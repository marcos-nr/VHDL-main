$date
  Tue Apr 23 20:11:56 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_tp2_1 $end
$var reg 1 ! clock $end
$var reg 1 " key $end
$var reg 1 # enable $end
$var reg 1 $ reset $end
$var reg 1 % led $end
$var reg 7 & segmentos[6:0] $end
$scope module uut $end
$var reg 1 ' clk $end
$var reg 1 ( key $end
$var reg 7 ) segmentos[6:0] $end
$var reg 1 * enable $end
$var reg 1 + reset $end
$var reg 1 , led $end
$var reg 1 - debounced_key $end
$var reg 4 . aux[3:0] $end
$scope module a $end
$var reg 1 / clk $end
$var reg 1 0 key $end
$var reg 1 1 debounced_key $end
$var reg 1 2 key_stable $end
$var reg 1 3 last_key $end
$upscope $end
$scope module b $end
$var reg 7 4 segmentos[6:0] $end
$var reg 4 5 bcd[3:0] $end
$var reg 1 6 enable $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
0"
1#
0$
0%
b1111110 &
0'
0(
b1111110 )
1*
0+
0,
U-
b0000 .
0/
00
U1
U2
U3
b1111110 4
b0000 5
16
#10000000
1!
1'
0-
1/
01
02
03
#20000000
0!
0'
0/
#30000000
1!
1'
1/
#40000000
0!
1"
0'
1(
0/
10
#50000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#60000000
0!
0'
0/
#70000000
1!
1'
1/
#80000000
0!
0'
0/
#90000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#100000000
0!
0'
0/
#110000000
1!
1'
1/
#120000000
0!
1"
0'
1(
0/
10
#130000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#140000000
0!
1$
0'
1+
0/
#150000000
1!
1'
1/
#160000000
0!
0'
0/
#170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#180000000
0!
0'
0/
#190000000
1!
1'
1/
#200000000
0!
0'
0/
#210000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#220000000
0!
0'
0/
#230000000
1!
1'
1/
#240000000
0!
0'
0/
#250000000
1!
1'
1/
#260000000
0!
0'
0/
#270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#280000000
0!
0'
0/
#290000000
1!
1'
1/
#300000000
0!
0'
0/
#310000000
1!
1'
1/
#320000000
0!
0'
0/
#330000000
1!
1'
1/
#340000000
0!
0'
0/
#350000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#360000000
0!
0'
0/
#370000000
1!
1'
1/
#380000000
0!
0'
0/
#390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#400000000
0!
0'
0/
#410000000
1!
1'
1/
#420000000
0!
0'
0/
#430000000
#440000000
1!
1'
1/
#450000000
0!
0'
0/
#460000000
1!
1'
1/
#470000000
0!
1"
0'
1(
0/
10
#480000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#490000000
0!
0'
0/
#500000000
1!
1'
1/
#510000000
0!
0'
0/
#520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#530000000
0!
0'
0/
#540000000
1!
1'
1/
#550000000
0!
1"
0'
1(
0/
10
#560000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#570000000
0!
1$
0'
1+
0/
#580000000
1!
1'
1/
#590000000
0!
0'
0/
#600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#610000000
0!
0'
0/
#620000000
1!
1'
1/
#630000000
0!
0'
0/
#640000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#650000000
0!
0'
0/
#660000000
1!
1'
1/
#670000000
0!
0'
0/
#680000000
1!
1'
1/
#690000000
0!
0'
0/
#700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#710000000
0!
0'
0/
#720000000
1!
1'
1/
#730000000
0!
0'
0/
#740000000
1!
1'
1/
#750000000
0!
0'
0/
#760000000
1!
1'
1/
#770000000
0!
0'
0/
#780000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#790000000
0!
0'
0/
#800000000
1!
1'
1/
#810000000
0!
0'
0/
#820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#830000000
0!
0'
0/
#840000000
1!
1'
1/
#850000000
0!
0'
0/
#860000000
#870000000
1!
1'
1/
#880000000
0!
0'
0/
#890000000
1!
1'
1/
#900000000
0!
1"
0'
1(
0/
10
#910000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#920000000
0!
0'
0/
#930000000
1!
1'
1/
#940000000
0!
0'
0/
#950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#960000000
0!
0'
0/
#970000000
1!
1'
1/
#980000000
0!
1"
0'
1(
0/
10
#990000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#1000000000
0!
1$
0'
1+
0/
#1010000000
1!
1'
1/
#1020000000
0!
0'
0/
#1030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#1040000000
0!
0'
0/
#1050000000
1!
1'
1/
#1060000000
0!
0'
0/
#1070000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#1080000000
0!
0'
0/
#1090000000
1!
1'
1/
#1100000000
0!
0'
0/
#1110000000
1!
1'
1/
#1120000000
0!
0'
0/
#1130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#1140000000
0!
0'
0/
#1150000000
1!
1'
1/
#1160000000
0!
0'
0/
#1170000000
1!
1'
1/
#1180000000
0!
0'
0/
#1190000000
1!
1'
1/
#1200000000
0!
0'
0/
#1210000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#1220000000
0!
0'
0/
#1230000000
1!
1'
1/
#1240000000
0!
0'
0/
#1250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#1260000000
0!
0'
0/
#1270000000
1!
1'
1/
#1280000000
0!
0'
0/
#1290000000
#1300000000
1!
1'
1/
#1310000000
0!
0'
0/
#1320000000
1!
1'
1/
#1330000000
0!
1"
0'
1(
0/
10
#1340000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#1350000000
0!
0'
0/
#1360000000
1!
1'
1/
#1370000000
0!
0'
0/
#1380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#1390000000
0!
0'
0/
#1400000000
1!
1'
1/
#1410000000
0!
1"
0'
1(
0/
10
#1420000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#1430000000
0!
1$
0'
1+
0/
#1440000000
1!
1'
1/
#1450000000
0!
0'
0/
#1460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#1470000000
0!
0'
0/
#1480000000
1!
1'
1/
#1490000000
0!
0'
0/
#1500000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#1510000000
0!
0'
0/
#1520000000
1!
1'
1/
#1530000000
0!
0'
0/
#1540000000
1!
1'
1/
#1550000000
0!
0'
0/
#1560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#1570000000
0!
0'
0/
#1580000000
1!
1'
1/
#1590000000
0!
0'
0/
#1600000000
1!
1'
1/
#1610000000
0!
0'
0/
#1620000000
1!
1'
1/
#1630000000
0!
0'
0/
#1640000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#1650000000
0!
0'
0/
#1660000000
1!
1'
1/
#1670000000
0!
0'
0/
#1680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#1690000000
0!
0'
0/
#1700000000
1!
1'
1/
#1710000000
0!
0'
0/
#1720000000
#1730000000
1!
1'
1/
#1740000000
0!
0'
0/
#1750000000
1!
1'
1/
#1760000000
0!
1"
0'
1(
0/
10
#1770000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#1780000000
0!
0'
0/
#1790000000
1!
1'
1/
#1800000000
0!
0'
0/
#1810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#1820000000
0!
0'
0/
#1830000000
1!
1'
1/
#1840000000
0!
1"
0'
1(
0/
10
#1850000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#1860000000
0!
1$
0'
1+
0/
#1870000000
1!
1'
1/
#1880000000
0!
0'
0/
#1890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#1900000000
0!
0'
0/
#1910000000
1!
1'
1/
#1920000000
0!
0'
0/
#1930000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#1940000000
0!
0'
0/
#1950000000
1!
1'
1/
#1960000000
0!
0'
0/
#1970000000
1!
1'
1/
#1980000000
0!
0'
0/
#1990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#2000000000
0!
0'
0/
#2010000000
1!
1'
1/
#2020000000
0!
0'
0/
#2030000000
1!
1'
1/
#2040000000
0!
0'
0/
#2050000000
1!
1'
1/
#2060000000
0!
0'
0/
#2070000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#2080000000
0!
0'
0/
#2090000000
1!
1'
1/
#2100000000
0!
0'
0/
#2110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#2120000000
0!
0'
0/
#2130000000
1!
1'
1/
#2140000000
0!
0'
0/
#2150000000
#2160000000
1!
1'
1/
#2170000000
0!
0'
0/
#2180000000
1!
1'
1/
#2190000000
0!
1"
0'
1(
0/
10
#2200000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#2210000000
0!
0'
0/
#2220000000
1!
1'
1/
#2230000000
0!
0'
0/
#2240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#2250000000
0!
0'
0/
#2260000000
1!
1'
1/
#2270000000
0!
1"
0'
1(
0/
10
#2280000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#2290000000
0!
1$
0'
1+
0/
#2300000000
1!
1'
1/
#2310000000
0!
0'
0/
#2320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#2330000000
0!
0'
0/
#2340000000
1!
1'
1/
#2350000000
0!
0'
0/
#2360000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#2370000000
0!
0'
0/
#2380000000
1!
1'
1/
#2390000000
0!
0'
0/
#2400000000
1!
1'
1/
#2410000000
0!
0'
0/
#2420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#2430000000
0!
0'
0/
#2440000000
1!
1'
1/
#2450000000
0!
0'
0/
#2460000000
1!
1'
1/
#2470000000
0!
0'
0/
#2480000000
1!
1'
1/
#2490000000
0!
0'
0/
#2500000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#2510000000
0!
0'
0/
#2520000000
1!
1'
1/
#2530000000
0!
0'
0/
#2540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#2550000000
0!
0'
0/
#2560000000
1!
1'
1/
#2570000000
0!
0'
0/
#2580000000
#2590000000
1!
1'
1/
#2600000000
0!
0'
0/
#2610000000
1!
1'
1/
#2620000000
0!
1"
0'
1(
0/
10
#2630000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#2640000000
0!
0'
0/
#2650000000
1!
1'
1/
#2660000000
0!
0'
0/
#2670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#2680000000
0!
0'
0/
#2690000000
1!
1'
1/
#2700000000
0!
1"
0'
1(
0/
10
#2710000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#2720000000
0!
1$
0'
1+
0/
#2730000000
1!
1'
1/
#2740000000
0!
0'
0/
#2750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#2760000000
0!
0'
0/
#2770000000
1!
1'
1/
#2780000000
0!
0'
0/
#2790000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#2800000000
0!
0'
0/
#2810000000
1!
1'
1/
#2820000000
0!
0'
0/
#2830000000
1!
1'
1/
#2840000000
0!
0'
0/
#2850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#2860000000
0!
0'
0/
#2870000000
1!
1'
1/
#2880000000
0!
0'
0/
#2890000000
1!
1'
1/
#2900000000
0!
0'
0/
#2910000000
1!
1'
1/
#2920000000
0!
0'
0/
#2930000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#2940000000
0!
0'
0/
#2950000000
1!
1'
1/
#2960000000
0!
0'
0/
#2970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#2980000000
0!
0'
0/
#2990000000
1!
1'
1/
#3000000000
0!
0'
0/
#3010000000
#3020000000
1!
1'
1/
#3030000000
0!
0'
0/
#3040000000
1!
1'
1/
#3050000000
0!
1"
0'
1(
0/
10
#3060000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#3070000000
0!
0'
0/
#3080000000
1!
1'
1/
#3090000000
0!
0'
0/
#3100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#3110000000
0!
0'
0/
#3120000000
1!
1'
1/
#3130000000
0!
1"
0'
1(
0/
10
#3140000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#3150000000
0!
1$
0'
1+
0/
#3160000000
1!
1'
1/
#3170000000
0!
0'
0/
#3180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#3190000000
0!
0'
0/
#3200000000
1!
1'
1/
#3210000000
0!
0'
0/
#3220000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#3230000000
0!
0'
0/
#3240000000
1!
1'
1/
#3250000000
0!
0'
0/
#3260000000
1!
1'
1/
#3270000000
0!
0'
0/
#3280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#3290000000
0!
0'
0/
#3300000000
1!
1'
1/
#3310000000
0!
0'
0/
#3320000000
1!
1'
1/
#3330000000
0!
0'
0/
#3340000000
1!
1'
1/
#3350000000
0!
0'
0/
#3360000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#3370000000
0!
0'
0/
#3380000000
1!
1'
1/
#3390000000
0!
0'
0/
#3400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#3410000000
0!
0'
0/
#3420000000
1!
1'
1/
#3430000000
0!
0'
0/
#3440000000
#3450000000
1!
1'
1/
#3460000000
0!
0'
0/
#3470000000
1!
1'
1/
#3480000000
0!
1"
0'
1(
0/
10
#3490000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#3500000000
0!
0'
0/
#3510000000
1!
1'
1/
#3520000000
0!
0'
0/
#3530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#3540000000
0!
0'
0/
#3550000000
1!
1'
1/
#3560000000
0!
1"
0'
1(
0/
10
#3570000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#3580000000
0!
1$
0'
1+
0/
#3590000000
1!
1'
1/
#3600000000
0!
0'
0/
#3610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#3620000000
0!
0'
0/
#3630000000
1!
1'
1/
#3640000000
0!
0'
0/
#3650000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#3660000000
0!
0'
0/
#3670000000
1!
1'
1/
#3680000000
0!
0'
0/
#3690000000
1!
1'
1/
#3700000000
0!
0'
0/
#3710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#3720000000
0!
0'
0/
#3730000000
1!
1'
1/
#3740000000
0!
0'
0/
#3750000000
1!
1'
1/
#3760000000
0!
0'
0/
#3770000000
1!
1'
1/
#3780000000
0!
0'
0/
#3790000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#3800000000
0!
0'
0/
#3810000000
1!
1'
1/
#3820000000
0!
0'
0/
#3830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#3840000000
0!
0'
0/
#3850000000
1!
1'
1/
#3860000000
0!
0'
0/
#3870000000
#3880000000
1!
1'
1/
#3890000000
0!
0'
0/
#3900000000
1!
1'
1/
#3910000000
0!
1"
0'
1(
0/
10
#3920000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#3930000000
0!
0'
0/
#3940000000
1!
1'
1/
#3950000000
0!
0'
0/
#3960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#3970000000
0!
0'
0/
#3980000000
1!
1'
1/
#3990000000
0!
1"
0'
1(
0/
10
#4000000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#4010000000
0!
1$
0'
1+
0/
#4020000000
1!
1'
1/
#4030000000
0!
0'
0/
#4040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#4050000000
0!
0'
0/
#4060000000
1!
1'
1/
#4070000000
0!
0'
0/
#4080000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#4090000000
0!
0'
0/
#4100000000
1!
1'
1/
#4110000000
0!
0'
0/
#4120000000
1!
1'
1/
#4130000000
0!
0'
0/
#4140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#4150000000
0!
0'
0/
#4160000000
1!
1'
1/
#4170000000
0!
0'
0/
#4180000000
1!
1'
1/
#4190000000
0!
0'
0/
#4200000000
1!
1'
1/
#4210000000
0!
0'
0/
#4220000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#4230000000
0!
0'
0/
#4240000000
1!
1'
1/
#4250000000
0!
0'
0/
#4260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#4270000000
0!
0'
0/
#4280000000
1!
1'
1/
#4290000000
0!
0'
0/
#4300000000
#4310000000
1!
1'
1/
#4320000000
0!
0'
0/
#4330000000
1!
1'
1/
#4340000000
0!
1"
0'
1(
0/
10
#4350000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#4360000000
0!
0'
0/
#4370000000
1!
1'
1/
#4380000000
0!
0'
0/
#4390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#4400000000
0!
0'
0/
#4410000000
1!
1'
1/
#4420000000
0!
1"
0'
1(
0/
10
#4430000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#4440000000
0!
1$
0'
1+
0/
#4450000000
1!
1'
1/
#4460000000
0!
0'
0/
#4470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#4480000000
0!
0'
0/
#4490000000
1!
1'
1/
#4500000000
0!
0'
0/
#4510000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#4520000000
0!
0'
0/
#4530000000
1!
1'
1/
#4540000000
0!
0'
0/
#4550000000
1!
1'
1/
#4560000000
0!
0'
0/
#4570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#4580000000
0!
0'
0/
#4590000000
1!
1'
1/
#4600000000
0!
0'
0/
#4610000000
1!
1'
1/
#4620000000
0!
0'
0/
#4630000000
1!
1'
1/
#4640000000
0!
0'
0/
#4650000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#4660000000
0!
0'
0/
#4670000000
1!
1'
1/
#4680000000
0!
0'
0/
#4690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#4700000000
0!
0'
0/
#4710000000
1!
1'
1/
#4720000000
0!
0'
0/
#4730000000
#4740000000
1!
1'
1/
#4750000000
0!
0'
0/
#4760000000
1!
1'
1/
#4770000000
0!
1"
0'
1(
0/
10
#4780000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#4790000000
0!
0'
0/
#4800000000
1!
1'
1/
#4810000000
0!
0'
0/
#4820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#4830000000
0!
0'
0/
#4840000000
1!
1'
1/
#4850000000
0!
1"
0'
1(
0/
10
#4860000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#4870000000
0!
1$
0'
1+
0/
#4880000000
1!
1'
1/
#4890000000
0!
0'
0/
#4900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#4910000000
0!
0'
0/
#4920000000
1!
1'
1/
#4930000000
0!
0'
0/
#4940000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#4950000000
0!
0'
0/
#4960000000
1!
1'
1/
#4970000000
0!
0'
0/
#4980000000
1!
1'
1/
#4990000000
0!
0'
0/
#5000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#5010000000
0!
0'
0/
#5020000000
1!
1'
1/
#5030000000
0!
0'
0/
#5040000000
1!
1'
1/
#5050000000
0!
0'
0/
#5060000000
1!
1'
1/
#5070000000
0!
0'
0/
#5080000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#5090000000
0!
0'
0/
#5100000000
1!
1'
1/
#5110000000
0!
0'
0/
#5120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#5130000000
0!
0'
0/
#5140000000
1!
1'
1/
#5150000000
0!
0'
0/
#5160000000
#5170000000
1!
1'
1/
#5180000000
0!
0'
0/
#5190000000
1!
1'
1/
#5200000000
0!
1"
0'
1(
0/
10
#5210000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#5220000000
0!
0'
0/
#5230000000
1!
1'
1/
#5240000000
0!
0'
0/
#5250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#5260000000
0!
0'
0/
#5270000000
1!
1'
1/
#5280000000
0!
1"
0'
1(
0/
10
#5290000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#5300000000
0!
1$
0'
1+
0/
#5310000000
1!
1'
1/
#5320000000
0!
0'
0/
#5330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#5340000000
0!
0'
0/
#5350000000
1!
1'
1/
#5360000000
0!
0'
0/
#5370000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#5380000000
0!
0'
0/
#5390000000
1!
1'
1/
#5400000000
0!
0'
0/
#5410000000
1!
1'
1/
#5420000000
0!
0'
0/
#5430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#5440000000
0!
0'
0/
#5450000000
1!
1'
1/
#5460000000
0!
0'
0/
#5470000000
1!
1'
1/
#5480000000
0!
0'
0/
#5490000000
1!
1'
1/
#5500000000
0!
0'
0/
#5510000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#5520000000
0!
0'
0/
#5530000000
1!
1'
1/
#5540000000
0!
0'
0/
#5550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#5560000000
0!
0'
0/
#5570000000
1!
1'
1/
#5580000000
0!
0'
0/
#5590000000
#5600000000
1!
1'
1/
#5610000000
0!
0'
0/
#5620000000
1!
1'
1/
#5630000000
0!
1"
0'
1(
0/
10
#5640000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#5650000000
0!
0'
0/
#5660000000
1!
1'
1/
#5670000000
0!
0'
0/
#5680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#5690000000
0!
0'
0/
#5700000000
1!
1'
1/
#5710000000
0!
1"
0'
1(
0/
10
#5720000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#5730000000
0!
1$
0'
1+
0/
#5740000000
1!
1'
1/
#5750000000
0!
0'
0/
#5760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#5770000000
0!
0'
0/
#5780000000
1!
1'
1/
#5790000000
0!
0'
0/
#5800000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#5810000000
0!
0'
0/
#5820000000
1!
1'
1/
#5830000000
0!
0'
0/
#5840000000
1!
1'
1/
#5850000000
0!
0'
0/
#5860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#5870000000
0!
0'
0/
#5880000000
1!
1'
1/
#5890000000
0!
0'
0/
#5900000000
1!
1'
1/
#5910000000
0!
0'
0/
#5920000000
1!
1'
1/
#5930000000
0!
0'
0/
#5940000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#5950000000
0!
0'
0/
#5960000000
1!
1'
1/
#5970000000
0!
0'
0/
#5980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#5990000000
0!
0'
0/
#6000000000
1!
1'
1/
#6010000000
0!
0'
0/
#6020000000
#6030000000
1!
1'
1/
#6040000000
0!
0'
0/
#6050000000
1!
1'
1/
#6060000000
0!
1"
0'
1(
0/
10
#6070000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#6080000000
0!
0'
0/
#6090000000
1!
1'
1/
#6100000000
0!
0'
0/
#6110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#6120000000
0!
0'
0/
#6130000000
1!
1'
1/
#6140000000
0!
1"
0'
1(
0/
10
#6150000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#6160000000
0!
1$
0'
1+
0/
#6170000000
1!
1'
1/
#6180000000
0!
0'
0/
#6190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#6200000000
0!
0'
0/
#6210000000
1!
1'
1/
#6220000000
0!
0'
0/
#6230000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#6240000000
0!
0'
0/
#6250000000
1!
1'
1/
#6260000000
0!
0'
0/
#6270000000
1!
1'
1/
#6280000000
0!
0'
0/
#6290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#6300000000
0!
0'
0/
#6310000000
1!
1'
1/
#6320000000
0!
0'
0/
#6330000000
1!
1'
1/
#6340000000
0!
0'
0/
#6350000000
1!
1'
1/
#6360000000
0!
0'
0/
#6370000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#6380000000
0!
0'
0/
#6390000000
1!
1'
1/
#6400000000
0!
0'
0/
#6410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#6420000000
0!
0'
0/
#6430000000
1!
1'
1/
#6440000000
0!
0'
0/
#6450000000
#6460000000
1!
1'
1/
#6470000000
0!
0'
0/
#6480000000
1!
1'
1/
#6490000000
0!
1"
0'
1(
0/
10
#6500000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#6510000000
0!
0'
0/
#6520000000
1!
1'
1/
#6530000000
0!
0'
0/
#6540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#6550000000
0!
0'
0/
#6560000000
1!
1'
1/
#6570000000
0!
1"
0'
1(
0/
10
#6580000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#6590000000
0!
1$
0'
1+
0/
#6600000000
1!
1'
1/
#6610000000
0!
0'
0/
#6620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#6630000000
0!
0'
0/
#6640000000
1!
1'
1/
#6650000000
0!
0'
0/
#6660000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#6670000000
0!
0'
0/
#6680000000
1!
1'
1/
#6690000000
0!
0'
0/
#6700000000
1!
1'
1/
#6710000000
0!
0'
0/
#6720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#6730000000
0!
0'
0/
#6740000000
1!
1'
1/
#6750000000
0!
0'
0/
#6760000000
1!
1'
1/
#6770000000
0!
0'
0/
#6780000000
1!
1'
1/
#6790000000
0!
0'
0/
#6800000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#6810000000
0!
0'
0/
#6820000000
1!
1'
1/
#6830000000
0!
0'
0/
#6840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#6850000000
0!
0'
0/
#6860000000
1!
1'
1/
#6870000000
0!
0'
0/
#6880000000
#6890000000
1!
1'
1/
#6900000000
0!
0'
0/
#6910000000
1!
1'
1/
#6920000000
0!
1"
0'
1(
0/
10
#6930000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#6940000000
0!
0'
0/
#6950000000
1!
1'
1/
#6960000000
0!
0'
0/
#6970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#6980000000
0!
0'
0/
#6990000000
1!
1'
1/
#7000000000
0!
1"
0'
1(
0/
10
#7010000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#7020000000
0!
1$
0'
1+
0/
#7030000000
1!
1'
1/
#7040000000
0!
0'
0/
#7050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#7060000000
0!
0'
0/
#7070000000
1!
1'
1/
#7080000000
0!
0'
0/
#7090000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#7100000000
0!
0'
0/
#7110000000
1!
1'
1/
#7120000000
0!
0'
0/
#7130000000
1!
1'
1/
#7140000000
0!
0'
0/
#7150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#7160000000
0!
0'
0/
#7170000000
1!
1'
1/
#7180000000
0!
0'
0/
#7190000000
1!
1'
1/
#7200000000
0!
0'
0/
#7210000000
1!
1'
1/
#7220000000
0!
0'
0/
#7230000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#7240000000
0!
0'
0/
#7250000000
1!
1'
1/
#7260000000
0!
0'
0/
#7270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#7280000000
0!
0'
0/
#7290000000
1!
1'
1/
#7300000000
0!
0'
0/
#7310000000
#7320000000
1!
1'
1/
#7330000000
0!
0'
0/
#7340000000
1!
1'
1/
#7350000000
0!
1"
0'
1(
0/
10
#7360000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#7370000000
0!
0'
0/
#7380000000
1!
1'
1/
#7390000000
0!
0'
0/
#7400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#7410000000
0!
0'
0/
#7420000000
1!
1'
1/
#7430000000
0!
1"
0'
1(
0/
10
#7440000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#7450000000
0!
1$
0'
1+
0/
#7460000000
1!
1'
1/
#7470000000
0!
0'
0/
#7480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#7490000000
0!
0'
0/
#7500000000
1!
1'
1/
#7510000000
0!
0'
0/
#7520000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#7530000000
0!
0'
0/
#7540000000
1!
1'
1/
#7550000000
0!
0'
0/
#7560000000
1!
1'
1/
#7570000000
0!
0'
0/
#7580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#7590000000
0!
0'
0/
#7600000000
1!
1'
1/
#7610000000
0!
0'
0/
#7620000000
1!
1'
1/
#7630000000
0!
0'
0/
#7640000000
1!
1'
1/
#7650000000
0!
0'
0/
#7660000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#7670000000
0!
0'
0/
#7680000000
1!
1'
1/
#7690000000
0!
0'
0/
#7700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#7710000000
0!
0'
0/
#7720000000
1!
1'
1/
#7730000000
0!
0'
0/
#7740000000
#7750000000
1!
1'
1/
#7760000000
0!
0'
0/
#7770000000
1!
1'
1/
#7780000000
0!
1"
0'
1(
0/
10
#7790000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#7800000000
0!
0'
0/
#7810000000
1!
1'
1/
#7820000000
0!
0'
0/
#7830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#7840000000
0!
0'
0/
#7850000000
1!
1'
1/
#7860000000
0!
1"
0'
1(
0/
10
#7870000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#7880000000
0!
1$
0'
1+
0/
#7890000000
1!
1'
1/
#7900000000
0!
0'
0/
#7910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#7920000000
0!
0'
0/
#7930000000
1!
1'
1/
#7940000000
0!
0'
0/
#7950000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#7960000000
0!
0'
0/
#7970000000
1!
1'
1/
#7980000000
0!
0'
0/
#7990000000
1!
1'
1/
#8000000000
0!
0'
0/
#8010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#8020000000
0!
0'
0/
#8030000000
1!
1'
1/
#8040000000
0!
0'
0/
#8050000000
1!
1'
1/
#8060000000
0!
0'
0/
#8070000000
1!
1'
1/
#8080000000
0!
0'
0/
#8090000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#8100000000
0!
0'
0/
#8110000000
1!
1'
1/
#8120000000
0!
0'
0/
#8130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#8140000000
0!
0'
0/
#8150000000
1!
1'
1/
#8160000000
0!
0'
0/
#8170000000
#8180000000
1!
1'
1/
#8190000000
0!
0'
0/
#8200000000
1!
1'
1/
#8210000000
0!
1"
0'
1(
0/
10
#8220000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#8230000000
0!
0'
0/
#8240000000
1!
1'
1/
#8250000000
0!
0'
0/
#8260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#8270000000
0!
0'
0/
#8280000000
1!
1'
1/
#8290000000
0!
1"
0'
1(
0/
10
#8300000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#8310000000
0!
1$
0'
1+
0/
#8320000000
1!
1'
1/
#8330000000
0!
0'
0/
#8340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#8350000000
0!
0'
0/
#8360000000
1!
1'
1/
#8370000000
0!
0'
0/
#8380000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#8390000000
0!
0'
0/
#8400000000
1!
1'
1/
#8410000000
0!
0'
0/
#8420000000
1!
1'
1/
#8430000000
0!
0'
0/
#8440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#8450000000
0!
0'
0/
#8460000000
1!
1'
1/
#8470000000
0!
0'
0/
#8480000000
1!
1'
1/
#8490000000
0!
0'
0/
#8500000000
1!
1'
1/
#8510000000
0!
0'
0/
#8520000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#8530000000
0!
0'
0/
#8540000000
1!
1'
1/
#8550000000
0!
0'
0/
#8560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#8570000000
0!
0'
0/
#8580000000
1!
1'
1/
#8590000000
0!
0'
0/
#8600000000
#8610000000
1!
1'
1/
#8620000000
0!
0'
0/
#8630000000
1!
1'
1/
#8640000000
0!
1"
0'
1(
0/
10
#8650000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#8660000000
0!
0'
0/
#8670000000
1!
1'
1/
#8680000000
0!
0'
0/
#8690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#8700000000
0!
0'
0/
#8710000000
1!
1'
1/
#8720000000
0!
1"
0'
1(
0/
10
#8730000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#8740000000
0!
1$
0'
1+
0/
#8750000000
1!
1'
1/
#8760000000
0!
0'
0/
#8770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#8780000000
0!
0'
0/
#8790000000
1!
1'
1/
#8800000000
0!
0'
0/
#8810000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#8820000000
0!
0'
0/
#8830000000
1!
1'
1/
#8840000000
0!
0'
0/
#8850000000
1!
1'
1/
#8860000000
0!
0'
0/
#8870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#8880000000
0!
0'
0/
#8890000000
1!
1'
1/
#8900000000
0!
0'
0/
#8910000000
1!
1'
1/
#8920000000
0!
0'
0/
#8930000000
1!
1'
1/
#8940000000
0!
0'
0/
#8950000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#8960000000
0!
0'
0/
#8970000000
1!
1'
1/
#8980000000
0!
0'
0/
#8990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#9000000000
0!
0'
0/
#9010000000
1!
1'
1/
#9020000000
0!
0'
0/
#9030000000
#9040000000
1!
1'
1/
#9050000000
0!
0'
0/
#9060000000
1!
1'
1/
#9070000000
0!
1"
0'
1(
0/
10
#9080000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#9090000000
0!
0'
0/
#9100000000
1!
1'
1/
#9110000000
0!
0'
0/
#9120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#9130000000
0!
0'
0/
#9140000000
1!
1'
1/
#9150000000
0!
1"
0'
1(
0/
10
#9160000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#9170000000
0!
1$
0'
1+
0/
#9180000000
1!
1'
1/
#9190000000
0!
0'
0/
#9200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#9210000000
0!
0'
0/
#9220000000
1!
1'
1/
#9230000000
0!
0'
0/
#9240000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#9250000000
0!
0'
0/
#9260000000
1!
1'
1/
#9270000000
0!
0'
0/
#9280000000
1!
1'
1/
#9290000000
0!
0'
0/
#9300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#9310000000
0!
0'
0/
#9320000000
1!
1'
1/
#9330000000
0!
0'
0/
#9340000000
1!
1'
1/
#9350000000
0!
0'
0/
#9360000000
1!
1'
1/
#9370000000
0!
0'
0/
#9380000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#9390000000
0!
0'
0/
#9400000000
1!
1'
1/
#9410000000
0!
0'
0/
#9420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#9430000000
0!
0'
0/
#9440000000
1!
1'
1/
#9450000000
0!
0'
0/
#9460000000
#9470000000
1!
1'
1/
#9480000000
0!
0'
0/
#9490000000
1!
1'
1/
#9500000000
0!
1"
0'
1(
0/
10
#9510000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#9520000000
0!
0'
0/
#9530000000
1!
1'
1/
#9540000000
0!
0'
0/
#9550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#9560000000
0!
0'
0/
#9570000000
1!
1'
1/
#9580000000
0!
1"
0'
1(
0/
10
#9590000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#9600000000
0!
1$
0'
1+
0/
#9610000000
1!
1'
1/
#9620000000
0!
0'
0/
#9630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#9640000000
0!
0'
0/
#9650000000
1!
1'
1/
#9660000000
0!
0'
0/
#9670000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#9680000000
0!
0'
0/
#9690000000
1!
1'
1/
#9700000000
0!
0'
0/
#9710000000
1!
1'
1/
#9720000000
0!
0'
0/
#9730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#9740000000
0!
0'
0/
#9750000000
1!
1'
1/
#9760000000
0!
0'
0/
#9770000000
1!
1'
1/
#9780000000
0!
0'
0/
#9790000000
1!
1'
1/
#9800000000
0!
0'
0/
#9810000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#9820000000
0!
0'
0/
#9830000000
1!
1'
1/
#9840000000
0!
0'
0/
#9850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#9860000000
0!
0'
0/
#9870000000
1!
1'
1/
#9880000000
0!
0'
0/
#9890000000
#9900000000
1!
1'
1/
#9910000000
0!
0'
0/
#9920000000
1!
1'
1/
#9930000000
0!
1"
0'
1(
0/
10
#9940000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#9950000000
0!
0'
0/
#9960000000
1!
1'
1/
#9970000000
0!
0'
0/
#9980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#9990000000
0!
0'
0/
#10000000000
1!
1'
1/
#10010000000
0!
1"
0'
1(
0/
10
#10020000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#10030000000
0!
1$
0'
1+
0/
#10040000000
1!
1'
1/
#10050000000
0!
0'
0/
#10060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#10070000000
0!
0'
0/
#10080000000
1!
1'
1/
#10090000000
0!
0'
0/
#10100000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#10110000000
0!
0'
0/
#10120000000
1!
1'
1/
#10130000000
0!
0'
0/
#10140000000
1!
1'
1/
#10150000000
0!
0'
0/
#10160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#10170000000
0!
0'
0/
#10180000000
1!
1'
1/
#10190000000
0!
0'
0/
#10200000000
1!
1'
1/
#10210000000
0!
0'
0/
#10220000000
1!
1'
1/
#10230000000
0!
0'
0/
#10240000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#10250000000
0!
0'
0/
#10260000000
1!
1'
1/
#10270000000
0!
0'
0/
#10280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#10290000000
0!
0'
0/
#10300000000
1!
1'
1/
#10310000000
0!
0'
0/
#10320000000
#10330000000
1!
1'
1/
#10340000000
0!
0'
0/
#10350000000
1!
1'
1/
#10360000000
0!
1"
0'
1(
0/
10
#10370000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#10380000000
0!
0'
0/
#10390000000
1!
1'
1/
#10400000000
0!
0'
0/
#10410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#10420000000
0!
0'
0/
#10430000000
1!
1'
1/
#10440000000
0!
1"
0'
1(
0/
10
#10450000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#10460000000
0!
1$
0'
1+
0/
#10470000000
1!
1'
1/
#10480000000
0!
0'
0/
#10490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#10500000000
0!
0'
0/
#10510000000
1!
1'
1/
#10520000000
0!
0'
0/
#10530000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#10540000000
0!
0'
0/
#10550000000
1!
1'
1/
#10560000000
0!
0'
0/
#10570000000
1!
1'
1/
#10580000000
0!
0'
0/
#10590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#10600000000
0!
0'
0/
#10610000000
1!
1'
1/
#10620000000
0!
0'
0/
#10630000000
1!
1'
1/
#10640000000
0!
0'
0/
#10650000000
1!
1'
1/
#10660000000
0!
0'
0/
#10670000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#10680000000
0!
0'
0/
#10690000000
1!
1'
1/
#10700000000
0!
0'
0/
#10710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#10720000000
0!
0'
0/
#10730000000
1!
1'
1/
#10740000000
0!
0'
0/
#10750000000
#10760000000
1!
1'
1/
#10770000000
0!
0'
0/
#10780000000
1!
1'
1/
#10790000000
0!
1"
0'
1(
0/
10
#10800000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#10810000000
0!
0'
0/
#10820000000
1!
1'
1/
#10830000000
0!
0'
0/
#10840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#10850000000
0!
0'
0/
#10860000000
1!
1'
1/
#10870000000
0!
1"
0'
1(
0/
10
#10880000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#10890000000
0!
1$
0'
1+
0/
#10900000000
1!
1'
1/
#10910000000
0!
0'
0/
#10920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#10930000000
0!
0'
0/
#10940000000
1!
1'
1/
#10950000000
0!
0'
0/
#10960000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#10970000000
0!
0'
0/
#10980000000
1!
1'
1/
#10990000000
0!
0'
0/
#11000000000
1!
1'
1/
#11010000000
0!
0'
0/
#11020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#11030000000
0!
0'
0/
#11040000000
1!
1'
1/
#11050000000
0!
0'
0/
#11060000000
1!
1'
1/
#11070000000
0!
0'
0/
#11080000000
1!
1'
1/
#11090000000
0!
0'
0/
#11100000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#11110000000
0!
0'
0/
#11120000000
1!
1'
1/
#11130000000
0!
0'
0/
#11140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#11150000000
0!
0'
0/
#11160000000
1!
1'
1/
#11170000000
0!
0'
0/
#11180000000
#11190000000
1!
1'
1/
#11200000000
0!
0'
0/
#11210000000
1!
1'
1/
#11220000000
0!
1"
0'
1(
0/
10
#11230000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#11240000000
0!
0'
0/
#11250000000
1!
1'
1/
#11260000000
0!
0'
0/
#11270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#11280000000
0!
0'
0/
#11290000000
1!
1'
1/
#11300000000
0!
1"
0'
1(
0/
10
#11310000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#11320000000
0!
1$
0'
1+
0/
#11330000000
1!
1'
1/
#11340000000
0!
0'
0/
#11350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#11360000000
0!
0'
0/
#11370000000
1!
1'
1/
#11380000000
0!
0'
0/
#11390000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#11400000000
0!
0'
0/
#11410000000
1!
1'
1/
#11420000000
0!
0'
0/
#11430000000
1!
1'
1/
#11440000000
0!
0'
0/
#11450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#11460000000
0!
0'
0/
#11470000000
1!
1'
1/
#11480000000
0!
0'
0/
#11490000000
1!
1'
1/
#11500000000
0!
0'
0/
#11510000000
1!
1'
1/
#11520000000
0!
0'
0/
#11530000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#11540000000
0!
0'
0/
#11550000000
1!
1'
1/
#11560000000
0!
0'
0/
#11570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#11580000000
0!
0'
0/
#11590000000
1!
1'
1/
#11600000000
0!
0'
0/
#11610000000
#11620000000
1!
1'
1/
#11630000000
0!
0'
0/
#11640000000
1!
1'
1/
#11650000000
0!
1"
0'
1(
0/
10
#11660000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#11670000000
0!
0'
0/
#11680000000
1!
1'
1/
#11690000000
0!
0'
0/
#11700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#11710000000
0!
0'
0/
#11720000000
1!
1'
1/
#11730000000
0!
1"
0'
1(
0/
10
#11740000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#11750000000
0!
1$
0'
1+
0/
#11760000000
1!
1'
1/
#11770000000
0!
0'
0/
#11780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#11790000000
0!
0'
0/
#11800000000
1!
1'
1/
#11810000000
0!
0'
0/
#11820000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#11830000000
0!
0'
0/
#11840000000
1!
1'
1/
#11850000000
0!
0'
0/
#11860000000
1!
1'
1/
#11870000000
0!
0'
0/
#11880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#11890000000
0!
0'
0/
#11900000000
1!
1'
1/
#11910000000
0!
0'
0/
#11920000000
1!
1'
1/
#11930000000
0!
0'
0/
#11940000000
1!
1'
1/
#11950000000
0!
0'
0/
#11960000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#11970000000
0!
0'
0/
#11980000000
1!
1'
1/
#11990000000
0!
0'
0/
#12000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#12010000000
0!
0'
0/
#12020000000
1!
1'
1/
#12030000000
0!
0'
0/
#12040000000
#12050000000
1!
1'
1/
#12060000000
0!
0'
0/
#12070000000
1!
1'
1/
#12080000000
0!
1"
0'
1(
0/
10
#12090000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#12100000000
0!
0'
0/
#12110000000
1!
1'
1/
#12120000000
0!
0'
0/
#12130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#12140000000
0!
0'
0/
#12150000000
1!
1'
1/
#12160000000
0!
1"
0'
1(
0/
10
#12170000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#12180000000
0!
1$
0'
1+
0/
#12190000000
1!
1'
1/
#12200000000
0!
0'
0/
#12210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#12220000000
0!
0'
0/
#12230000000
1!
1'
1/
#12240000000
0!
0'
0/
#12250000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#12260000000
0!
0'
0/
#12270000000
1!
1'
1/
#12280000000
0!
0'
0/
#12290000000
1!
1'
1/
#12300000000
0!
0'
0/
#12310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#12320000000
0!
0'
0/
#12330000000
1!
1'
1/
#12340000000
0!
0'
0/
#12350000000
1!
1'
1/
#12360000000
0!
0'
0/
#12370000000
1!
1'
1/
#12380000000
0!
0'
0/
#12390000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#12400000000
0!
0'
0/
#12410000000
1!
1'
1/
#12420000000
0!
0'
0/
#12430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#12440000000
0!
0'
0/
#12450000000
1!
1'
1/
#12460000000
0!
0'
0/
#12470000000
#12480000000
1!
1'
1/
#12490000000
0!
0'
0/
#12500000000
1!
1'
1/
#12510000000
0!
1"
0'
1(
0/
10
#12520000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#12530000000
0!
0'
0/
#12540000000
1!
1'
1/
#12550000000
0!
0'
0/
#12560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#12570000000
0!
0'
0/
#12580000000
1!
1'
1/
#12590000000
0!
1"
0'
1(
0/
10
#12600000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#12610000000
0!
1$
0'
1+
0/
#12620000000
1!
1'
1/
#12630000000
0!
0'
0/
#12640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#12650000000
0!
0'
0/
#12660000000
1!
1'
1/
#12670000000
0!
0'
0/
#12680000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#12690000000
0!
0'
0/
#12700000000
1!
1'
1/
#12710000000
0!
0'
0/
#12720000000
1!
1'
1/
#12730000000
0!
0'
0/
#12740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#12750000000
0!
0'
0/
#12760000000
1!
1'
1/
#12770000000
0!
0'
0/
#12780000000
1!
1'
1/
#12790000000
0!
0'
0/
#12800000000
1!
1'
1/
#12810000000
0!
0'
0/
#12820000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#12830000000
0!
0'
0/
#12840000000
1!
1'
1/
#12850000000
0!
0'
0/
#12860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#12870000000
0!
0'
0/
#12880000000
1!
1'
1/
#12890000000
0!
0'
0/
#12900000000
#12910000000
1!
1'
1/
#12920000000
0!
0'
0/
#12930000000
1!
1'
1/
#12940000000
0!
1"
0'
1(
0/
10
#12950000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#12960000000
0!
0'
0/
#12970000000
1!
1'
1/
#12980000000
0!
0'
0/
#12990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#13000000000
0!
0'
0/
#13010000000
1!
1'
1/
#13020000000
0!
1"
0'
1(
0/
10
#13030000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#13040000000
0!
1$
0'
1+
0/
#13050000000
1!
1'
1/
#13060000000
0!
0'
0/
#13070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#13080000000
0!
0'
0/
#13090000000
1!
1'
1/
#13100000000
0!
0'
0/
#13110000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#13120000000
0!
0'
0/
#13130000000
1!
1'
1/
#13140000000
0!
0'
0/
#13150000000
1!
1'
1/
#13160000000
0!
0'
0/
#13170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#13180000000
0!
0'
0/
#13190000000
1!
1'
1/
#13200000000
0!
0'
0/
#13210000000
1!
1'
1/
#13220000000
0!
0'
0/
#13230000000
1!
1'
1/
#13240000000
0!
0'
0/
#13250000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#13260000000
0!
0'
0/
#13270000000
1!
1'
1/
#13280000000
0!
0'
0/
#13290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#13300000000
0!
0'
0/
#13310000000
1!
1'
1/
#13320000000
0!
0'
0/
#13330000000
#13340000000
1!
1'
1/
#13350000000
0!
0'
0/
#13360000000
1!
1'
1/
#13370000000
0!
1"
0'
1(
0/
10
#13380000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#13390000000
0!
0'
0/
#13400000000
1!
1'
1/
#13410000000
0!
0'
0/
#13420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#13430000000
0!
0'
0/
#13440000000
1!
1'
1/
#13450000000
0!
1"
0'
1(
0/
10
#13460000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#13470000000
0!
1$
0'
1+
0/
#13480000000
1!
1'
1/
#13490000000
0!
0'
0/
#13500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#13510000000
0!
0'
0/
#13520000000
1!
1'
1/
#13530000000
0!
0'
0/
#13540000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#13550000000
0!
0'
0/
#13560000000
1!
1'
1/
#13570000000
0!
0'
0/
#13580000000
1!
1'
1/
#13590000000
0!
0'
0/
#13600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#13610000000
0!
0'
0/
#13620000000
1!
1'
1/
#13630000000
0!
0'
0/
#13640000000
1!
1'
1/
#13650000000
0!
0'
0/
#13660000000
1!
1'
1/
#13670000000
0!
0'
0/
#13680000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#13690000000
0!
0'
0/
#13700000000
1!
1'
1/
#13710000000
0!
0'
0/
#13720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#13730000000
0!
0'
0/
#13740000000
1!
1'
1/
#13750000000
0!
0'
0/
#13760000000
#13770000000
1!
1'
1/
#13780000000
0!
0'
0/
#13790000000
1!
1'
1/
#13800000000
0!
1"
0'
1(
0/
10
#13810000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#13820000000
0!
0'
0/
#13830000000
1!
1'
1/
#13840000000
0!
0'
0/
#13850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#13860000000
0!
0'
0/
#13870000000
1!
1'
1/
#13880000000
0!
1"
0'
1(
0/
10
#13890000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#13900000000
0!
1$
0'
1+
0/
#13910000000
1!
1'
1/
#13920000000
0!
0'
0/
#13930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#13940000000
0!
0'
0/
#13950000000
1!
1'
1/
#13960000000
0!
0'
0/
#13970000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#13980000000
0!
0'
0/
#13990000000
1!
1'
1/
#14000000000
0!
0'
0/
#14010000000
1!
1'
1/
#14020000000
0!
0'
0/
#14030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#14040000000
0!
0'
0/
#14050000000
1!
1'
1/
#14060000000
0!
0'
0/
#14070000000
1!
1'
1/
#14080000000
0!
0'
0/
#14090000000
1!
1'
1/
#14100000000
0!
0'
0/
#14110000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#14120000000
0!
0'
0/
#14130000000
1!
1'
1/
#14140000000
0!
0'
0/
#14150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#14160000000
0!
0'
0/
#14170000000
1!
1'
1/
#14180000000
0!
0'
0/
#14190000000
#14200000000
1!
1'
1/
#14210000000
0!
0'
0/
#14220000000
1!
1'
1/
#14230000000
0!
1"
0'
1(
0/
10
#14240000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#14250000000
0!
0'
0/
#14260000000
1!
1'
1/
#14270000000
0!
0'
0/
#14280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#14290000000
0!
0'
0/
#14300000000
1!
1'
1/
#14310000000
0!
1"
0'
1(
0/
10
#14320000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#14330000000
0!
1$
0'
1+
0/
#14340000000
1!
1'
1/
#14350000000
0!
0'
0/
#14360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#14370000000
0!
0'
0/
#14380000000
1!
1'
1/
#14390000000
0!
0'
0/
#14400000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#14410000000
0!
0'
0/
#14420000000
1!
1'
1/
#14430000000
0!
0'
0/
#14440000000
1!
1'
1/
#14450000000
0!
0'
0/
#14460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#14470000000
0!
0'
0/
#14480000000
1!
1'
1/
#14490000000
0!
0'
0/
#14500000000
1!
1'
1/
#14510000000
0!
0'
0/
#14520000000
1!
1'
1/
#14530000000
0!
0'
0/
#14540000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#14550000000
0!
0'
0/
#14560000000
1!
1'
1/
#14570000000
0!
0'
0/
#14580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#14590000000
0!
0'
0/
#14600000000
1!
1'
1/
#14610000000
0!
0'
0/
#14620000000
#14630000000
1!
1'
1/
#14640000000
0!
0'
0/
#14650000000
1!
1'
1/
#14660000000
0!
1"
0'
1(
0/
10
#14670000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#14680000000
0!
0'
0/
#14690000000
1!
1'
1/
#14700000000
0!
0'
0/
#14710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#14720000000
0!
0'
0/
#14730000000
1!
1'
1/
#14740000000
0!
1"
0'
1(
0/
10
#14750000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#14760000000
0!
1$
0'
1+
0/
#14770000000
1!
1'
1/
#14780000000
0!
0'
0/
#14790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#14800000000
0!
0'
0/
#14810000000
1!
1'
1/
#14820000000
0!
0'
0/
#14830000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#14840000000
0!
0'
0/
#14850000000
1!
1'
1/
#14860000000
0!
0'
0/
#14870000000
1!
1'
1/
#14880000000
0!
0'
0/
#14890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#14900000000
0!
0'
0/
#14910000000
1!
1'
1/
#14920000000
0!
0'
0/
#14930000000
1!
1'
1/
#14940000000
0!
0'
0/
#14950000000
1!
1'
1/
#14960000000
0!
0'
0/
#14970000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#14980000000
0!
0'
0/
#14990000000
1!
1'
1/
#15000000000
0!
0'
0/
#15010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#15020000000
0!
0'
0/
#15030000000
1!
1'
1/
#15040000000
0!
0'
0/
#15050000000
#15060000000
1!
1'
1/
#15070000000
0!
0'
0/
#15080000000
1!
1'
1/
#15090000000
0!
1"
0'
1(
0/
10
#15100000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#15110000000
0!
0'
0/
#15120000000
1!
1'
1/
#15130000000
0!
0'
0/
#15140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#15150000000
0!
0'
0/
#15160000000
1!
1'
1/
#15170000000
0!
1"
0'
1(
0/
10
#15180000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#15190000000
0!
1$
0'
1+
0/
#15200000000
1!
1'
1/
#15210000000
0!
0'
0/
#15220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#15230000000
0!
0'
0/
#15240000000
1!
1'
1/
#15250000000
0!
0'
0/
#15260000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#15270000000
0!
0'
0/
#15280000000
1!
1'
1/
#15290000000
0!
0'
0/
#15300000000
1!
1'
1/
#15310000000
0!
0'
0/
#15320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#15330000000
0!
0'
0/
#15340000000
1!
1'
1/
#15350000000
0!
0'
0/
#15360000000
1!
1'
1/
#15370000000
0!
0'
0/
#15380000000
1!
1'
1/
#15390000000
0!
0'
0/
#15400000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#15410000000
0!
0'
0/
#15420000000
1!
1'
1/
#15430000000
0!
0'
0/
#15440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#15450000000
0!
0'
0/
#15460000000
1!
1'
1/
#15470000000
0!
0'
0/
#15480000000
#15490000000
1!
1'
1/
#15500000000
0!
0'
0/
#15510000000
1!
1'
1/
#15520000000
0!
1"
0'
1(
0/
10
#15530000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#15540000000
0!
0'
0/
#15550000000
1!
1'
1/
#15560000000
0!
0'
0/
#15570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#15580000000
0!
0'
0/
#15590000000
1!
1'
1/
#15600000000
0!
1"
0'
1(
0/
10
#15610000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#15620000000
0!
1$
0'
1+
0/
#15630000000
1!
1'
1/
#15640000000
0!
0'
0/
#15650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#15660000000
0!
0'
0/
#15670000000
1!
1'
1/
#15680000000
0!
0'
0/
#15690000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#15700000000
0!
0'
0/
#15710000000
1!
1'
1/
#15720000000
0!
0'
0/
#15730000000
1!
1'
1/
#15740000000
0!
0'
0/
#15750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#15760000000
0!
0'
0/
#15770000000
1!
1'
1/
#15780000000
0!
0'
0/
#15790000000
1!
1'
1/
#15800000000
0!
0'
0/
#15810000000
1!
1'
1/
#15820000000
0!
0'
0/
#15830000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#15840000000
0!
0'
0/
#15850000000
1!
1'
1/
#15860000000
0!
0'
0/
#15870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#15880000000
0!
0'
0/
#15890000000
1!
1'
1/
#15900000000
0!
0'
0/
#15910000000
#15920000000
1!
1'
1/
#15930000000
0!
0'
0/
#15940000000
1!
1'
1/
#15950000000
0!
1"
0'
1(
0/
10
#15960000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#15970000000
0!
0'
0/
#15980000000
1!
1'
1/
#15990000000
0!
0'
0/
#16000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#16010000000
0!
0'
0/
#16020000000
1!
1'
1/
#16030000000
0!
1"
0'
1(
0/
10
#16040000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#16050000000
0!
1$
0'
1+
0/
#16060000000
1!
1'
1/
#16070000000
0!
0'
0/
#16080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#16090000000
0!
0'
0/
#16100000000
1!
1'
1/
#16110000000
0!
0'
0/
#16120000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#16130000000
0!
0'
0/
#16140000000
1!
1'
1/
#16150000000
0!
0'
0/
#16160000000
1!
1'
1/
#16170000000
0!
0'
0/
#16180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#16190000000
0!
0'
0/
#16200000000
1!
1'
1/
#16210000000
0!
0'
0/
#16220000000
1!
1'
1/
#16230000000
0!
0'
0/
#16240000000
1!
1'
1/
#16250000000
0!
0'
0/
#16260000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#16270000000
0!
0'
0/
#16280000000
1!
1'
1/
#16290000000
0!
0'
0/
#16300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#16310000000
0!
0'
0/
#16320000000
1!
1'
1/
#16330000000
0!
0'
0/
#16340000000
#16350000000
1!
1'
1/
#16360000000
0!
0'
0/
#16370000000
1!
1'
1/
#16380000000
0!
1"
0'
1(
0/
10
#16390000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#16400000000
0!
0'
0/
#16410000000
1!
1'
1/
#16420000000
0!
0'
0/
#16430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#16440000000
0!
0'
0/
#16450000000
1!
1'
1/
#16460000000
0!
1"
0'
1(
0/
10
#16470000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#16480000000
0!
1$
0'
1+
0/
#16490000000
1!
1'
1/
#16500000000
0!
0'
0/
#16510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#16520000000
0!
0'
0/
#16530000000
1!
1'
1/
#16540000000
0!
0'
0/
#16550000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#16560000000
0!
0'
0/
#16570000000
1!
1'
1/
#16580000000
0!
0'
0/
#16590000000
1!
1'
1/
#16600000000
0!
0'
0/
#16610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#16620000000
0!
0'
0/
#16630000000
1!
1'
1/
#16640000000
0!
0'
0/
#16650000000
1!
1'
1/
#16660000000
0!
0'
0/
#16670000000
1!
1'
1/
#16680000000
0!
0'
0/
#16690000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#16700000000
0!
0'
0/
#16710000000
1!
1'
1/
#16720000000
0!
0'
0/
#16730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#16740000000
0!
0'
0/
#16750000000
1!
1'
1/
#16760000000
0!
0'
0/
#16770000000
#16780000000
1!
1'
1/
#16790000000
0!
0'
0/
#16800000000
1!
1'
1/
#16810000000
0!
1"
0'
1(
0/
10
#16820000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#16830000000
0!
0'
0/
#16840000000
1!
1'
1/
#16850000000
0!
0'
0/
#16860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#16870000000
0!
0'
0/
#16880000000
1!
1'
1/
#16890000000
0!
1"
0'
1(
0/
10
#16900000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#16910000000
0!
1$
0'
1+
0/
#16920000000
1!
1'
1/
#16930000000
0!
0'
0/
#16940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#16950000000
0!
0'
0/
#16960000000
1!
1'
1/
#16970000000
0!
0'
0/
#16980000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#16990000000
0!
0'
0/
#17000000000
1!
1'
1/
#17010000000
0!
0'
0/
#17020000000
1!
1'
1/
#17030000000
0!
0'
0/
#17040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#17050000000
0!
0'
0/
#17060000000
1!
1'
1/
#17070000000
0!
0'
0/
#17080000000
1!
1'
1/
#17090000000
0!
0'
0/
#17100000000
1!
1'
1/
#17110000000
0!
0'
0/
#17120000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#17130000000
0!
0'
0/
#17140000000
1!
1'
1/
#17150000000
0!
0'
0/
#17160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#17170000000
0!
0'
0/
#17180000000
1!
1'
1/
#17190000000
0!
0'
0/
#17200000000
#17210000000
1!
1'
1/
#17220000000
0!
0'
0/
#17230000000
1!
1'
1/
#17240000000
0!
1"
0'
1(
0/
10
#17250000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#17260000000
0!
0'
0/
#17270000000
1!
1'
1/
#17280000000
0!
0'
0/
#17290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#17300000000
0!
0'
0/
#17310000000
1!
1'
1/
#17320000000
0!
1"
0'
1(
0/
10
#17330000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#17340000000
0!
1$
0'
1+
0/
#17350000000
1!
1'
1/
#17360000000
0!
0'
0/
#17370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#17380000000
0!
0'
0/
#17390000000
1!
1'
1/
#17400000000
0!
0'
0/
#17410000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#17420000000
0!
0'
0/
#17430000000
1!
1'
1/
#17440000000
0!
0'
0/
#17450000000
1!
1'
1/
#17460000000
0!
0'
0/
#17470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#17480000000
0!
0'
0/
#17490000000
1!
1'
1/
#17500000000
0!
0'
0/
#17510000000
1!
1'
1/
#17520000000
0!
0'
0/
#17530000000
1!
1'
1/
#17540000000
0!
0'
0/
#17550000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#17560000000
0!
0'
0/
#17570000000
1!
1'
1/
#17580000000
0!
0'
0/
#17590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#17600000000
0!
0'
0/
#17610000000
1!
1'
1/
#17620000000
0!
0'
0/
#17630000000
#17640000000
1!
1'
1/
#17650000000
0!
0'
0/
#17660000000
1!
1'
1/
#17670000000
0!
1"
0'
1(
0/
10
#17680000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#17690000000
0!
0'
0/
#17700000000
1!
1'
1/
#17710000000
0!
0'
0/
#17720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#17730000000
0!
0'
0/
#17740000000
1!
1'
1/
#17750000000
0!
1"
0'
1(
0/
10
#17760000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#17770000000
0!
1$
0'
1+
0/
#17780000000
1!
1'
1/
#17790000000
0!
0'
0/
#17800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#17810000000
0!
0'
0/
#17820000000
1!
1'
1/
#17830000000
0!
0'
0/
#17840000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#17850000000
0!
0'
0/
#17860000000
1!
1'
1/
#17870000000
0!
0'
0/
#17880000000
1!
1'
1/
#17890000000
0!
0'
0/
#17900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#17910000000
0!
0'
0/
#17920000000
1!
1'
1/
#17930000000
0!
0'
0/
#17940000000
1!
1'
1/
#17950000000
0!
0'
0/
#17960000000
1!
1'
1/
#17970000000
0!
0'
0/
#17980000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#17990000000
0!
0'
0/
#18000000000
1!
1'
1/
#18010000000
0!
0'
0/
#18020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#18030000000
0!
0'
0/
#18040000000
1!
1'
1/
#18050000000
0!
0'
0/
#18060000000
#18070000000
1!
1'
1/
#18080000000
0!
0'
0/
#18090000000
1!
1'
1/
#18100000000
0!
1"
0'
1(
0/
10
#18110000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#18120000000
0!
0'
0/
#18130000000
1!
1'
1/
#18140000000
0!
0'
0/
#18150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#18160000000
0!
0'
0/
#18170000000
1!
1'
1/
#18180000000
0!
1"
0'
1(
0/
10
#18190000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#18200000000
0!
1$
0'
1+
0/
#18210000000
1!
1'
1/
#18220000000
0!
0'
0/
#18230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#18240000000
0!
0'
0/
#18250000000
1!
1'
1/
#18260000000
0!
0'
0/
#18270000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#18280000000
0!
0'
0/
#18290000000
1!
1'
1/
#18300000000
0!
0'
0/
#18310000000
1!
1'
1/
#18320000000
0!
0'
0/
#18330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#18340000000
0!
0'
0/
#18350000000
1!
1'
1/
#18360000000
0!
0'
0/
#18370000000
1!
1'
1/
#18380000000
0!
0'
0/
#18390000000
1!
1'
1/
#18400000000
0!
0'
0/
#18410000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#18420000000
0!
0'
0/
#18430000000
1!
1'
1/
#18440000000
0!
0'
0/
#18450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#18460000000
0!
0'
0/
#18470000000
1!
1'
1/
#18480000000
0!
0'
0/
#18490000000
#18500000000
1!
1'
1/
#18510000000
0!
0'
0/
#18520000000
1!
1'
1/
#18530000000
0!
1"
0'
1(
0/
10
#18540000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#18550000000
0!
0'
0/
#18560000000
1!
1'
1/
#18570000000
0!
0'
0/
#18580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#18590000000
0!
0'
0/
#18600000000
1!
1'
1/
#18610000000
0!
1"
0'
1(
0/
10
#18620000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#18630000000
0!
1$
0'
1+
0/
#18640000000
1!
1'
1/
#18650000000
0!
0'
0/
#18660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#18670000000
0!
0'
0/
#18680000000
1!
1'
1/
#18690000000
0!
0'
0/
#18700000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#18710000000
0!
0'
0/
#18720000000
1!
1'
1/
#18730000000
0!
0'
0/
#18740000000
1!
1'
1/
#18750000000
0!
0'
0/
#18760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#18770000000
0!
0'
0/
#18780000000
1!
1'
1/
#18790000000
0!
0'
0/
#18800000000
1!
1'
1/
#18810000000
0!
0'
0/
#18820000000
1!
1'
1/
#18830000000
0!
0'
0/
#18840000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#18850000000
0!
0'
0/
#18860000000
1!
1'
1/
#18870000000
0!
0'
0/
#18880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#18890000000
0!
0'
0/
#18900000000
1!
1'
1/
#18910000000
0!
0'
0/
#18920000000
#18930000000
1!
1'
1/
#18940000000
0!
0'
0/
#18950000000
1!
1'
1/
#18960000000
0!
1"
0'
1(
0/
10
#18970000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#18980000000
0!
0'
0/
#18990000000
1!
1'
1/
#19000000000
0!
0'
0/
#19010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#19020000000
0!
0'
0/
#19030000000
1!
1'
1/
#19040000000
0!
1"
0'
1(
0/
10
#19050000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#19060000000
0!
1$
0'
1+
0/
#19070000000
1!
1'
1/
#19080000000
0!
0'
0/
#19090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#19100000000
0!
0'
0/
#19110000000
1!
1'
1/
#19120000000
0!
0'
0/
#19130000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#19140000000
0!
0'
0/
#19150000000
1!
1'
1/
#19160000000
0!
0'
0/
#19170000000
1!
1'
1/
#19180000000
0!
0'
0/
#19190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#19200000000
0!
0'
0/
#19210000000
1!
1'
1/
#19220000000
0!
0'
0/
#19230000000
1!
1'
1/
#19240000000
0!
0'
0/
#19250000000
1!
1'
1/
#19260000000
0!
0'
0/
#19270000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#19280000000
0!
0'
0/
#19290000000
1!
1'
1/
#19300000000
0!
0'
0/
#19310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#19320000000
0!
0'
0/
#19330000000
1!
1'
1/
#19340000000
0!
0'
0/
#19350000000
#19360000000
1!
1'
1/
#19370000000
0!
0'
0/
#19380000000
1!
1'
1/
#19390000000
0!
1"
0'
1(
0/
10
#19400000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#19410000000
0!
0'
0/
#19420000000
1!
1'
1/
#19430000000
0!
0'
0/
#19440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#19450000000
0!
0'
0/
#19460000000
1!
1'
1/
#19470000000
0!
1"
0'
1(
0/
10
#19480000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#19490000000
0!
1$
0'
1+
0/
#19500000000
1!
1'
1/
#19510000000
0!
0'
0/
#19520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#19530000000
0!
0'
0/
#19540000000
1!
1'
1/
#19550000000
0!
0'
0/
#19560000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#19570000000
0!
0'
0/
#19580000000
1!
1'
1/
#19590000000
0!
0'
0/
#19600000000
1!
1'
1/
#19610000000
0!
0'
0/
#19620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#19630000000
0!
0'
0/
#19640000000
1!
1'
1/
#19650000000
0!
0'
0/
#19660000000
1!
1'
1/
#19670000000
0!
0'
0/
#19680000000
1!
1'
1/
#19690000000
0!
0'
0/
#19700000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#19710000000
0!
0'
0/
#19720000000
1!
1'
1/
#19730000000
0!
0'
0/
#19740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#19750000000
0!
0'
0/
#19760000000
1!
1'
1/
#19770000000
0!
0'
0/
#19780000000
#19790000000
1!
1'
1/
#19800000000
0!
0'
0/
#19810000000
1!
1'
1/
#19820000000
0!
1"
0'
1(
0/
10
#19830000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#19840000000
0!
0'
0/
#19850000000
1!
1'
1/
#19860000000
0!
0'
0/
#19870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#19880000000
0!
0'
0/
#19890000000
1!
1'
1/
#19900000000
0!
1"
0'
1(
0/
10
#19910000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#19920000000
0!
1$
0'
1+
0/
#19930000000
1!
1'
1/
#19940000000
0!
0'
0/
#19950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#19960000000
0!
0'
0/
#19970000000
1!
1'
1/
#19980000000
0!
0'
0/
#19990000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#20000000000
0!
0'
0/
#20010000000
1!
1'
1/
#20020000000
0!
0'
0/
#20030000000
1!
1'
1/
#20040000000
0!
0'
0/
#20050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#20060000000
0!
0'
0/
#20070000000
1!
1'
1/
#20080000000
0!
0'
0/
#20090000000
1!
1'
1/
#20100000000
0!
0'
0/
#20110000000
1!
1'
1/
#20120000000
0!
0'
0/
#20130000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#20140000000
0!
0'
0/
#20150000000
1!
1'
1/
#20160000000
0!
0'
0/
#20170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#20180000000
0!
0'
0/
#20190000000
1!
1'
1/
#20200000000
0!
0'
0/
#20210000000
#20220000000
1!
1'
1/
#20230000000
0!
0'
0/
#20240000000
1!
1'
1/
#20250000000
0!
1"
0'
1(
0/
10
#20260000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#20270000000
0!
0'
0/
#20280000000
1!
1'
1/
#20290000000
0!
0'
0/
#20300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#20310000000
0!
0'
0/
#20320000000
1!
1'
1/
#20330000000
0!
1"
0'
1(
0/
10
#20340000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#20350000000
0!
1$
0'
1+
0/
#20360000000
1!
1'
1/
#20370000000
0!
0'
0/
#20380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#20390000000
0!
0'
0/
#20400000000
1!
1'
1/
#20410000000
0!
0'
0/
#20420000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#20430000000
0!
0'
0/
#20440000000
1!
1'
1/
#20450000000
0!
0'
0/
#20460000000
1!
1'
1/
#20470000000
0!
0'
0/
#20480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#20490000000
0!
0'
0/
#20500000000
1!
1'
1/
#20510000000
0!
0'
0/
#20520000000
1!
1'
1/
#20530000000
0!
0'
0/
#20540000000
1!
1'
1/
#20550000000
0!
0'
0/
#20560000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#20570000000
0!
0'
0/
#20580000000
1!
1'
1/
#20590000000
0!
0'
0/
#20600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#20610000000
0!
0'
0/
#20620000000
1!
1'
1/
#20630000000
0!
0'
0/
#20640000000
#20650000000
1!
1'
1/
#20660000000
0!
0'
0/
#20670000000
1!
1'
1/
#20680000000
0!
1"
0'
1(
0/
10
#20690000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#20700000000
0!
0'
0/
#20710000000
1!
1'
1/
#20720000000
0!
0'
0/
#20730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#20740000000
0!
0'
0/
#20750000000
1!
1'
1/
#20760000000
0!
1"
0'
1(
0/
10
#20770000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#20780000000
0!
1$
0'
1+
0/
#20790000000
1!
1'
1/
#20800000000
0!
0'
0/
#20810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#20820000000
0!
0'
0/
#20830000000
1!
1'
1/
#20840000000
0!
0'
0/
#20850000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#20860000000
0!
0'
0/
#20870000000
1!
1'
1/
#20880000000
0!
0'
0/
#20890000000
1!
1'
1/
#20900000000
0!
0'
0/
#20910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#20920000000
0!
0'
0/
#20930000000
1!
1'
1/
#20940000000
0!
0'
0/
#20950000000
1!
1'
1/
#20960000000
0!
0'
0/
#20970000000
1!
1'
1/
#20980000000
0!
0'
0/
#20990000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#21000000000
0!
0'
0/
#21010000000
1!
1'
1/
#21020000000
0!
0'
0/
#21030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#21040000000
0!
0'
0/
#21050000000
1!
1'
1/
#21060000000
0!
0'
0/
#21070000000
#21080000000
1!
1'
1/
#21090000000
0!
0'
0/
#21100000000
1!
1'
1/
#21110000000
0!
1"
0'
1(
0/
10
#21120000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#21130000000
0!
0'
0/
#21140000000
1!
1'
1/
#21150000000
0!
0'
0/
#21160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#21170000000
0!
0'
0/
#21180000000
1!
1'
1/
#21190000000
0!
1"
0'
1(
0/
10
#21200000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#21210000000
0!
1$
0'
1+
0/
#21220000000
1!
1'
1/
#21230000000
0!
0'
0/
#21240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#21250000000
0!
0'
0/
#21260000000
1!
1'
1/
#21270000000
0!
0'
0/
#21280000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#21290000000
0!
0'
0/
#21300000000
1!
1'
1/
#21310000000
0!
0'
0/
#21320000000
1!
1'
1/
#21330000000
0!
0'
0/
#21340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#21350000000
0!
0'
0/
#21360000000
1!
1'
1/
#21370000000
0!
0'
0/
#21380000000
1!
1'
1/
#21390000000
0!
0'
0/
#21400000000
1!
1'
1/
#21410000000
0!
0'
0/
#21420000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#21430000000
0!
0'
0/
#21440000000
1!
1'
1/
#21450000000
0!
0'
0/
#21460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#21470000000
0!
0'
0/
#21480000000
1!
1'
1/
#21490000000
0!
0'
0/
#21500000000
#21510000000
1!
1'
1/
#21520000000
0!
0'
0/
#21530000000
1!
1'
1/
#21540000000
0!
1"
0'
1(
0/
10
#21550000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#21560000000
0!
0'
0/
#21570000000
1!
1'
1/
#21580000000
0!
0'
0/
#21590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#21600000000
0!
0'
0/
#21610000000
1!
1'
1/
#21620000000
0!
1"
0'
1(
0/
10
#21630000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#21640000000
0!
1$
0'
1+
0/
#21650000000
1!
1'
1/
#21660000000
0!
0'
0/
#21670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#21680000000
0!
0'
0/
#21690000000
1!
1'
1/
#21700000000
0!
0'
0/
#21710000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#21720000000
0!
0'
0/
#21730000000
1!
1'
1/
#21740000000
0!
0'
0/
#21750000000
1!
1'
1/
#21760000000
0!
0'
0/
#21770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#21780000000
0!
0'
0/
#21790000000
1!
1'
1/
#21800000000
0!
0'
0/
#21810000000
1!
1'
1/
#21820000000
0!
0'
0/
#21830000000
1!
1'
1/
#21840000000
0!
0'
0/
#21850000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#21860000000
0!
0'
0/
#21870000000
1!
1'
1/
#21880000000
0!
0'
0/
#21890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#21900000000
0!
0'
0/
#21910000000
1!
1'
1/
#21920000000
0!
0'
0/
#21930000000
#21940000000
1!
1'
1/
#21950000000
0!
0'
0/
#21960000000
1!
1'
1/
#21970000000
0!
1"
0'
1(
0/
10
#21980000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#21990000000
0!
0'
0/
#22000000000
1!
1'
1/
#22010000000
0!
0'
0/
#22020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#22030000000
0!
0'
0/
#22040000000
1!
1'
1/
#22050000000
0!
1"
0'
1(
0/
10
#22060000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#22070000000
0!
1$
0'
1+
0/
#22080000000
1!
1'
1/
#22090000000
0!
0'
0/
#22100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#22110000000
0!
0'
0/
#22120000000
1!
1'
1/
#22130000000
0!
0'
0/
#22140000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#22150000000
0!
0'
0/
#22160000000
1!
1'
1/
#22170000000
0!
0'
0/
#22180000000
1!
1'
1/
#22190000000
0!
0'
0/
#22200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#22210000000
0!
0'
0/
#22220000000
1!
1'
1/
#22230000000
0!
0'
0/
#22240000000
1!
1'
1/
#22250000000
0!
0'
0/
#22260000000
1!
1'
1/
#22270000000
0!
0'
0/
#22280000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#22290000000
0!
0'
0/
#22300000000
1!
1'
1/
#22310000000
0!
0'
0/
#22320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#22330000000
0!
0'
0/
#22340000000
1!
1'
1/
#22350000000
0!
0'
0/
#22360000000
#22370000000
1!
1'
1/
#22380000000
0!
0'
0/
#22390000000
1!
1'
1/
#22400000000
0!
1"
0'
1(
0/
10
#22410000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#22420000000
0!
0'
0/
#22430000000
1!
1'
1/
#22440000000
0!
0'
0/
#22450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#22460000000
0!
0'
0/
#22470000000
1!
1'
1/
#22480000000
0!
1"
0'
1(
0/
10
#22490000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#22500000000
0!
1$
0'
1+
0/
#22510000000
1!
1'
1/
#22520000000
0!
0'
0/
#22530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#22540000000
0!
0'
0/
#22550000000
1!
1'
1/
#22560000000
0!
0'
0/
#22570000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#22580000000
0!
0'
0/
#22590000000
1!
1'
1/
#22600000000
0!
0'
0/
#22610000000
1!
1'
1/
#22620000000
0!
0'
0/
#22630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#22640000000
0!
0'
0/
#22650000000
1!
1'
1/
#22660000000
0!
0'
0/
#22670000000
1!
1'
1/
#22680000000
0!
0'
0/
#22690000000
1!
1'
1/
#22700000000
0!
0'
0/
#22710000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#22720000000
0!
0'
0/
#22730000000
1!
1'
1/
#22740000000
0!
0'
0/
#22750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#22760000000
0!
0'
0/
#22770000000
1!
1'
1/
#22780000000
0!
0'
0/
#22790000000
#22800000000
1!
1'
1/
#22810000000
0!
0'
0/
#22820000000
1!
1'
1/
#22830000000
0!
1"
0'
1(
0/
10
#22840000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#22850000000
0!
0'
0/
#22860000000
1!
1'
1/
#22870000000
0!
0'
0/
#22880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#22890000000
0!
0'
0/
#22900000000
1!
1'
1/
#22910000000
0!
1"
0'
1(
0/
10
#22920000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#22930000000
0!
1$
0'
1+
0/
#22940000000
1!
1'
1/
#22950000000
0!
0'
0/
#22960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#22970000000
0!
0'
0/
#22980000000
1!
1'
1/
#22990000000
0!
0'
0/
#23000000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#23010000000
0!
0'
0/
#23020000000
1!
1'
1/
#23030000000
0!
0'
0/
#23040000000
1!
1'
1/
#23050000000
0!
0'
0/
#23060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#23070000000
0!
0'
0/
#23080000000
1!
1'
1/
#23090000000
0!
0'
0/
#23100000000
1!
1'
1/
#23110000000
0!
0'
0/
#23120000000
1!
1'
1/
#23130000000
0!
0'
0/
#23140000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#23150000000
0!
0'
0/
#23160000000
1!
1'
1/
#23170000000
0!
0'
0/
#23180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#23190000000
0!
0'
0/
#23200000000
1!
1'
1/
#23210000000
0!
0'
0/
#23220000000
#23230000000
1!
1'
1/
#23240000000
0!
0'
0/
#23250000000
1!
1'
1/
#23260000000
0!
1"
0'
1(
0/
10
#23270000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#23280000000
0!
0'
0/
#23290000000
1!
1'
1/
#23300000000
0!
0'
0/
#23310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#23320000000
0!
0'
0/
#23330000000
1!
1'
1/
#23340000000
0!
1"
0'
1(
0/
10
#23350000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#23360000000
0!
1$
0'
1+
0/
#23370000000
1!
1'
1/
#23380000000
0!
0'
0/
#23390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#23400000000
0!
0'
0/
#23410000000
1!
1'
1/
#23420000000
0!
0'
0/
#23430000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#23440000000
0!
0'
0/
#23450000000
1!
1'
1/
#23460000000
0!
0'
0/
#23470000000
1!
1'
1/
#23480000000
0!
0'
0/
#23490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#23500000000
0!
0'
0/
#23510000000
1!
1'
1/
#23520000000
0!
0'
0/
#23530000000
1!
1'
1/
#23540000000
0!
0'
0/
#23550000000
1!
1'
1/
#23560000000
0!
0'
0/
#23570000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#23580000000
0!
0'
0/
#23590000000
1!
1'
1/
#23600000000
0!
0'
0/
#23610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#23620000000
0!
0'
0/
#23630000000
1!
1'
1/
#23640000000
0!
0'
0/
#23650000000
#23660000000
1!
1'
1/
#23670000000
0!
0'
0/
#23680000000
1!
1'
1/
#23690000000
0!
1"
0'
1(
0/
10
#23700000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#23710000000
0!
0'
0/
#23720000000
1!
1'
1/
#23730000000
0!
0'
0/
#23740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#23750000000
0!
0'
0/
#23760000000
1!
1'
1/
#23770000000
0!
1"
0'
1(
0/
10
#23780000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#23790000000
0!
1$
0'
1+
0/
#23800000000
1!
1'
1/
#23810000000
0!
0'
0/
#23820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#23830000000
0!
0'
0/
#23840000000
1!
1'
1/
#23850000000
0!
0'
0/
#23860000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#23870000000
0!
0'
0/
#23880000000
1!
1'
1/
#23890000000
0!
0'
0/
#23900000000
1!
1'
1/
#23910000000
0!
0'
0/
#23920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#23930000000
0!
0'
0/
#23940000000
1!
1'
1/
#23950000000
0!
0'
0/
#23960000000
1!
1'
1/
#23970000000
0!
0'
0/
#23980000000
1!
1'
1/
#23990000000
0!
0'
0/
#24000000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#24010000000
0!
0'
0/
#24020000000
1!
1'
1/
#24030000000
0!
0'
0/
#24040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#24050000000
0!
0'
0/
#24060000000
1!
1'
1/
#24070000000
0!
0'
0/
#24080000000
#24090000000
1!
1'
1/
#24100000000
0!
0'
0/
#24110000000
1!
1'
1/
#24120000000
0!
1"
0'
1(
0/
10
#24130000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#24140000000
0!
0'
0/
#24150000000
1!
1'
1/
#24160000000
0!
0'
0/
#24170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#24180000000
0!
0'
0/
#24190000000
1!
1'
1/
#24200000000
0!
1"
0'
1(
0/
10
#24210000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#24220000000
0!
1$
0'
1+
0/
#24230000000
1!
1'
1/
#24240000000
0!
0'
0/
#24250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#24260000000
0!
0'
0/
#24270000000
1!
1'
1/
#24280000000
0!
0'
0/
#24290000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#24300000000
0!
0'
0/
#24310000000
1!
1'
1/
#24320000000
0!
0'
0/
#24330000000
1!
1'
1/
#24340000000
0!
0'
0/
#24350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#24360000000
0!
0'
0/
#24370000000
1!
1'
1/
#24380000000
0!
0'
0/
#24390000000
1!
1'
1/
#24400000000
0!
0'
0/
#24410000000
1!
1'
1/
#24420000000
0!
0'
0/
#24430000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#24440000000
0!
0'
0/
#24450000000
1!
1'
1/
#24460000000
0!
0'
0/
#24470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#24480000000
0!
0'
0/
#24490000000
1!
1'
1/
#24500000000
0!
0'
0/
#24510000000
#24520000000
1!
1'
1/
#24530000000
0!
0'
0/
#24540000000
1!
1'
1/
#24550000000
0!
1"
0'
1(
0/
10
#24560000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#24570000000
0!
0'
0/
#24580000000
1!
1'
1/
#24590000000
0!
0'
0/
#24600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#24610000000
0!
0'
0/
#24620000000
1!
1'
1/
#24630000000
0!
1"
0'
1(
0/
10
#24640000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#24650000000
0!
1$
0'
1+
0/
#24660000000
1!
1'
1/
#24670000000
0!
0'
0/
#24680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#24690000000
0!
0'
0/
#24700000000
1!
1'
1/
#24710000000
0!
0'
0/
#24720000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#24730000000
0!
0'
0/
#24740000000
1!
1'
1/
#24750000000
0!
0'
0/
#24760000000
1!
1'
1/
#24770000000
0!
0'
0/
#24780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#24790000000
0!
0'
0/
#24800000000
1!
1'
1/
#24810000000
0!
0'
0/
#24820000000
1!
1'
1/
#24830000000
0!
0'
0/
#24840000000
1!
1'
1/
#24850000000
0!
0'
0/
#24860000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#24870000000
0!
0'
0/
#24880000000
1!
1'
1/
#24890000000
0!
0'
0/
#24900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#24910000000
0!
0'
0/
#24920000000
1!
1'
1/
#24930000000
0!
0'
0/
#24940000000
#24950000000
1!
1'
1/
#24960000000
0!
0'
0/
#24970000000
1!
1'
1/
#24980000000
0!
1"
0'
1(
0/
10
#24990000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#25000000000
0!
0'
0/
#25010000000
1!
1'
1/
#25020000000
0!
0'
0/
#25030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#25040000000
0!
0'
0/
#25050000000
1!
1'
1/
#25060000000
0!
1"
0'
1(
0/
10
#25070000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#25080000000
0!
1$
0'
1+
0/
#25090000000
1!
1'
1/
#25100000000
0!
0'
0/
#25110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#25120000000
0!
0'
0/
#25130000000
1!
1'
1/
#25140000000
0!
0'
0/
#25150000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#25160000000
0!
0'
0/
#25170000000
1!
1'
1/
#25180000000
0!
0'
0/
#25190000000
1!
1'
1/
#25200000000
0!
0'
0/
#25210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#25220000000
0!
0'
0/
#25230000000
1!
1'
1/
#25240000000
0!
0'
0/
#25250000000
1!
1'
1/
#25260000000
0!
0'
0/
#25270000000
1!
1'
1/
#25280000000
0!
0'
0/
#25290000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#25300000000
0!
0'
0/
#25310000000
1!
1'
1/
#25320000000
0!
0'
0/
#25330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#25340000000
0!
0'
0/
#25350000000
1!
1'
1/
#25360000000
0!
0'
0/
#25370000000
#25380000000
1!
1'
1/
#25390000000
0!
0'
0/
#25400000000
1!
1'
1/
#25410000000
0!
1"
0'
1(
0/
10
#25420000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#25430000000
0!
0'
0/
#25440000000
1!
1'
1/
#25450000000
0!
0'
0/
#25460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#25470000000
0!
0'
0/
#25480000000
1!
1'
1/
#25490000000
0!
1"
0'
1(
0/
10
#25500000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#25510000000
0!
1$
0'
1+
0/
#25520000000
1!
1'
1/
#25530000000
0!
0'
0/
#25540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#25550000000
0!
0'
0/
#25560000000
1!
1'
1/
#25570000000
0!
0'
0/
#25580000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#25590000000
0!
0'
0/
#25600000000
1!
1'
1/
#25610000000
0!
0'
0/
#25620000000
1!
1'
1/
#25630000000
0!
0'
0/
#25640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#25650000000
0!
0'
0/
#25660000000
1!
1'
1/
#25670000000
0!
0'
0/
#25680000000
1!
1'
1/
#25690000000
0!
0'
0/
#25700000000
1!
1'
1/
#25710000000
0!
0'
0/
#25720000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#25730000000
0!
0'
0/
#25740000000
1!
1'
1/
#25750000000
0!
0'
0/
#25760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#25770000000
0!
0'
0/
#25780000000
1!
1'
1/
#25790000000
0!
0'
0/
#25800000000
#25810000000
1!
1'
1/
#25820000000
0!
0'
0/
#25830000000
1!
1'
1/
#25840000000
0!
1"
0'
1(
0/
10
#25850000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#25860000000
0!
0'
0/
#25870000000
1!
1'
1/
#25880000000
0!
0'
0/
#25890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#25900000000
0!
0'
0/
#25910000000
1!
1'
1/
#25920000000
0!
1"
0'
1(
0/
10
#25930000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#25940000000
0!
1$
0'
1+
0/
#25950000000
1!
1'
1/
#25960000000
0!
0'
0/
#25970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#25980000000
0!
0'
0/
#25990000000
1!
1'
1/
#26000000000
0!
0'
0/
#26010000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#26020000000
0!
0'
0/
#26030000000
1!
1'
1/
#26040000000
0!
0'
0/
#26050000000
1!
1'
1/
#26060000000
0!
0'
0/
#26070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#26080000000
0!
0'
0/
#26090000000
1!
1'
1/
#26100000000
0!
0'
0/
#26110000000
1!
1'
1/
#26120000000
0!
0'
0/
#26130000000
1!
1'
1/
#26140000000
0!
0'
0/
#26150000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#26160000000
0!
0'
0/
#26170000000
1!
1'
1/
#26180000000
0!
0'
0/
#26190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#26200000000
0!
0'
0/
#26210000000
1!
1'
1/
#26220000000
0!
0'
0/
#26230000000
#26240000000
1!
1'
1/
#26250000000
0!
0'
0/
#26260000000
1!
1'
1/
#26270000000
0!
1"
0'
1(
0/
10
#26280000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#26290000000
0!
0'
0/
#26300000000
1!
1'
1/
#26310000000
0!
0'
0/
#26320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#26330000000
0!
0'
0/
#26340000000
1!
1'
1/
#26350000000
0!
1"
0'
1(
0/
10
#26360000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#26370000000
0!
1$
0'
1+
0/
#26380000000
1!
1'
1/
#26390000000
0!
0'
0/
#26400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#26410000000
0!
0'
0/
#26420000000
1!
1'
1/
#26430000000
0!
0'
0/
#26440000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#26450000000
0!
0'
0/
#26460000000
1!
1'
1/
#26470000000
0!
0'
0/
#26480000000
1!
1'
1/
#26490000000
0!
0'
0/
#26500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#26510000000
0!
0'
0/
#26520000000
1!
1'
1/
#26530000000
0!
0'
0/
#26540000000
1!
1'
1/
#26550000000
0!
0'
0/
#26560000000
1!
1'
1/
#26570000000
0!
0'
0/
#26580000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#26590000000
0!
0'
0/
#26600000000
1!
1'
1/
#26610000000
0!
0'
0/
#26620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#26630000000
0!
0'
0/
#26640000000
1!
1'
1/
#26650000000
0!
0'
0/
#26660000000
#26670000000
1!
1'
1/
#26680000000
0!
0'
0/
#26690000000
1!
1'
1/
#26700000000
0!
1"
0'
1(
0/
10
#26710000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#26720000000
0!
0'
0/
#26730000000
1!
1'
1/
#26740000000
0!
0'
0/
#26750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#26760000000
0!
0'
0/
#26770000000
1!
1'
1/
#26780000000
0!
1"
0'
1(
0/
10
#26790000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#26800000000
0!
1$
0'
1+
0/
#26810000000
1!
1'
1/
#26820000000
0!
0'
0/
#26830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#26840000000
0!
0'
0/
#26850000000
1!
1'
1/
#26860000000
0!
0'
0/
#26870000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#26880000000
0!
0'
0/
#26890000000
1!
1'
1/
#26900000000
0!
0'
0/
#26910000000
1!
1'
1/
#26920000000
0!
0'
0/
#26930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#26940000000
0!
0'
0/
#26950000000
1!
1'
1/
#26960000000
0!
0'
0/
#26970000000
1!
1'
1/
#26980000000
0!
0'
0/
#26990000000
1!
1'
1/
#27000000000
0!
0'
0/
#27010000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#27020000000
0!
0'
0/
#27030000000
1!
1'
1/
#27040000000
0!
0'
0/
#27050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#27060000000
0!
0'
0/
#27070000000
1!
1'
1/
#27080000000
0!
0'
0/
#27090000000
#27100000000
1!
1'
1/
#27110000000
0!
0'
0/
#27120000000
1!
1'
1/
#27130000000
0!
1"
0'
1(
0/
10
#27140000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#27150000000
0!
0'
0/
#27160000000
1!
1'
1/
#27170000000
0!
0'
0/
#27180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#27190000000
0!
0'
0/
#27200000000
1!
1'
1/
#27210000000
0!
1"
0'
1(
0/
10
#27220000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#27230000000
0!
1$
0'
1+
0/
#27240000000
1!
1'
1/
#27250000000
0!
0'
0/
#27260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#27270000000
0!
0'
0/
#27280000000
1!
1'
1/
#27290000000
0!
0'
0/
#27300000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#27310000000
0!
0'
0/
#27320000000
1!
1'
1/
#27330000000
0!
0'
0/
#27340000000
1!
1'
1/
#27350000000
0!
0'
0/
#27360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#27370000000
0!
0'
0/
#27380000000
1!
1'
1/
#27390000000
0!
0'
0/
#27400000000
1!
1'
1/
#27410000000
0!
0'
0/
#27420000000
1!
1'
1/
#27430000000
0!
0'
0/
#27440000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#27450000000
0!
0'
0/
#27460000000
1!
1'
1/
#27470000000
0!
0'
0/
#27480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#27490000000
0!
0'
0/
#27500000000
1!
1'
1/
#27510000000
0!
0'
0/
#27520000000
#27530000000
1!
1'
1/
#27540000000
0!
0'
0/
#27550000000
1!
1'
1/
#27560000000
0!
1"
0'
1(
0/
10
#27570000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#27580000000
0!
0'
0/
#27590000000
1!
1'
1/
#27600000000
0!
0'
0/
#27610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#27620000000
0!
0'
0/
#27630000000
1!
1'
1/
#27640000000
0!
1"
0'
1(
0/
10
#27650000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#27660000000
0!
1$
0'
1+
0/
#27670000000
1!
1'
1/
#27680000000
0!
0'
0/
#27690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#27700000000
0!
0'
0/
#27710000000
1!
1'
1/
#27720000000
0!
0'
0/
#27730000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#27740000000
0!
0'
0/
#27750000000
1!
1'
1/
#27760000000
0!
0'
0/
#27770000000
1!
1'
1/
#27780000000
0!
0'
0/
#27790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#27800000000
0!
0'
0/
#27810000000
1!
1'
1/
#27820000000
0!
0'
0/
#27830000000
1!
1'
1/
#27840000000
0!
0'
0/
#27850000000
1!
1'
1/
#27860000000
0!
0'
0/
#27870000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#27880000000
0!
0'
0/
#27890000000
1!
1'
1/
#27900000000
0!
0'
0/
#27910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#27920000000
0!
0'
0/
#27930000000
1!
1'
1/
#27940000000
0!
0'
0/
#27950000000
#27960000000
1!
1'
1/
#27970000000
0!
0'
0/
#27980000000
1!
1'
1/
#27990000000
0!
1"
0'
1(
0/
10
#28000000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#28010000000
0!
0'
0/
#28020000000
1!
1'
1/
#28030000000
0!
0'
0/
#28040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#28050000000
0!
0'
0/
#28060000000
1!
1'
1/
#28070000000
0!
1"
0'
1(
0/
10
#28080000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#28090000000
0!
1$
0'
1+
0/
#28100000000
1!
1'
1/
#28110000000
0!
0'
0/
#28120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#28130000000
0!
0'
0/
#28140000000
1!
1'
1/
#28150000000
0!
0'
0/
#28160000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#28170000000
0!
0'
0/
#28180000000
1!
1'
1/
#28190000000
0!
0'
0/
#28200000000
1!
1'
1/
#28210000000
0!
0'
0/
#28220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#28230000000
0!
0'
0/
#28240000000
1!
1'
1/
#28250000000
0!
0'
0/
#28260000000
1!
1'
1/
#28270000000
0!
0'
0/
#28280000000
1!
1'
1/
#28290000000
0!
0'
0/
#28300000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#28310000000
0!
0'
0/
#28320000000
1!
1'
1/
#28330000000
0!
0'
0/
#28340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#28350000000
0!
0'
0/
#28360000000
1!
1'
1/
#28370000000
0!
0'
0/
#28380000000
#28390000000
1!
1'
1/
#28400000000
0!
0'
0/
#28410000000
1!
1'
1/
#28420000000
0!
1"
0'
1(
0/
10
#28430000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#28440000000
0!
0'
0/
#28450000000
1!
1'
1/
#28460000000
0!
0'
0/
#28470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#28480000000
0!
0'
0/
#28490000000
1!
1'
1/
#28500000000
0!
1"
0'
1(
0/
10
#28510000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#28520000000
0!
1$
0'
1+
0/
#28530000000
1!
1'
1/
#28540000000
0!
0'
0/
#28550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#28560000000
0!
0'
0/
#28570000000
1!
1'
1/
#28580000000
0!
0'
0/
#28590000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#28600000000
0!
0'
0/
#28610000000
1!
1'
1/
#28620000000
0!
0'
0/
#28630000000
1!
1'
1/
#28640000000
0!
0'
0/
#28650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#28660000000
0!
0'
0/
#28670000000
1!
1'
1/
#28680000000
0!
0'
0/
#28690000000
1!
1'
1/
#28700000000
0!
0'
0/
#28710000000
1!
1'
1/
#28720000000
0!
0'
0/
#28730000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#28740000000
0!
0'
0/
#28750000000
1!
1'
1/
#28760000000
0!
0'
0/
#28770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#28780000000
0!
0'
0/
#28790000000
1!
1'
1/
#28800000000
0!
0'
0/
#28810000000
#28820000000
1!
1'
1/
#28830000000
0!
0'
0/
#28840000000
1!
1'
1/
#28850000000
0!
1"
0'
1(
0/
10
#28860000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#28870000000
0!
0'
0/
#28880000000
1!
1'
1/
#28890000000
0!
0'
0/
#28900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#28910000000
0!
0'
0/
#28920000000
1!
1'
1/
#28930000000
0!
1"
0'
1(
0/
10
#28940000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#28950000000
0!
1$
0'
1+
0/
#28960000000
1!
1'
1/
#28970000000
0!
0'
0/
#28980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#28990000000
0!
0'
0/
#29000000000
1!
1'
1/
#29010000000
0!
0'
0/
#29020000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#29030000000
0!
0'
0/
#29040000000
1!
1'
1/
#29050000000
0!
0'
0/
#29060000000
1!
1'
1/
#29070000000
0!
0'
0/
#29080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#29090000000
0!
0'
0/
#29100000000
1!
1'
1/
#29110000000
0!
0'
0/
#29120000000
1!
1'
1/
#29130000000
0!
0'
0/
#29140000000
1!
1'
1/
#29150000000
0!
0'
0/
#29160000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#29170000000
0!
0'
0/
#29180000000
1!
1'
1/
#29190000000
0!
0'
0/
#29200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#29210000000
0!
0'
0/
#29220000000
1!
1'
1/
#29230000000
0!
0'
0/
#29240000000
#29250000000
1!
1'
1/
#29260000000
0!
0'
0/
#29270000000
1!
1'
1/
#29280000000
0!
1"
0'
1(
0/
10
#29290000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#29300000000
0!
0'
0/
#29310000000
1!
1'
1/
#29320000000
0!
0'
0/
#29330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#29340000000
0!
0'
0/
#29350000000
1!
1'
1/
#29360000000
0!
1"
0'
1(
0/
10
#29370000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#29380000000
0!
1$
0'
1+
0/
#29390000000
1!
1'
1/
#29400000000
0!
0'
0/
#29410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#29420000000
0!
0'
0/
#29430000000
1!
1'
1/
#29440000000
0!
0'
0/
#29450000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#29460000000
0!
0'
0/
#29470000000
1!
1'
1/
#29480000000
0!
0'
0/
#29490000000
1!
1'
1/
#29500000000
0!
0'
0/
#29510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#29520000000
0!
0'
0/
#29530000000
1!
1'
1/
#29540000000
0!
0'
0/
#29550000000
1!
1'
1/
#29560000000
0!
0'
0/
#29570000000
1!
1'
1/
#29580000000
0!
0'
0/
#29590000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#29600000000
0!
0'
0/
#29610000000
1!
1'
1/
#29620000000
0!
0'
0/
#29630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#29640000000
0!
0'
0/
#29650000000
1!
1'
1/
#29660000000
0!
0'
0/
#29670000000
#29680000000
1!
1'
1/
#29690000000
0!
0'
0/
#29700000000
1!
1'
1/
#29710000000
0!
1"
0'
1(
0/
10
#29720000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#29730000000
0!
0'
0/
#29740000000
1!
1'
1/
#29750000000
0!
0'
0/
#29760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#29770000000
0!
0'
0/
#29780000000
1!
1'
1/
#29790000000
0!
1"
0'
1(
0/
10
#29800000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#29810000000
0!
1$
0'
1+
0/
#29820000000
1!
1'
1/
#29830000000
0!
0'
0/
#29840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#29850000000
0!
0'
0/
#29860000000
1!
1'
1/
#29870000000
0!
0'
0/
#29880000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#29890000000
0!
0'
0/
#29900000000
1!
1'
1/
#29910000000
0!
0'
0/
#29920000000
1!
1'
1/
#29930000000
0!
0'
0/
#29940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#29950000000
0!
0'
0/
#29960000000
1!
1'
1/
#29970000000
0!
0'
0/
#29980000000
1!
1'
1/
#29990000000
0!
0'
0/
#30000000000
1!
1'
1/
#30010000000
0!
0'
0/
#30020000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#30030000000
0!
0'
0/
#30040000000
1!
1'
1/
#30050000000
0!
0'
0/
#30060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#30070000000
0!
0'
0/
#30080000000
1!
1'
1/
#30090000000
0!
0'
0/
#30100000000
#30110000000
1!
1'
1/
#30120000000
0!
0'
0/
#30130000000
1!
1'
1/
#30140000000
0!
1"
0'
1(
0/
10
#30150000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#30160000000
0!
0'
0/
#30170000000
1!
1'
1/
#30180000000
0!
0'
0/
#30190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#30200000000
0!
0'
0/
#30210000000
1!
1'
1/
#30220000000
0!
1"
0'
1(
0/
10
#30230000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#30240000000
0!
1$
0'
1+
0/
#30250000000
1!
1'
1/
#30260000000
0!
0'
0/
#30270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#30280000000
0!
0'
0/
#30290000000
1!
1'
1/
#30300000000
0!
0'
0/
#30310000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#30320000000
0!
0'
0/
#30330000000
1!
1'
1/
#30340000000
0!
0'
0/
#30350000000
1!
1'
1/
#30360000000
0!
0'
0/
#30370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#30380000000
0!
0'
0/
#30390000000
1!
1'
1/
#30400000000
0!
0'
0/
#30410000000
1!
1'
1/
#30420000000
0!
0'
0/
#30430000000
1!
1'
1/
#30440000000
0!
0'
0/
#30450000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#30460000000
0!
0'
0/
#30470000000
1!
1'
1/
#30480000000
0!
0'
0/
#30490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#30500000000
0!
0'
0/
#30510000000
1!
1'
1/
#30520000000
0!
0'
0/
#30530000000
#30540000000
1!
1'
1/
#30550000000
0!
0'
0/
#30560000000
1!
1'
1/
#30570000000
0!
1"
0'
1(
0/
10
#30580000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#30590000000
0!
0'
0/
#30600000000
1!
1'
1/
#30610000000
0!
0'
0/
#30620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#30630000000
0!
0'
0/
#30640000000
1!
1'
1/
#30650000000
0!
1"
0'
1(
0/
10
#30660000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#30670000000
0!
1$
0'
1+
0/
#30680000000
1!
1'
1/
#30690000000
0!
0'
0/
#30700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#30710000000
0!
0'
0/
#30720000000
1!
1'
1/
#30730000000
0!
0'
0/
#30740000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#30750000000
0!
0'
0/
#30760000000
1!
1'
1/
#30770000000
0!
0'
0/
#30780000000
1!
1'
1/
#30790000000
0!
0'
0/
#30800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#30810000000
0!
0'
0/
#30820000000
1!
1'
1/
#30830000000
0!
0'
0/
#30840000000
1!
1'
1/
#30850000000
0!
0'
0/
#30860000000
1!
1'
1/
#30870000000
0!
0'
0/
#30880000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#30890000000
0!
0'
0/
#30900000000
1!
1'
1/
#30910000000
0!
0'
0/
#30920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#30930000000
0!
0'
0/
#30940000000
1!
1'
1/
#30950000000
0!
0'
0/
#30960000000
#30970000000
1!
1'
1/
#30980000000
0!
0'
0/
#30990000000
1!
1'
1/
#31000000000
0!
1"
0'
1(
0/
10
#31010000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#31020000000
0!
0'
0/
#31030000000
1!
1'
1/
#31040000000
0!
0'
0/
#31050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#31060000000
0!
0'
0/
#31070000000
1!
1'
1/
#31080000000
0!
1"
0'
1(
0/
10
#31090000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#31100000000
0!
1$
0'
1+
0/
#31110000000
1!
1'
1/
#31120000000
0!
0'
0/
#31130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#31140000000
0!
0'
0/
#31150000000
1!
1'
1/
#31160000000
0!
0'
0/
#31170000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#31180000000
0!
0'
0/
#31190000000
1!
1'
1/
#31200000000
0!
0'
0/
#31210000000
1!
1'
1/
#31220000000
0!
0'
0/
#31230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#31240000000
0!
0'
0/
#31250000000
1!
1'
1/
#31260000000
0!
0'
0/
#31270000000
1!
1'
1/
#31280000000
0!
0'
0/
#31290000000
1!
1'
1/
#31300000000
0!
0'
0/
#31310000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#31320000000
0!
0'
0/
#31330000000
1!
1'
1/
#31340000000
0!
0'
0/
#31350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#31360000000
0!
0'
0/
#31370000000
1!
1'
1/
#31380000000
0!
0'
0/
#31390000000
#31400000000
1!
1'
1/
#31410000000
0!
0'
0/
#31420000000
1!
1'
1/
#31430000000
0!
1"
0'
1(
0/
10
#31440000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#31450000000
0!
0'
0/
#31460000000
1!
1'
1/
#31470000000
0!
0'
0/
#31480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#31490000000
0!
0'
0/
#31500000000
1!
1'
1/
#31510000000
0!
1"
0'
1(
0/
10
#31520000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#31530000000
0!
1$
0'
1+
0/
#31540000000
1!
1'
1/
#31550000000
0!
0'
0/
#31560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#31570000000
0!
0'
0/
#31580000000
1!
1'
1/
#31590000000
0!
0'
0/
#31600000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#31610000000
0!
0'
0/
#31620000000
1!
1'
1/
#31630000000
0!
0'
0/
#31640000000
1!
1'
1/
#31650000000
0!
0'
0/
#31660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#31670000000
0!
0'
0/
#31680000000
1!
1'
1/
#31690000000
0!
0'
0/
#31700000000
1!
1'
1/
#31710000000
0!
0'
0/
#31720000000
1!
1'
1/
#31730000000
0!
0'
0/
#31740000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#31750000000
0!
0'
0/
#31760000000
1!
1'
1/
#31770000000
0!
0'
0/
#31780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#31790000000
0!
0'
0/
#31800000000
1!
1'
1/
#31810000000
0!
0'
0/
#31820000000
#31830000000
1!
1'
1/
#31840000000
0!
0'
0/
#31850000000
1!
1'
1/
#31860000000
0!
1"
0'
1(
0/
10
#31870000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#31880000000
0!
0'
0/
#31890000000
1!
1'
1/
#31900000000
0!
0'
0/
#31910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#31920000000
0!
0'
0/
#31930000000
1!
1'
1/
#31940000000
0!
1"
0'
1(
0/
10
#31950000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#31960000000
0!
1$
0'
1+
0/
#31970000000
1!
1'
1/
#31980000000
0!
0'
0/
#31990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#32000000000
0!
0'
0/
#32010000000
1!
1'
1/
#32020000000
0!
0'
0/
#32030000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#32040000000
0!
0'
0/
#32050000000
1!
1'
1/
#32060000000
0!
0'
0/
#32070000000
1!
1'
1/
#32080000000
0!
0'
0/
#32090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#32100000000
0!
0'
0/
#32110000000
1!
1'
1/
#32120000000
0!
0'
0/
#32130000000
1!
1'
1/
#32140000000
0!
0'
0/
#32150000000
1!
1'
1/
#32160000000
0!
0'
0/
#32170000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#32180000000
0!
0'
0/
#32190000000
1!
1'
1/
#32200000000
0!
0'
0/
#32210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#32220000000
0!
0'
0/
#32230000000
1!
1'
1/
#32240000000
0!
0'
0/
#32250000000
#32260000000
1!
1'
1/
#32270000000
0!
0'
0/
#32280000000
1!
1'
1/
#32290000000
0!
1"
0'
1(
0/
10
#32300000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#32310000000
0!
0'
0/
#32320000000
1!
1'
1/
#32330000000
0!
0'
0/
#32340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#32350000000
0!
0'
0/
#32360000000
1!
1'
1/
#32370000000
0!
1"
0'
1(
0/
10
#32380000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#32390000000
0!
1$
0'
1+
0/
#32400000000
1!
1'
1/
#32410000000
0!
0'
0/
#32420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#32430000000
0!
0'
0/
#32440000000
1!
1'
1/
#32450000000
0!
0'
0/
#32460000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#32470000000
0!
0'
0/
#32480000000
1!
1'
1/
#32490000000
0!
0'
0/
#32500000000
1!
1'
1/
#32510000000
0!
0'
0/
#32520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#32530000000
0!
0'
0/
#32540000000
1!
1'
1/
#32550000000
0!
0'
0/
#32560000000
1!
1'
1/
#32570000000
0!
0'
0/
#32580000000
1!
1'
1/
#32590000000
0!
0'
0/
#32600000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#32610000000
0!
0'
0/
#32620000000
1!
1'
1/
#32630000000
0!
0'
0/
#32640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#32650000000
0!
0'
0/
#32660000000
1!
1'
1/
#32670000000
0!
0'
0/
#32680000000
#32690000000
1!
1'
1/
#32700000000
0!
0'
0/
#32710000000
1!
1'
1/
#32720000000
0!
1"
0'
1(
0/
10
#32730000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#32740000000
0!
0'
0/
#32750000000
1!
1'
1/
#32760000000
0!
0'
0/
#32770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#32780000000
0!
0'
0/
#32790000000
1!
1'
1/
#32800000000
0!
1"
0'
1(
0/
10
#32810000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#32820000000
0!
1$
0'
1+
0/
#32830000000
1!
1'
1/
#32840000000
0!
0'
0/
#32850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#32860000000
0!
0'
0/
#32870000000
1!
1'
1/
#32880000000
0!
0'
0/
#32890000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#32900000000
0!
0'
0/
#32910000000
1!
1'
1/
#32920000000
0!
0'
0/
#32930000000
1!
1'
1/
#32940000000
0!
0'
0/
#32950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#32960000000
0!
0'
0/
#32970000000
1!
1'
1/
#32980000000
0!
0'
0/
#32990000000
1!
1'
1/
#33000000000
0!
0'
0/
#33010000000
1!
1'
1/
#33020000000
0!
0'
0/
#33030000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#33040000000
0!
0'
0/
#33050000000
1!
1'
1/
#33060000000
0!
0'
0/
#33070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#33080000000
0!
0'
0/
#33090000000
1!
1'
1/
#33100000000
0!
0'
0/
#33110000000
#33120000000
1!
1'
1/
#33130000000
0!
0'
0/
#33140000000
1!
1'
1/
#33150000000
0!
1"
0'
1(
0/
10
#33160000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#33170000000
0!
0'
0/
#33180000000
1!
1'
1/
#33190000000
0!
0'
0/
#33200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#33210000000
0!
0'
0/
#33220000000
1!
1'
1/
#33230000000
0!
1"
0'
1(
0/
10
#33240000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#33250000000
0!
1$
0'
1+
0/
#33260000000
1!
1'
1/
#33270000000
0!
0'
0/
#33280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#33290000000
0!
0'
0/
#33300000000
1!
1'
1/
#33310000000
0!
0'
0/
#33320000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#33330000000
0!
0'
0/
#33340000000
1!
1'
1/
#33350000000
0!
0'
0/
#33360000000
1!
1'
1/
#33370000000
0!
0'
0/
#33380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#33390000000
0!
0'
0/
#33400000000
1!
1'
1/
#33410000000
0!
0'
0/
#33420000000
1!
1'
1/
#33430000000
0!
0'
0/
#33440000000
1!
1'
1/
#33450000000
0!
0'
0/
#33460000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#33470000000
0!
0'
0/
#33480000000
1!
1'
1/
#33490000000
0!
0'
0/
#33500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#33510000000
0!
0'
0/
#33520000000
1!
1'
1/
#33530000000
0!
0'
0/
#33540000000
#33550000000
1!
1'
1/
#33560000000
0!
0'
0/
#33570000000
1!
1'
1/
#33580000000
0!
1"
0'
1(
0/
10
#33590000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#33600000000
0!
0'
0/
#33610000000
1!
1'
1/
#33620000000
0!
0'
0/
#33630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#33640000000
0!
0'
0/
#33650000000
1!
1'
1/
#33660000000
0!
1"
0'
1(
0/
10
#33670000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#33680000000
0!
1$
0'
1+
0/
#33690000000
1!
1'
1/
#33700000000
0!
0'
0/
#33710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#33720000000
0!
0'
0/
#33730000000
1!
1'
1/
#33740000000
0!
0'
0/
#33750000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#33760000000
0!
0'
0/
#33770000000
1!
1'
1/
#33780000000
0!
0'
0/
#33790000000
1!
1'
1/
#33800000000
0!
0'
0/
#33810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#33820000000
0!
0'
0/
#33830000000
1!
1'
1/
#33840000000
0!
0'
0/
#33850000000
1!
1'
1/
#33860000000
0!
0'
0/
#33870000000
1!
1'
1/
#33880000000
0!
0'
0/
#33890000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#33900000000
0!
0'
0/
#33910000000
1!
1'
1/
#33920000000
0!
0'
0/
#33930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#33940000000
0!
0'
0/
#33950000000
1!
1'
1/
#33960000000
0!
0'
0/
#33970000000
#33980000000
1!
1'
1/
#33990000000
0!
0'
0/
#34000000000
1!
1'
1/
#34010000000
0!
1"
0'
1(
0/
10
#34020000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#34030000000
0!
0'
0/
#34040000000
1!
1'
1/
#34050000000
0!
0'
0/
#34060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#34070000000
0!
0'
0/
#34080000000
1!
1'
1/
#34090000000
0!
1"
0'
1(
0/
10
#34100000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#34110000000
0!
1$
0'
1+
0/
#34120000000
1!
1'
1/
#34130000000
0!
0'
0/
#34140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#34150000000
0!
0'
0/
#34160000000
1!
1'
1/
#34170000000
0!
0'
0/
#34180000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#34190000000
0!
0'
0/
#34200000000
1!
1'
1/
#34210000000
0!
0'
0/
#34220000000
1!
1'
1/
#34230000000
0!
0'
0/
#34240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#34250000000
0!
0'
0/
#34260000000
1!
1'
1/
#34270000000
0!
0'
0/
#34280000000
1!
1'
1/
#34290000000
0!
0'
0/
#34300000000
1!
1'
1/
#34310000000
0!
0'
0/
#34320000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#34330000000
0!
0'
0/
#34340000000
1!
1'
1/
#34350000000
0!
0'
0/
#34360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#34370000000
0!
0'
0/
#34380000000
1!
1'
1/
#34390000000
0!
0'
0/
#34400000000
#34410000000
1!
1'
1/
#34420000000
0!
0'
0/
#34430000000
1!
1'
1/
#34440000000
0!
1"
0'
1(
0/
10
#34450000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#34460000000
0!
0'
0/
#34470000000
1!
1'
1/
#34480000000
0!
0'
0/
#34490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#34500000000
0!
0'
0/
#34510000000
1!
1'
1/
#34520000000
0!
1"
0'
1(
0/
10
#34530000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#34540000000
0!
1$
0'
1+
0/
#34550000000
1!
1'
1/
#34560000000
0!
0'
0/
#34570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#34580000000
0!
0'
0/
#34590000000
1!
1'
1/
#34600000000
0!
0'
0/
#34610000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#34620000000
0!
0'
0/
#34630000000
1!
1'
1/
#34640000000
0!
0'
0/
#34650000000
1!
1'
1/
#34660000000
0!
0'
0/
#34670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#34680000000
0!
0'
0/
#34690000000
1!
1'
1/
#34700000000
0!
0'
0/
#34710000000
1!
1'
1/
#34720000000
0!
0'
0/
#34730000000
1!
1'
1/
#34740000000
0!
0'
0/
#34750000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#34760000000
0!
0'
0/
#34770000000
1!
1'
1/
#34780000000
0!
0'
0/
#34790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#34800000000
0!
0'
0/
#34810000000
1!
1'
1/
#34820000000
0!
0'
0/
#34830000000
#34840000000
1!
1'
1/
#34850000000
0!
0'
0/
#34860000000
1!
1'
1/
#34870000000
0!
1"
0'
1(
0/
10
#34880000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#34890000000
0!
0'
0/
#34900000000
1!
1'
1/
#34910000000
0!
0'
0/
#34920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#34930000000
0!
0'
0/
#34940000000
1!
1'
1/
#34950000000
0!
1"
0'
1(
0/
10
#34960000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#34970000000
0!
1$
0'
1+
0/
#34980000000
1!
1'
1/
#34990000000
0!
0'
0/
#35000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#35010000000
0!
0'
0/
#35020000000
1!
1'
1/
#35030000000
0!
0'
0/
#35040000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#35050000000
0!
0'
0/
#35060000000
1!
1'
1/
#35070000000
0!
0'
0/
#35080000000
1!
1'
1/
#35090000000
0!
0'
0/
#35100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#35110000000
0!
0'
0/
#35120000000
1!
1'
1/
#35130000000
0!
0'
0/
#35140000000
1!
1'
1/
#35150000000
0!
0'
0/
#35160000000
1!
1'
1/
#35170000000
0!
0'
0/
#35180000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#35190000000
0!
0'
0/
#35200000000
1!
1'
1/
#35210000000
0!
0'
0/
#35220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#35230000000
0!
0'
0/
#35240000000
1!
1'
1/
#35250000000
0!
0'
0/
#35260000000
#35270000000
1!
1'
1/
#35280000000
0!
0'
0/
#35290000000
1!
1'
1/
#35300000000
0!
1"
0'
1(
0/
10
#35310000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#35320000000
0!
0'
0/
#35330000000
1!
1'
1/
#35340000000
0!
0'
0/
#35350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#35360000000
0!
0'
0/
#35370000000
1!
1'
1/
#35380000000
0!
1"
0'
1(
0/
10
#35390000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#35400000000
0!
1$
0'
1+
0/
#35410000000
1!
1'
1/
#35420000000
0!
0'
0/
#35430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#35440000000
0!
0'
0/
#35450000000
1!
1'
1/
#35460000000
0!
0'
0/
#35470000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#35480000000
0!
0'
0/
#35490000000
1!
1'
1/
#35500000000
0!
0'
0/
#35510000000
1!
1'
1/
#35520000000
0!
0'
0/
#35530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#35540000000
0!
0'
0/
#35550000000
1!
1'
1/
#35560000000
0!
0'
0/
#35570000000
1!
1'
1/
#35580000000
0!
0'
0/
#35590000000
1!
1'
1/
#35600000000
0!
0'
0/
#35610000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#35620000000
0!
0'
0/
#35630000000
1!
1'
1/
#35640000000
0!
0'
0/
#35650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#35660000000
0!
0'
0/
#35670000000
1!
1'
1/
#35680000000
0!
0'
0/
#35690000000
#35700000000
1!
1'
1/
#35710000000
0!
0'
0/
#35720000000
1!
1'
1/
#35730000000
0!
1"
0'
1(
0/
10
#35740000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#35750000000
0!
0'
0/
#35760000000
1!
1'
1/
#35770000000
0!
0'
0/
#35780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#35790000000
0!
0'
0/
#35800000000
1!
1'
1/
#35810000000
0!
1"
0'
1(
0/
10
#35820000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#35830000000
0!
1$
0'
1+
0/
#35840000000
1!
1'
1/
#35850000000
0!
0'
0/
#35860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#35870000000
0!
0'
0/
#35880000000
1!
1'
1/
#35890000000
0!
0'
0/
#35900000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#35910000000
0!
0'
0/
#35920000000
1!
1'
1/
#35930000000
0!
0'
0/
#35940000000
1!
1'
1/
#35950000000
0!
0'
0/
#35960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#35970000000
0!
0'
0/
#35980000000
1!
1'
1/
#35990000000
0!
0'
0/
#36000000000
1!
1'
1/
#36010000000
0!
0'
0/
#36020000000
1!
1'
1/
#36030000000
0!
0'
0/
#36040000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#36050000000
0!
0'
0/
#36060000000
1!
1'
1/
#36070000000
0!
0'
0/
#36080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#36090000000
0!
0'
0/
#36100000000
1!
1'
1/
#36110000000
0!
0'
0/
#36120000000
#36130000000
1!
1'
1/
#36140000000
0!
0'
0/
#36150000000
1!
1'
1/
#36160000000
0!
1"
0'
1(
0/
10
#36170000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#36180000000
0!
0'
0/
#36190000000
1!
1'
1/
#36200000000
0!
0'
0/
#36210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#36220000000
0!
0'
0/
#36230000000
1!
1'
1/
#36240000000
0!
1"
0'
1(
0/
10
#36250000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#36260000000
0!
1$
0'
1+
0/
#36270000000
1!
1'
1/
#36280000000
0!
0'
0/
#36290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#36300000000
0!
0'
0/
#36310000000
1!
1'
1/
#36320000000
0!
0'
0/
#36330000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#36340000000
0!
0'
0/
#36350000000
1!
1'
1/
#36360000000
0!
0'
0/
#36370000000
1!
1'
1/
#36380000000
0!
0'
0/
#36390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#36400000000
0!
0'
0/
#36410000000
1!
1'
1/
#36420000000
0!
0'
0/
#36430000000
1!
1'
1/
#36440000000
0!
0'
0/
#36450000000
1!
1'
1/
#36460000000
0!
0'
0/
#36470000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#36480000000
0!
0'
0/
#36490000000
1!
1'
1/
#36500000000
0!
0'
0/
#36510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#36520000000
0!
0'
0/
#36530000000
1!
1'
1/
#36540000000
0!
0'
0/
#36550000000
#36560000000
1!
1'
1/
#36570000000
0!
0'
0/
#36580000000
1!
1'
1/
#36590000000
0!
1"
0'
1(
0/
10
#36600000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#36610000000
0!
0'
0/
#36620000000
1!
1'
1/
#36630000000
0!
0'
0/
#36640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#36650000000
0!
0'
0/
#36660000000
1!
1'
1/
#36670000000
0!
1"
0'
1(
0/
10
#36680000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#36690000000
0!
1$
0'
1+
0/
#36700000000
1!
1'
1/
#36710000000
0!
0'
0/
#36720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#36730000000
0!
0'
0/
#36740000000
1!
1'
1/
#36750000000
0!
0'
0/
#36760000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#36770000000
0!
0'
0/
#36780000000
1!
1'
1/
#36790000000
0!
0'
0/
#36800000000
1!
1'
1/
#36810000000
0!
0'
0/
#36820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#36830000000
0!
0'
0/
#36840000000
1!
1'
1/
#36850000000
0!
0'
0/
#36860000000
1!
1'
1/
#36870000000
0!
0'
0/
#36880000000
1!
1'
1/
#36890000000
0!
0'
0/
#36900000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#36910000000
0!
0'
0/
#36920000000
1!
1'
1/
#36930000000
0!
0'
0/
#36940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#36950000000
0!
0'
0/
#36960000000
1!
1'
1/
#36970000000
0!
0'
0/
#36980000000
#36990000000
1!
1'
1/
#37000000000
0!
0'
0/
#37010000000
1!
1'
1/
#37020000000
0!
1"
0'
1(
0/
10
#37030000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#37040000000
0!
0'
0/
#37050000000
1!
1'
1/
#37060000000
0!
0'
0/
#37070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#37080000000
0!
0'
0/
#37090000000
1!
1'
1/
#37100000000
0!
1"
0'
1(
0/
10
#37110000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#37120000000
0!
1$
0'
1+
0/
#37130000000
1!
1'
1/
#37140000000
0!
0'
0/
#37150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#37160000000
0!
0'
0/
#37170000000
1!
1'
1/
#37180000000
0!
0'
0/
#37190000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#37200000000
0!
0'
0/
#37210000000
1!
1'
1/
#37220000000
0!
0'
0/
#37230000000
1!
1'
1/
#37240000000
0!
0'
0/
#37250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#37260000000
0!
0'
0/
#37270000000
1!
1'
1/
#37280000000
0!
0'
0/
#37290000000
1!
1'
1/
#37300000000
0!
0'
0/
#37310000000
1!
1'
1/
#37320000000
0!
0'
0/
#37330000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#37340000000
0!
0'
0/
#37350000000
1!
1'
1/
#37360000000
0!
0'
0/
#37370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#37380000000
0!
0'
0/
#37390000000
1!
1'
1/
#37400000000
0!
0'
0/
#37410000000
#37420000000
1!
1'
1/
#37430000000
0!
0'
0/
#37440000000
1!
1'
1/
#37450000000
0!
1"
0'
1(
0/
10
#37460000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#37470000000
0!
0'
0/
#37480000000
1!
1'
1/
#37490000000
0!
0'
0/
#37500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#37510000000
0!
0'
0/
#37520000000
1!
1'
1/
#37530000000
0!
1"
0'
1(
0/
10
#37540000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#37550000000
0!
1$
0'
1+
0/
#37560000000
1!
1'
1/
#37570000000
0!
0'
0/
#37580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#37590000000
0!
0'
0/
#37600000000
1!
1'
1/
#37610000000
0!
0'
0/
#37620000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#37630000000
0!
0'
0/
#37640000000
1!
1'
1/
#37650000000
0!
0'
0/
#37660000000
1!
1'
1/
#37670000000
0!
0'
0/
#37680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#37690000000
0!
0'
0/
#37700000000
1!
1'
1/
#37710000000
0!
0'
0/
#37720000000
1!
1'
1/
#37730000000
0!
0'
0/
#37740000000
1!
1'
1/
#37750000000
0!
0'
0/
#37760000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#37770000000
0!
0'
0/
#37780000000
1!
1'
1/
#37790000000
0!
0'
0/
#37800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#37810000000
0!
0'
0/
#37820000000
1!
1'
1/
#37830000000
0!
0'
0/
#37840000000
#37850000000
1!
1'
1/
#37860000000
0!
0'
0/
#37870000000
1!
1'
1/
#37880000000
0!
1"
0'
1(
0/
10
#37890000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#37900000000
0!
0'
0/
#37910000000
1!
1'
1/
#37920000000
0!
0'
0/
#37930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#37940000000
0!
0'
0/
#37950000000
1!
1'
1/
#37960000000
0!
1"
0'
1(
0/
10
#37970000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#37980000000
0!
1$
0'
1+
0/
#37990000000
1!
1'
1/
#38000000000
0!
0'
0/
#38010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#38020000000
0!
0'
0/
#38030000000
1!
1'
1/
#38040000000
0!
0'
0/
#38050000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#38060000000
0!
0'
0/
#38070000000
1!
1'
1/
#38080000000
0!
0'
0/
#38090000000
1!
1'
1/
#38100000000
0!
0'
0/
#38110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#38120000000
0!
0'
0/
#38130000000
1!
1'
1/
#38140000000
0!
0'
0/
#38150000000
1!
1'
1/
#38160000000
0!
0'
0/
#38170000000
1!
1'
1/
#38180000000
0!
0'
0/
#38190000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#38200000000
0!
0'
0/
#38210000000
1!
1'
1/
#38220000000
0!
0'
0/
#38230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#38240000000
0!
0'
0/
#38250000000
1!
1'
1/
#38260000000
0!
0'
0/
#38270000000
#38280000000
1!
1'
1/
#38290000000
0!
0'
0/
#38300000000
1!
1'
1/
#38310000000
0!
1"
0'
1(
0/
10
#38320000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#38330000000
0!
0'
0/
#38340000000
1!
1'
1/
#38350000000
0!
0'
0/
#38360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#38370000000
0!
0'
0/
#38380000000
1!
1'
1/
#38390000000
0!
1"
0'
1(
0/
10
#38400000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#38410000000
0!
1$
0'
1+
0/
#38420000000
1!
1'
1/
#38430000000
0!
0'
0/
#38440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#38450000000
0!
0'
0/
#38460000000
1!
1'
1/
#38470000000
0!
0'
0/
#38480000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#38490000000
0!
0'
0/
#38500000000
1!
1'
1/
#38510000000
0!
0'
0/
#38520000000
1!
1'
1/
#38530000000
0!
0'
0/
#38540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#38550000000
0!
0'
0/
#38560000000
1!
1'
1/
#38570000000
0!
0'
0/
#38580000000
1!
1'
1/
#38590000000
0!
0'
0/
#38600000000
1!
1'
1/
#38610000000
0!
0'
0/
#38620000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#38630000000
0!
0'
0/
#38640000000
1!
1'
1/
#38650000000
0!
0'
0/
#38660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#38670000000
0!
0'
0/
#38680000000
1!
1'
1/
#38690000000
0!
0'
0/
#38700000000
#38710000000
1!
1'
1/
#38720000000
0!
0'
0/
#38730000000
1!
1'
1/
#38740000000
0!
1"
0'
1(
0/
10
#38750000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#38760000000
0!
0'
0/
#38770000000
1!
1'
1/
#38780000000
0!
0'
0/
#38790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#38800000000
0!
0'
0/
#38810000000
1!
1'
1/
#38820000000
0!
1"
0'
1(
0/
10
#38830000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#38840000000
0!
1$
0'
1+
0/
#38850000000
1!
1'
1/
#38860000000
0!
0'
0/
#38870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#38880000000
0!
0'
0/
#38890000000
1!
1'
1/
#38900000000
0!
0'
0/
#38910000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#38920000000
0!
0'
0/
#38930000000
1!
1'
1/
#38940000000
0!
0'
0/
#38950000000
1!
1'
1/
#38960000000
0!
0'
0/
#38970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#38980000000
0!
0'
0/
#38990000000
1!
1'
1/
#39000000000
0!
0'
0/
#39010000000
1!
1'
1/
#39020000000
0!
0'
0/
#39030000000
1!
1'
1/
#39040000000
0!
0'
0/
#39050000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#39060000000
0!
0'
0/
#39070000000
1!
1'
1/
#39080000000
0!
0'
0/
#39090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#39100000000
0!
0'
0/
#39110000000
1!
1'
1/
#39120000000
0!
0'
0/
#39130000000
#39140000000
1!
1'
1/
#39150000000
0!
0'
0/
#39160000000
1!
1'
1/
#39170000000
0!
1"
0'
1(
0/
10
#39180000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#39190000000
0!
0'
0/
#39200000000
1!
1'
1/
#39210000000
0!
0'
0/
#39220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#39230000000
0!
0'
0/
#39240000000
1!
1'
1/
#39250000000
0!
1"
0'
1(
0/
10
#39260000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#39270000000
0!
1$
0'
1+
0/
#39280000000
1!
1'
1/
#39290000000
0!
0'
0/
#39300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#39310000000
0!
0'
0/
#39320000000
1!
1'
1/
#39330000000
0!
0'
0/
#39340000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#39350000000
0!
0'
0/
#39360000000
1!
1'
1/
#39370000000
0!
0'
0/
#39380000000
1!
1'
1/
#39390000000
0!
0'
0/
#39400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#39410000000
0!
0'
0/
#39420000000
1!
1'
1/
#39430000000
0!
0'
0/
#39440000000
1!
1'
1/
#39450000000
0!
0'
0/
#39460000000
1!
1'
1/
#39470000000
0!
0'
0/
#39480000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#39490000000
0!
0'
0/
#39500000000
1!
1'
1/
#39510000000
0!
0'
0/
#39520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#39530000000
0!
0'
0/
#39540000000
1!
1'
1/
#39550000000
0!
0'
0/
#39560000000
#39570000000
1!
1'
1/
#39580000000
0!
0'
0/
#39590000000
1!
1'
1/
#39600000000
0!
1"
0'
1(
0/
10
#39610000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#39620000000
0!
0'
0/
#39630000000
1!
1'
1/
#39640000000
0!
0'
0/
#39650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#39660000000
0!
0'
0/
#39670000000
1!
1'
1/
#39680000000
0!
1"
0'
1(
0/
10
#39690000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#39700000000
0!
1$
0'
1+
0/
#39710000000
1!
1'
1/
#39720000000
0!
0'
0/
#39730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#39740000000
0!
0'
0/
#39750000000
1!
1'
1/
#39760000000
0!
0'
0/
#39770000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#39780000000
0!
0'
0/
#39790000000
1!
1'
1/
#39800000000
0!
0'
0/
#39810000000
1!
1'
1/
#39820000000
0!
0'
0/
#39830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#39840000000
0!
0'
0/
#39850000000
1!
1'
1/
#39860000000
0!
0'
0/
#39870000000
1!
1'
1/
#39880000000
0!
0'
0/
#39890000000
1!
1'
1/
#39900000000
0!
0'
0/
#39910000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#39920000000
0!
0'
0/
#39930000000
1!
1'
1/
#39940000000
0!
0'
0/
#39950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#39960000000
0!
0'
0/
#39970000000
1!
1'
1/
#39980000000
0!
0'
0/
#39990000000
#40000000000
1!
1'
1/
#40010000000
0!
0'
0/
#40020000000
1!
1'
1/
#40030000000
0!
1"
0'
1(
0/
10
#40040000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#40050000000
0!
0'
0/
#40060000000
1!
1'
1/
#40070000000
0!
0'
0/
#40080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#40090000000
0!
0'
0/
#40100000000
1!
1'
1/
#40110000000
0!
1"
0'
1(
0/
10
#40120000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#40130000000
0!
1$
0'
1+
0/
#40140000000
1!
1'
1/
#40150000000
0!
0'
0/
#40160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#40170000000
0!
0'
0/
#40180000000
1!
1'
1/
#40190000000
0!
0'
0/
#40200000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#40210000000
0!
0'
0/
#40220000000
1!
1'
1/
#40230000000
0!
0'
0/
#40240000000
1!
1'
1/
#40250000000
0!
0'
0/
#40260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#40270000000
0!
0'
0/
#40280000000
1!
1'
1/
#40290000000
0!
0'
0/
#40300000000
1!
1'
1/
#40310000000
0!
0'
0/
#40320000000
1!
1'
1/
#40330000000
0!
0'
0/
#40340000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#40350000000
0!
0'
0/
#40360000000
1!
1'
1/
#40370000000
0!
0'
0/
#40380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#40390000000
0!
0'
0/
#40400000000
1!
1'
1/
#40410000000
0!
0'
0/
#40420000000
#40430000000
1!
1'
1/
#40440000000
0!
0'
0/
#40450000000
1!
1'
1/
#40460000000
0!
1"
0'
1(
0/
10
#40470000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#40480000000
0!
0'
0/
#40490000000
1!
1'
1/
#40500000000
0!
0'
0/
#40510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#40520000000
0!
0'
0/
#40530000000
1!
1'
1/
#40540000000
0!
1"
0'
1(
0/
10
#40550000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#40560000000
0!
1$
0'
1+
0/
#40570000000
1!
1'
1/
#40580000000
0!
0'
0/
#40590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#40600000000
0!
0'
0/
#40610000000
1!
1'
1/
#40620000000
0!
0'
0/
#40630000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#40640000000
0!
0'
0/
#40650000000
1!
1'
1/
#40660000000
0!
0'
0/
#40670000000
1!
1'
1/
#40680000000
0!
0'
0/
#40690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#40700000000
0!
0'
0/
#40710000000
1!
1'
1/
#40720000000
0!
0'
0/
#40730000000
1!
1'
1/
#40740000000
0!
0'
0/
#40750000000
1!
1'
1/
#40760000000
0!
0'
0/
#40770000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#40780000000
0!
0'
0/
#40790000000
1!
1'
1/
#40800000000
0!
0'
0/
#40810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#40820000000
0!
0'
0/
#40830000000
1!
1'
1/
#40840000000
0!
0'
0/
#40850000000
#40860000000
1!
1'
1/
#40870000000
0!
0'
0/
#40880000000
1!
1'
1/
#40890000000
0!
1"
0'
1(
0/
10
#40900000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#40910000000
0!
0'
0/
#40920000000
1!
1'
1/
#40930000000
0!
0'
0/
#40940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#40950000000
0!
0'
0/
#40960000000
1!
1'
1/
#40970000000
0!
1"
0'
1(
0/
10
#40980000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#40990000000
0!
1$
0'
1+
0/
#41000000000
1!
1'
1/
#41010000000
0!
0'
0/
#41020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#41030000000
0!
0'
0/
#41040000000
1!
1'
1/
#41050000000
0!
0'
0/
#41060000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#41070000000
0!
0'
0/
#41080000000
1!
1'
1/
#41090000000
0!
0'
0/
#41100000000
1!
1'
1/
#41110000000
0!
0'
0/
#41120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#41130000000
0!
0'
0/
#41140000000
1!
1'
1/
#41150000000
0!
0'
0/
#41160000000
1!
1'
1/
#41170000000
0!
0'
0/
#41180000000
1!
1'
1/
#41190000000
0!
0'
0/
#41200000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#41210000000
0!
0'
0/
#41220000000
1!
1'
1/
#41230000000
0!
0'
0/
#41240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#41250000000
0!
0'
0/
#41260000000
1!
1'
1/
#41270000000
0!
0'
0/
#41280000000
#41290000000
1!
1'
1/
#41300000000
0!
0'
0/
#41310000000
1!
1'
1/
#41320000000
0!
1"
0'
1(
0/
10
#41330000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#41340000000
0!
0'
0/
#41350000000
1!
1'
1/
#41360000000
0!
0'
0/
#41370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#41380000000
0!
0'
0/
#41390000000
1!
1'
1/
#41400000000
0!
1"
0'
1(
0/
10
#41410000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#41420000000
0!
1$
0'
1+
0/
#41430000000
1!
1'
1/
#41440000000
0!
0'
0/
#41450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#41460000000
0!
0'
0/
#41470000000
1!
1'
1/
#41480000000
0!
0'
0/
#41490000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#41500000000
0!
0'
0/
#41510000000
1!
1'
1/
#41520000000
0!
0'
0/
#41530000000
1!
1'
1/
#41540000000
0!
0'
0/
#41550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#41560000000
0!
0'
0/
#41570000000
1!
1'
1/
#41580000000
0!
0'
0/
#41590000000
1!
1'
1/
#41600000000
0!
0'
0/
#41610000000
1!
1'
1/
#41620000000
0!
0'
0/
#41630000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#41640000000
0!
0'
0/
#41650000000
1!
1'
1/
#41660000000
0!
0'
0/
#41670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#41680000000
0!
0'
0/
#41690000000
1!
1'
1/
#41700000000
0!
0'
0/
#41710000000
#41720000000
1!
1'
1/
#41730000000
0!
0'
0/
#41740000000
1!
1'
1/
#41750000000
0!
1"
0'
1(
0/
10
#41760000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#41770000000
0!
0'
0/
#41780000000
1!
1'
1/
#41790000000
0!
0'
0/
#41800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#41810000000
0!
0'
0/
#41820000000
1!
1'
1/
#41830000000
0!
1"
0'
1(
0/
10
#41840000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#41850000000
0!
1$
0'
1+
0/
#41860000000
1!
1'
1/
#41870000000
0!
0'
0/
#41880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#41890000000
0!
0'
0/
#41900000000
1!
1'
1/
#41910000000
0!
0'
0/
#41920000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#41930000000
0!
0'
0/
#41940000000
1!
1'
1/
#41950000000
0!
0'
0/
#41960000000
1!
1'
1/
#41970000000
0!
0'
0/
#41980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#41990000000
0!
0'
0/
#42000000000
1!
1'
1/
#42010000000
0!
0'
0/
#42020000000
1!
1'
1/
#42030000000
0!
0'
0/
#42040000000
1!
1'
1/
#42050000000
0!
0'
0/
#42060000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#42070000000
0!
0'
0/
#42080000000
1!
1'
1/
#42090000000
0!
0'
0/
#42100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#42110000000
0!
0'
0/
#42120000000
1!
1'
1/
#42130000000
0!
0'
0/
#42140000000
#42150000000
1!
1'
1/
#42160000000
0!
0'
0/
#42170000000
1!
1'
1/
#42180000000
0!
1"
0'
1(
0/
10
#42190000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#42200000000
0!
0'
0/
#42210000000
1!
1'
1/
#42220000000
0!
0'
0/
#42230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#42240000000
0!
0'
0/
#42250000000
1!
1'
1/
#42260000000
0!
1"
0'
1(
0/
10
#42270000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#42280000000
0!
1$
0'
1+
0/
#42290000000
1!
1'
1/
#42300000000
0!
0'
0/
#42310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#42320000000
0!
0'
0/
#42330000000
1!
1'
1/
#42340000000
0!
0'
0/
#42350000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#42360000000
0!
0'
0/
#42370000000
1!
1'
1/
#42380000000
0!
0'
0/
#42390000000
1!
1'
1/
#42400000000
0!
0'
0/
#42410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#42420000000
0!
0'
0/
#42430000000
1!
1'
1/
#42440000000
0!
0'
0/
#42450000000
1!
1'
1/
#42460000000
0!
0'
0/
#42470000000
1!
1'
1/
#42480000000
0!
0'
0/
#42490000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#42500000000
0!
0'
0/
#42510000000
1!
1'
1/
#42520000000
0!
0'
0/
#42530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#42540000000
0!
0'
0/
#42550000000
1!
1'
1/
#42560000000
0!
0'
0/
#42570000000
#42580000000
1!
1'
1/
#42590000000
0!
0'
0/
#42600000000
1!
1'
1/
#42610000000
0!
1"
0'
1(
0/
10
#42620000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#42630000000
0!
0'
0/
#42640000000
1!
1'
1/
#42650000000
0!
0'
0/
#42660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#42670000000
0!
0'
0/
#42680000000
1!
1'
1/
#42690000000
0!
1"
0'
1(
0/
10
#42700000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#42710000000
0!
1$
0'
1+
0/
#42720000000
1!
1'
1/
#42730000000
0!
0'
0/
#42740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#42750000000
0!
0'
0/
#42760000000
1!
1'
1/
#42770000000
0!
0'
0/
#42780000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#42790000000
0!
0'
0/
#42800000000
1!
1'
1/
#42810000000
0!
0'
0/
#42820000000
1!
1'
1/
#42830000000
0!
0'
0/
#42840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#42850000000
0!
0'
0/
#42860000000
1!
1'
1/
#42870000000
0!
0'
0/
#42880000000
1!
1'
1/
#42890000000
0!
0'
0/
#42900000000
1!
1'
1/
#42910000000
0!
0'
0/
#42920000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#42930000000
0!
0'
0/
#42940000000
1!
1'
1/
#42950000000
0!
0'
0/
#42960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#42970000000
0!
0'
0/
#42980000000
1!
1'
1/
#42990000000
0!
0'
0/
#43000000000
#43010000000
1!
1'
1/
#43020000000
0!
0'
0/
#43030000000
1!
1'
1/
#43040000000
0!
1"
0'
1(
0/
10
#43050000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#43060000000
0!
0'
0/
#43070000000
1!
1'
1/
#43080000000
0!
0'
0/
#43090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#43100000000
0!
0'
0/
#43110000000
1!
1'
1/
#43120000000
0!
1"
0'
1(
0/
10
#43130000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#43140000000
0!
1$
0'
1+
0/
#43150000000
1!
1'
1/
#43160000000
0!
0'
0/
#43170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#43180000000
0!
0'
0/
#43190000000
1!
1'
1/
#43200000000
0!
0'
0/
#43210000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#43220000000
0!
0'
0/
#43230000000
1!
1'
1/
#43240000000
0!
0'
0/
#43250000000
1!
1'
1/
#43260000000
0!
0'
0/
#43270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#43280000000
0!
0'
0/
#43290000000
1!
1'
1/
#43300000000
0!
0'
0/
#43310000000
1!
1'
1/
#43320000000
0!
0'
0/
#43330000000
1!
1'
1/
#43340000000
0!
0'
0/
#43350000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#43360000000
0!
0'
0/
#43370000000
1!
1'
1/
#43380000000
0!
0'
0/
#43390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#43400000000
0!
0'
0/
#43410000000
1!
1'
1/
#43420000000
0!
0'
0/
#43430000000
#43440000000
1!
1'
1/
#43450000000
0!
0'
0/
#43460000000
1!
1'
1/
#43470000000
0!
1"
0'
1(
0/
10
#43480000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#43490000000
0!
0'
0/
#43500000000
1!
1'
1/
#43510000000
0!
0'
0/
#43520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#43530000000
0!
0'
0/
#43540000000
1!
1'
1/
#43550000000
0!
1"
0'
1(
0/
10
#43560000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#43570000000
0!
1$
0'
1+
0/
#43580000000
1!
1'
1/
#43590000000
0!
0'
0/
#43600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#43610000000
0!
0'
0/
#43620000000
1!
1'
1/
#43630000000
0!
0'
0/
#43640000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#43650000000
0!
0'
0/
#43660000000
1!
1'
1/
#43670000000
0!
0'
0/
#43680000000
1!
1'
1/
#43690000000
0!
0'
0/
#43700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#43710000000
0!
0'
0/
#43720000000
1!
1'
1/
#43730000000
0!
0'
0/
#43740000000
1!
1'
1/
#43750000000
0!
0'
0/
#43760000000
1!
1'
1/
#43770000000
0!
0'
0/
#43780000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#43790000000
0!
0'
0/
#43800000000
1!
1'
1/
#43810000000
0!
0'
0/
#43820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#43830000000
0!
0'
0/
#43840000000
1!
1'
1/
#43850000000
0!
0'
0/
#43860000000
#43870000000
1!
1'
1/
#43880000000
0!
0'
0/
#43890000000
1!
1'
1/
#43900000000
0!
1"
0'
1(
0/
10
#43910000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#43920000000
0!
0'
0/
#43930000000
1!
1'
1/
#43940000000
0!
0'
0/
#43950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#43960000000
0!
0'
0/
#43970000000
1!
1'
1/
#43980000000
0!
1"
0'
1(
0/
10
#43990000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#44000000000
0!
1$
0'
1+
0/
#44010000000
1!
1'
1/
#44020000000
0!
0'
0/
#44030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#44040000000
0!
0'
0/
#44050000000
1!
1'
1/
#44060000000
0!
0'
0/
#44070000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#44080000000
0!
0'
0/
#44090000000
1!
1'
1/
#44100000000
0!
0'
0/
#44110000000
1!
1'
1/
#44120000000
0!
0'
0/
#44130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#44140000000
0!
0'
0/
#44150000000
1!
1'
1/
#44160000000
0!
0'
0/
#44170000000
1!
1'
1/
#44180000000
0!
0'
0/
#44190000000
1!
1'
1/
#44200000000
0!
0'
0/
#44210000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#44220000000
0!
0'
0/
#44230000000
1!
1'
1/
#44240000000
0!
0'
0/
#44250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#44260000000
0!
0'
0/
#44270000000
1!
1'
1/
#44280000000
0!
0'
0/
#44290000000
#44300000000
1!
1'
1/
#44310000000
0!
0'
0/
#44320000000
1!
1'
1/
#44330000000
0!
1"
0'
1(
0/
10
#44340000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#44350000000
0!
0'
0/
#44360000000
1!
1'
1/
#44370000000
0!
0'
0/
#44380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#44390000000
0!
0'
0/
#44400000000
1!
1'
1/
#44410000000
0!
1"
0'
1(
0/
10
#44420000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#44430000000
0!
1$
0'
1+
0/
#44440000000
1!
1'
1/
#44450000000
0!
0'
0/
#44460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#44470000000
0!
0'
0/
#44480000000
1!
1'
1/
#44490000000
0!
0'
0/
#44500000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#44510000000
0!
0'
0/
#44520000000
1!
1'
1/
#44530000000
0!
0'
0/
#44540000000
1!
1'
1/
#44550000000
0!
0'
0/
#44560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#44570000000
0!
0'
0/
#44580000000
1!
1'
1/
#44590000000
0!
0'
0/
#44600000000
1!
1'
1/
#44610000000
0!
0'
0/
#44620000000
1!
1'
1/
#44630000000
0!
0'
0/
#44640000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#44650000000
0!
0'
0/
#44660000000
1!
1'
1/
#44670000000
0!
0'
0/
#44680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#44690000000
0!
0'
0/
#44700000000
1!
1'
1/
#44710000000
0!
0'
0/
#44720000000
#44730000000
1!
1'
1/
#44740000000
0!
0'
0/
#44750000000
1!
1'
1/
#44760000000
0!
1"
0'
1(
0/
10
#44770000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#44780000000
0!
0'
0/
#44790000000
1!
1'
1/
#44800000000
0!
0'
0/
#44810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#44820000000
0!
0'
0/
#44830000000
1!
1'
1/
#44840000000
0!
1"
0'
1(
0/
10
#44850000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#44860000000
0!
1$
0'
1+
0/
#44870000000
1!
1'
1/
#44880000000
0!
0'
0/
#44890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#44900000000
0!
0'
0/
#44910000000
1!
1'
1/
#44920000000
0!
0'
0/
#44930000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#44940000000
0!
0'
0/
#44950000000
1!
1'
1/
#44960000000
0!
0'
0/
#44970000000
1!
1'
1/
#44980000000
0!
0'
0/
#44990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#45000000000
0!
0'
0/
#45010000000
1!
1'
1/
#45020000000
0!
0'
0/
#45030000000
1!
1'
1/
#45040000000
0!
0'
0/
#45050000000
1!
1'
1/
#45060000000
0!
0'
0/
#45070000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#45080000000
0!
0'
0/
#45090000000
1!
1'
1/
#45100000000
0!
0'
0/
#45110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#45120000000
0!
0'
0/
#45130000000
1!
1'
1/
#45140000000
0!
0'
0/
#45150000000
#45160000000
1!
1'
1/
#45170000000
0!
0'
0/
#45180000000
1!
1'
1/
#45190000000
0!
1"
0'
1(
0/
10
#45200000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#45210000000
0!
0'
0/
#45220000000
1!
1'
1/
#45230000000
0!
0'
0/
#45240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#45250000000
0!
0'
0/
#45260000000
1!
1'
1/
#45270000000
0!
1"
0'
1(
0/
10
#45280000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#45290000000
0!
1$
0'
1+
0/
#45300000000
1!
1'
1/
#45310000000
0!
0'
0/
#45320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#45330000000
0!
0'
0/
#45340000000
1!
1'
1/
#45350000000
0!
0'
0/
#45360000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#45370000000
0!
0'
0/
#45380000000
1!
1'
1/
#45390000000
0!
0'
0/
#45400000000
1!
1'
1/
#45410000000
0!
0'
0/
#45420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#45430000000
0!
0'
0/
#45440000000
1!
1'
1/
#45450000000
0!
0'
0/
#45460000000
1!
1'
1/
#45470000000
0!
0'
0/
#45480000000
1!
1'
1/
#45490000000
0!
0'
0/
#45500000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#45510000000
0!
0'
0/
#45520000000
1!
1'
1/
#45530000000
0!
0'
0/
#45540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#45550000000
0!
0'
0/
#45560000000
1!
1'
1/
#45570000000
0!
0'
0/
#45580000000
#45590000000
1!
1'
1/
#45600000000
0!
0'
0/
#45610000000
1!
1'
1/
#45620000000
0!
1"
0'
1(
0/
10
#45630000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#45640000000
0!
0'
0/
#45650000000
1!
1'
1/
#45660000000
0!
0'
0/
#45670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#45680000000
0!
0'
0/
#45690000000
1!
1'
1/
#45700000000
0!
1"
0'
1(
0/
10
#45710000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#45720000000
0!
1$
0'
1+
0/
#45730000000
1!
1'
1/
#45740000000
0!
0'
0/
#45750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#45760000000
0!
0'
0/
#45770000000
1!
1'
1/
#45780000000
0!
0'
0/
#45790000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#45800000000
0!
0'
0/
#45810000000
1!
1'
1/
#45820000000
0!
0'
0/
#45830000000
1!
1'
1/
#45840000000
0!
0'
0/
#45850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#45860000000
0!
0'
0/
#45870000000
1!
1'
1/
#45880000000
0!
0'
0/
#45890000000
1!
1'
1/
#45900000000
0!
0'
0/
#45910000000
1!
1'
1/
#45920000000
0!
0'
0/
#45930000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#45940000000
0!
0'
0/
#45950000000
1!
1'
1/
#45960000000
0!
0'
0/
#45970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#45980000000
0!
0'
0/
#45990000000
1!
1'
1/
#46000000000
0!
0'
0/
#46010000000
#46020000000
1!
1'
1/
#46030000000
0!
0'
0/
#46040000000
1!
1'
1/
#46050000000
0!
1"
0'
1(
0/
10
#46060000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#46070000000
0!
0'
0/
#46080000000
1!
1'
1/
#46090000000
0!
0'
0/
#46100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#46110000000
0!
0'
0/
#46120000000
1!
1'
1/
#46130000000
0!
1"
0'
1(
0/
10
#46140000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#46150000000
0!
1$
0'
1+
0/
#46160000000
1!
1'
1/
#46170000000
0!
0'
0/
#46180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#46190000000
0!
0'
0/
#46200000000
1!
1'
1/
#46210000000
0!
0'
0/
#46220000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#46230000000
0!
0'
0/
#46240000000
1!
1'
1/
#46250000000
0!
0'
0/
#46260000000
1!
1'
1/
#46270000000
0!
0'
0/
#46280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#46290000000
0!
0'
0/
#46300000000
1!
1'
1/
#46310000000
0!
0'
0/
#46320000000
1!
1'
1/
#46330000000
0!
0'
0/
#46340000000
1!
1'
1/
#46350000000
0!
0'
0/
#46360000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#46370000000
0!
0'
0/
#46380000000
1!
1'
1/
#46390000000
0!
0'
0/
#46400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#46410000000
0!
0'
0/
#46420000000
1!
1'
1/
#46430000000
0!
0'
0/
#46440000000
#46450000000
1!
1'
1/
#46460000000
0!
0'
0/
#46470000000
1!
1'
1/
#46480000000
0!
1"
0'
1(
0/
10
#46490000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#46500000000
0!
0'
0/
#46510000000
1!
1'
1/
#46520000000
0!
0'
0/
#46530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#46540000000
0!
0'
0/
#46550000000
1!
1'
1/
#46560000000
0!
1"
0'
1(
0/
10
#46570000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#46580000000
0!
1$
0'
1+
0/
#46590000000
1!
1'
1/
#46600000000
0!
0'
0/
#46610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#46620000000
0!
0'
0/
#46630000000
1!
1'
1/
#46640000000
0!
0'
0/
#46650000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#46660000000
0!
0'
0/
#46670000000
1!
1'
1/
#46680000000
0!
0'
0/
#46690000000
1!
1'
1/
#46700000000
0!
0'
0/
#46710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#46720000000
0!
0'
0/
#46730000000
1!
1'
1/
#46740000000
0!
0'
0/
#46750000000
1!
1'
1/
#46760000000
0!
0'
0/
#46770000000
1!
1'
1/
#46780000000
0!
0'
0/
#46790000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#46800000000
0!
0'
0/
#46810000000
1!
1'
1/
#46820000000
0!
0'
0/
#46830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#46840000000
0!
0'
0/
#46850000000
1!
1'
1/
#46860000000
0!
0'
0/
#46870000000
#46880000000
1!
1'
1/
#46890000000
0!
0'
0/
#46900000000
1!
1'
1/
#46910000000
0!
1"
0'
1(
0/
10
#46920000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#46930000000
0!
0'
0/
#46940000000
1!
1'
1/
#46950000000
0!
0'
0/
#46960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#46970000000
0!
0'
0/
#46980000000
1!
1'
1/
#46990000000
0!
1"
0'
1(
0/
10
#47000000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#47010000000
0!
1$
0'
1+
0/
#47020000000
1!
1'
1/
#47030000000
0!
0'
0/
#47040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#47050000000
0!
0'
0/
#47060000000
1!
1'
1/
#47070000000
0!
0'
0/
#47080000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#47090000000
0!
0'
0/
#47100000000
1!
1'
1/
#47110000000
0!
0'
0/
#47120000000
1!
1'
1/
#47130000000
0!
0'
0/
#47140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#47150000000
0!
0'
0/
#47160000000
1!
1'
1/
#47170000000
0!
0'
0/
#47180000000
1!
1'
1/
#47190000000
0!
0'
0/
#47200000000
1!
1'
1/
#47210000000
0!
0'
0/
#47220000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#47230000000
0!
0'
0/
#47240000000
1!
1'
1/
#47250000000
0!
0'
0/
#47260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#47270000000
0!
0'
0/
#47280000000
1!
1'
1/
#47290000000
0!
0'
0/
#47300000000
#47310000000
1!
1'
1/
#47320000000
0!
0'
0/
#47330000000
1!
1'
1/
#47340000000
0!
1"
0'
1(
0/
10
#47350000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#47360000000
0!
0'
0/
#47370000000
1!
1'
1/
#47380000000
0!
0'
0/
#47390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#47400000000
0!
0'
0/
#47410000000
1!
1'
1/
#47420000000
0!
1"
0'
1(
0/
10
#47430000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#47440000000
0!
1$
0'
1+
0/
#47450000000
1!
1'
1/
#47460000000
0!
0'
0/
#47470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#47480000000
0!
0'
0/
#47490000000
1!
1'
1/
#47500000000
0!
0'
0/
#47510000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#47520000000
0!
0'
0/
#47530000000
1!
1'
1/
#47540000000
0!
0'
0/
#47550000000
1!
1'
1/
#47560000000
0!
0'
0/
#47570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#47580000000
0!
0'
0/
#47590000000
1!
1'
1/
#47600000000
0!
0'
0/
#47610000000
1!
1'
1/
#47620000000
0!
0'
0/
#47630000000
1!
1'
1/
#47640000000
0!
0'
0/
#47650000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#47660000000
0!
0'
0/
#47670000000
1!
1'
1/
#47680000000
0!
0'
0/
#47690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#47700000000
0!
0'
0/
#47710000000
1!
1'
1/
#47720000000
0!
0'
0/
#47730000000
#47740000000
1!
1'
1/
#47750000000
0!
0'
0/
#47760000000
1!
1'
1/
#47770000000
0!
1"
0'
1(
0/
10
#47780000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#47790000000
0!
0'
0/
#47800000000
1!
1'
1/
#47810000000
0!
0'
0/
#47820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#47830000000
0!
0'
0/
#47840000000
1!
1'
1/
#47850000000
0!
1"
0'
1(
0/
10
#47860000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#47870000000
0!
1$
0'
1+
0/
#47880000000
1!
1'
1/
#47890000000
0!
0'
0/
#47900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#47910000000
0!
0'
0/
#47920000000
1!
1'
1/
#47930000000
0!
0'
0/
#47940000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#47950000000
0!
0'
0/
#47960000000
1!
1'
1/
#47970000000
0!
0'
0/
#47980000000
1!
1'
1/
#47990000000
0!
0'
0/
#48000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#48010000000
0!
0'
0/
#48020000000
1!
1'
1/
#48030000000
0!
0'
0/
#48040000000
1!
1'
1/
#48050000000
0!
0'
0/
#48060000000
1!
1'
1/
#48070000000
0!
0'
0/
#48080000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#48090000000
0!
0'
0/
#48100000000
1!
1'
1/
#48110000000
0!
0'
0/
#48120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#48130000000
0!
0'
0/
#48140000000
1!
1'
1/
#48150000000
0!
0'
0/
#48160000000
#48170000000
1!
1'
1/
#48180000000
0!
0'
0/
#48190000000
1!
1'
1/
#48200000000
0!
1"
0'
1(
0/
10
#48210000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#48220000000
0!
0'
0/
#48230000000
1!
1'
1/
#48240000000
0!
0'
0/
#48250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#48260000000
0!
0'
0/
#48270000000
1!
1'
1/
#48280000000
0!
1"
0'
1(
0/
10
#48290000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#48300000000
0!
1$
0'
1+
0/
#48310000000
1!
1'
1/
#48320000000
0!
0'
0/
#48330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#48340000000
0!
0'
0/
#48350000000
1!
1'
1/
#48360000000
0!
0'
0/
#48370000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#48380000000
0!
0'
0/
#48390000000
1!
1'
1/
#48400000000
0!
0'
0/
#48410000000
1!
1'
1/
#48420000000
0!
0'
0/
#48430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#48440000000
0!
0'
0/
#48450000000
1!
1'
1/
#48460000000
0!
0'
0/
#48470000000
1!
1'
1/
#48480000000
0!
0'
0/
#48490000000
1!
1'
1/
#48500000000
0!
0'
0/
#48510000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#48520000000
0!
0'
0/
#48530000000
1!
1'
1/
#48540000000
0!
0'
0/
#48550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#48560000000
0!
0'
0/
#48570000000
1!
1'
1/
#48580000000
0!
0'
0/
#48590000000
#48600000000
1!
1'
1/
#48610000000
0!
0'
0/
#48620000000
1!
1'
1/
#48630000000
0!
1"
0'
1(
0/
10
#48640000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#48650000000
0!
0'
0/
#48660000000
1!
1'
1/
#48670000000
0!
0'
0/
#48680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#48690000000
0!
0'
0/
#48700000000
1!
1'
1/
#48710000000
0!
1"
0'
1(
0/
10
#48720000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#48730000000
0!
1$
0'
1+
0/
#48740000000
1!
1'
1/
#48750000000
0!
0'
0/
#48760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#48770000000
0!
0'
0/
#48780000000
1!
1'
1/
#48790000000
0!
0'
0/
#48800000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#48810000000
0!
0'
0/
#48820000000
1!
1'
1/
#48830000000
0!
0'
0/
#48840000000
1!
1'
1/
#48850000000
0!
0'
0/
#48860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#48870000000
0!
0'
0/
#48880000000
1!
1'
1/
#48890000000
0!
0'
0/
#48900000000
1!
1'
1/
#48910000000
0!
0'
0/
#48920000000
1!
1'
1/
#48930000000
0!
0'
0/
#48940000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#48950000000
0!
0'
0/
#48960000000
1!
1'
1/
#48970000000
0!
0'
0/
#48980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#48990000000
0!
0'
0/
#49000000000
1!
1'
1/
#49010000000
0!
0'
0/
#49020000000
#49030000000
1!
1'
1/
#49040000000
0!
0'
0/
#49050000000
1!
1'
1/
#49060000000
0!
1"
0'
1(
0/
10
#49070000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#49080000000
0!
0'
0/
#49090000000
1!
1'
1/
#49100000000
0!
0'
0/
#49110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#49120000000
0!
0'
0/
#49130000000
1!
1'
1/
#49140000000
0!
1"
0'
1(
0/
10
#49150000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#49160000000
0!
1$
0'
1+
0/
#49170000000
1!
1'
1/
#49180000000
0!
0'
0/
#49190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#49200000000
0!
0'
0/
#49210000000
1!
1'
1/
#49220000000
0!
0'
0/
#49230000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#49240000000
0!
0'
0/
#49250000000
1!
1'
1/
#49260000000
0!
0'
0/
#49270000000
1!
1'
1/
#49280000000
0!
0'
0/
#49290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#49300000000
0!
0'
0/
#49310000000
1!
1'
1/
#49320000000
0!
0'
0/
#49330000000
1!
1'
1/
#49340000000
0!
0'
0/
#49350000000
1!
1'
1/
#49360000000
0!
0'
0/
#49370000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#49380000000
0!
0'
0/
#49390000000
1!
1'
1/
#49400000000
0!
0'
0/
#49410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#49420000000
0!
0'
0/
#49430000000
1!
1'
1/
#49440000000
0!
0'
0/
#49450000000
#49460000000
1!
1'
1/
#49470000000
0!
0'
0/
#49480000000
1!
1'
1/
#49490000000
0!
1"
0'
1(
0/
10
#49500000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#49510000000
0!
0'
0/
#49520000000
1!
1'
1/
#49530000000
0!
0'
0/
#49540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#49550000000
0!
0'
0/
#49560000000
1!
1'
1/
#49570000000
0!
1"
0'
1(
0/
10
#49580000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#49590000000
0!
1$
0'
1+
0/
#49600000000
1!
1'
1/
#49610000000
0!
0'
0/
#49620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#49630000000
0!
0'
0/
#49640000000
1!
1'
1/
#49650000000
0!
0'
0/
#49660000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#49670000000
0!
0'
0/
#49680000000
1!
1'
1/
#49690000000
0!
0'
0/
#49700000000
1!
1'
1/
#49710000000
0!
0'
0/
#49720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#49730000000
0!
0'
0/
#49740000000
1!
1'
1/
#49750000000
0!
0'
0/
#49760000000
1!
1'
1/
#49770000000
0!
0'
0/
#49780000000
1!
1'
1/
#49790000000
0!
0'
0/
#49800000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#49810000000
0!
0'
0/
#49820000000
1!
1'
1/
#49830000000
0!
0'
0/
#49840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#49850000000
0!
0'
0/
#49860000000
1!
1'
1/
#49870000000
0!
0'
0/
#49880000000
#49890000000
1!
1'
1/
#49900000000
0!
0'
0/
#49910000000
1!
1'
1/
#49920000000
0!
1"
0'
1(
0/
10
#49930000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#49940000000
0!
0'
0/
#49950000000
1!
1'
1/
#49960000000
0!
0'
0/
#49970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#49980000000
0!
0'
0/
#49990000000
1!
1'
1/
#50000000000
0!
1"
0'
1(
0/
10
#50010000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#50020000000
0!
1$
0'
1+
0/
#50030000000
1!
1'
1/
#50040000000
0!
0'
0/
#50050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#50060000000
0!
0'
0/
#50070000000
1!
1'
1/
#50080000000
0!
0'
0/
#50090000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#50100000000
0!
0'
0/
#50110000000
1!
1'
1/
#50120000000
0!
0'
0/
#50130000000
1!
1'
1/
#50140000000
0!
0'
0/
#50150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#50160000000
0!
0'
0/
#50170000000
1!
1'
1/
#50180000000
0!
0'
0/
#50190000000
1!
1'
1/
#50200000000
0!
0'
0/
#50210000000
1!
1'
1/
#50220000000
0!
0'
0/
#50230000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#50240000000
0!
0'
0/
#50250000000
1!
1'
1/
#50260000000
0!
0'
0/
#50270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#50280000000
0!
0'
0/
#50290000000
1!
1'
1/
#50300000000
0!
0'
0/
#50310000000
#50320000000
1!
1'
1/
#50330000000
0!
0'
0/
#50340000000
1!
1'
1/
#50350000000
0!
1"
0'
1(
0/
10
#50360000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#50370000000
0!
0'
0/
#50380000000
1!
1'
1/
#50390000000
0!
0'
0/
#50400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#50410000000
0!
0'
0/
#50420000000
1!
1'
1/
#50430000000
0!
1"
0'
1(
0/
10
#50440000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#50450000000
0!
1$
0'
1+
0/
#50460000000
1!
1'
1/
#50470000000
0!
0'
0/
#50480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#50490000000
0!
0'
0/
#50500000000
1!
1'
1/
#50510000000
0!
0'
0/
#50520000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#50530000000
0!
0'
0/
#50540000000
1!
1'
1/
#50550000000
0!
0'
0/
#50560000000
1!
1'
1/
#50570000000
0!
0'
0/
#50580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#50590000000
0!
0'
0/
#50600000000
1!
1'
1/
#50610000000
0!
0'
0/
#50620000000
1!
1'
1/
#50630000000
0!
0'
0/
#50640000000
1!
1'
1/
#50650000000
0!
0'
0/
#50660000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#50670000000
0!
0'
0/
#50680000000
1!
1'
1/
#50690000000
0!
0'
0/
#50700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#50710000000
0!
0'
0/
#50720000000
1!
1'
1/
#50730000000
0!
0'
0/
#50740000000
#50750000000
1!
1'
1/
#50760000000
0!
0'
0/
#50770000000
1!
1'
1/
#50780000000
0!
1"
0'
1(
0/
10
#50790000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#50800000000
0!
0'
0/
#50810000000
1!
1'
1/
#50820000000
0!
0'
0/
#50830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#50840000000
0!
0'
0/
#50850000000
1!
1'
1/
#50860000000
0!
1"
0'
1(
0/
10
#50870000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#50880000000
0!
1$
0'
1+
0/
#50890000000
1!
1'
1/
#50900000000
0!
0'
0/
#50910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#50920000000
0!
0'
0/
#50930000000
1!
1'
1/
#50940000000
0!
0'
0/
#50950000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#50960000000
0!
0'
0/
#50970000000
1!
1'
1/
#50980000000
0!
0'
0/
#50990000000
1!
1'
1/
#51000000000
0!
0'
0/
#51010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#51020000000
0!
0'
0/
#51030000000
1!
1'
1/
#51040000000
0!
0'
0/
#51050000000
1!
1'
1/
#51060000000
0!
0'
0/
#51070000000
1!
1'
1/
#51080000000
0!
0'
0/
#51090000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#51100000000
0!
0'
0/
#51110000000
1!
1'
1/
#51120000000
0!
0'
0/
#51130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#51140000000
0!
0'
0/
#51150000000
1!
1'
1/
#51160000000
0!
0'
0/
#51170000000
#51180000000
1!
1'
1/
#51190000000
0!
0'
0/
#51200000000
1!
1'
1/
#51210000000
0!
1"
0'
1(
0/
10
#51220000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#51230000000
0!
0'
0/
#51240000000
1!
1'
1/
#51250000000
0!
0'
0/
#51260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#51270000000
0!
0'
0/
#51280000000
1!
1'
1/
#51290000000
0!
1"
0'
1(
0/
10
#51300000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#51310000000
0!
1$
0'
1+
0/
#51320000000
1!
1'
1/
#51330000000
0!
0'
0/
#51340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#51350000000
0!
0'
0/
#51360000000
1!
1'
1/
#51370000000
0!
0'
0/
#51380000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#51390000000
0!
0'
0/
#51400000000
1!
1'
1/
#51410000000
0!
0'
0/
#51420000000
1!
1'
1/
#51430000000
0!
0'
0/
#51440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#51450000000
0!
0'
0/
#51460000000
1!
1'
1/
#51470000000
0!
0'
0/
#51480000000
1!
1'
1/
#51490000000
0!
0'
0/
#51500000000
1!
1'
1/
#51510000000
0!
0'
0/
#51520000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#51530000000
0!
0'
0/
#51540000000
1!
1'
1/
#51550000000
0!
0'
0/
#51560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#51570000000
0!
0'
0/
#51580000000
1!
1'
1/
#51590000000
0!
0'
0/
#51600000000
#51610000000
1!
1'
1/
#51620000000
0!
0'
0/
#51630000000
1!
1'
1/
#51640000000
0!
1"
0'
1(
0/
10
#51650000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#51660000000
0!
0'
0/
#51670000000
1!
1'
1/
#51680000000
0!
0'
0/
#51690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#51700000000
0!
0'
0/
#51710000000
1!
1'
1/
#51720000000
0!
1"
0'
1(
0/
10
#51730000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#51740000000
0!
1$
0'
1+
0/
#51750000000
1!
1'
1/
#51760000000
0!
0'
0/
#51770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#51780000000
0!
0'
0/
#51790000000
1!
1'
1/
#51800000000
0!
0'
0/
#51810000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#51820000000
0!
0'
0/
#51830000000
1!
1'
1/
#51840000000
0!
0'
0/
#51850000000
1!
1'
1/
#51860000000
0!
0'
0/
#51870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#51880000000
0!
0'
0/
#51890000000
1!
1'
1/
#51900000000
0!
0'
0/
#51910000000
1!
1'
1/
#51920000000
0!
0'
0/
#51930000000
1!
1'
1/
#51940000000
0!
0'
0/
#51950000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#51960000000
0!
0'
0/
#51970000000
1!
1'
1/
#51980000000
0!
0'
0/
#51990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#52000000000
0!
0'
0/
#52010000000
1!
1'
1/
#52020000000
0!
0'
0/
#52030000000
#52040000000
1!
1'
1/
#52050000000
0!
0'
0/
#52060000000
1!
1'
1/
#52070000000
0!
1"
0'
1(
0/
10
#52080000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#52090000000
0!
0'
0/
#52100000000
1!
1'
1/
#52110000000
0!
0'
0/
#52120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#52130000000
0!
0'
0/
#52140000000
1!
1'
1/
#52150000000
0!
1"
0'
1(
0/
10
#52160000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#52170000000
0!
1$
0'
1+
0/
#52180000000
1!
1'
1/
#52190000000
0!
0'
0/
#52200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#52210000000
0!
0'
0/
#52220000000
1!
1'
1/
#52230000000
0!
0'
0/
#52240000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#52250000000
0!
0'
0/
#52260000000
1!
1'
1/
#52270000000
0!
0'
0/
#52280000000
1!
1'
1/
#52290000000
0!
0'
0/
#52300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#52310000000
0!
0'
0/
#52320000000
1!
1'
1/
#52330000000
0!
0'
0/
#52340000000
1!
1'
1/
#52350000000
0!
0'
0/
#52360000000
1!
1'
1/
#52370000000
0!
0'
0/
#52380000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#52390000000
0!
0'
0/
#52400000000
1!
1'
1/
#52410000000
0!
0'
0/
#52420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#52430000000
0!
0'
0/
#52440000000
1!
1'
1/
#52450000000
0!
0'
0/
#52460000000
#52470000000
1!
1'
1/
#52480000000
0!
0'
0/
#52490000000
1!
1'
1/
#52500000000
0!
1"
0'
1(
0/
10
#52510000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#52520000000
0!
0'
0/
#52530000000
1!
1'
1/
#52540000000
0!
0'
0/
#52550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#52560000000
0!
0'
0/
#52570000000
1!
1'
1/
#52580000000
0!
1"
0'
1(
0/
10
#52590000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#52600000000
0!
1$
0'
1+
0/
#52610000000
1!
1'
1/
#52620000000
0!
0'
0/
#52630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#52640000000
0!
0'
0/
#52650000000
1!
1'
1/
#52660000000
0!
0'
0/
#52670000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#52680000000
0!
0'
0/
#52690000000
1!
1'
1/
#52700000000
0!
0'
0/
#52710000000
1!
1'
1/
#52720000000
0!
0'
0/
#52730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#52740000000
0!
0'
0/
#52750000000
1!
1'
1/
#52760000000
0!
0'
0/
#52770000000
1!
1'
1/
#52780000000
0!
0'
0/
#52790000000
1!
1'
1/
#52800000000
0!
0'
0/
#52810000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#52820000000
0!
0'
0/
#52830000000
1!
1'
1/
#52840000000
0!
0'
0/
#52850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#52860000000
0!
0'
0/
#52870000000
1!
1'
1/
#52880000000
0!
0'
0/
#52890000000
#52900000000
1!
1'
1/
#52910000000
0!
0'
0/
#52920000000
1!
1'
1/
#52930000000
0!
1"
0'
1(
0/
10
#52940000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#52950000000
0!
0'
0/
#52960000000
1!
1'
1/
#52970000000
0!
0'
0/
#52980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#52990000000
0!
0'
0/
#53000000000
1!
1'
1/
#53010000000
0!
1"
0'
1(
0/
10
#53020000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#53030000000
0!
1$
0'
1+
0/
#53040000000
1!
1'
1/
#53050000000
0!
0'
0/
#53060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#53070000000
0!
0'
0/
#53080000000
1!
1'
1/
#53090000000
0!
0'
0/
#53100000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#53110000000
0!
0'
0/
#53120000000
1!
1'
1/
#53130000000
0!
0'
0/
#53140000000
1!
1'
1/
#53150000000
0!
0'
0/
#53160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#53170000000
0!
0'
0/
#53180000000
1!
1'
1/
#53190000000
0!
0'
0/
#53200000000
1!
1'
1/
#53210000000
0!
0'
0/
#53220000000
1!
1'
1/
#53230000000
0!
0'
0/
#53240000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#53250000000
0!
0'
0/
#53260000000
1!
1'
1/
#53270000000
0!
0'
0/
#53280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#53290000000
0!
0'
0/
#53300000000
1!
1'
1/
#53310000000
0!
0'
0/
#53320000000
#53330000000
1!
1'
1/
#53340000000
0!
0'
0/
#53350000000
1!
1'
1/
#53360000000
0!
1"
0'
1(
0/
10
#53370000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#53380000000
0!
0'
0/
#53390000000
1!
1'
1/
#53400000000
0!
0'
0/
#53410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#53420000000
0!
0'
0/
#53430000000
1!
1'
1/
#53440000000
0!
1"
0'
1(
0/
10
#53450000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#53460000000
0!
1$
0'
1+
0/
#53470000000
1!
1'
1/
#53480000000
0!
0'
0/
#53490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#53500000000
0!
0'
0/
#53510000000
1!
1'
1/
#53520000000
0!
0'
0/
#53530000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#53540000000
0!
0'
0/
#53550000000
1!
1'
1/
#53560000000
0!
0'
0/
#53570000000
1!
1'
1/
#53580000000
0!
0'
0/
#53590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#53600000000
0!
0'
0/
#53610000000
1!
1'
1/
#53620000000
0!
0'
0/
#53630000000
1!
1'
1/
#53640000000
0!
0'
0/
#53650000000
1!
1'
1/
#53660000000
0!
0'
0/
#53670000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#53680000000
0!
0'
0/
#53690000000
1!
1'
1/
#53700000000
0!
0'
0/
#53710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#53720000000
0!
0'
0/
#53730000000
1!
1'
1/
#53740000000
0!
0'
0/
#53750000000
#53760000000
1!
1'
1/
#53770000000
0!
0'
0/
#53780000000
1!
1'
1/
#53790000000
0!
1"
0'
1(
0/
10
#53800000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#53810000000
0!
0'
0/
#53820000000
1!
1'
1/
#53830000000
0!
0'
0/
#53840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#53850000000
0!
0'
0/
#53860000000
1!
1'
1/
#53870000000
0!
1"
0'
1(
0/
10
#53880000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#53890000000
0!
1$
0'
1+
0/
#53900000000
1!
1'
1/
#53910000000
0!
0'
0/
#53920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#53930000000
0!
0'
0/
#53940000000
1!
1'
1/
#53950000000
0!
0'
0/
#53960000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#53970000000
0!
0'
0/
#53980000000
1!
1'
1/
#53990000000
0!
0'
0/
#54000000000
1!
1'
1/
#54010000000
0!
0'
0/
#54020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#54030000000
0!
0'
0/
#54040000000
1!
1'
1/
#54050000000
0!
0'
0/
#54060000000
1!
1'
1/
#54070000000
0!
0'
0/
#54080000000
1!
1'
1/
#54090000000
0!
0'
0/
#54100000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#54110000000
0!
0'
0/
#54120000000
1!
1'
1/
#54130000000
0!
0'
0/
#54140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#54150000000
0!
0'
0/
#54160000000
1!
1'
1/
#54170000000
0!
0'
0/
#54180000000
#54190000000
1!
1'
1/
#54200000000
0!
0'
0/
#54210000000
1!
1'
1/
#54220000000
0!
1"
0'
1(
0/
10
#54230000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#54240000000
0!
0'
0/
#54250000000
1!
1'
1/
#54260000000
0!
0'
0/
#54270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#54280000000
0!
0'
0/
#54290000000
1!
1'
1/
#54300000000
0!
1"
0'
1(
0/
10
#54310000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#54320000000
0!
1$
0'
1+
0/
#54330000000
1!
1'
1/
#54340000000
0!
0'
0/
#54350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#54360000000
0!
0'
0/
#54370000000
1!
1'
1/
#54380000000
0!
0'
0/
#54390000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#54400000000
0!
0'
0/
#54410000000
1!
1'
1/
#54420000000
0!
0'
0/
#54430000000
1!
1'
1/
#54440000000
0!
0'
0/
#54450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#54460000000
0!
0'
0/
#54470000000
1!
1'
1/
#54480000000
0!
0'
0/
#54490000000
1!
1'
1/
#54500000000
0!
0'
0/
#54510000000
1!
1'
1/
#54520000000
0!
0'
0/
#54530000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#54540000000
0!
0'
0/
#54550000000
1!
1'
1/
#54560000000
0!
0'
0/
#54570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#54580000000
0!
0'
0/
#54590000000
1!
1'
1/
#54600000000
0!
0'
0/
#54610000000
#54620000000
1!
1'
1/
#54630000000
0!
0'
0/
#54640000000
1!
1'
1/
#54650000000
0!
1"
0'
1(
0/
10
#54660000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#54670000000
0!
0'
0/
#54680000000
1!
1'
1/
#54690000000
0!
0'
0/
#54700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#54710000000
0!
0'
0/
#54720000000
1!
1'
1/
#54730000000
0!
1"
0'
1(
0/
10
#54740000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#54750000000
0!
1$
0'
1+
0/
#54760000000
1!
1'
1/
#54770000000
0!
0'
0/
#54780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#54790000000
0!
0'
0/
#54800000000
1!
1'
1/
#54810000000
0!
0'
0/
#54820000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#54830000000
0!
0'
0/
#54840000000
1!
1'
1/
#54850000000
0!
0'
0/
#54860000000
1!
1'
1/
#54870000000
0!
0'
0/
#54880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#54890000000
0!
0'
0/
#54900000000
1!
1'
1/
#54910000000
0!
0'
0/
#54920000000
1!
1'
1/
#54930000000
0!
0'
0/
#54940000000
1!
1'
1/
#54950000000
0!
0'
0/
#54960000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#54970000000
0!
0'
0/
#54980000000
1!
1'
1/
#54990000000
0!
0'
0/
#55000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#55010000000
0!
0'
0/
#55020000000
1!
1'
1/
#55030000000
0!
0'
0/
#55040000000
#55050000000
1!
1'
1/
#55060000000
0!
0'
0/
#55070000000
1!
1'
1/
#55080000000
0!
1"
0'
1(
0/
10
#55090000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#55100000000
0!
0'
0/
#55110000000
1!
1'
1/
#55120000000
0!
0'
0/
#55130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#55140000000
0!
0'
0/
#55150000000
1!
1'
1/
#55160000000
0!
1"
0'
1(
0/
10
#55170000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#55180000000
0!
1$
0'
1+
0/
#55190000000
1!
1'
1/
#55200000000
0!
0'
0/
#55210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#55220000000
0!
0'
0/
#55230000000
1!
1'
1/
#55240000000
0!
0'
0/
#55250000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#55260000000
0!
0'
0/
#55270000000
1!
1'
1/
#55280000000
0!
0'
0/
#55290000000
1!
1'
1/
#55300000000
0!
0'
0/
#55310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#55320000000
0!
0'
0/
#55330000000
1!
1'
1/
#55340000000
0!
0'
0/
#55350000000
1!
1'
1/
#55360000000
0!
0'
0/
#55370000000
1!
1'
1/
#55380000000
0!
0'
0/
#55390000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#55400000000
0!
0'
0/
#55410000000
1!
1'
1/
#55420000000
0!
0'
0/
#55430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#55440000000
0!
0'
0/
#55450000000
1!
1'
1/
#55460000000
0!
0'
0/
#55470000000
#55480000000
1!
1'
1/
#55490000000
0!
0'
0/
#55500000000
1!
1'
1/
#55510000000
0!
1"
0'
1(
0/
10
#55520000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#55530000000
0!
0'
0/
#55540000000
1!
1'
1/
#55550000000
0!
0'
0/
#55560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#55570000000
0!
0'
0/
#55580000000
1!
1'
1/
#55590000000
0!
1"
0'
1(
0/
10
#55600000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#55610000000
0!
1$
0'
1+
0/
#55620000000
1!
1'
1/
#55630000000
0!
0'
0/
#55640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#55650000000
0!
0'
0/
#55660000000
1!
1'
1/
#55670000000
0!
0'
0/
#55680000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#55690000000
0!
0'
0/
#55700000000
1!
1'
1/
#55710000000
0!
0'
0/
#55720000000
1!
1'
1/
#55730000000
0!
0'
0/
#55740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#55750000000
0!
0'
0/
#55760000000
1!
1'
1/
#55770000000
0!
0'
0/
#55780000000
1!
1'
1/
#55790000000
0!
0'
0/
#55800000000
1!
1'
1/
#55810000000
0!
0'
0/
#55820000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#55830000000
0!
0'
0/
#55840000000
1!
1'
1/
#55850000000
0!
0'
0/
#55860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#55870000000
0!
0'
0/
#55880000000
1!
1'
1/
#55890000000
0!
0'
0/
#55900000000
#55910000000
1!
1'
1/
#55920000000
0!
0'
0/
#55930000000
1!
1'
1/
#55940000000
0!
1"
0'
1(
0/
10
#55950000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#55960000000
0!
0'
0/
#55970000000
1!
1'
1/
#55980000000
0!
0'
0/
#55990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#56000000000
0!
0'
0/
#56010000000
1!
1'
1/
#56020000000
0!
1"
0'
1(
0/
10
#56030000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#56040000000
0!
1$
0'
1+
0/
#56050000000
1!
1'
1/
#56060000000
0!
0'
0/
#56070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#56080000000
0!
0'
0/
#56090000000
1!
1'
1/
#56100000000
0!
0'
0/
#56110000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#56120000000
0!
0'
0/
#56130000000
1!
1'
1/
#56140000000
0!
0'
0/
#56150000000
1!
1'
1/
#56160000000
0!
0'
0/
#56170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#56180000000
0!
0'
0/
#56190000000
1!
1'
1/
#56200000000
0!
0'
0/
#56210000000
1!
1'
1/
#56220000000
0!
0'
0/
#56230000000
1!
1'
1/
#56240000000
0!
0'
0/
#56250000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#56260000000
0!
0'
0/
#56270000000
1!
1'
1/
#56280000000
0!
0'
0/
#56290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#56300000000
0!
0'
0/
#56310000000
1!
1'
1/
#56320000000
0!
0'
0/
#56330000000
#56340000000
1!
1'
1/
#56350000000
0!
0'
0/
#56360000000
1!
1'
1/
#56370000000
0!
1"
0'
1(
0/
10
#56380000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#56390000000
0!
0'
0/
#56400000000
1!
1'
1/
#56410000000
0!
0'
0/
#56420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#56430000000
0!
0'
0/
#56440000000
1!
1'
1/
#56450000000
0!
1"
0'
1(
0/
10
#56460000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#56470000000
0!
1$
0'
1+
0/
#56480000000
1!
1'
1/
#56490000000
0!
0'
0/
#56500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#56510000000
0!
0'
0/
#56520000000
1!
1'
1/
#56530000000
0!
0'
0/
#56540000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#56550000000
0!
0'
0/
#56560000000
1!
1'
1/
#56570000000
0!
0'
0/
#56580000000
1!
1'
1/
#56590000000
0!
0'
0/
#56600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#56610000000
0!
0'
0/
#56620000000
1!
1'
1/
#56630000000
0!
0'
0/
#56640000000
1!
1'
1/
#56650000000
0!
0'
0/
#56660000000
1!
1'
1/
#56670000000
0!
0'
0/
#56680000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#56690000000
0!
0'
0/
#56700000000
1!
1'
1/
#56710000000
0!
0'
0/
#56720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#56730000000
0!
0'
0/
#56740000000
1!
1'
1/
#56750000000
0!
0'
0/
#56760000000
#56770000000
1!
1'
1/
#56780000000
0!
0'
0/
#56790000000
1!
1'
1/
#56800000000
0!
1"
0'
1(
0/
10
#56810000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#56820000000
0!
0'
0/
#56830000000
1!
1'
1/
#56840000000
0!
0'
0/
#56850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#56860000000
0!
0'
0/
#56870000000
1!
1'
1/
#56880000000
0!
1"
0'
1(
0/
10
#56890000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#56900000000
0!
1$
0'
1+
0/
#56910000000
1!
1'
1/
#56920000000
0!
0'
0/
#56930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#56940000000
0!
0'
0/
#56950000000
1!
1'
1/
#56960000000
0!
0'
0/
#56970000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#56980000000
0!
0'
0/
#56990000000
1!
1'
1/
#57000000000
0!
0'
0/
#57010000000
1!
1'
1/
#57020000000
0!
0'
0/
#57030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#57040000000
0!
0'
0/
#57050000000
1!
1'
1/
#57060000000
0!
0'
0/
#57070000000
1!
1'
1/
#57080000000
0!
0'
0/
#57090000000
1!
1'
1/
#57100000000
0!
0'
0/
#57110000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#57120000000
0!
0'
0/
#57130000000
1!
1'
1/
#57140000000
0!
0'
0/
#57150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#57160000000
0!
0'
0/
#57170000000
1!
1'
1/
#57180000000
0!
0'
0/
#57190000000
#57200000000
1!
1'
1/
#57210000000
0!
0'
0/
#57220000000
1!
1'
1/
#57230000000
0!
1"
0'
1(
0/
10
#57240000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#57250000000
0!
0'
0/
#57260000000
1!
1'
1/
#57270000000
0!
0'
0/
#57280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#57290000000
0!
0'
0/
#57300000000
1!
1'
1/
#57310000000
0!
1"
0'
1(
0/
10
#57320000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#57330000000
0!
1$
0'
1+
0/
#57340000000
1!
1'
1/
#57350000000
0!
0'
0/
#57360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#57370000000
0!
0'
0/
#57380000000
1!
1'
1/
#57390000000
0!
0'
0/
#57400000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#57410000000
0!
0'
0/
#57420000000
1!
1'
1/
#57430000000
0!
0'
0/
#57440000000
1!
1'
1/
#57450000000
0!
0'
0/
#57460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#57470000000
0!
0'
0/
#57480000000
1!
1'
1/
#57490000000
0!
0'
0/
#57500000000
1!
1'
1/
#57510000000
0!
0'
0/
#57520000000
1!
1'
1/
#57530000000
0!
0'
0/
#57540000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#57550000000
0!
0'
0/
#57560000000
1!
1'
1/
#57570000000
0!
0'
0/
#57580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#57590000000
0!
0'
0/
#57600000000
1!
1'
1/
#57610000000
0!
0'
0/
#57620000000
#57630000000
1!
1'
1/
#57640000000
0!
0'
0/
#57650000000
1!
1'
1/
#57660000000
0!
1"
0'
1(
0/
10
#57670000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#57680000000
0!
0'
0/
#57690000000
1!
1'
1/
#57700000000
0!
0'
0/
#57710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#57720000000
0!
0'
0/
#57730000000
1!
1'
1/
#57740000000
0!
1"
0'
1(
0/
10
#57750000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#57760000000
0!
1$
0'
1+
0/
#57770000000
1!
1'
1/
#57780000000
0!
0'
0/
#57790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#57800000000
0!
0'
0/
#57810000000
1!
1'
1/
#57820000000
0!
0'
0/
#57830000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#57840000000
0!
0'
0/
#57850000000
1!
1'
1/
#57860000000
0!
0'
0/
#57870000000
1!
1'
1/
#57880000000
0!
0'
0/
#57890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#57900000000
0!
0'
0/
#57910000000
1!
1'
1/
#57920000000
0!
0'
0/
#57930000000
1!
1'
1/
#57940000000
0!
0'
0/
#57950000000
1!
1'
1/
#57960000000
0!
0'
0/
#57970000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#57980000000
0!
0'
0/
#57990000000
1!
1'
1/
#58000000000
0!
0'
0/
#58010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#58020000000
0!
0'
0/
#58030000000
1!
1'
1/
#58040000000
0!
0'
0/
#58050000000
#58060000000
1!
1'
1/
#58070000000
0!
0'
0/
#58080000000
1!
1'
1/
#58090000000
0!
1"
0'
1(
0/
10
#58100000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#58110000000
0!
0'
0/
#58120000000
1!
1'
1/
#58130000000
0!
0'
0/
#58140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#58150000000
0!
0'
0/
#58160000000
1!
1'
1/
#58170000000
0!
1"
0'
1(
0/
10
#58180000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#58190000000
0!
1$
0'
1+
0/
#58200000000
1!
1'
1/
#58210000000
0!
0'
0/
#58220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#58230000000
0!
0'
0/
#58240000000
1!
1'
1/
#58250000000
0!
0'
0/
#58260000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#58270000000
0!
0'
0/
#58280000000
1!
1'
1/
#58290000000
0!
0'
0/
#58300000000
1!
1'
1/
#58310000000
0!
0'
0/
#58320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#58330000000
0!
0'
0/
#58340000000
1!
1'
1/
#58350000000
0!
0'
0/
#58360000000
1!
1'
1/
#58370000000
0!
0'
0/
#58380000000
1!
1'
1/
#58390000000
0!
0'
0/
#58400000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#58410000000
0!
0'
0/
#58420000000
1!
1'
1/
#58430000000
0!
0'
0/
#58440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#58450000000
0!
0'
0/
#58460000000
1!
1'
1/
#58470000000
0!
0'
0/
#58480000000
#58490000000
1!
1'
1/
#58500000000
0!
0'
0/
#58510000000
1!
1'
1/
#58520000000
0!
1"
0'
1(
0/
10
#58530000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#58540000000
0!
0'
0/
#58550000000
1!
1'
1/
#58560000000
0!
0'
0/
#58570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#58580000000
0!
0'
0/
#58590000000
1!
1'
1/
#58600000000
0!
1"
0'
1(
0/
10
#58610000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#58620000000
0!
1$
0'
1+
0/
#58630000000
1!
1'
1/
#58640000000
0!
0'
0/
#58650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#58660000000
0!
0'
0/
#58670000000
1!
1'
1/
#58680000000
0!
0'
0/
#58690000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#58700000000
0!
0'
0/
#58710000000
1!
1'
1/
#58720000000
0!
0'
0/
#58730000000
1!
1'
1/
#58740000000
0!
0'
0/
#58750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#58760000000
0!
0'
0/
#58770000000
1!
1'
1/
#58780000000
0!
0'
0/
#58790000000
1!
1'
1/
#58800000000
0!
0'
0/
#58810000000
1!
1'
1/
#58820000000
0!
0'
0/
#58830000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#58840000000
0!
0'
0/
#58850000000
1!
1'
1/
#58860000000
0!
0'
0/
#58870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#58880000000
0!
0'
0/
#58890000000
1!
1'
1/
#58900000000
0!
0'
0/
#58910000000
#58920000000
1!
1'
1/
#58930000000
0!
0'
0/
#58940000000
1!
1'
1/
#58950000000
0!
1"
0'
1(
0/
10
#58960000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#58970000000
0!
0'
0/
#58980000000
1!
1'
1/
#58990000000
0!
0'
0/
#59000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#59010000000
0!
0'
0/
#59020000000
1!
1'
1/
#59030000000
0!
1"
0'
1(
0/
10
#59040000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#59050000000
0!
1$
0'
1+
0/
#59060000000
1!
1'
1/
#59070000000
0!
0'
0/
#59080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#59090000000
0!
0'
0/
#59100000000
1!
1'
1/
#59110000000
0!
0'
0/
#59120000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#59130000000
0!
0'
0/
#59140000000
1!
1'
1/
#59150000000
0!
0'
0/
#59160000000
1!
1'
1/
#59170000000
0!
0'
0/
#59180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#59190000000
0!
0'
0/
#59200000000
1!
1'
1/
#59210000000
0!
0'
0/
#59220000000
1!
1'
1/
#59230000000
0!
0'
0/
#59240000000
1!
1'
1/
#59250000000
0!
0'
0/
#59260000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#59270000000
0!
0'
0/
#59280000000
1!
1'
1/
#59290000000
0!
0'
0/
#59300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#59310000000
0!
0'
0/
#59320000000
1!
1'
1/
#59330000000
0!
0'
0/
#59340000000
#59350000000
1!
1'
1/
#59360000000
0!
0'
0/
#59370000000
1!
1'
1/
#59380000000
0!
1"
0'
1(
0/
10
#59390000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#59400000000
0!
0'
0/
#59410000000
1!
1'
1/
#59420000000
0!
0'
0/
#59430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#59440000000
0!
0'
0/
#59450000000
1!
1'
1/
#59460000000
0!
1"
0'
1(
0/
10
#59470000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#59480000000
0!
1$
0'
1+
0/
#59490000000
1!
1'
1/
#59500000000
0!
0'
0/
#59510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#59520000000
0!
0'
0/
#59530000000
1!
1'
1/
#59540000000
0!
0'
0/
#59550000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#59560000000
0!
0'
0/
#59570000000
1!
1'
1/
#59580000000
0!
0'
0/
#59590000000
1!
1'
1/
#59600000000
0!
0'
0/
#59610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#59620000000
0!
0'
0/
#59630000000
1!
1'
1/
#59640000000
0!
0'
0/
#59650000000
1!
1'
1/
#59660000000
0!
0'
0/
#59670000000
1!
1'
1/
#59680000000
0!
0'
0/
#59690000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#59700000000
0!
0'
0/
#59710000000
1!
1'
1/
#59720000000
0!
0'
0/
#59730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#59740000000
0!
0'
0/
#59750000000
1!
1'
1/
#59760000000
0!
0'
0/
#59770000000
#59780000000
1!
1'
1/
#59790000000
0!
0'
0/
#59800000000
1!
1'
1/
#59810000000
0!
1"
0'
1(
0/
10
#59820000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#59830000000
0!
0'
0/
#59840000000
1!
1'
1/
#59850000000
0!
0'
0/
#59860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#59870000000
0!
0'
0/
#59880000000
1!
1'
1/
#59890000000
0!
1"
0'
1(
0/
10
#59900000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#59910000000
0!
1$
0'
1+
0/
#59920000000
1!
1'
1/
#59930000000
0!
0'
0/
#59940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#59950000000
0!
0'
0/
#59960000000
1!
1'
1/
#59970000000
0!
0'
0/
#59980000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#59990000000
0!
0'
0/
#60000000000
1!
1'
1/
#60010000000
0!
0'
0/
#60020000000
1!
1'
1/
#60030000000
0!
0'
0/
#60040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#60050000000
0!
0'
0/
#60060000000
1!
1'
1/
#60070000000
0!
0'
0/
#60080000000
1!
1'
1/
#60090000000
0!
0'
0/
#60100000000
1!
1'
1/
#60110000000
0!
0'
0/
#60120000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#60130000000
0!
0'
0/
#60140000000
1!
1'
1/
#60150000000
0!
0'
0/
#60160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#60170000000
0!
0'
0/
#60180000000
1!
1'
1/
#60190000000
0!
0'
0/
#60200000000
#60210000000
1!
1'
1/
#60220000000
0!
0'
0/
#60230000000
1!
1'
1/
#60240000000
0!
1"
0'
1(
0/
10
#60250000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#60260000000
0!
0'
0/
#60270000000
1!
1'
1/
#60280000000
0!
0'
0/
#60290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#60300000000
0!
0'
0/
#60310000000
1!
1'
1/
#60320000000
0!
1"
0'
1(
0/
10
#60330000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#60340000000
0!
1$
0'
1+
0/
#60350000000
1!
1'
1/
#60360000000
0!
0'
0/
#60370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#60380000000
0!
0'
0/
#60390000000
1!
1'
1/
#60400000000
0!
0'
0/
#60410000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#60420000000
0!
0'
0/
#60430000000
1!
1'
1/
#60440000000
0!
0'
0/
#60450000000
1!
1'
1/
#60460000000
0!
0'
0/
#60470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#60480000000
0!
0'
0/
#60490000000
1!
1'
1/
#60500000000
0!
0'
0/
#60510000000
1!
1'
1/
#60520000000
0!
0'
0/
#60530000000
1!
1'
1/
#60540000000
0!
0'
0/
#60550000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#60560000000
0!
0'
0/
#60570000000
1!
1'
1/
#60580000000
0!
0'
0/
#60590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#60600000000
0!
0'
0/
#60610000000
1!
1'
1/
#60620000000
0!
0'
0/
#60630000000
#60640000000
1!
1'
1/
#60650000000
0!
0'
0/
#60660000000
1!
1'
1/
#60670000000
0!
1"
0'
1(
0/
10
#60680000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#60690000000
0!
0'
0/
#60700000000
1!
1'
1/
#60710000000
0!
0'
0/
#60720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#60730000000
0!
0'
0/
#60740000000
1!
1'
1/
#60750000000
0!
1"
0'
1(
0/
10
#60760000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#60770000000
0!
1$
0'
1+
0/
#60780000000
1!
1'
1/
#60790000000
0!
0'
0/
#60800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#60810000000
0!
0'
0/
#60820000000
1!
1'
1/
#60830000000
0!
0'
0/
#60840000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#60850000000
0!
0'
0/
#60860000000
1!
1'
1/
#60870000000
0!
0'
0/
#60880000000
1!
1'
1/
#60890000000
0!
0'
0/
#60900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#60910000000
0!
0'
0/
#60920000000
1!
1'
1/
#60930000000
0!
0'
0/
#60940000000
1!
1'
1/
#60950000000
0!
0'
0/
#60960000000
1!
1'
1/
#60970000000
0!
0'
0/
#60980000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#60990000000
0!
0'
0/
#61000000000
1!
1'
1/
#61010000000
0!
0'
0/
#61020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#61030000000
0!
0'
0/
#61040000000
1!
1'
1/
#61050000000
0!
0'
0/
#61060000000
#61070000000
1!
1'
1/
#61080000000
0!
0'
0/
#61090000000
1!
1'
1/
#61100000000
0!
1"
0'
1(
0/
10
#61110000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#61120000000
0!
0'
0/
#61130000000
1!
1'
1/
#61140000000
0!
0'
0/
#61150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#61160000000
0!
0'
0/
#61170000000
1!
1'
1/
#61180000000
0!
1"
0'
1(
0/
10
#61190000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#61200000000
0!
1$
0'
1+
0/
#61210000000
1!
1'
1/
#61220000000
0!
0'
0/
#61230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#61240000000
0!
0'
0/
#61250000000
1!
1'
1/
#61260000000
0!
0'
0/
#61270000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#61280000000
0!
0'
0/
#61290000000
1!
1'
1/
#61300000000
0!
0'
0/
#61310000000
1!
1'
1/
#61320000000
0!
0'
0/
#61330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#61340000000
0!
0'
0/
#61350000000
1!
1'
1/
#61360000000
0!
0'
0/
#61370000000
1!
1'
1/
#61380000000
0!
0'
0/
#61390000000
1!
1'
1/
#61400000000
0!
0'
0/
#61410000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#61420000000
0!
0'
0/
#61430000000
1!
1'
1/
#61440000000
0!
0'
0/
#61450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#61460000000
0!
0'
0/
#61470000000
1!
1'
1/
#61480000000
0!
0'
0/
#61490000000
#61500000000
1!
1'
1/
#61510000000
0!
0'
0/
#61520000000
1!
1'
1/
#61530000000
0!
1"
0'
1(
0/
10
#61540000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#61550000000
0!
0'
0/
#61560000000
1!
1'
1/
#61570000000
0!
0'
0/
#61580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#61590000000
0!
0'
0/
#61600000000
1!
1'
1/
#61610000000
0!
1"
0'
1(
0/
10
#61620000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#61630000000
0!
1$
0'
1+
0/
#61640000000
1!
1'
1/
#61650000000
0!
0'
0/
#61660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#61670000000
0!
0'
0/
#61680000000
1!
1'
1/
#61690000000
0!
0'
0/
#61700000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#61710000000
0!
0'
0/
#61720000000
1!
1'
1/
#61730000000
0!
0'
0/
#61740000000
1!
1'
1/
#61750000000
0!
0'
0/
#61760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#61770000000
0!
0'
0/
#61780000000
1!
1'
1/
#61790000000
0!
0'
0/
#61800000000
1!
1'
1/
#61810000000
0!
0'
0/
#61820000000
1!
1'
1/
#61830000000
0!
0'
0/
#61840000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#61850000000
0!
0'
0/
#61860000000
1!
1'
1/
#61870000000
0!
0'
0/
#61880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#61890000000
0!
0'
0/
#61900000000
1!
1'
1/
#61910000000
0!
0'
0/
#61920000000
#61930000000
1!
1'
1/
#61940000000
0!
0'
0/
#61950000000
1!
1'
1/
#61960000000
0!
1"
0'
1(
0/
10
#61970000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#61980000000
0!
0'
0/
#61990000000
1!
1'
1/
#62000000000
0!
0'
0/
#62010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#62020000000
0!
0'
0/
#62030000000
1!
1'
1/
#62040000000
0!
1"
0'
1(
0/
10
#62050000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#62060000000
0!
1$
0'
1+
0/
#62070000000
1!
1'
1/
#62080000000
0!
0'
0/
#62090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#62100000000
0!
0'
0/
#62110000000
1!
1'
1/
#62120000000
0!
0'
0/
#62130000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#62140000000
0!
0'
0/
#62150000000
1!
1'
1/
#62160000000
0!
0'
0/
#62170000000
1!
1'
1/
#62180000000
0!
0'
0/
#62190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#62200000000
0!
0'
0/
#62210000000
1!
1'
1/
#62220000000
0!
0'
0/
#62230000000
1!
1'
1/
#62240000000
0!
0'
0/
#62250000000
1!
1'
1/
#62260000000
0!
0'
0/
#62270000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#62280000000
0!
0'
0/
#62290000000
1!
1'
1/
#62300000000
0!
0'
0/
#62310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#62320000000
0!
0'
0/
#62330000000
1!
1'
1/
#62340000000
0!
0'
0/
#62350000000
#62360000000
1!
1'
1/
#62370000000
0!
0'
0/
#62380000000
1!
1'
1/
#62390000000
0!
1"
0'
1(
0/
10
#62400000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#62410000000
0!
0'
0/
#62420000000
1!
1'
1/
#62430000000
0!
0'
0/
#62440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#62450000000
0!
0'
0/
#62460000000
1!
1'
1/
#62470000000
0!
1"
0'
1(
0/
10
#62480000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#62490000000
0!
1$
0'
1+
0/
#62500000000
1!
1'
1/
#62510000000
0!
0'
0/
#62520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#62530000000
0!
0'
0/
#62540000000
1!
1'
1/
#62550000000
0!
0'
0/
#62560000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#62570000000
0!
0'
0/
#62580000000
1!
1'
1/
#62590000000
0!
0'
0/
#62600000000
1!
1'
1/
#62610000000
0!
0'
0/
#62620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#62630000000
0!
0'
0/
#62640000000
1!
1'
1/
#62650000000
0!
0'
0/
#62660000000
1!
1'
1/
#62670000000
0!
0'
0/
#62680000000
1!
1'
1/
#62690000000
0!
0'
0/
#62700000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#62710000000
0!
0'
0/
#62720000000
1!
1'
1/
#62730000000
0!
0'
0/
#62740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#62750000000
0!
0'
0/
#62760000000
1!
1'
1/
#62770000000
0!
0'
0/
#62780000000
#62790000000
1!
1'
1/
#62800000000
0!
0'
0/
#62810000000
1!
1'
1/
#62820000000
0!
1"
0'
1(
0/
10
#62830000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#62840000000
0!
0'
0/
#62850000000
1!
1'
1/
#62860000000
0!
0'
0/
#62870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#62880000000
0!
0'
0/
#62890000000
1!
1'
1/
#62900000000
0!
1"
0'
1(
0/
10
#62910000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#62920000000
0!
1$
0'
1+
0/
#62930000000
1!
1'
1/
#62940000000
0!
0'
0/
#62950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#62960000000
0!
0'
0/
#62970000000
1!
1'
1/
#62980000000
0!
0'
0/
#62990000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#63000000000
0!
0'
0/
#63010000000
1!
1'
1/
#63020000000
0!
0'
0/
#63030000000
1!
1'
1/
#63040000000
0!
0'
0/
#63050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#63060000000
0!
0'
0/
#63070000000
1!
1'
1/
#63080000000
0!
0'
0/
#63090000000
1!
1'
1/
#63100000000
0!
0'
0/
#63110000000
1!
1'
1/
#63120000000
0!
0'
0/
#63130000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#63140000000
0!
0'
0/
#63150000000
1!
1'
1/
#63160000000
0!
0'
0/
#63170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#63180000000
0!
0'
0/
#63190000000
1!
1'
1/
#63200000000
0!
0'
0/
#63210000000
#63220000000
1!
1'
1/
#63230000000
0!
0'
0/
#63240000000
1!
1'
1/
#63250000000
0!
1"
0'
1(
0/
10
#63260000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#63270000000
0!
0'
0/
#63280000000
1!
1'
1/
#63290000000
0!
0'
0/
#63300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#63310000000
0!
0'
0/
#63320000000
1!
1'
1/
#63330000000
0!
1"
0'
1(
0/
10
#63340000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#63350000000
0!
1$
0'
1+
0/
#63360000000
1!
1'
1/
#63370000000
0!
0'
0/
#63380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#63390000000
0!
0'
0/
#63400000000
1!
1'
1/
#63410000000
0!
0'
0/
#63420000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#63430000000
0!
0'
0/
#63440000000
1!
1'
1/
#63450000000
0!
0'
0/
#63460000000
1!
1'
1/
#63470000000
0!
0'
0/
#63480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#63490000000
0!
0'
0/
#63500000000
1!
1'
1/
#63510000000
0!
0'
0/
#63520000000
1!
1'
1/
#63530000000
0!
0'
0/
#63540000000
1!
1'
1/
#63550000000
0!
0'
0/
#63560000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#63570000000
0!
0'
0/
#63580000000
1!
1'
1/
#63590000000
0!
0'
0/
#63600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#63610000000
0!
0'
0/
#63620000000
1!
1'
1/
#63630000000
0!
0'
0/
#63640000000
#63650000000
1!
1'
1/
#63660000000
0!
0'
0/
#63670000000
1!
1'
1/
#63680000000
0!
1"
0'
1(
0/
10
#63690000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#63700000000
0!
0'
0/
#63710000000
1!
1'
1/
#63720000000
0!
0'
0/
#63730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#63740000000
0!
0'
0/
#63750000000
1!
1'
1/
#63760000000
0!
1"
0'
1(
0/
10
#63770000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#63780000000
0!
1$
0'
1+
0/
#63790000000
1!
1'
1/
#63800000000
0!
0'
0/
#63810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#63820000000
0!
0'
0/
#63830000000
1!
1'
1/
#63840000000
0!
0'
0/
#63850000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#63860000000
0!
0'
0/
#63870000000
1!
1'
1/
#63880000000
0!
0'
0/
#63890000000
1!
1'
1/
#63900000000
0!
0'
0/
#63910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#63920000000
0!
0'
0/
#63930000000
1!
1'
1/
#63940000000
0!
0'
0/
#63950000000
1!
1'
1/
#63960000000
0!
0'
0/
#63970000000
1!
1'
1/
#63980000000
0!
0'
0/
#63990000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#64000000000
0!
0'
0/
#64010000000
1!
1'
1/
#64020000000
0!
0'
0/
#64030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#64040000000
0!
0'
0/
#64050000000
1!
1'
1/
#64060000000
0!
0'
0/
#64070000000
#64080000000
1!
1'
1/
#64090000000
0!
0'
0/
#64100000000
1!
1'
1/
#64110000000
0!
1"
0'
1(
0/
10
#64120000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#64130000000
0!
0'
0/
#64140000000
1!
1'
1/
#64150000000
0!
0'
0/
#64160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#64170000000
0!
0'
0/
#64180000000
1!
1'
1/
#64190000000
0!
1"
0'
1(
0/
10
#64200000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#64210000000
0!
1$
0'
1+
0/
#64220000000
1!
1'
1/
#64230000000
0!
0'
0/
#64240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#64250000000
0!
0'
0/
#64260000000
1!
1'
1/
#64270000000
0!
0'
0/
#64280000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#64290000000
0!
0'
0/
#64300000000
1!
1'
1/
#64310000000
0!
0'
0/
#64320000000
1!
1'
1/
#64330000000
0!
0'
0/
#64340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#64350000000
0!
0'
0/
#64360000000
1!
1'
1/
#64370000000
0!
0'
0/
#64380000000
1!
1'
1/
#64390000000
0!
0'
0/
#64400000000
1!
1'
1/
#64410000000
0!
0'
0/
#64420000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#64430000000
0!
0'
0/
#64440000000
1!
1'
1/
#64450000000
0!
0'
0/
#64460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#64470000000
0!
0'
0/
#64480000000
1!
1'
1/
#64490000000
0!
0'
0/
#64500000000
#64510000000
1!
1'
1/
#64520000000
0!
0'
0/
#64530000000
1!
1'
1/
#64540000000
0!
1"
0'
1(
0/
10
#64550000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#64560000000
0!
0'
0/
#64570000000
1!
1'
1/
#64580000000
0!
0'
0/
#64590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#64600000000
0!
0'
0/
#64610000000
1!
1'
1/
#64620000000
0!
1"
0'
1(
0/
10
#64630000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#64640000000
0!
1$
0'
1+
0/
#64650000000
1!
1'
1/
#64660000000
0!
0'
0/
#64670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#64680000000
0!
0'
0/
#64690000000
1!
1'
1/
#64700000000
0!
0'
0/
#64710000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#64720000000
0!
0'
0/
#64730000000
1!
1'
1/
#64740000000
0!
0'
0/
#64750000000
1!
1'
1/
#64760000000
0!
0'
0/
#64770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#64780000000
0!
0'
0/
#64790000000
1!
1'
1/
#64800000000
0!
0'
0/
#64810000000
1!
1'
1/
#64820000000
0!
0'
0/
#64830000000
1!
1'
1/
#64840000000
0!
0'
0/
#64850000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#64860000000
0!
0'
0/
#64870000000
1!
1'
1/
#64880000000
0!
0'
0/
#64890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#64900000000
0!
0'
0/
#64910000000
1!
1'
1/
#64920000000
0!
0'
0/
#64930000000
#64940000000
1!
1'
1/
#64950000000
0!
0'
0/
#64960000000
1!
1'
1/
#64970000000
0!
1"
0'
1(
0/
10
#64980000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#64990000000
0!
0'
0/
#65000000000
1!
1'
1/
#65010000000
0!
0'
0/
#65020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#65030000000
0!
0'
0/
#65040000000
1!
1'
1/
#65050000000
0!
1"
0'
1(
0/
10
#65060000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#65070000000
0!
1$
0'
1+
0/
#65080000000
1!
1'
1/
#65090000000
0!
0'
0/
#65100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#65110000000
0!
0'
0/
#65120000000
1!
1'
1/
#65130000000
0!
0'
0/
#65140000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#65150000000
0!
0'
0/
#65160000000
1!
1'
1/
#65170000000
0!
0'
0/
#65180000000
1!
1'
1/
#65190000000
0!
0'
0/
#65200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#65210000000
0!
0'
0/
#65220000000
1!
1'
1/
#65230000000
0!
0'
0/
#65240000000
1!
1'
1/
#65250000000
0!
0'
0/
#65260000000
1!
1'
1/
#65270000000
0!
0'
0/
#65280000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#65290000000
0!
0'
0/
#65300000000
1!
1'
1/
#65310000000
0!
0'
0/
#65320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#65330000000
0!
0'
0/
#65340000000
1!
1'
1/
#65350000000
0!
0'
0/
#65360000000
#65370000000
1!
1'
1/
#65380000000
0!
0'
0/
#65390000000
1!
1'
1/
#65400000000
0!
1"
0'
1(
0/
10
#65410000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#65420000000
0!
0'
0/
#65430000000
1!
1'
1/
#65440000000
0!
0'
0/
#65450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#65460000000
0!
0'
0/
#65470000000
1!
1'
1/
#65480000000
0!
1"
0'
1(
0/
10
#65490000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#65500000000
0!
1$
0'
1+
0/
#65510000000
1!
1'
1/
#65520000000
0!
0'
0/
#65530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#65540000000
0!
0'
0/
#65550000000
1!
1'
1/
#65560000000
0!
0'
0/
#65570000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#65580000000
0!
0'
0/
#65590000000
1!
1'
1/
#65600000000
0!
0'
0/
#65610000000
1!
1'
1/
#65620000000
0!
0'
0/
#65630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#65640000000
0!
0'
0/
#65650000000
1!
1'
1/
#65660000000
0!
0'
0/
#65670000000
1!
1'
1/
#65680000000
0!
0'
0/
#65690000000
1!
1'
1/
#65700000000
0!
0'
0/
#65710000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#65720000000
0!
0'
0/
#65730000000
1!
1'
1/
#65740000000
0!
0'
0/
#65750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#65760000000
0!
0'
0/
#65770000000
1!
1'
1/
#65780000000
0!
0'
0/
#65790000000
#65800000000
1!
1'
1/
#65810000000
0!
0'
0/
#65820000000
1!
1'
1/
#65830000000
0!
1"
0'
1(
0/
10
#65840000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#65850000000
0!
0'
0/
#65860000000
1!
1'
1/
#65870000000
0!
0'
0/
#65880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#65890000000
0!
0'
0/
#65900000000
1!
1'
1/
#65910000000
0!
1"
0'
1(
0/
10
#65920000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#65930000000
0!
1$
0'
1+
0/
#65940000000
1!
1'
1/
#65950000000
0!
0'
0/
#65960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#65970000000
0!
0'
0/
#65980000000
1!
1'
1/
#65990000000
0!
0'
0/
#66000000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#66010000000
0!
0'
0/
#66020000000
1!
1'
1/
#66030000000
0!
0'
0/
#66040000000
1!
1'
1/
#66050000000
0!
0'
0/
#66060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#66070000000
0!
0'
0/
#66080000000
1!
1'
1/
#66090000000
0!
0'
0/
#66100000000
1!
1'
1/
#66110000000
0!
0'
0/
#66120000000
1!
1'
1/
#66130000000
0!
0'
0/
#66140000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#66150000000
0!
0'
0/
#66160000000
1!
1'
1/
#66170000000
0!
0'
0/
#66180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#66190000000
0!
0'
0/
#66200000000
1!
1'
1/
#66210000000
0!
0'
0/
#66220000000
#66230000000
1!
1'
1/
#66240000000
0!
0'
0/
#66250000000
1!
1'
1/
#66260000000
0!
1"
0'
1(
0/
10
#66270000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#66280000000
0!
0'
0/
#66290000000
1!
1'
1/
#66300000000
0!
0'
0/
#66310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#66320000000
0!
0'
0/
#66330000000
1!
1'
1/
#66340000000
0!
1"
0'
1(
0/
10
#66350000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#66360000000
0!
1$
0'
1+
0/
#66370000000
1!
1'
1/
#66380000000
0!
0'
0/
#66390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#66400000000
0!
0'
0/
#66410000000
1!
1'
1/
#66420000000
0!
0'
0/
#66430000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#66440000000
0!
0'
0/
#66450000000
1!
1'
1/
#66460000000
0!
0'
0/
#66470000000
1!
1'
1/
#66480000000
0!
0'
0/
#66490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#66500000000
0!
0'
0/
#66510000000
1!
1'
1/
#66520000000
0!
0'
0/
#66530000000
1!
1'
1/
#66540000000
0!
0'
0/
#66550000000
1!
1'
1/
#66560000000
0!
0'
0/
#66570000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#66580000000
0!
0'
0/
#66590000000
1!
1'
1/
#66600000000
0!
0'
0/
#66610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#66620000000
0!
0'
0/
#66630000000
1!
1'
1/
#66640000000
0!
0'
0/
#66650000000
#66660000000
1!
1'
1/
#66670000000
0!
0'
0/
#66680000000
1!
1'
1/
#66690000000
0!
1"
0'
1(
0/
10
#66700000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#66710000000
0!
0'
0/
#66720000000
1!
1'
1/
#66730000000
0!
0'
0/
#66740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#66750000000
0!
0'
0/
#66760000000
1!
1'
1/
#66770000000
0!
1"
0'
1(
0/
10
#66780000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#66790000000
0!
1$
0'
1+
0/
#66800000000
1!
1'
1/
#66810000000
0!
0'
0/
#66820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#66830000000
0!
0'
0/
#66840000000
1!
1'
1/
#66850000000
0!
0'
0/
#66860000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#66870000000
0!
0'
0/
#66880000000
1!
1'
1/
#66890000000
0!
0'
0/
#66900000000
1!
1'
1/
#66910000000
0!
0'
0/
#66920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#66930000000
0!
0'
0/
#66940000000
1!
1'
1/
#66950000000
0!
0'
0/
#66960000000
1!
1'
1/
#66970000000
0!
0'
0/
#66980000000
1!
1'
1/
#66990000000
0!
0'
0/
#67000000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#67010000000
0!
0'
0/
#67020000000
1!
1'
1/
#67030000000
0!
0'
0/
#67040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#67050000000
0!
0'
0/
#67060000000
1!
1'
1/
#67070000000
0!
0'
0/
#67080000000
#67090000000
1!
1'
1/
#67100000000
0!
0'
0/
#67110000000
1!
1'
1/
#67120000000
0!
1"
0'
1(
0/
10
#67130000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#67140000000
0!
0'
0/
#67150000000
1!
1'
1/
#67160000000
0!
0'
0/
#67170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#67180000000
0!
0'
0/
#67190000000
1!
1'
1/
#67200000000
0!
1"
0'
1(
0/
10
#67210000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#67220000000
0!
1$
0'
1+
0/
#67230000000
1!
1'
1/
#67240000000
0!
0'
0/
#67250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#67260000000
0!
0'
0/
#67270000000
1!
1'
1/
#67280000000
0!
0'
0/
#67290000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#67300000000
0!
0'
0/
#67310000000
1!
1'
1/
#67320000000
0!
0'
0/
#67330000000
1!
1'
1/
#67340000000
0!
0'
0/
#67350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#67360000000
0!
0'
0/
#67370000000
1!
1'
1/
#67380000000
0!
0'
0/
#67390000000
1!
1'
1/
#67400000000
0!
0'
0/
#67410000000
1!
1'
1/
#67420000000
0!
0'
0/
#67430000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#67440000000
0!
0'
0/
#67450000000
1!
1'
1/
#67460000000
0!
0'
0/
#67470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#67480000000
0!
0'
0/
#67490000000
1!
1'
1/
#67500000000
0!
0'
0/
#67510000000
#67520000000
1!
1'
1/
#67530000000
0!
0'
0/
#67540000000
1!
1'
1/
#67550000000
0!
1"
0'
1(
0/
10
#67560000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#67570000000
0!
0'
0/
#67580000000
1!
1'
1/
#67590000000
0!
0'
0/
#67600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#67610000000
0!
0'
0/
#67620000000
1!
1'
1/
#67630000000
0!
1"
0'
1(
0/
10
#67640000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#67650000000
0!
1$
0'
1+
0/
#67660000000
1!
1'
1/
#67670000000
0!
0'
0/
#67680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#67690000000
0!
0'
0/
#67700000000
1!
1'
1/
#67710000000
0!
0'
0/
#67720000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#67730000000
0!
0'
0/
#67740000000
1!
1'
1/
#67750000000
0!
0'
0/
#67760000000
1!
1'
1/
#67770000000
0!
0'
0/
#67780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#67790000000
0!
0'
0/
#67800000000
1!
1'
1/
#67810000000
0!
0'
0/
#67820000000
1!
1'
1/
#67830000000
0!
0'
0/
#67840000000
1!
1'
1/
#67850000000
0!
0'
0/
#67860000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#67870000000
0!
0'
0/
#67880000000
1!
1'
1/
#67890000000
0!
0'
0/
#67900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#67910000000
0!
0'
0/
#67920000000
1!
1'
1/
#67930000000
0!
0'
0/
#67940000000
#67950000000
1!
1'
1/
#67960000000
0!
0'
0/
#67970000000
1!
1'
1/
#67980000000
0!
1"
0'
1(
0/
10
#67990000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#68000000000
0!
0'
0/
#68010000000
1!
1'
1/
#68020000000
0!
0'
0/
#68030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#68040000000
0!
0'
0/
#68050000000
1!
1'
1/
#68060000000
0!
1"
0'
1(
0/
10
#68070000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#68080000000
0!
1$
0'
1+
0/
#68090000000
1!
1'
1/
#68100000000
0!
0'
0/
#68110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#68120000000
0!
0'
0/
#68130000000
1!
1'
1/
#68140000000
0!
0'
0/
#68150000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#68160000000
0!
0'
0/
#68170000000
1!
1'
1/
#68180000000
0!
0'
0/
#68190000000
1!
1'
1/
#68200000000
0!
0'
0/
#68210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#68220000000
0!
0'
0/
#68230000000
1!
1'
1/
#68240000000
0!
0'
0/
#68250000000
1!
1'
1/
#68260000000
0!
0'
0/
#68270000000
1!
1'
1/
#68280000000
0!
0'
0/
#68290000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#68300000000
0!
0'
0/
#68310000000
1!
1'
1/
#68320000000
0!
0'
0/
#68330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#68340000000
0!
0'
0/
#68350000000
1!
1'
1/
#68360000000
0!
0'
0/
#68370000000
#68380000000
1!
1'
1/
#68390000000
0!
0'
0/
#68400000000
1!
1'
1/
#68410000000
0!
1"
0'
1(
0/
10
#68420000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#68430000000
0!
0'
0/
#68440000000
1!
1'
1/
#68450000000
0!
0'
0/
#68460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#68470000000
0!
0'
0/
#68480000000
1!
1'
1/
#68490000000
0!
1"
0'
1(
0/
10
#68500000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#68510000000
0!
1$
0'
1+
0/
#68520000000
1!
1'
1/
#68530000000
0!
0'
0/
#68540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#68550000000
0!
0'
0/
#68560000000
1!
1'
1/
#68570000000
0!
0'
0/
#68580000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#68590000000
0!
0'
0/
#68600000000
1!
1'
1/
#68610000000
0!
0'
0/
#68620000000
1!
1'
1/
#68630000000
0!
0'
0/
#68640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#68650000000
0!
0'
0/
#68660000000
1!
1'
1/
#68670000000
0!
0'
0/
#68680000000
1!
1'
1/
#68690000000
0!
0'
0/
#68700000000
1!
1'
1/
#68710000000
0!
0'
0/
#68720000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#68730000000
0!
0'
0/
#68740000000
1!
1'
1/
#68750000000
0!
0'
0/
#68760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#68770000000
0!
0'
0/
#68780000000
1!
1'
1/
#68790000000
0!
0'
0/
#68800000000
#68810000000
1!
1'
1/
#68820000000
0!
0'
0/
#68830000000
1!
1'
1/
#68840000000
0!
1"
0'
1(
0/
10
#68850000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#68860000000
0!
0'
0/
#68870000000
1!
1'
1/
#68880000000
0!
0'
0/
#68890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#68900000000
0!
0'
0/
#68910000000
1!
1'
1/
#68920000000
0!
1"
0'
1(
0/
10
#68930000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#68940000000
0!
1$
0'
1+
0/
#68950000000
1!
1'
1/
#68960000000
0!
0'
0/
#68970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#68980000000
0!
0'
0/
#68990000000
1!
1'
1/
#69000000000
0!
0'
0/
#69010000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#69020000000
0!
0'
0/
#69030000000
1!
1'
1/
#69040000000
0!
0'
0/
#69050000000
1!
1'
1/
#69060000000
0!
0'
0/
#69070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#69080000000
0!
0'
0/
#69090000000
1!
1'
1/
#69100000000
0!
0'
0/
#69110000000
1!
1'
1/
#69120000000
0!
0'
0/
#69130000000
1!
1'
1/
#69140000000
0!
0'
0/
#69150000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#69160000000
0!
0'
0/
#69170000000
1!
1'
1/
#69180000000
0!
0'
0/
#69190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#69200000000
0!
0'
0/
#69210000000
1!
1'
1/
#69220000000
0!
0'
0/
#69230000000
#69240000000
1!
1'
1/
#69250000000
0!
0'
0/
#69260000000
1!
1'
1/
#69270000000
0!
1"
0'
1(
0/
10
#69280000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#69290000000
0!
0'
0/
#69300000000
1!
1'
1/
#69310000000
0!
0'
0/
#69320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#69330000000
0!
0'
0/
#69340000000
1!
1'
1/
#69350000000
0!
1"
0'
1(
0/
10
#69360000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#69370000000
0!
1$
0'
1+
0/
#69380000000
1!
1'
1/
#69390000000
0!
0'
0/
#69400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#69410000000
0!
0'
0/
#69420000000
1!
1'
1/
#69430000000
0!
0'
0/
#69440000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#69450000000
0!
0'
0/
#69460000000
1!
1'
1/
#69470000000
0!
0'
0/
#69480000000
1!
1'
1/
#69490000000
0!
0'
0/
#69500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#69510000000
0!
0'
0/
#69520000000
1!
1'
1/
#69530000000
0!
0'
0/
#69540000000
1!
1'
1/
#69550000000
0!
0'
0/
#69560000000
1!
1'
1/
#69570000000
0!
0'
0/
#69580000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#69590000000
0!
0'
0/
#69600000000
1!
1'
1/
#69610000000
0!
0'
0/
#69620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#69630000000
0!
0'
0/
#69640000000
1!
1'
1/
#69650000000
0!
0'
0/
#69660000000
#69670000000
1!
1'
1/
#69680000000
0!
0'
0/
#69690000000
1!
1'
1/
#69700000000
0!
1"
0'
1(
0/
10
#69710000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#69720000000
0!
0'
0/
#69730000000
1!
1'
1/
#69740000000
0!
0'
0/
#69750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#69760000000
0!
0'
0/
#69770000000
1!
1'
1/
#69780000000
0!
1"
0'
1(
0/
10
#69790000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#69800000000
0!
1$
0'
1+
0/
#69810000000
1!
1'
1/
#69820000000
0!
0'
0/
#69830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#69840000000
0!
0'
0/
#69850000000
1!
1'
1/
#69860000000
0!
0'
0/
#69870000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#69880000000
0!
0'
0/
#69890000000
1!
1'
1/
#69900000000
0!
0'
0/
#69910000000
1!
1'
1/
#69920000000
0!
0'
0/
#69930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#69940000000
0!
0'
0/
#69950000000
1!
1'
1/
#69960000000
0!
0'
0/
#69970000000
1!
1'
1/
#69980000000
0!
0'
0/
#69990000000
1!
1'
1/
#70000000000
0!
0'
0/
#70010000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#70020000000
0!
0'
0/
#70030000000
1!
1'
1/
#70040000000
0!
0'
0/
#70050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#70060000000
0!
0'
0/
#70070000000
1!
1'
1/
#70080000000
0!
0'
0/
#70090000000
#70100000000
1!
1'
1/
#70110000000
0!
0'
0/
#70120000000
1!
1'
1/
#70130000000
0!
1"
0'
1(
0/
10
#70140000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#70150000000
0!
0'
0/
#70160000000
1!
1'
1/
#70170000000
0!
0'
0/
#70180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#70190000000
0!
0'
0/
#70200000000
1!
1'
1/
#70210000000
0!
1"
0'
1(
0/
10
#70220000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#70230000000
0!
1$
0'
1+
0/
#70240000000
1!
1'
1/
#70250000000
0!
0'
0/
#70260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#70270000000
0!
0'
0/
#70280000000
1!
1'
1/
#70290000000
0!
0'
0/
#70300000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#70310000000
0!
0'
0/
#70320000000
1!
1'
1/
#70330000000
0!
0'
0/
#70340000000
1!
1'
1/
#70350000000
0!
0'
0/
#70360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#70370000000
0!
0'
0/
#70380000000
1!
1'
1/
#70390000000
0!
0'
0/
#70400000000
1!
1'
1/
#70410000000
0!
0'
0/
#70420000000
1!
1'
1/
#70430000000
0!
0'
0/
#70440000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#70450000000
0!
0'
0/
#70460000000
1!
1'
1/
#70470000000
0!
0'
0/
#70480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#70490000000
0!
0'
0/
#70500000000
1!
1'
1/
#70510000000
0!
0'
0/
#70520000000
#70530000000
1!
1'
1/
#70540000000
0!
0'
0/
#70550000000
1!
1'
1/
#70560000000
0!
1"
0'
1(
0/
10
#70570000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#70580000000
0!
0'
0/
#70590000000
1!
1'
1/
#70600000000
0!
0'
0/
#70610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#70620000000
0!
0'
0/
#70630000000
1!
1'
1/
#70640000000
0!
1"
0'
1(
0/
10
#70650000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#70660000000
0!
1$
0'
1+
0/
#70670000000
1!
1'
1/
#70680000000
0!
0'
0/
#70690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#70700000000
0!
0'
0/
#70710000000
1!
1'
1/
#70720000000
0!
0'
0/
#70730000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#70740000000
0!
0'
0/
#70750000000
1!
1'
1/
#70760000000
0!
0'
0/
#70770000000
1!
1'
1/
#70780000000
0!
0'
0/
#70790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#70800000000
0!
0'
0/
#70810000000
1!
1'
1/
#70820000000
0!
0'
0/
#70830000000
1!
1'
1/
#70840000000
0!
0'
0/
#70850000000
1!
1'
1/
#70860000000
0!
0'
0/
#70870000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#70880000000
0!
0'
0/
#70890000000
1!
1'
1/
#70900000000
0!
0'
0/
#70910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#70920000000
0!
0'
0/
#70930000000
1!
1'
1/
#70940000000
0!
0'
0/
#70950000000
#70960000000
1!
1'
1/
#70970000000
0!
0'
0/
#70980000000
1!
1'
1/
#70990000000
0!
1"
0'
1(
0/
10
#71000000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#71010000000
0!
0'
0/
#71020000000
1!
1'
1/
#71030000000
0!
0'
0/
#71040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#71050000000
0!
0'
0/
#71060000000
1!
1'
1/
#71070000000
0!
1"
0'
1(
0/
10
#71080000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#71090000000
0!
1$
0'
1+
0/
#71100000000
1!
1'
1/
#71110000000
0!
0'
0/
#71120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#71130000000
0!
0'
0/
#71140000000
1!
1'
1/
#71150000000
0!
0'
0/
#71160000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#71170000000
0!
0'
0/
#71180000000
1!
1'
1/
#71190000000
0!
0'
0/
#71200000000
1!
1'
1/
#71210000000
0!
0'
0/
#71220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#71230000000
0!
0'
0/
#71240000000
1!
1'
1/
#71250000000
0!
0'
0/
#71260000000
1!
1'
1/
#71270000000
0!
0'
0/
#71280000000
1!
1'
1/
#71290000000
0!
0'
0/
#71300000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#71310000000
0!
0'
0/
#71320000000
1!
1'
1/
#71330000000
0!
0'
0/
#71340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#71350000000
0!
0'
0/
#71360000000
1!
1'
1/
#71370000000
0!
0'
0/
#71380000000
#71390000000
1!
1'
1/
#71400000000
0!
0'
0/
#71410000000
1!
1'
1/
#71420000000
0!
1"
0'
1(
0/
10
#71430000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#71440000000
0!
0'
0/
#71450000000
1!
1'
1/
#71460000000
0!
0'
0/
#71470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#71480000000
0!
0'
0/
#71490000000
1!
1'
1/
#71500000000
0!
1"
0'
1(
0/
10
#71510000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#71520000000
0!
1$
0'
1+
0/
#71530000000
1!
1'
1/
#71540000000
0!
0'
0/
#71550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#71560000000
0!
0'
0/
#71570000000
1!
1'
1/
#71580000000
0!
0'
0/
#71590000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#71600000000
0!
0'
0/
#71610000000
1!
1'
1/
#71620000000
0!
0'
0/
#71630000000
1!
1'
1/
#71640000000
0!
0'
0/
#71650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#71660000000
0!
0'
0/
#71670000000
1!
1'
1/
#71680000000
0!
0'
0/
#71690000000
1!
1'
1/
#71700000000
0!
0'
0/
#71710000000
1!
1'
1/
#71720000000
0!
0'
0/
#71730000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#71740000000
0!
0'
0/
#71750000000
1!
1'
1/
#71760000000
0!
0'
0/
#71770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#71780000000
0!
0'
0/
#71790000000
1!
1'
1/
#71800000000
0!
0'
0/
#71810000000
#71820000000
1!
1'
1/
#71830000000
0!
0'
0/
#71840000000
1!
1'
1/
#71850000000
0!
1"
0'
1(
0/
10
#71860000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#71870000000
0!
0'
0/
#71880000000
1!
1'
1/
#71890000000
0!
0'
0/
#71900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#71910000000
0!
0'
0/
#71920000000
1!
1'
1/
#71930000000
0!
1"
0'
1(
0/
10
#71940000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#71950000000
0!
1$
0'
1+
0/
#71960000000
1!
1'
1/
#71970000000
0!
0'
0/
#71980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#71990000000
0!
0'
0/
#72000000000
1!
1'
1/
#72010000000
0!
0'
0/
#72020000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#72030000000
0!
0'
0/
#72040000000
1!
1'
1/
#72050000000
0!
0'
0/
#72060000000
1!
1'
1/
#72070000000
0!
0'
0/
#72080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#72090000000
0!
0'
0/
#72100000000
1!
1'
1/
#72110000000
0!
0'
0/
#72120000000
1!
1'
1/
#72130000000
0!
0'
0/
#72140000000
1!
1'
1/
#72150000000
0!
0'
0/
#72160000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#72170000000
0!
0'
0/
#72180000000
1!
1'
1/
#72190000000
0!
0'
0/
#72200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#72210000000
0!
0'
0/
#72220000000
1!
1'
1/
#72230000000
0!
0'
0/
#72240000000
#72250000000
1!
1'
1/
#72260000000
0!
0'
0/
#72270000000
1!
1'
1/
#72280000000
0!
1"
0'
1(
0/
10
#72290000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#72300000000
0!
0'
0/
#72310000000
1!
1'
1/
#72320000000
0!
0'
0/
#72330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#72340000000
0!
0'
0/
#72350000000
1!
1'
1/
#72360000000
0!
1"
0'
1(
0/
10
#72370000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#72380000000
0!
1$
0'
1+
0/
#72390000000
1!
1'
1/
#72400000000
0!
0'
0/
#72410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#72420000000
0!
0'
0/
#72430000000
1!
1'
1/
#72440000000
0!
0'
0/
#72450000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#72460000000
0!
0'
0/
#72470000000
1!
1'
1/
#72480000000
0!
0'
0/
#72490000000
1!
1'
1/
#72500000000
0!
0'
0/
#72510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#72520000000
0!
0'
0/
#72530000000
1!
1'
1/
#72540000000
0!
0'
0/
#72550000000
1!
1'
1/
#72560000000
0!
0'
0/
#72570000000
1!
1'
1/
#72580000000
0!
0'
0/
#72590000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#72600000000
0!
0'
0/
#72610000000
1!
1'
1/
#72620000000
0!
0'
0/
#72630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#72640000000
0!
0'
0/
#72650000000
1!
1'
1/
#72660000000
0!
0'
0/
#72670000000
#72680000000
1!
1'
1/
#72690000000
0!
0'
0/
#72700000000
1!
1'
1/
#72710000000
0!
1"
0'
1(
0/
10
#72720000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#72730000000
0!
0'
0/
#72740000000
1!
1'
1/
#72750000000
0!
0'
0/
#72760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#72770000000
0!
0'
0/
#72780000000
1!
1'
1/
#72790000000
0!
1"
0'
1(
0/
10
#72800000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#72810000000
0!
1$
0'
1+
0/
#72820000000
1!
1'
1/
#72830000000
0!
0'
0/
#72840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#72850000000
0!
0'
0/
#72860000000
1!
1'
1/
#72870000000
0!
0'
0/
#72880000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#72890000000
0!
0'
0/
#72900000000
1!
1'
1/
#72910000000
0!
0'
0/
#72920000000
1!
1'
1/
#72930000000
0!
0'
0/
#72940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#72950000000
0!
0'
0/
#72960000000
1!
1'
1/
#72970000000
0!
0'
0/
#72980000000
1!
1'
1/
#72990000000
0!
0'
0/
#73000000000
1!
1'
1/
#73010000000
0!
0'
0/
#73020000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#73030000000
0!
0'
0/
#73040000000
1!
1'
1/
#73050000000
0!
0'
0/
#73060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#73070000000
0!
0'
0/
#73080000000
1!
1'
1/
#73090000000
0!
0'
0/
#73100000000
#73110000000
1!
1'
1/
#73120000000
0!
0'
0/
#73130000000
1!
1'
1/
#73140000000
0!
1"
0'
1(
0/
10
#73150000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#73160000000
0!
0'
0/
#73170000000
1!
1'
1/
#73180000000
0!
0'
0/
#73190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#73200000000
0!
0'
0/
#73210000000
1!
1'
1/
#73220000000
0!
1"
0'
1(
0/
10
#73230000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#73240000000
0!
1$
0'
1+
0/
#73250000000
1!
1'
1/
#73260000000
0!
0'
0/
#73270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#73280000000
0!
0'
0/
#73290000000
1!
1'
1/
#73300000000
0!
0'
0/
#73310000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#73320000000
0!
0'
0/
#73330000000
1!
1'
1/
#73340000000
0!
0'
0/
#73350000000
1!
1'
1/
#73360000000
0!
0'
0/
#73370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#73380000000
0!
0'
0/
#73390000000
1!
1'
1/
#73400000000
0!
0'
0/
#73410000000
1!
1'
1/
#73420000000
0!
0'
0/
#73430000000
1!
1'
1/
#73440000000
0!
0'
0/
#73450000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#73460000000
0!
0'
0/
#73470000000
1!
1'
1/
#73480000000
0!
0'
0/
#73490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#73500000000
0!
0'
0/
#73510000000
1!
1'
1/
#73520000000
0!
0'
0/
#73530000000
#73540000000
1!
1'
1/
#73550000000
0!
0'
0/
#73560000000
1!
1'
1/
#73570000000
0!
1"
0'
1(
0/
10
#73580000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#73590000000
0!
0'
0/
#73600000000
1!
1'
1/
#73610000000
0!
0'
0/
#73620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#73630000000
0!
0'
0/
#73640000000
1!
1'
1/
#73650000000
0!
1"
0'
1(
0/
10
#73660000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#73670000000
0!
1$
0'
1+
0/
#73680000000
1!
1'
1/
#73690000000
0!
0'
0/
#73700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#73710000000
0!
0'
0/
#73720000000
1!
1'
1/
#73730000000
0!
0'
0/
#73740000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#73750000000
0!
0'
0/
#73760000000
1!
1'
1/
#73770000000
0!
0'
0/
#73780000000
1!
1'
1/
#73790000000
0!
0'
0/
#73800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#73810000000
0!
0'
0/
#73820000000
1!
1'
1/
#73830000000
0!
0'
0/
#73840000000
1!
1'
1/
#73850000000
0!
0'
0/
#73860000000
1!
1'
1/
#73870000000
0!
0'
0/
#73880000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#73890000000
0!
0'
0/
#73900000000
1!
1'
1/
#73910000000
0!
0'
0/
#73920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#73930000000
0!
0'
0/
#73940000000
1!
1'
1/
#73950000000
0!
0'
0/
#73960000000
#73970000000
1!
1'
1/
#73980000000
0!
0'
0/
#73990000000
1!
1'
1/
#74000000000
0!
1"
0'
1(
0/
10
#74010000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#74020000000
0!
0'
0/
#74030000000
1!
1'
1/
#74040000000
0!
0'
0/
#74050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#74060000000
0!
0'
0/
#74070000000
1!
1'
1/
#74080000000
0!
1"
0'
1(
0/
10
#74090000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#74100000000
0!
1$
0'
1+
0/
#74110000000
1!
1'
1/
#74120000000
0!
0'
0/
#74130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#74140000000
0!
0'
0/
#74150000000
1!
1'
1/
#74160000000
0!
0'
0/
#74170000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#74180000000
0!
0'
0/
#74190000000
1!
1'
1/
#74200000000
0!
0'
0/
#74210000000
1!
1'
1/
#74220000000
0!
0'
0/
#74230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#74240000000
0!
0'
0/
#74250000000
1!
1'
1/
#74260000000
0!
0'
0/
#74270000000
1!
1'
1/
#74280000000
0!
0'
0/
#74290000000
1!
1'
1/
#74300000000
0!
0'
0/
#74310000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#74320000000
0!
0'
0/
#74330000000
1!
1'
1/
#74340000000
0!
0'
0/
#74350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#74360000000
0!
0'
0/
#74370000000
1!
1'
1/
#74380000000
0!
0'
0/
#74390000000
#74400000000
1!
1'
1/
#74410000000
0!
0'
0/
#74420000000
1!
1'
1/
#74430000000
0!
1"
0'
1(
0/
10
#74440000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#74450000000
0!
0'
0/
#74460000000
1!
1'
1/
#74470000000
0!
0'
0/
#74480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#74490000000
0!
0'
0/
#74500000000
1!
1'
1/
#74510000000
0!
1"
0'
1(
0/
10
#74520000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#74530000000
0!
1$
0'
1+
0/
#74540000000
1!
1'
1/
#74550000000
0!
0'
0/
#74560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#74570000000
0!
0'
0/
#74580000000
1!
1'
1/
#74590000000
0!
0'
0/
#74600000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#74610000000
0!
0'
0/
#74620000000
1!
1'
1/
#74630000000
0!
0'
0/
#74640000000
1!
1'
1/
#74650000000
0!
0'
0/
#74660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#74670000000
0!
0'
0/
#74680000000
1!
1'
1/
#74690000000
0!
0'
0/
#74700000000
1!
1'
1/
#74710000000
0!
0'
0/
#74720000000
1!
1'
1/
#74730000000
0!
0'
0/
#74740000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#74750000000
0!
0'
0/
#74760000000
1!
1'
1/
#74770000000
0!
0'
0/
#74780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#74790000000
0!
0'
0/
#74800000000
1!
1'
1/
#74810000000
0!
0'
0/
#74820000000
#74830000000
1!
1'
1/
#74840000000
0!
0'
0/
#74850000000
1!
1'
1/
#74860000000
0!
1"
0'
1(
0/
10
#74870000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#74880000000
0!
0'
0/
#74890000000
1!
1'
1/
#74900000000
0!
0'
0/
#74910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#74920000000
0!
0'
0/
#74930000000
1!
1'
1/
#74940000000
0!
1"
0'
1(
0/
10
#74950000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#74960000000
0!
1$
0'
1+
0/
#74970000000
1!
1'
1/
#74980000000
0!
0'
0/
#74990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#75000000000
0!
0'
0/
#75010000000
1!
1'
1/
#75020000000
0!
0'
0/
#75030000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#75040000000
0!
0'
0/
#75050000000
1!
1'
1/
#75060000000
0!
0'
0/
#75070000000
1!
1'
1/
#75080000000
0!
0'
0/
#75090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#75100000000
0!
0'
0/
#75110000000
1!
1'
1/
#75120000000
0!
0'
0/
#75130000000
1!
1'
1/
#75140000000
0!
0'
0/
#75150000000
1!
1'
1/
#75160000000
0!
0'
0/
#75170000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#75180000000
0!
0'
0/
#75190000000
1!
1'
1/
#75200000000
0!
0'
0/
#75210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#75220000000
0!
0'
0/
#75230000000
1!
1'
1/
#75240000000
0!
0'
0/
#75250000000
#75260000000
1!
1'
1/
#75270000000
0!
0'
0/
#75280000000
1!
1'
1/
#75290000000
0!
1"
0'
1(
0/
10
#75300000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#75310000000
0!
0'
0/
#75320000000
1!
1'
1/
#75330000000
0!
0'
0/
#75340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#75350000000
0!
0'
0/
#75360000000
1!
1'
1/
#75370000000
0!
1"
0'
1(
0/
10
#75380000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#75390000000
0!
1$
0'
1+
0/
#75400000000
1!
1'
1/
#75410000000
0!
0'
0/
#75420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#75430000000
0!
0'
0/
#75440000000
1!
1'
1/
#75450000000
0!
0'
0/
#75460000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#75470000000
0!
0'
0/
#75480000000
1!
1'
1/
#75490000000
0!
0'
0/
#75500000000
1!
1'
1/
#75510000000
0!
0'
0/
#75520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#75530000000
0!
0'
0/
#75540000000
1!
1'
1/
#75550000000
0!
0'
0/
#75560000000
1!
1'
1/
#75570000000
0!
0'
0/
#75580000000
1!
1'
1/
#75590000000
0!
0'
0/
#75600000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#75610000000
0!
0'
0/
#75620000000
1!
1'
1/
#75630000000
0!
0'
0/
#75640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#75650000000
0!
0'
0/
#75660000000
1!
1'
1/
#75670000000
0!
0'
0/
#75680000000
#75690000000
1!
1'
1/
#75700000000
0!
0'
0/
#75710000000
1!
1'
1/
#75720000000
0!
1"
0'
1(
0/
10
#75730000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#75740000000
0!
0'
0/
#75750000000
1!
1'
1/
#75760000000
0!
0'
0/
#75770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#75780000000
0!
0'
0/
#75790000000
1!
1'
1/
#75800000000
0!
1"
0'
1(
0/
10
#75810000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#75820000000
0!
1$
0'
1+
0/
#75830000000
1!
1'
1/
#75840000000
0!
0'
0/
#75850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#75860000000
0!
0'
0/
#75870000000
1!
1'
1/
#75880000000
0!
0'
0/
#75890000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#75900000000
0!
0'
0/
#75910000000
1!
1'
1/
#75920000000
0!
0'
0/
#75930000000
1!
1'
1/
#75940000000
0!
0'
0/
#75950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#75960000000
0!
0'
0/
#75970000000
1!
1'
1/
#75980000000
0!
0'
0/
#75990000000
1!
1'
1/
#76000000000
0!
0'
0/
#76010000000
1!
1'
1/
#76020000000
0!
0'
0/
#76030000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#76040000000
0!
0'
0/
#76050000000
1!
1'
1/
#76060000000
0!
0'
0/
#76070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#76080000000
0!
0'
0/
#76090000000
1!
1'
1/
#76100000000
0!
0'
0/
#76110000000
#76120000000
1!
1'
1/
#76130000000
0!
0'
0/
#76140000000
1!
1'
1/
#76150000000
0!
1"
0'
1(
0/
10
#76160000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#76170000000
0!
0'
0/
#76180000000
1!
1'
1/
#76190000000
0!
0'
0/
#76200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#76210000000
0!
0'
0/
#76220000000
1!
1'
1/
#76230000000
0!
1"
0'
1(
0/
10
#76240000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#76250000000
0!
1$
0'
1+
0/
#76260000000
1!
1'
1/
#76270000000
0!
0'
0/
#76280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#76290000000
0!
0'
0/
#76300000000
1!
1'
1/
#76310000000
0!
0'
0/
#76320000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#76330000000
0!
0'
0/
#76340000000
1!
1'
1/
#76350000000
0!
0'
0/
#76360000000
1!
1'
1/
#76370000000
0!
0'
0/
#76380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#76390000000
0!
0'
0/
#76400000000
1!
1'
1/
#76410000000
0!
0'
0/
#76420000000
1!
1'
1/
#76430000000
0!
0'
0/
#76440000000
1!
1'
1/
#76450000000
0!
0'
0/
#76460000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#76470000000
0!
0'
0/
#76480000000
1!
1'
1/
#76490000000
0!
0'
0/
#76500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#76510000000
0!
0'
0/
#76520000000
1!
1'
1/
#76530000000
0!
0'
0/
#76540000000
#76550000000
1!
1'
1/
#76560000000
0!
0'
0/
#76570000000
1!
1'
1/
#76580000000
0!
1"
0'
1(
0/
10
#76590000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#76600000000
0!
0'
0/
#76610000000
1!
1'
1/
#76620000000
0!
0'
0/
#76630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#76640000000
0!
0'
0/
#76650000000
1!
1'
1/
#76660000000
0!
1"
0'
1(
0/
10
#76670000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#76680000000
0!
1$
0'
1+
0/
#76690000000
1!
1'
1/
#76700000000
0!
0'
0/
#76710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#76720000000
0!
0'
0/
#76730000000
1!
1'
1/
#76740000000
0!
0'
0/
#76750000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#76760000000
0!
0'
0/
#76770000000
1!
1'
1/
#76780000000
0!
0'
0/
#76790000000
1!
1'
1/
#76800000000
0!
0'
0/
#76810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#76820000000
0!
0'
0/
#76830000000
1!
1'
1/
#76840000000
0!
0'
0/
#76850000000
1!
1'
1/
#76860000000
0!
0'
0/
#76870000000
1!
1'
1/
#76880000000
0!
0'
0/
#76890000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#76900000000
0!
0'
0/
#76910000000
1!
1'
1/
#76920000000
0!
0'
0/
#76930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#76940000000
0!
0'
0/
#76950000000
1!
1'
1/
#76960000000
0!
0'
0/
#76970000000
#76980000000
1!
1'
1/
#76990000000
0!
0'
0/
#77000000000
1!
1'
1/
#77010000000
0!
1"
0'
1(
0/
10
#77020000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#77030000000
0!
0'
0/
#77040000000
1!
1'
1/
#77050000000
0!
0'
0/
#77060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#77070000000
0!
0'
0/
#77080000000
1!
1'
1/
#77090000000
0!
1"
0'
1(
0/
10
#77100000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#77110000000
0!
1$
0'
1+
0/
#77120000000
1!
1'
1/
#77130000000
0!
0'
0/
#77140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#77150000000
0!
0'
0/
#77160000000
1!
1'
1/
#77170000000
0!
0'
0/
#77180000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#77190000000
0!
0'
0/
#77200000000
1!
1'
1/
#77210000000
0!
0'
0/
#77220000000
1!
1'
1/
#77230000000
0!
0'
0/
#77240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#77250000000
0!
0'
0/
#77260000000
1!
1'
1/
#77270000000
0!
0'
0/
#77280000000
1!
1'
1/
#77290000000
0!
0'
0/
#77300000000
1!
1'
1/
#77310000000
0!
0'
0/
#77320000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#77330000000
0!
0'
0/
#77340000000
1!
1'
1/
#77350000000
0!
0'
0/
#77360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#77370000000
0!
0'
0/
#77380000000
1!
1'
1/
#77390000000
0!
0'
0/
#77400000000
#77410000000
1!
1'
1/
#77420000000
0!
0'
0/
#77430000000
1!
1'
1/
#77440000000
0!
1"
0'
1(
0/
10
#77450000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#77460000000
0!
0'
0/
#77470000000
1!
1'
1/
#77480000000
0!
0'
0/
#77490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#77500000000
0!
0'
0/
#77510000000
1!
1'
1/
#77520000000
0!
1"
0'
1(
0/
10
#77530000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#77540000000
0!
1$
0'
1+
0/
#77550000000
1!
1'
1/
#77560000000
0!
0'
0/
#77570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#77580000000
0!
0'
0/
#77590000000
1!
1'
1/
#77600000000
0!
0'
0/
#77610000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#77620000000
0!
0'
0/
#77630000000
1!
1'
1/
#77640000000
0!
0'
0/
#77650000000
1!
1'
1/
#77660000000
0!
0'
0/
#77670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#77680000000
0!
0'
0/
#77690000000
1!
1'
1/
#77700000000
0!
0'
0/
#77710000000
1!
1'
1/
#77720000000
0!
0'
0/
#77730000000
1!
1'
1/
#77740000000
0!
0'
0/
#77750000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#77760000000
0!
0'
0/
#77770000000
1!
1'
1/
#77780000000
0!
0'
0/
#77790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#77800000000
0!
0'
0/
#77810000000
1!
1'
1/
#77820000000
0!
0'
0/
#77830000000
#77840000000
1!
1'
1/
#77850000000
0!
0'
0/
#77860000000
1!
1'
1/
#77870000000
0!
1"
0'
1(
0/
10
#77880000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#77890000000
0!
0'
0/
#77900000000
1!
1'
1/
#77910000000
0!
0'
0/
#77920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#77930000000
0!
0'
0/
#77940000000
1!
1'
1/
#77950000000
0!
1"
0'
1(
0/
10
#77960000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#77970000000
0!
1$
0'
1+
0/
#77980000000
1!
1'
1/
#77990000000
0!
0'
0/
#78000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#78010000000
0!
0'
0/
#78020000000
1!
1'
1/
#78030000000
0!
0'
0/
#78040000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#78050000000
0!
0'
0/
#78060000000
1!
1'
1/
#78070000000
0!
0'
0/
#78080000000
1!
1'
1/
#78090000000
0!
0'
0/
#78100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#78110000000
0!
0'
0/
#78120000000
1!
1'
1/
#78130000000
0!
0'
0/
#78140000000
1!
1'
1/
#78150000000
0!
0'
0/
#78160000000
1!
1'
1/
#78170000000
0!
0'
0/
#78180000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#78190000000
0!
0'
0/
#78200000000
1!
1'
1/
#78210000000
0!
0'
0/
#78220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#78230000000
0!
0'
0/
#78240000000
1!
1'
1/
#78250000000
0!
0'
0/
#78260000000
#78270000000
1!
1'
1/
#78280000000
0!
0'
0/
#78290000000
1!
1'
1/
#78300000000
0!
1"
0'
1(
0/
10
#78310000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#78320000000
0!
0'
0/
#78330000000
1!
1'
1/
#78340000000
0!
0'
0/
#78350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#78360000000
0!
0'
0/
#78370000000
1!
1'
1/
#78380000000
0!
1"
0'
1(
0/
10
#78390000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#78400000000
0!
1$
0'
1+
0/
#78410000000
1!
1'
1/
#78420000000
0!
0'
0/
#78430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#78440000000
0!
0'
0/
#78450000000
1!
1'
1/
#78460000000
0!
0'
0/
#78470000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#78480000000
0!
0'
0/
#78490000000
1!
1'
1/
#78500000000
0!
0'
0/
#78510000000
1!
1'
1/
#78520000000
0!
0'
0/
#78530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#78540000000
0!
0'
0/
#78550000000
1!
1'
1/
#78560000000
0!
0'
0/
#78570000000
1!
1'
1/
#78580000000
0!
0'
0/
#78590000000
1!
1'
1/
#78600000000
0!
0'
0/
#78610000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#78620000000
0!
0'
0/
#78630000000
1!
1'
1/
#78640000000
0!
0'
0/
#78650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#78660000000
0!
0'
0/
#78670000000
1!
1'
1/
#78680000000
0!
0'
0/
#78690000000
#78700000000
1!
1'
1/
#78710000000
0!
0'
0/
#78720000000
1!
1'
1/
#78730000000
0!
1"
0'
1(
0/
10
#78740000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#78750000000
0!
0'
0/
#78760000000
1!
1'
1/
#78770000000
0!
0'
0/
#78780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#78790000000
0!
0'
0/
#78800000000
1!
1'
1/
#78810000000
0!
1"
0'
1(
0/
10
#78820000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#78830000000
0!
1$
0'
1+
0/
#78840000000
1!
1'
1/
#78850000000
0!
0'
0/
#78860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#78870000000
0!
0'
0/
#78880000000
1!
1'
1/
#78890000000
0!
0'
0/
#78900000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#78910000000
0!
0'
0/
#78920000000
1!
1'
1/
#78930000000
0!
0'
0/
#78940000000
1!
1'
1/
#78950000000
0!
0'
0/
#78960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#78970000000
0!
0'
0/
#78980000000
1!
1'
1/
#78990000000
0!
0'
0/
#79000000000
1!
1'
1/
#79010000000
0!
0'
0/
#79020000000
1!
1'
1/
#79030000000
0!
0'
0/
#79040000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#79050000000
0!
0'
0/
#79060000000
1!
1'
1/
#79070000000
0!
0'
0/
#79080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#79090000000
0!
0'
0/
#79100000000
1!
1'
1/
#79110000000
0!
0'
0/
#79120000000
#79130000000
1!
1'
1/
#79140000000
0!
0'
0/
#79150000000
1!
1'
1/
#79160000000
0!
1"
0'
1(
0/
10
#79170000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#79180000000
0!
0'
0/
#79190000000
1!
1'
1/
#79200000000
0!
0'
0/
#79210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#79220000000
0!
0'
0/
#79230000000
1!
1'
1/
#79240000000
0!
1"
0'
1(
0/
10
#79250000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#79260000000
0!
1$
0'
1+
0/
#79270000000
1!
1'
1/
#79280000000
0!
0'
0/
#79290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#79300000000
0!
0'
0/
#79310000000
1!
1'
1/
#79320000000
0!
0'
0/
#79330000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#79340000000
0!
0'
0/
#79350000000
1!
1'
1/
#79360000000
0!
0'
0/
#79370000000
1!
1'
1/
#79380000000
0!
0'
0/
#79390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#79400000000
0!
0'
0/
#79410000000
1!
1'
1/
#79420000000
0!
0'
0/
#79430000000
1!
1'
1/
#79440000000
0!
0'
0/
#79450000000
1!
1'
1/
#79460000000
0!
0'
0/
#79470000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#79480000000
0!
0'
0/
#79490000000
1!
1'
1/
#79500000000
0!
0'
0/
#79510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#79520000000
0!
0'
0/
#79530000000
1!
1'
1/
#79540000000
0!
0'
0/
#79550000000
#79560000000
1!
1'
1/
#79570000000
0!
0'
0/
#79580000000
1!
1'
1/
#79590000000
0!
1"
0'
1(
0/
10
#79600000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#79610000000
0!
0'
0/
#79620000000
1!
1'
1/
#79630000000
0!
0'
0/
#79640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#79650000000
0!
0'
0/
#79660000000
1!
1'
1/
#79670000000
0!
1"
0'
1(
0/
10
#79680000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#79690000000
0!
1$
0'
1+
0/
#79700000000
1!
1'
1/
#79710000000
0!
0'
0/
#79720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#79730000000
0!
0'
0/
#79740000000
1!
1'
1/
#79750000000
0!
0'
0/
#79760000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#79770000000
0!
0'
0/
#79780000000
1!
1'
1/
#79790000000
0!
0'
0/
#79800000000
1!
1'
1/
#79810000000
0!
0'
0/
#79820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#79830000000
0!
0'
0/
#79840000000
1!
1'
1/
#79850000000
0!
0'
0/
#79860000000
1!
1'
1/
#79870000000
0!
0'
0/
#79880000000
1!
1'
1/
#79890000000
0!
0'
0/
#79900000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#79910000000
0!
0'
0/
#79920000000
1!
1'
1/
#79930000000
0!
0'
0/
#79940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#79950000000
0!
0'
0/
#79960000000
1!
1'
1/
#79970000000
0!
0'
0/
#79980000000
#79990000000
1!
1'
1/
#80000000000
0!
0'
0/
#80010000000
1!
1'
1/
#80020000000
0!
1"
0'
1(
0/
10
#80030000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#80040000000
0!
0'
0/
#80050000000
1!
1'
1/
#80060000000
0!
0'
0/
#80070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#80080000000
0!
0'
0/
#80090000000
1!
1'
1/
#80100000000
0!
1"
0'
1(
0/
10
#80110000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#80120000000
0!
1$
0'
1+
0/
#80130000000
1!
1'
1/
#80140000000
0!
0'
0/
#80150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#80160000000
0!
0'
0/
#80170000000
1!
1'
1/
#80180000000
0!
0'
0/
#80190000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#80200000000
0!
0'
0/
#80210000000
1!
1'
1/
#80220000000
0!
0'
0/
#80230000000
1!
1'
1/
#80240000000
0!
0'
0/
#80250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#80260000000
0!
0'
0/
#80270000000
1!
1'
1/
#80280000000
0!
0'
0/
#80290000000
1!
1'
1/
#80300000000
0!
0'
0/
#80310000000
1!
1'
1/
#80320000000
0!
0'
0/
#80330000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#80340000000
0!
0'
0/
#80350000000
1!
1'
1/
#80360000000
0!
0'
0/
#80370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#80380000000
0!
0'
0/
#80390000000
1!
1'
1/
#80400000000
0!
0'
0/
#80410000000
#80420000000
1!
1'
1/
#80430000000
0!
0'
0/
#80440000000
1!
1'
1/
#80450000000
0!
1"
0'
1(
0/
10
#80460000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#80470000000
0!
0'
0/
#80480000000
1!
1'
1/
#80490000000
0!
0'
0/
#80500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#80510000000
0!
0'
0/
#80520000000
1!
1'
1/
#80530000000
0!
1"
0'
1(
0/
10
#80540000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#80550000000
0!
1$
0'
1+
0/
#80560000000
1!
1'
1/
#80570000000
0!
0'
0/
#80580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#80590000000
0!
0'
0/
#80600000000
1!
1'
1/
#80610000000
0!
0'
0/
#80620000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#80630000000
0!
0'
0/
#80640000000
1!
1'
1/
#80650000000
0!
0'
0/
#80660000000
1!
1'
1/
#80670000000
0!
0'
0/
#80680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#80690000000
0!
0'
0/
#80700000000
1!
1'
1/
#80710000000
0!
0'
0/
#80720000000
1!
1'
1/
#80730000000
0!
0'
0/
#80740000000
1!
1'
1/
#80750000000
0!
0'
0/
#80760000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#80770000000
0!
0'
0/
#80780000000
1!
1'
1/
#80790000000
0!
0'
0/
#80800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#80810000000
0!
0'
0/
#80820000000
1!
1'
1/
#80830000000
0!
0'
0/
#80840000000
#80850000000
1!
1'
1/
#80860000000
0!
0'
0/
#80870000000
1!
1'
1/
#80880000000
0!
1"
0'
1(
0/
10
#80890000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#80900000000
0!
0'
0/
#80910000000
1!
1'
1/
#80920000000
0!
0'
0/
#80930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#80940000000
0!
0'
0/
#80950000000
1!
1'
1/
#80960000000
0!
1"
0'
1(
0/
10
#80970000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#80980000000
0!
1$
0'
1+
0/
#80990000000
1!
1'
1/
#81000000000
0!
0'
0/
#81010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#81020000000
0!
0'
0/
#81030000000
1!
1'
1/
#81040000000
0!
0'
0/
#81050000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#81060000000
0!
0'
0/
#81070000000
1!
1'
1/
#81080000000
0!
0'
0/
#81090000000
1!
1'
1/
#81100000000
0!
0'
0/
#81110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#81120000000
0!
0'
0/
#81130000000
1!
1'
1/
#81140000000
0!
0'
0/
#81150000000
1!
1'
1/
#81160000000
0!
0'
0/
#81170000000
1!
1'
1/
#81180000000
0!
0'
0/
#81190000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#81200000000
0!
0'
0/
#81210000000
1!
1'
1/
#81220000000
0!
0'
0/
#81230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#81240000000
0!
0'
0/
#81250000000
1!
1'
1/
#81260000000
0!
0'
0/
#81270000000
#81280000000
1!
1'
1/
#81290000000
0!
0'
0/
#81300000000
1!
1'
1/
#81310000000
0!
1"
0'
1(
0/
10
#81320000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#81330000000
0!
0'
0/
#81340000000
1!
1'
1/
#81350000000
0!
0'
0/
#81360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#81370000000
0!
0'
0/
#81380000000
1!
1'
1/
#81390000000
0!
1"
0'
1(
0/
10
#81400000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#81410000000
0!
1$
0'
1+
0/
#81420000000
1!
1'
1/
#81430000000
0!
0'
0/
#81440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#81450000000
0!
0'
0/
#81460000000
1!
1'
1/
#81470000000
0!
0'
0/
#81480000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#81490000000
0!
0'
0/
#81500000000
1!
1'
1/
#81510000000
0!
0'
0/
#81520000000
1!
1'
1/
#81530000000
0!
0'
0/
#81540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#81550000000
0!
0'
0/
#81560000000
1!
1'
1/
#81570000000
0!
0'
0/
#81580000000
1!
1'
1/
#81590000000
0!
0'
0/
#81600000000
1!
1'
1/
#81610000000
0!
0'
0/
#81620000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#81630000000
0!
0'
0/
#81640000000
1!
1'
1/
#81650000000
0!
0'
0/
#81660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#81670000000
0!
0'
0/
#81680000000
1!
1'
1/
#81690000000
0!
0'
0/
#81700000000
#81710000000
1!
1'
1/
#81720000000
0!
0'
0/
#81730000000
1!
1'
1/
#81740000000
0!
1"
0'
1(
0/
10
#81750000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#81760000000
0!
0'
0/
#81770000000
1!
1'
1/
#81780000000
0!
0'
0/
#81790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#81800000000
0!
0'
0/
#81810000000
1!
1'
1/
#81820000000
0!
1"
0'
1(
0/
10
#81830000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#81840000000
0!
1$
0'
1+
0/
#81850000000
1!
1'
1/
#81860000000
0!
0'
0/
#81870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#81880000000
0!
0'
0/
#81890000000
1!
1'
1/
#81900000000
0!
0'
0/
#81910000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#81920000000
0!
0'
0/
#81930000000
1!
1'
1/
#81940000000
0!
0'
0/
#81950000000
1!
1'
1/
#81960000000
0!
0'
0/
#81970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#81980000000
0!
0'
0/
#81990000000
1!
1'
1/
#82000000000
0!
0'
0/
#82010000000
1!
1'
1/
#82020000000
0!
0'
0/
#82030000000
1!
1'
1/
#82040000000
0!
0'
0/
#82050000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#82060000000
0!
0'
0/
#82070000000
1!
1'
1/
#82080000000
0!
0'
0/
#82090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#82100000000
0!
0'
0/
#82110000000
1!
1'
1/
#82120000000
0!
0'
0/
#82130000000
#82140000000
1!
1'
1/
#82150000000
0!
0'
0/
#82160000000
1!
1'
1/
#82170000000
0!
1"
0'
1(
0/
10
#82180000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#82190000000
0!
0'
0/
#82200000000
1!
1'
1/
#82210000000
0!
0'
0/
#82220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#82230000000
0!
0'
0/
#82240000000
1!
1'
1/
#82250000000
0!
1"
0'
1(
0/
10
#82260000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#82270000000
0!
1$
0'
1+
0/
#82280000000
1!
1'
1/
#82290000000
0!
0'
0/
#82300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#82310000000
0!
0'
0/
#82320000000
1!
1'
1/
#82330000000
0!
0'
0/
#82340000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#82350000000
0!
0'
0/
#82360000000
1!
1'
1/
#82370000000
0!
0'
0/
#82380000000
1!
1'
1/
#82390000000
0!
0'
0/
#82400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#82410000000
0!
0'
0/
#82420000000
1!
1'
1/
#82430000000
0!
0'
0/
#82440000000
1!
1'
1/
#82450000000
0!
0'
0/
#82460000000
1!
1'
1/
#82470000000
0!
0'
0/
#82480000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#82490000000
0!
0'
0/
#82500000000
1!
1'
1/
#82510000000
0!
0'
0/
#82520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#82530000000
0!
0'
0/
#82540000000
1!
1'
1/
#82550000000
0!
0'
0/
#82560000000
#82570000000
1!
1'
1/
#82580000000
0!
0'
0/
#82590000000
1!
1'
1/
#82600000000
0!
1"
0'
1(
0/
10
#82610000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#82620000000
0!
0'
0/
#82630000000
1!
1'
1/
#82640000000
0!
0'
0/
#82650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#82660000000
0!
0'
0/
#82670000000
1!
1'
1/
#82680000000
0!
1"
0'
1(
0/
10
#82690000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#82700000000
0!
1$
0'
1+
0/
#82710000000
1!
1'
1/
#82720000000
0!
0'
0/
#82730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#82740000000
0!
0'
0/
#82750000000
1!
1'
1/
#82760000000
0!
0'
0/
#82770000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#82780000000
0!
0'
0/
#82790000000
1!
1'
1/
#82800000000
0!
0'
0/
#82810000000
1!
1'
1/
#82820000000
0!
0'
0/
#82830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#82840000000
0!
0'
0/
#82850000000
1!
1'
1/
#82860000000
0!
0'
0/
#82870000000
1!
1'
1/
#82880000000
0!
0'
0/
#82890000000
1!
1'
1/
#82900000000
0!
0'
0/
#82910000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#82920000000
0!
0'
0/
#82930000000
1!
1'
1/
#82940000000
0!
0'
0/
#82950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#82960000000
0!
0'
0/
#82970000000
1!
1'
1/
#82980000000
0!
0'
0/
#82990000000
#83000000000
1!
1'
1/
#83010000000
0!
0'
0/
#83020000000
1!
1'
1/
#83030000000
0!
1"
0'
1(
0/
10
#83040000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#83050000000
0!
0'
0/
#83060000000
1!
1'
1/
#83070000000
0!
0'
0/
#83080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#83090000000
0!
0'
0/
#83100000000
1!
1'
1/
#83110000000
0!
1"
0'
1(
0/
10
#83120000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#83130000000
0!
1$
0'
1+
0/
#83140000000
1!
1'
1/
#83150000000
0!
0'
0/
#83160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#83170000000
0!
0'
0/
#83180000000
1!
1'
1/
#83190000000
0!
0'
0/
#83200000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#83210000000
0!
0'
0/
#83220000000
1!
1'
1/
#83230000000
0!
0'
0/
#83240000000
1!
1'
1/
#83250000000
0!
0'
0/
#83260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#83270000000
0!
0'
0/
#83280000000
1!
1'
1/
#83290000000
0!
0'
0/
#83300000000
1!
1'
1/
#83310000000
0!
0'
0/
#83320000000
1!
1'
1/
#83330000000
0!
0'
0/
#83340000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#83350000000
0!
0'
0/
#83360000000
1!
1'
1/
#83370000000
0!
0'
0/
#83380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#83390000000
0!
0'
0/
#83400000000
1!
1'
1/
#83410000000
0!
0'
0/
#83420000000
#83430000000
1!
1'
1/
#83440000000
0!
0'
0/
#83450000000
1!
1'
1/
#83460000000
0!
1"
0'
1(
0/
10
#83470000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#83480000000
0!
0'
0/
#83490000000
1!
1'
1/
#83500000000
0!
0'
0/
#83510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#83520000000
0!
0'
0/
#83530000000
1!
1'
1/
#83540000000
0!
1"
0'
1(
0/
10
#83550000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#83560000000
0!
1$
0'
1+
0/
#83570000000
1!
1'
1/
#83580000000
0!
0'
0/
#83590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#83600000000
0!
0'
0/
#83610000000
1!
1'
1/
#83620000000
0!
0'
0/
#83630000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#83640000000
0!
0'
0/
#83650000000
1!
1'
1/
#83660000000
0!
0'
0/
#83670000000
1!
1'
1/
#83680000000
0!
0'
0/
#83690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#83700000000
0!
0'
0/
#83710000000
1!
1'
1/
#83720000000
0!
0'
0/
#83730000000
1!
1'
1/
#83740000000
0!
0'
0/
#83750000000
1!
1'
1/
#83760000000
0!
0'
0/
#83770000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#83780000000
0!
0'
0/
#83790000000
1!
1'
1/
#83800000000
0!
0'
0/
#83810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#83820000000
0!
0'
0/
#83830000000
1!
1'
1/
#83840000000
0!
0'
0/
#83850000000
#83860000000
1!
1'
1/
#83870000000
0!
0'
0/
#83880000000
1!
1'
1/
#83890000000
0!
1"
0'
1(
0/
10
#83900000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#83910000000
0!
0'
0/
#83920000000
1!
1'
1/
#83930000000
0!
0'
0/
#83940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#83950000000
0!
0'
0/
#83960000000
1!
1'
1/
#83970000000
0!
1"
0'
1(
0/
10
#83980000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#83990000000
0!
1$
0'
1+
0/
#84000000000
1!
1'
1/
#84010000000
0!
0'
0/
#84020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#84030000000
0!
0'
0/
#84040000000
1!
1'
1/
#84050000000
0!
0'
0/
#84060000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#84070000000
0!
0'
0/
#84080000000
1!
1'
1/
#84090000000
0!
0'
0/
#84100000000
1!
1'
1/
#84110000000
0!
0'
0/
#84120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#84130000000
0!
0'
0/
#84140000000
1!
1'
1/
#84150000000
0!
0'
0/
#84160000000
1!
1'
1/
#84170000000
0!
0'
0/
#84180000000
1!
1'
1/
#84190000000
0!
0'
0/
#84200000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#84210000000
0!
0'
0/
#84220000000
1!
1'
1/
#84230000000
0!
0'
0/
#84240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#84250000000
0!
0'
0/
#84260000000
1!
1'
1/
#84270000000
0!
0'
0/
#84280000000
#84290000000
1!
1'
1/
#84300000000
0!
0'
0/
#84310000000
1!
1'
1/
#84320000000
0!
1"
0'
1(
0/
10
#84330000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#84340000000
0!
0'
0/
#84350000000
1!
1'
1/
#84360000000
0!
0'
0/
#84370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#84380000000
0!
0'
0/
#84390000000
1!
1'
1/
#84400000000
0!
1"
0'
1(
0/
10
#84410000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#84420000000
0!
1$
0'
1+
0/
#84430000000
1!
1'
1/
#84440000000
0!
0'
0/
#84450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#84460000000
0!
0'
0/
#84470000000
1!
1'
1/
#84480000000
0!
0'
0/
#84490000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#84500000000
0!
0'
0/
#84510000000
1!
1'
1/
#84520000000
0!
0'
0/
#84530000000
1!
1'
1/
#84540000000
0!
0'
0/
#84550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#84560000000
0!
0'
0/
#84570000000
1!
1'
1/
#84580000000
0!
0'
0/
#84590000000
1!
1'
1/
#84600000000
0!
0'
0/
#84610000000
1!
1'
1/
#84620000000
0!
0'
0/
#84630000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#84640000000
0!
0'
0/
#84650000000
1!
1'
1/
#84660000000
0!
0'
0/
#84670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#84680000000
0!
0'
0/
#84690000000
1!
1'
1/
#84700000000
0!
0'
0/
#84710000000
#84720000000
1!
1'
1/
#84730000000
0!
0'
0/
#84740000000
1!
1'
1/
#84750000000
0!
1"
0'
1(
0/
10
#84760000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#84770000000
0!
0'
0/
#84780000000
1!
1'
1/
#84790000000
0!
0'
0/
#84800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#84810000000
0!
0'
0/
#84820000000
1!
1'
1/
#84830000000
0!
1"
0'
1(
0/
10
#84840000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#84850000000
0!
1$
0'
1+
0/
#84860000000
1!
1'
1/
#84870000000
0!
0'
0/
#84880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#84890000000
0!
0'
0/
#84900000000
1!
1'
1/
#84910000000
0!
0'
0/
#84920000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#84930000000
0!
0'
0/
#84940000000
1!
1'
1/
#84950000000
0!
0'
0/
#84960000000
1!
1'
1/
#84970000000
0!
0'
0/
#84980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#84990000000
0!
0'
0/
#85000000000
1!
1'
1/
#85010000000
0!
0'
0/
#85020000000
1!
1'
1/
#85030000000
0!
0'
0/
#85040000000
1!
1'
1/
#85050000000
0!
0'
0/
#85060000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#85070000000
0!
0'
0/
#85080000000
1!
1'
1/
#85090000000
0!
0'
0/
#85100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#85110000000
0!
0'
0/
#85120000000
1!
1'
1/
#85130000000
0!
0'
0/
#85140000000
#85150000000
1!
1'
1/
#85160000000
0!
0'
0/
#85170000000
1!
1'
1/
#85180000000
0!
1"
0'
1(
0/
10
#85190000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#85200000000
0!
0'
0/
#85210000000
1!
1'
1/
#85220000000
0!
0'
0/
#85230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#85240000000
0!
0'
0/
#85250000000
1!
1'
1/
#85260000000
0!
1"
0'
1(
0/
10
#85270000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#85280000000
0!
1$
0'
1+
0/
#85290000000
1!
1'
1/
#85300000000
0!
0'
0/
#85310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#85320000000
0!
0'
0/
#85330000000
1!
1'
1/
#85340000000
0!
0'
0/
#85350000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#85360000000
0!
0'
0/
#85370000000
1!
1'
1/
#85380000000
0!
0'
0/
#85390000000
1!
1'
1/
#85400000000
0!
0'
0/
#85410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#85420000000
0!
0'
0/
#85430000000
1!
1'
1/
#85440000000
0!
0'
0/
#85450000000
1!
1'
1/
#85460000000
0!
0'
0/
#85470000000
1!
1'
1/
#85480000000
0!
0'
0/
#85490000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#85500000000
0!
0'
0/
#85510000000
1!
1'
1/
#85520000000
0!
0'
0/
#85530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#85540000000
0!
0'
0/
#85550000000
1!
1'
1/
#85560000000
0!
0'
0/
#85570000000
#85580000000
1!
1'
1/
#85590000000
0!
0'
0/
#85600000000
1!
1'
1/
#85610000000
0!
1"
0'
1(
0/
10
#85620000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#85630000000
0!
0'
0/
#85640000000
1!
1'
1/
#85650000000
0!
0'
0/
#85660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#85670000000
0!
0'
0/
#85680000000
1!
1'
1/
#85690000000
0!
1"
0'
1(
0/
10
#85700000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#85710000000
0!
1$
0'
1+
0/
#85720000000
1!
1'
1/
#85730000000
0!
0'
0/
#85740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#85750000000
0!
0'
0/
#85760000000
1!
1'
1/
#85770000000
0!
0'
0/
#85780000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#85790000000
0!
0'
0/
#85800000000
1!
1'
1/
#85810000000
0!
0'
0/
#85820000000
1!
1'
1/
#85830000000
0!
0'
0/
#85840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#85850000000
0!
0'
0/
#85860000000
1!
1'
1/
#85870000000
0!
0'
0/
#85880000000
1!
1'
1/
#85890000000
0!
0'
0/
#85900000000
1!
1'
1/
#85910000000
0!
0'
0/
#85920000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#85930000000
0!
0'
0/
#85940000000
1!
1'
1/
#85950000000
0!
0'
0/
#85960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#85970000000
0!
0'
0/
#85980000000
1!
1'
1/
#85990000000
0!
0'
0/
#86000000000
#86010000000
1!
1'
1/
#86020000000
0!
0'
0/
#86030000000
1!
1'
1/
#86040000000
0!
1"
0'
1(
0/
10
#86050000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#86060000000
0!
0'
0/
#86070000000
1!
1'
1/
#86080000000
0!
0'
0/
#86090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#86100000000
0!
0'
0/
#86110000000
1!
1'
1/
#86120000000
0!
1"
0'
1(
0/
10
#86130000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#86140000000
0!
1$
0'
1+
0/
#86150000000
1!
1'
1/
#86160000000
0!
0'
0/
#86170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#86180000000
0!
0'
0/
#86190000000
1!
1'
1/
#86200000000
0!
0'
0/
#86210000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#86220000000
0!
0'
0/
#86230000000
1!
1'
1/
#86240000000
0!
0'
0/
#86250000000
1!
1'
1/
#86260000000
0!
0'
0/
#86270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#86280000000
0!
0'
0/
#86290000000
1!
1'
1/
#86300000000
0!
0'
0/
#86310000000
1!
1'
1/
#86320000000
0!
0'
0/
#86330000000
1!
1'
1/
#86340000000
0!
0'
0/
#86350000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#86360000000
0!
0'
0/
#86370000000
1!
1'
1/
#86380000000
0!
0'
0/
#86390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#86400000000
0!
0'
0/
#86410000000
1!
1'
1/
#86420000000
0!
0'
0/
#86430000000
#86440000000
1!
1'
1/
#86450000000
0!
0'
0/
#86460000000
1!
1'
1/
#86470000000
0!
1"
0'
1(
0/
10
#86480000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#86490000000
0!
0'
0/
#86500000000
1!
1'
1/
#86510000000
0!
0'
0/
#86520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#86530000000
0!
0'
0/
#86540000000
1!
1'
1/
#86550000000
0!
1"
0'
1(
0/
10
#86560000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#86570000000
0!
1$
0'
1+
0/
#86580000000
1!
1'
1/
#86590000000
0!
0'
0/
#86600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#86610000000
0!
0'
0/
#86620000000
1!
1'
1/
#86630000000
0!
0'
0/
#86640000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#86650000000
0!
0'
0/
#86660000000
1!
1'
1/
#86670000000
0!
0'
0/
#86680000000
1!
1'
1/
#86690000000
0!
0'
0/
#86700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#86710000000
0!
0'
0/
#86720000000
1!
1'
1/
#86730000000
0!
0'
0/
#86740000000
1!
1'
1/
#86750000000
0!
0'
0/
#86760000000
1!
1'
1/
#86770000000
0!
0'
0/
#86780000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#86790000000
0!
0'
0/
#86800000000
1!
1'
1/
#86810000000
0!
0'
0/
#86820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#86830000000
0!
0'
0/
#86840000000
1!
1'
1/
#86850000000
0!
0'
0/
#86860000000
#86870000000
1!
1'
1/
#86880000000
0!
0'
0/
#86890000000
1!
1'
1/
#86900000000
0!
1"
0'
1(
0/
10
#86910000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#86920000000
0!
0'
0/
#86930000000
1!
1'
1/
#86940000000
0!
0'
0/
#86950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#86960000000
0!
0'
0/
#86970000000
1!
1'
1/
#86980000000
0!
1"
0'
1(
0/
10
#86990000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#87000000000
0!
1$
0'
1+
0/
#87010000000
1!
1'
1/
#87020000000
0!
0'
0/
#87030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#87040000000
0!
0'
0/
#87050000000
1!
1'
1/
#87060000000
0!
0'
0/
#87070000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#87080000000
0!
0'
0/
#87090000000
1!
1'
1/
#87100000000
0!
0'
0/
#87110000000
1!
1'
1/
#87120000000
0!
0'
0/
#87130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#87140000000
0!
0'
0/
#87150000000
1!
1'
1/
#87160000000
0!
0'
0/
#87170000000
1!
1'
1/
#87180000000
0!
0'
0/
#87190000000
1!
1'
1/
#87200000000
0!
0'
0/
#87210000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#87220000000
0!
0'
0/
#87230000000
1!
1'
1/
#87240000000
0!
0'
0/
#87250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#87260000000
0!
0'
0/
#87270000000
1!
1'
1/
#87280000000
0!
0'
0/
#87290000000
#87300000000
1!
1'
1/
#87310000000
0!
0'
0/
#87320000000
1!
1'
1/
#87330000000
0!
1"
0'
1(
0/
10
#87340000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#87350000000
0!
0'
0/
#87360000000
1!
1'
1/
#87370000000
0!
0'
0/
#87380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#87390000000
0!
0'
0/
#87400000000
1!
1'
1/
#87410000000
0!
1"
0'
1(
0/
10
#87420000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#87430000000
0!
1$
0'
1+
0/
#87440000000
1!
1'
1/
#87450000000
0!
0'
0/
#87460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#87470000000
0!
0'
0/
#87480000000
1!
1'
1/
#87490000000
0!
0'
0/
#87500000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#87510000000
0!
0'
0/
#87520000000
1!
1'
1/
#87530000000
0!
0'
0/
#87540000000
1!
1'
1/
#87550000000
0!
0'
0/
#87560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#87570000000
0!
0'
0/
#87580000000
1!
1'
1/
#87590000000
0!
0'
0/
#87600000000
1!
1'
1/
#87610000000
0!
0'
0/
#87620000000
1!
1'
1/
#87630000000
0!
0'
0/
#87640000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#87650000000
0!
0'
0/
#87660000000
1!
1'
1/
#87670000000
0!
0'
0/
#87680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#87690000000
0!
0'
0/
#87700000000
1!
1'
1/
#87710000000
0!
0'
0/
#87720000000
#87730000000
1!
1'
1/
#87740000000
0!
0'
0/
#87750000000
1!
1'
1/
#87760000000
0!
1"
0'
1(
0/
10
#87770000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#87780000000
0!
0'
0/
#87790000000
1!
1'
1/
#87800000000
0!
0'
0/
#87810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#87820000000
0!
0'
0/
#87830000000
1!
1'
1/
#87840000000
0!
1"
0'
1(
0/
10
#87850000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#87860000000
0!
1$
0'
1+
0/
#87870000000
1!
1'
1/
#87880000000
0!
0'
0/
#87890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#87900000000
0!
0'
0/
#87910000000
1!
1'
1/
#87920000000
0!
0'
0/
#87930000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#87940000000
0!
0'
0/
#87950000000
1!
1'
1/
#87960000000
0!
0'
0/
#87970000000
1!
1'
1/
#87980000000
0!
0'
0/
#87990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#88000000000
0!
0'
0/
#88010000000
1!
1'
1/
#88020000000
0!
0'
0/
#88030000000
1!
1'
1/
#88040000000
0!
0'
0/
#88050000000
1!
1'
1/
#88060000000
0!
0'
0/
#88070000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#88080000000
0!
0'
0/
#88090000000
1!
1'
1/
#88100000000
0!
0'
0/
#88110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#88120000000
0!
0'
0/
#88130000000
1!
1'
1/
#88140000000
0!
0'
0/
#88150000000
#88160000000
1!
1'
1/
#88170000000
0!
0'
0/
#88180000000
1!
1'
1/
#88190000000
0!
1"
0'
1(
0/
10
#88200000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#88210000000
0!
0'
0/
#88220000000
1!
1'
1/
#88230000000
0!
0'
0/
#88240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#88250000000
0!
0'
0/
#88260000000
1!
1'
1/
#88270000000
0!
1"
0'
1(
0/
10
#88280000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#88290000000
0!
1$
0'
1+
0/
#88300000000
1!
1'
1/
#88310000000
0!
0'
0/
#88320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#88330000000
0!
0'
0/
#88340000000
1!
1'
1/
#88350000000
0!
0'
0/
#88360000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#88370000000
0!
0'
0/
#88380000000
1!
1'
1/
#88390000000
0!
0'
0/
#88400000000
1!
1'
1/
#88410000000
0!
0'
0/
#88420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#88430000000
0!
0'
0/
#88440000000
1!
1'
1/
#88450000000
0!
0'
0/
#88460000000
1!
1'
1/
#88470000000
0!
0'
0/
#88480000000
1!
1'
1/
#88490000000
0!
0'
0/
#88500000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#88510000000
0!
0'
0/
#88520000000
1!
1'
1/
#88530000000
0!
0'
0/
#88540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#88550000000
0!
0'
0/
#88560000000
1!
1'
1/
#88570000000
0!
0'
0/
#88580000000
#88590000000
1!
1'
1/
#88600000000
0!
0'
0/
#88610000000
1!
1'
1/
#88620000000
0!
1"
0'
1(
0/
10
#88630000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#88640000000
0!
0'
0/
#88650000000
1!
1'
1/
#88660000000
0!
0'
0/
#88670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#88680000000
0!
0'
0/
#88690000000
1!
1'
1/
#88700000000
0!
1"
0'
1(
0/
10
#88710000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#88720000000
0!
1$
0'
1+
0/
#88730000000
1!
1'
1/
#88740000000
0!
0'
0/
#88750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#88760000000
0!
0'
0/
#88770000000
1!
1'
1/
#88780000000
0!
0'
0/
#88790000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#88800000000
0!
0'
0/
#88810000000
1!
1'
1/
#88820000000
0!
0'
0/
#88830000000
1!
1'
1/
#88840000000
0!
0'
0/
#88850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#88860000000
0!
0'
0/
#88870000000
1!
1'
1/
#88880000000
0!
0'
0/
#88890000000
1!
1'
1/
#88900000000
0!
0'
0/
#88910000000
1!
1'
1/
#88920000000
0!
0'
0/
#88930000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#88940000000
0!
0'
0/
#88950000000
1!
1'
1/
#88960000000
0!
0'
0/
#88970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#88980000000
0!
0'
0/
#88990000000
1!
1'
1/
#89000000000
0!
0'
0/
#89010000000
#89020000000
1!
1'
1/
#89030000000
0!
0'
0/
#89040000000
1!
1'
1/
#89050000000
0!
1"
0'
1(
0/
10
#89060000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#89070000000
0!
0'
0/
#89080000000
1!
1'
1/
#89090000000
0!
0'
0/
#89100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#89110000000
0!
0'
0/
#89120000000
1!
1'
1/
#89130000000
0!
1"
0'
1(
0/
10
#89140000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#89150000000
0!
1$
0'
1+
0/
#89160000000
1!
1'
1/
#89170000000
0!
0'
0/
#89180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#89190000000
0!
0'
0/
#89200000000
1!
1'
1/
#89210000000
0!
0'
0/
#89220000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#89230000000
0!
0'
0/
#89240000000
1!
1'
1/
#89250000000
0!
0'
0/
#89260000000
1!
1'
1/
#89270000000
0!
0'
0/
#89280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#89290000000
0!
0'
0/
#89300000000
1!
1'
1/
#89310000000
0!
0'
0/
#89320000000
1!
1'
1/
#89330000000
0!
0'
0/
#89340000000
1!
1'
1/
#89350000000
0!
0'
0/
#89360000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#89370000000
0!
0'
0/
#89380000000
1!
1'
1/
#89390000000
0!
0'
0/
#89400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#89410000000
0!
0'
0/
#89420000000
1!
1'
1/
#89430000000
0!
0'
0/
#89440000000
#89450000000
1!
1'
1/
#89460000000
0!
0'
0/
#89470000000
1!
1'
1/
#89480000000
0!
1"
0'
1(
0/
10
#89490000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#89500000000
0!
0'
0/
#89510000000
1!
1'
1/
#89520000000
0!
0'
0/
#89530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#89540000000
0!
0'
0/
#89550000000
1!
1'
1/
#89560000000
0!
1"
0'
1(
0/
10
#89570000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#89580000000
0!
1$
0'
1+
0/
#89590000000
1!
1'
1/
#89600000000
0!
0'
0/
#89610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#89620000000
0!
0'
0/
#89630000000
1!
1'
1/
#89640000000
0!
0'
0/
#89650000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#89660000000
0!
0'
0/
#89670000000
1!
1'
1/
#89680000000
0!
0'
0/
#89690000000
1!
1'
1/
#89700000000
0!
0'
0/
#89710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#89720000000
0!
0'
0/
#89730000000
1!
1'
1/
#89740000000
0!
0'
0/
#89750000000
1!
1'
1/
#89760000000
0!
0'
0/
#89770000000
1!
1'
1/
#89780000000
0!
0'
0/
#89790000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#89800000000
0!
0'
0/
#89810000000
1!
1'
1/
#89820000000
0!
0'
0/
#89830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#89840000000
0!
0'
0/
#89850000000
1!
1'
1/
#89860000000
0!
0'
0/
#89870000000
#89880000000
1!
1'
1/
#89890000000
0!
0'
0/
#89900000000
1!
1'
1/
#89910000000
0!
1"
0'
1(
0/
10
#89920000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#89930000000
0!
0'
0/
#89940000000
1!
1'
1/
#89950000000
0!
0'
0/
#89960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#89970000000
0!
0'
0/
#89980000000
1!
1'
1/
#89990000000
0!
1"
0'
1(
0/
10
#90000000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#90010000000
0!
1$
0'
1+
0/
#90020000000
1!
1'
1/
#90030000000
0!
0'
0/
#90040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#90050000000
0!
0'
0/
#90060000000
1!
1'
1/
#90070000000
0!
0'
0/
#90080000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#90090000000
0!
0'
0/
#90100000000
1!
1'
1/
#90110000000
0!
0'
0/
#90120000000
1!
1'
1/
#90130000000
0!
0'
0/
#90140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#90150000000
0!
0'
0/
#90160000000
1!
1'
1/
#90170000000
0!
0'
0/
#90180000000
1!
1'
1/
#90190000000
0!
0'
0/
#90200000000
1!
1'
1/
#90210000000
0!
0'
0/
#90220000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#90230000000
0!
0'
0/
#90240000000
1!
1'
1/
#90250000000
0!
0'
0/
#90260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#90270000000
0!
0'
0/
#90280000000
1!
1'
1/
#90290000000
0!
0'
0/
#90300000000
#90310000000
1!
1'
1/
#90320000000
0!
0'
0/
#90330000000
1!
1'
1/
#90340000000
0!
1"
0'
1(
0/
10
#90350000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#90360000000
0!
0'
0/
#90370000000
1!
1'
1/
#90380000000
0!
0'
0/
#90390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#90400000000
0!
0'
0/
#90410000000
1!
1'
1/
#90420000000
0!
1"
0'
1(
0/
10
#90430000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#90440000000
0!
1$
0'
1+
0/
#90450000000
1!
1'
1/
#90460000000
0!
0'
0/
#90470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#90480000000
0!
0'
0/
#90490000000
1!
1'
1/
#90500000000
0!
0'
0/
#90510000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#90520000000
0!
0'
0/
#90530000000
1!
1'
1/
#90540000000
0!
0'
0/
#90550000000
1!
1'
1/
#90560000000
0!
0'
0/
#90570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#90580000000
0!
0'
0/
#90590000000
1!
1'
1/
#90600000000
0!
0'
0/
#90610000000
1!
1'
1/
#90620000000
0!
0'
0/
#90630000000
1!
1'
1/
#90640000000
0!
0'
0/
#90650000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#90660000000
0!
0'
0/
#90670000000
1!
1'
1/
#90680000000
0!
0'
0/
#90690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#90700000000
0!
0'
0/
#90710000000
1!
1'
1/
#90720000000
0!
0'
0/
#90730000000
#90740000000
1!
1'
1/
#90750000000
0!
0'
0/
#90760000000
1!
1'
1/
#90770000000
0!
1"
0'
1(
0/
10
#90780000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#90790000000
0!
0'
0/
#90800000000
1!
1'
1/
#90810000000
0!
0'
0/
#90820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#90830000000
0!
0'
0/
#90840000000
1!
1'
1/
#90850000000
0!
1"
0'
1(
0/
10
#90860000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#90870000000
0!
1$
0'
1+
0/
#90880000000
1!
1'
1/
#90890000000
0!
0'
0/
#90900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#90910000000
0!
0'
0/
#90920000000
1!
1'
1/
#90930000000
0!
0'
0/
#90940000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#90950000000
0!
0'
0/
#90960000000
1!
1'
1/
#90970000000
0!
0'
0/
#90980000000
1!
1'
1/
#90990000000
0!
0'
0/
#91000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#91010000000
0!
0'
0/
#91020000000
1!
1'
1/
#91030000000
0!
0'
0/
#91040000000
1!
1'
1/
#91050000000
0!
0'
0/
#91060000000
1!
1'
1/
#91070000000
0!
0'
0/
#91080000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#91090000000
0!
0'
0/
#91100000000
1!
1'
1/
#91110000000
0!
0'
0/
#91120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#91130000000
0!
0'
0/
#91140000000
1!
1'
1/
#91150000000
0!
0'
0/
#91160000000
#91170000000
1!
1'
1/
#91180000000
0!
0'
0/
#91190000000
1!
1'
1/
#91200000000
0!
1"
0'
1(
0/
10
#91210000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#91220000000
0!
0'
0/
#91230000000
1!
1'
1/
#91240000000
0!
0'
0/
#91250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#91260000000
0!
0'
0/
#91270000000
1!
1'
1/
#91280000000
0!
1"
0'
1(
0/
10
#91290000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#91300000000
0!
1$
0'
1+
0/
#91310000000
1!
1'
1/
#91320000000
0!
0'
0/
#91330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#91340000000
0!
0'
0/
#91350000000
1!
1'
1/
#91360000000
0!
0'
0/
#91370000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#91380000000
0!
0'
0/
#91390000000
1!
1'
1/
#91400000000
0!
0'
0/
#91410000000
1!
1'
1/
#91420000000
0!
0'
0/
#91430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#91440000000
0!
0'
0/
#91450000000
1!
1'
1/
#91460000000
0!
0'
0/
#91470000000
1!
1'
1/
#91480000000
0!
0'
0/
#91490000000
1!
1'
1/
#91500000000
0!
0'
0/
#91510000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#91520000000
0!
0'
0/
#91530000000
1!
1'
1/
#91540000000
0!
0'
0/
#91550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#91560000000
0!
0'
0/
#91570000000
1!
1'
1/
#91580000000
0!
0'
0/
#91590000000
#91600000000
1!
1'
1/
#91610000000
0!
0'
0/
#91620000000
1!
1'
1/
#91630000000
0!
1"
0'
1(
0/
10
#91640000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#91650000000
0!
0'
0/
#91660000000
1!
1'
1/
#91670000000
0!
0'
0/
#91680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#91690000000
0!
0'
0/
#91700000000
1!
1'
1/
#91710000000
0!
1"
0'
1(
0/
10
#91720000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#91730000000
0!
1$
0'
1+
0/
#91740000000
1!
1'
1/
#91750000000
0!
0'
0/
#91760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#91770000000
0!
0'
0/
#91780000000
1!
1'
1/
#91790000000
0!
0'
0/
#91800000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#91810000000
0!
0'
0/
#91820000000
1!
1'
1/
#91830000000
0!
0'
0/
#91840000000
1!
1'
1/
#91850000000
0!
0'
0/
#91860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#91870000000
0!
0'
0/
#91880000000
1!
1'
1/
#91890000000
0!
0'
0/
#91900000000
1!
1'
1/
#91910000000
0!
0'
0/
#91920000000
1!
1'
1/
#91930000000
0!
0'
0/
#91940000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#91950000000
0!
0'
0/
#91960000000
1!
1'
1/
#91970000000
0!
0'
0/
#91980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#91990000000
0!
0'
0/
#92000000000
1!
1'
1/
#92010000000
0!
0'
0/
#92020000000
#92030000000
1!
1'
1/
#92040000000
0!
0'
0/
#92050000000
1!
1'
1/
#92060000000
0!
1"
0'
1(
0/
10
#92070000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#92080000000
0!
0'
0/
#92090000000
1!
1'
1/
#92100000000
0!
0'
0/
#92110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#92120000000
0!
0'
0/
#92130000000
1!
1'
1/
#92140000000
0!
1"
0'
1(
0/
10
#92150000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#92160000000
0!
1$
0'
1+
0/
#92170000000
1!
1'
1/
#92180000000
0!
0'
0/
#92190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#92200000000
0!
0'
0/
#92210000000
1!
1'
1/
#92220000000
0!
0'
0/
#92230000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#92240000000
0!
0'
0/
#92250000000
1!
1'
1/
#92260000000
0!
0'
0/
#92270000000
1!
1'
1/
#92280000000
0!
0'
0/
#92290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#92300000000
0!
0'
0/
#92310000000
1!
1'
1/
#92320000000
0!
0'
0/
#92330000000
1!
1'
1/
#92340000000
0!
0'
0/
#92350000000
1!
1'
1/
#92360000000
0!
0'
0/
#92370000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#92380000000
0!
0'
0/
#92390000000
1!
1'
1/
#92400000000
0!
0'
0/
#92410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#92420000000
0!
0'
0/
#92430000000
1!
1'
1/
#92440000000
0!
0'
0/
#92450000000
#92460000000
1!
1'
1/
#92470000000
0!
0'
0/
#92480000000
1!
1'
1/
#92490000000
0!
1"
0'
1(
0/
10
#92500000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#92510000000
0!
0'
0/
#92520000000
1!
1'
1/
#92530000000
0!
0'
0/
#92540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#92550000000
0!
0'
0/
#92560000000
1!
1'
1/
#92570000000
0!
1"
0'
1(
0/
10
#92580000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#92590000000
0!
1$
0'
1+
0/
#92600000000
1!
1'
1/
#92610000000
0!
0'
0/
#92620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#92630000000
0!
0'
0/
#92640000000
1!
1'
1/
#92650000000
0!
0'
0/
#92660000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#92670000000
0!
0'
0/
#92680000000
1!
1'
1/
#92690000000
0!
0'
0/
#92700000000
1!
1'
1/
#92710000000
0!
0'
0/
#92720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#92730000000
0!
0'
0/
#92740000000
1!
1'
1/
#92750000000
0!
0'
0/
#92760000000
1!
1'
1/
#92770000000
0!
0'
0/
#92780000000
1!
1'
1/
#92790000000
0!
0'
0/
#92800000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#92810000000
0!
0'
0/
#92820000000
1!
1'
1/
#92830000000
0!
0'
0/
#92840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#92850000000
0!
0'
0/
#92860000000
1!
1'
1/
#92870000000
0!
0'
0/
#92880000000
#92890000000
1!
1'
1/
#92900000000
0!
0'
0/
#92910000000
1!
1'
1/
#92920000000
0!
1"
0'
1(
0/
10
#92930000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#92940000000
0!
0'
0/
#92950000000
1!
1'
1/
#92960000000
0!
0'
0/
#92970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#92980000000
0!
0'
0/
#92990000000
1!
1'
1/
#93000000000
0!
1"
0'
1(
0/
10
#93010000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#93020000000
0!
1$
0'
1+
0/
#93030000000
1!
1'
1/
#93040000000
0!
0'
0/
#93050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#93060000000
0!
0'
0/
#93070000000
1!
1'
1/
#93080000000
0!
0'
0/
#93090000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#93100000000
0!
0'
0/
#93110000000
1!
1'
1/
#93120000000
0!
0'
0/
#93130000000
1!
1'
1/
#93140000000
0!
0'
0/
#93150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#93160000000
0!
0'
0/
#93170000000
1!
1'
1/
#93180000000
0!
0'
0/
#93190000000
1!
1'
1/
#93200000000
0!
0'
0/
#93210000000
1!
1'
1/
#93220000000
0!
0'
0/
#93230000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#93240000000
0!
0'
0/
#93250000000
1!
1'
1/
#93260000000
0!
0'
0/
#93270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#93280000000
0!
0'
0/
#93290000000
1!
1'
1/
#93300000000
0!
0'
0/
#93310000000
#93320000000
1!
1'
1/
#93330000000
0!
0'
0/
#93340000000
1!
1'
1/
#93350000000
0!
1"
0'
1(
0/
10
#93360000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#93370000000
0!
0'
0/
#93380000000
1!
1'
1/
#93390000000
0!
0'
0/
#93400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#93410000000
0!
0'
0/
#93420000000
1!
1'
1/
#93430000000
0!
1"
0'
1(
0/
10
#93440000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#93450000000
0!
1$
0'
1+
0/
#93460000000
1!
1'
1/
#93470000000
0!
0'
0/
#93480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#93490000000
0!
0'
0/
#93500000000
1!
1'
1/
#93510000000
0!
0'
0/
#93520000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#93530000000
0!
0'
0/
#93540000000
1!
1'
1/
#93550000000
0!
0'
0/
#93560000000
1!
1'
1/
#93570000000
0!
0'
0/
#93580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#93590000000
0!
0'
0/
#93600000000
1!
1'
1/
#93610000000
0!
0'
0/
#93620000000
1!
1'
1/
#93630000000
0!
0'
0/
#93640000000
1!
1'
1/
#93650000000
0!
0'
0/
#93660000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#93670000000
0!
0'
0/
#93680000000
1!
1'
1/
#93690000000
0!
0'
0/
#93700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#93710000000
0!
0'
0/
#93720000000
1!
1'
1/
#93730000000
0!
0'
0/
#93740000000
#93750000000
1!
1'
1/
#93760000000
0!
0'
0/
#93770000000
1!
1'
1/
#93780000000
0!
1"
0'
1(
0/
10
#93790000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#93800000000
0!
0'
0/
#93810000000
1!
1'
1/
#93820000000
0!
0'
0/
#93830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#93840000000
0!
0'
0/
#93850000000
1!
1'
1/
#93860000000
0!
1"
0'
1(
0/
10
#93870000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#93880000000
0!
1$
0'
1+
0/
#93890000000
1!
1'
1/
#93900000000
0!
0'
0/
#93910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#93920000000
0!
0'
0/
#93930000000
1!
1'
1/
#93940000000
0!
0'
0/
#93950000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#93960000000
0!
0'
0/
#93970000000
1!
1'
1/
#93980000000
0!
0'
0/
#93990000000
1!
1'
1/
#94000000000
0!
0'
0/
#94010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#94020000000
0!
0'
0/
#94030000000
1!
1'
1/
#94040000000
0!
0'
0/
#94050000000
1!
1'
1/
#94060000000
0!
0'
0/
#94070000000
1!
1'
1/
#94080000000
0!
0'
0/
#94090000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#94100000000
0!
0'
0/
#94110000000
1!
1'
1/
#94120000000
0!
0'
0/
#94130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#94140000000
0!
0'
0/
#94150000000
1!
1'
1/
#94160000000
0!
0'
0/
#94170000000
#94180000000
1!
1'
1/
#94190000000
0!
0'
0/
#94200000000
1!
1'
1/
#94210000000
0!
1"
0'
1(
0/
10
#94220000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#94230000000
0!
0'
0/
#94240000000
1!
1'
1/
#94250000000
0!
0'
0/
#94260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#94270000000
0!
0'
0/
#94280000000
1!
1'
1/
#94290000000
0!
1"
0'
1(
0/
10
#94300000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#94310000000
0!
1$
0'
1+
0/
#94320000000
1!
1'
1/
#94330000000
0!
0'
0/
#94340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#94350000000
0!
0'
0/
#94360000000
1!
1'
1/
#94370000000
0!
0'
0/
#94380000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#94390000000
0!
0'
0/
#94400000000
1!
1'
1/
#94410000000
0!
0'
0/
#94420000000
1!
1'
1/
#94430000000
0!
0'
0/
#94440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#94450000000
0!
0'
0/
#94460000000
1!
1'
1/
#94470000000
0!
0'
0/
#94480000000
1!
1'
1/
#94490000000
0!
0'
0/
#94500000000
1!
1'
1/
#94510000000
0!
0'
0/
#94520000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#94530000000
0!
0'
0/
#94540000000
1!
1'
1/
#94550000000
0!
0'
0/
#94560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#94570000000
0!
0'
0/
#94580000000
1!
1'
1/
#94590000000
0!
0'
0/
#94600000000
#94610000000
1!
1'
1/
#94620000000
0!
0'
0/
#94630000000
1!
1'
1/
#94640000000
0!
1"
0'
1(
0/
10
#94650000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#94660000000
0!
0'
0/
#94670000000
1!
1'
1/
#94680000000
0!
0'
0/
#94690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#94700000000
0!
0'
0/
#94710000000
1!
1'
1/
#94720000000
0!
1"
0'
1(
0/
10
#94730000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#94740000000
0!
1$
0'
1+
0/
#94750000000
1!
1'
1/
#94760000000
0!
0'
0/
#94770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#94780000000
0!
0'
0/
#94790000000
1!
1'
1/
#94800000000
0!
0'
0/
#94810000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#94820000000
0!
0'
0/
#94830000000
1!
1'
1/
#94840000000
0!
0'
0/
#94850000000
1!
1'
1/
#94860000000
0!
0'
0/
#94870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#94880000000
0!
0'
0/
#94890000000
1!
1'
1/
#94900000000
0!
0'
0/
#94910000000
1!
1'
1/
#94920000000
0!
0'
0/
#94930000000
1!
1'
1/
#94940000000
0!
0'
0/
#94950000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#94960000000
0!
0'
0/
#94970000000
1!
1'
1/
#94980000000
0!
0'
0/
#94990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#95000000000
0!
0'
0/
#95010000000
1!
1'
1/
#95020000000
0!
0'
0/
#95030000000
#95040000000
1!
1'
1/
#95050000000
0!
0'
0/
#95060000000
1!
1'
1/
#95070000000
0!
1"
0'
1(
0/
10
#95080000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#95090000000
0!
0'
0/
#95100000000
1!
1'
1/
#95110000000
0!
0'
0/
#95120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#95130000000
0!
0'
0/
#95140000000
1!
1'
1/
#95150000000
0!
1"
0'
1(
0/
10
#95160000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#95170000000
0!
1$
0'
1+
0/
#95180000000
1!
1'
1/
#95190000000
0!
0'
0/
#95200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#95210000000
0!
0'
0/
#95220000000
1!
1'
1/
#95230000000
0!
0'
0/
#95240000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#95250000000
0!
0'
0/
#95260000000
1!
1'
1/
#95270000000
0!
0'
0/
#95280000000
1!
1'
1/
#95290000000
0!
0'
0/
#95300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#95310000000
0!
0'
0/
#95320000000
1!
1'
1/
#95330000000
0!
0'
0/
#95340000000
1!
1'
1/
#95350000000
0!
0'
0/
#95360000000
1!
1'
1/
#95370000000
0!
0'
0/
#95380000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#95390000000
0!
0'
0/
#95400000000
1!
1'
1/
#95410000000
0!
0'
0/
#95420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#95430000000
0!
0'
0/
#95440000000
1!
1'
1/
#95450000000
0!
0'
0/
#95460000000
#95470000000
1!
1'
1/
#95480000000
0!
0'
0/
#95490000000
1!
1'
1/
#95500000000
0!
1"
0'
1(
0/
10
#95510000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#95520000000
0!
0'
0/
#95530000000
1!
1'
1/
#95540000000
0!
0'
0/
#95550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#95560000000
0!
0'
0/
#95570000000
1!
1'
1/
#95580000000
0!
1"
0'
1(
0/
10
#95590000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#95600000000
0!
1$
0'
1+
0/
#95610000000
1!
1'
1/
#95620000000
0!
0'
0/
#95630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#95640000000
0!
0'
0/
#95650000000
1!
1'
1/
#95660000000
0!
0'
0/
#95670000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#95680000000
0!
0'
0/
#95690000000
1!
1'
1/
#95700000000
0!
0'
0/
#95710000000
1!
1'
1/
#95720000000
0!
0'
0/
#95730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#95740000000
0!
0'
0/
#95750000000
1!
1'
1/
#95760000000
0!
0'
0/
#95770000000
1!
1'
1/
#95780000000
0!
0'
0/
#95790000000
1!
1'
1/
#95800000000
0!
0'
0/
#95810000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#95820000000
0!
0'
0/
#95830000000
1!
1'
1/
#95840000000
0!
0'
0/
#95850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#95860000000
0!
0'
0/
#95870000000
1!
1'
1/
#95880000000
0!
0'
0/
#95890000000
#95900000000
1!
1'
1/
#95910000000
0!
0'
0/
#95920000000
1!
1'
1/
#95930000000
0!
1"
0'
1(
0/
10
#95940000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#95950000000
0!
0'
0/
#95960000000
1!
1'
1/
#95970000000
0!
0'
0/
#95980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#95990000000
0!
0'
0/
#96000000000
1!
1'
1/
#96010000000
0!
1"
0'
1(
0/
10
#96020000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#96030000000
0!
1$
0'
1+
0/
#96040000000
1!
1'
1/
#96050000000
0!
0'
0/
#96060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#96070000000
0!
0'
0/
#96080000000
1!
1'
1/
#96090000000
0!
0'
0/
#96100000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#96110000000
0!
0'
0/
#96120000000
1!
1'
1/
#96130000000
0!
0'
0/
#96140000000
1!
1'
1/
#96150000000
0!
0'
0/
#96160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#96170000000
0!
0'
0/
#96180000000
1!
1'
1/
#96190000000
0!
0'
0/
#96200000000
1!
1'
1/
#96210000000
0!
0'
0/
#96220000000
1!
1'
1/
#96230000000
0!
0'
0/
#96240000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#96250000000
0!
0'
0/
#96260000000
1!
1'
1/
#96270000000
0!
0'
0/
#96280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#96290000000
0!
0'
0/
#96300000000
1!
1'
1/
#96310000000
0!
0'
0/
#96320000000
#96330000000
1!
1'
1/
#96340000000
0!
0'
0/
#96350000000
1!
1'
1/
#96360000000
0!
1"
0'
1(
0/
10
#96370000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#96380000000
0!
0'
0/
#96390000000
1!
1'
1/
#96400000000
0!
0'
0/
#96410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#96420000000
0!
0'
0/
#96430000000
1!
1'
1/
#96440000000
0!
1"
0'
1(
0/
10
#96450000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#96460000000
0!
1$
0'
1+
0/
#96470000000
1!
1'
1/
#96480000000
0!
0'
0/
#96490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#96500000000
0!
0'
0/
#96510000000
1!
1'
1/
#96520000000
0!
0'
0/
#96530000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#96540000000
0!
0'
0/
#96550000000
1!
1'
1/
#96560000000
0!
0'
0/
#96570000000
1!
1'
1/
#96580000000
0!
0'
0/
#96590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#96600000000
0!
0'
0/
#96610000000
1!
1'
1/
#96620000000
0!
0'
0/
#96630000000
1!
1'
1/
#96640000000
0!
0'
0/
#96650000000
1!
1'
1/
#96660000000
0!
0'
0/
#96670000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#96680000000
0!
0'
0/
#96690000000
1!
1'
1/
#96700000000
0!
0'
0/
#96710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#96720000000
0!
0'
0/
#96730000000
1!
1'
1/
#96740000000
0!
0'
0/
#96750000000
#96760000000
1!
1'
1/
#96770000000
0!
0'
0/
#96780000000
1!
1'
1/
#96790000000
0!
1"
0'
1(
0/
10
#96800000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#96810000000
0!
0'
0/
#96820000000
1!
1'
1/
#96830000000
0!
0'
0/
#96840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#96850000000
0!
0'
0/
#96860000000
1!
1'
1/
#96870000000
0!
1"
0'
1(
0/
10
#96880000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#96890000000
0!
1$
0'
1+
0/
#96900000000
1!
1'
1/
#96910000000
0!
0'
0/
#96920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#96930000000
0!
0'
0/
#96940000000
1!
1'
1/
#96950000000
0!
0'
0/
#96960000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#96970000000
0!
0'
0/
#96980000000
1!
1'
1/
#96990000000
0!
0'
0/
#97000000000
1!
1'
1/
#97010000000
0!
0'
0/
#97020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#97030000000
0!
0'
0/
#97040000000
1!
1'
1/
#97050000000
0!
0'
0/
#97060000000
1!
1'
1/
#97070000000
0!
0'
0/
#97080000000
1!
1'
1/
#97090000000
0!
0'
0/
#97100000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#97110000000
0!
0'
0/
#97120000000
1!
1'
1/
#97130000000
0!
0'
0/
#97140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#97150000000
0!
0'
0/
#97160000000
1!
1'
1/
#97170000000
0!
0'
0/
#97180000000
#97190000000
1!
1'
1/
#97200000000
0!
0'
0/
#97210000000
1!
1'
1/
#97220000000
0!
1"
0'
1(
0/
10
#97230000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#97240000000
0!
0'
0/
#97250000000
1!
1'
1/
#97260000000
0!
0'
0/
#97270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#97280000000
0!
0'
0/
#97290000000
1!
1'
1/
#97300000000
0!
1"
0'
1(
0/
10
#97310000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#97320000000
0!
1$
0'
1+
0/
#97330000000
1!
1'
1/
#97340000000
0!
0'
0/
#97350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#97360000000
0!
0'
0/
#97370000000
1!
1'
1/
#97380000000
0!
0'
0/
#97390000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#97400000000
0!
0'
0/
#97410000000
1!
1'
1/
#97420000000
0!
0'
0/
#97430000000
1!
1'
1/
#97440000000
0!
0'
0/
#97450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#97460000000
0!
0'
0/
#97470000000
1!
1'
1/
#97480000000
0!
0'
0/
#97490000000
1!
1'
1/
#97500000000
0!
0'
0/
#97510000000
1!
1'
1/
#97520000000
0!
0'
0/
#97530000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#97540000000
0!
0'
0/
#97550000000
1!
1'
1/
#97560000000
0!
0'
0/
#97570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#97580000000
0!
0'
0/
#97590000000
1!
1'
1/
#97600000000
0!
0'
0/
#97610000000
#97620000000
1!
1'
1/
#97630000000
0!
0'
0/
#97640000000
1!
1'
1/
#97650000000
0!
1"
0'
1(
0/
10
#97660000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#97670000000
0!
0'
0/
#97680000000
1!
1'
1/
#97690000000
0!
0'
0/
#97700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#97710000000
0!
0'
0/
#97720000000
1!
1'
1/
#97730000000
0!
1"
0'
1(
0/
10
#97740000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#97750000000
0!
1$
0'
1+
0/
#97760000000
1!
1'
1/
#97770000000
0!
0'
0/
#97780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#97790000000
0!
0'
0/
#97800000000
1!
1'
1/
#97810000000
0!
0'
0/
#97820000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#97830000000
0!
0'
0/
#97840000000
1!
1'
1/
#97850000000
0!
0'
0/
#97860000000
1!
1'
1/
#97870000000
0!
0'
0/
#97880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#97890000000
0!
0'
0/
#97900000000
1!
1'
1/
#97910000000
0!
0'
0/
#97920000000
1!
1'
1/
#97930000000
0!
0'
0/
#97940000000
1!
1'
1/
#97950000000
0!
0'
0/
#97960000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#97970000000
0!
0'
0/
#97980000000
1!
1'
1/
#97990000000
0!
0'
0/
#98000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#98010000000
0!
0'
0/
#98020000000
1!
1'
1/
#98030000000
0!
0'
0/
#98040000000
#98050000000
1!
1'
1/
#98060000000
0!
0'
0/
#98070000000
1!
1'
1/
#98080000000
0!
1"
0'
1(
0/
10
#98090000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#98100000000
0!
0'
0/
#98110000000
1!
1'
1/
#98120000000
0!
0'
0/
#98130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#98140000000
0!
0'
0/
#98150000000
1!
1'
1/
#98160000000
0!
1"
0'
1(
0/
10
#98170000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#98180000000
0!
1$
0'
1+
0/
#98190000000
1!
1'
1/
#98200000000
0!
0'
0/
#98210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#98220000000
0!
0'
0/
#98230000000
1!
1'
1/
#98240000000
0!
0'
0/
#98250000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#98260000000
0!
0'
0/
#98270000000
1!
1'
1/
#98280000000
0!
0'
0/
#98290000000
1!
1'
1/
#98300000000
0!
0'
0/
#98310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#98320000000
0!
0'
0/
#98330000000
1!
1'
1/
#98340000000
0!
0'
0/
#98350000000
1!
1'
1/
#98360000000
0!
0'
0/
#98370000000
1!
1'
1/
#98380000000
0!
0'
0/
#98390000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#98400000000
0!
0'
0/
#98410000000
1!
1'
1/
#98420000000
0!
0'
0/
#98430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#98440000000
0!
0'
0/
#98450000000
1!
1'
1/
#98460000000
0!
0'
0/
#98470000000
#98480000000
1!
1'
1/
#98490000000
0!
0'
0/
#98500000000
1!
1'
1/
#98510000000
0!
1"
0'
1(
0/
10
#98520000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#98530000000
0!
0'
0/
#98540000000
1!
1'
1/
#98550000000
0!
0'
0/
#98560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#98570000000
0!
0'
0/
#98580000000
1!
1'
1/
#98590000000
0!
1"
0'
1(
0/
10
#98600000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#98610000000
0!
1$
0'
1+
0/
#98620000000
1!
1'
1/
#98630000000
0!
0'
0/
#98640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#98650000000
0!
0'
0/
#98660000000
1!
1'
1/
#98670000000
0!
0'
0/
#98680000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#98690000000
0!
0'
0/
#98700000000
1!
1'
1/
#98710000000
0!
0'
0/
#98720000000
1!
1'
1/
#98730000000
0!
0'
0/
#98740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#98750000000
0!
0'
0/
#98760000000
1!
1'
1/
#98770000000
0!
0'
0/
#98780000000
1!
1'
1/
#98790000000
0!
0'
0/
#98800000000
1!
1'
1/
#98810000000
0!
0'
0/
#98820000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#98830000000
0!
0'
0/
#98840000000
1!
1'
1/
#98850000000
0!
0'
0/
#98860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#98870000000
0!
0'
0/
#98880000000
1!
1'
1/
#98890000000
0!
0'
0/
#98900000000
#98910000000
1!
1'
1/
#98920000000
0!
0'
0/
#98930000000
1!
1'
1/
#98940000000
0!
1"
0'
1(
0/
10
#98950000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#98960000000
0!
0'
0/
#98970000000
1!
1'
1/
#98980000000
0!
0'
0/
#98990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#99000000000
0!
0'
0/
#99010000000
1!
1'
1/
#99020000000
0!
1"
0'
1(
0/
10
#99030000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#99040000000
0!
1$
0'
1+
0/
#99050000000
1!
1'
1/
#99060000000
0!
0'
0/
#99070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#99080000000
0!
0'
0/
#99090000000
1!
1'
1/
#99100000000
0!
0'
0/
#99110000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#99120000000
0!
0'
0/
#99130000000
1!
1'
1/
#99140000000
0!
0'
0/
#99150000000
1!
1'
1/
#99160000000
0!
0'
0/
#99170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#99180000000
0!
0'
0/
#99190000000
1!
1'
1/
#99200000000
0!
0'
0/
#99210000000
1!
1'
1/
#99220000000
0!
0'
0/
#99230000000
1!
1'
1/
#99240000000
0!
0'
0/
#99250000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#99260000000
0!
0'
0/
#99270000000
1!
1'
1/
#99280000000
0!
0'
0/
#99290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#99300000000
0!
0'
0/
#99310000000
1!
1'
1/
#99320000000
0!
0'
0/
#99330000000
#99340000000
1!
1'
1/
#99350000000
0!
0'
0/
#99360000000
1!
1'
1/
#99370000000
0!
1"
0'
1(
0/
10
#99380000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#99390000000
0!
0'
0/
#99400000000
1!
1'
1/
#99410000000
0!
0'
0/
#99420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#99430000000
0!
0'
0/
#99440000000
1!
1'
1/
#99450000000
0!
1"
0'
1(
0/
10
#99460000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#99470000000
0!
1$
0'
1+
0/
#99480000000
1!
1'
1/
#99490000000
0!
0'
0/
#99500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#99510000000
0!
0'
0/
#99520000000
1!
1'
1/
#99530000000
0!
0'
0/
#99540000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#99550000000
0!
0'
0/
#99560000000
1!
1'
1/
#99570000000
0!
0'
0/
#99580000000
1!
1'
1/
#99590000000
0!
0'
0/
#99600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#99610000000
0!
0'
0/
#99620000000
1!
1'
1/
#99630000000
0!
0'
0/
#99640000000
1!
1'
1/
#99650000000
0!
0'
0/
#99660000000
1!
1'
1/
#99670000000
0!
0'
0/
#99680000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#99690000000
0!
0'
0/
#99700000000
1!
1'
1/
#99710000000
0!
0'
0/
#99720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#99730000000
0!
0'
0/
#99740000000
1!
1'
1/
#99750000000
0!
0'
0/
#99760000000
#99770000000
1!
1'
1/
#99780000000
0!
0'
0/
#99790000000
1!
1'
1/
#99800000000
0!
1"
0'
1(
0/
10
#99810000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#99820000000
0!
0'
0/
#99830000000
1!
1'
1/
#99840000000
0!
0'
0/
#99850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#99860000000
0!
0'
0/
#99870000000
1!
1'
1/
#99880000000
0!
1"
0'
1(
0/
10
#99890000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#99900000000
0!
1$
0'
1+
0/
#99910000000
1!
1'
1/
#99920000000
0!
0'
0/
#99930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#99940000000
0!
0'
0/
#99950000000
1!
1'
1/
#99960000000
0!
0'
0/
#99970000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#99980000000
0!
0'
0/
#99990000000
1!
1'
1/
#100000000000
0!
0'
0/
#100010000000
1!
1'
1/
#100020000000
0!
0'
0/
#100030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#100040000000
0!
0'
0/
#100050000000
1!
1'
1/
#100060000000
0!
0'
0/
#100070000000
1!
1'
1/
#100080000000
0!
0'
0/
#100090000000
1!
1'
1/
#100100000000
0!
0'
0/
#100110000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#100120000000
0!
0'
0/
#100130000000
1!
1'
1/
#100140000000
0!
0'
0/
#100150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#100160000000
0!
0'
0/
#100170000000
1!
1'
1/
#100180000000
0!
0'
0/
#100190000000
#100200000000
1!
1'
1/
#100210000000
0!
0'
0/
#100220000000
1!
1'
1/
#100230000000
0!
1"
0'
1(
0/
10
#100240000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#100250000000
0!
0'
0/
#100260000000
1!
1'
1/
#100270000000
0!
0'
0/
#100280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#100290000000
0!
0'
0/
#100300000000
1!
1'
1/
#100310000000
0!
1"
0'
1(
0/
10
#100320000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#100330000000
0!
1$
0'
1+
0/
#100340000000
1!
1'
1/
#100350000000
0!
0'
0/
#100360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#100370000000
0!
0'
0/
#100380000000
1!
1'
1/
#100390000000
0!
0'
0/
#100400000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#100410000000
0!
0'
0/
#100420000000
1!
1'
1/
#100430000000
0!
0'
0/
#100440000000
1!
1'
1/
#100450000000
0!
0'
0/
#100460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#100470000000
0!
0'
0/
#100480000000
1!
1'
1/
#100490000000
0!
0'
0/
#100500000000
1!
1'
1/
#100510000000
0!
0'
0/
#100520000000
1!
1'
1/
#100530000000
0!
0'
0/
#100540000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#100550000000
0!
0'
0/
#100560000000
1!
1'
1/
#100570000000
0!
0'
0/
#100580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#100590000000
0!
0'
0/
#100600000000
1!
1'
1/
#100610000000
0!
0'
0/
#100620000000
#100630000000
1!
1'
1/
#100640000000
0!
0'
0/
#100650000000
1!
1'
1/
#100660000000
0!
1"
0'
1(
0/
10
#100670000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#100680000000
0!
0'
0/
#100690000000
1!
1'
1/
#100700000000
0!
0'
0/
#100710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#100720000000
0!
0'
0/
#100730000000
1!
1'
1/
#100740000000
0!
1"
0'
1(
0/
10
#100750000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#100760000000
0!
1$
0'
1+
0/
#100770000000
1!
1'
1/
#100780000000
0!
0'
0/
#100790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#100800000000
0!
0'
0/
#100810000000
1!
1'
1/
#100820000000
0!
0'
0/
#100830000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#100840000000
0!
0'
0/
#100850000000
1!
1'
1/
#100860000000
0!
0'
0/
#100870000000
1!
1'
1/
#100880000000
0!
0'
0/
#100890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#100900000000
0!
0'
0/
#100910000000
1!
1'
1/
#100920000000
0!
0'
0/
#100930000000
1!
1'
1/
#100940000000
0!
0'
0/
#100950000000
1!
1'
1/
#100960000000
0!
0'
0/
#100970000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#100980000000
0!
0'
0/
#100990000000
1!
1'
1/
#101000000000
0!
0'
0/
#101010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#101020000000
0!
0'
0/
#101030000000
1!
1'
1/
#101040000000
0!
0'
0/
#101050000000
#101060000000
1!
1'
1/
#101070000000
0!
0'
0/
#101080000000
1!
1'
1/
#101090000000
0!
1"
0'
1(
0/
10
#101100000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#101110000000
0!
0'
0/
#101120000000
1!
1'
1/
#101130000000
0!
0'
0/
#101140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#101150000000
0!
0'
0/
#101160000000
1!
1'
1/
#101170000000
0!
1"
0'
1(
0/
10
#101180000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#101190000000
0!
1$
0'
1+
0/
#101200000000
1!
1'
1/
#101210000000
0!
0'
0/
#101220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#101230000000
0!
0'
0/
#101240000000
1!
1'
1/
#101250000000
0!
0'
0/
#101260000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#101270000000
0!
0'
0/
#101280000000
1!
1'
1/
#101290000000
0!
0'
0/
#101300000000
1!
1'
1/
#101310000000
0!
0'
0/
#101320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#101330000000
0!
0'
0/
#101340000000
1!
1'
1/
#101350000000
0!
0'
0/
#101360000000
1!
1'
1/
#101370000000
0!
0'
0/
#101380000000
1!
1'
1/
#101390000000
0!
0'
0/
#101400000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#101410000000
0!
0'
0/
#101420000000
1!
1'
1/
#101430000000
0!
0'
0/
#101440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#101450000000
0!
0'
0/
#101460000000
1!
1'
1/
#101470000000
0!
0'
0/
#101480000000
#101490000000
1!
1'
1/
#101500000000
0!
0'
0/
#101510000000
1!
1'
1/
#101520000000
0!
1"
0'
1(
0/
10
#101530000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#101540000000
0!
0'
0/
#101550000000
1!
1'
1/
#101560000000
0!
0'
0/
#101570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#101580000000
0!
0'
0/
#101590000000
1!
1'
1/
#101600000000
0!
1"
0'
1(
0/
10
#101610000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#101620000000
0!
1$
0'
1+
0/
#101630000000
1!
1'
1/
#101640000000
0!
0'
0/
#101650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#101660000000
0!
0'
0/
#101670000000
1!
1'
1/
#101680000000
0!
0'
0/
#101690000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#101700000000
0!
0'
0/
#101710000000
1!
1'
1/
#101720000000
0!
0'
0/
#101730000000
1!
1'
1/
#101740000000
0!
0'
0/
#101750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#101760000000
0!
0'
0/
#101770000000
1!
1'
1/
#101780000000
0!
0'
0/
#101790000000
1!
1'
1/
#101800000000
0!
0'
0/
#101810000000
1!
1'
1/
#101820000000
0!
0'
0/
#101830000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#101840000000
0!
0'
0/
#101850000000
1!
1'
1/
#101860000000
0!
0'
0/
#101870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#101880000000
0!
0'
0/
#101890000000
1!
1'
1/
#101900000000
0!
0'
0/
#101910000000
#101920000000
1!
1'
1/
#101930000000
0!
0'
0/
#101940000000
1!
1'
1/
#101950000000
0!
1"
0'
1(
0/
10
#101960000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#101970000000
0!
0'
0/
#101980000000
1!
1'
1/
#101990000000
0!
0'
0/
#102000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#102010000000
0!
0'
0/
#102020000000
1!
1'
1/
#102030000000
0!
1"
0'
1(
0/
10
#102040000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#102050000000
0!
1$
0'
1+
0/
#102060000000
1!
1'
1/
#102070000000
0!
0'
0/
#102080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#102090000000
0!
0'
0/
#102100000000
1!
1'
1/
#102110000000
0!
0'
0/
#102120000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#102130000000
0!
0'
0/
#102140000000
1!
1'
1/
#102150000000
0!
0'
0/
#102160000000
1!
1'
1/
#102170000000
0!
0'
0/
#102180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#102190000000
0!
0'
0/
#102200000000
1!
1'
1/
#102210000000
0!
0'
0/
#102220000000
1!
1'
1/
#102230000000
0!
0'
0/
#102240000000
1!
1'
1/
#102250000000
0!
0'
0/
#102260000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#102270000000
0!
0'
0/
#102280000000
1!
1'
1/
#102290000000
0!
0'
0/
#102300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#102310000000
0!
0'
0/
#102320000000
1!
1'
1/
#102330000000
0!
0'
0/
#102340000000
#102350000000
1!
1'
1/
#102360000000
0!
0'
0/
#102370000000
1!
1'
1/
#102380000000
0!
1"
0'
1(
0/
10
#102390000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#102400000000
0!
0'
0/
#102410000000
1!
1'
1/
#102420000000
0!
0'
0/
#102430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#102440000000
0!
0'
0/
#102450000000
1!
1'
1/
#102460000000
0!
1"
0'
1(
0/
10
#102470000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#102480000000
0!
1$
0'
1+
0/
#102490000000
1!
1'
1/
#102500000000
0!
0'
0/
#102510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#102520000000
0!
0'
0/
#102530000000
1!
1'
1/
#102540000000
0!
0'
0/
#102550000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#102560000000
0!
0'
0/
#102570000000
1!
1'
1/
#102580000000
0!
0'
0/
#102590000000
1!
1'
1/
#102600000000
0!
0'
0/
#102610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#102620000000
0!
0'
0/
#102630000000
1!
1'
1/
#102640000000
0!
0'
0/
#102650000000
1!
1'
1/
#102660000000
0!
0'
0/
#102670000000
1!
1'
1/
#102680000000
0!
0'
0/
#102690000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#102700000000
0!
0'
0/
#102710000000
1!
1'
1/
#102720000000
0!
0'
0/
#102730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#102740000000
0!
0'
0/
#102750000000
1!
1'
1/
#102760000000
0!
0'
0/
#102770000000
#102780000000
1!
1'
1/
#102790000000
0!
0'
0/
#102800000000
1!
1'
1/
#102810000000
0!
1"
0'
1(
0/
10
#102820000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#102830000000
0!
0'
0/
#102840000000
1!
1'
1/
#102850000000
0!
0'
0/
#102860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#102870000000
0!
0'
0/
#102880000000
1!
1'
1/
#102890000000
0!
1"
0'
1(
0/
10
#102900000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#102910000000
0!
1$
0'
1+
0/
#102920000000
1!
1'
1/
#102930000000
0!
0'
0/
#102940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#102950000000
0!
0'
0/
#102960000000
1!
1'
1/
#102970000000
0!
0'
0/
#102980000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#102990000000
0!
0'
0/
#103000000000
1!
1'
1/
#103010000000
0!
0'
0/
#103020000000
1!
1'
1/
#103030000000
0!
0'
0/
#103040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#103050000000
0!
0'
0/
#103060000000
1!
1'
1/
#103070000000
0!
0'
0/
#103080000000
1!
1'
1/
#103090000000
0!
0'
0/
#103100000000
1!
1'
1/
#103110000000
0!
0'
0/
#103120000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#103130000000
0!
0'
0/
#103140000000
1!
1'
1/
#103150000000
0!
0'
0/
#103160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#103170000000
0!
0'
0/
#103180000000
1!
1'
1/
#103190000000
0!
0'
0/
#103200000000
#103210000000
1!
1'
1/
#103220000000
0!
0'
0/
#103230000000
1!
1'
1/
#103240000000
0!
1"
0'
1(
0/
10
#103250000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#103260000000
0!
0'
0/
#103270000000
1!
1'
1/
#103280000000
0!
0'
0/
#103290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#103300000000
0!
0'
0/
#103310000000
1!
1'
1/
#103320000000
0!
1"
0'
1(
0/
10
#103330000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#103340000000
0!
1$
0'
1+
0/
#103350000000
1!
1'
1/
#103360000000
0!
0'
0/
#103370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#103380000000
0!
0'
0/
#103390000000
1!
1'
1/
#103400000000
0!
0'
0/
#103410000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#103420000000
0!
0'
0/
#103430000000
1!
1'
1/
#103440000000
0!
0'
0/
#103450000000
1!
1'
1/
#103460000000
0!
0'
0/
#103470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#103480000000
0!
0'
0/
#103490000000
1!
1'
1/
#103500000000
0!
0'
0/
#103510000000
1!
1'
1/
#103520000000
0!
0'
0/
#103530000000
1!
1'
1/
#103540000000
0!
0'
0/
#103550000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#103560000000
0!
0'
0/
#103570000000
1!
1'
1/
#103580000000
0!
0'
0/
#103590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#103600000000
0!
0'
0/
#103610000000
1!
1'
1/
#103620000000
0!
0'
0/
#103630000000
#103640000000
1!
1'
1/
#103650000000
0!
0'
0/
#103660000000
1!
1'
1/
#103670000000
0!
1"
0'
1(
0/
10
#103680000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#103690000000
0!
0'
0/
#103700000000
1!
1'
1/
#103710000000
0!
0'
0/
#103720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#103730000000
0!
0'
0/
#103740000000
1!
1'
1/
#103750000000
0!
1"
0'
1(
0/
10
#103760000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#103770000000
0!
1$
0'
1+
0/
#103780000000
1!
1'
1/
#103790000000
0!
0'
0/
#103800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#103810000000
0!
0'
0/
#103820000000
1!
1'
1/
#103830000000
0!
0'
0/
#103840000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#103850000000
0!
0'
0/
#103860000000
1!
1'
1/
#103870000000
0!
0'
0/
#103880000000
1!
1'
1/
#103890000000
0!
0'
0/
#103900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#103910000000
0!
0'
0/
#103920000000
1!
1'
1/
#103930000000
0!
0'
0/
#103940000000
1!
1'
1/
#103950000000
0!
0'
0/
#103960000000
1!
1'
1/
#103970000000
0!
0'
0/
#103980000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#103990000000
0!
0'
0/
#104000000000
1!
1'
1/
#104010000000
0!
0'
0/
#104020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#104030000000
0!
0'
0/
#104040000000
1!
1'
1/
#104050000000
0!
0'
0/
#104060000000
#104070000000
1!
1'
1/
#104080000000
0!
0'
0/
#104090000000
1!
1'
1/
#104100000000
0!
1"
0'
1(
0/
10
#104110000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#104120000000
0!
0'
0/
#104130000000
1!
1'
1/
#104140000000
0!
0'
0/
#104150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#104160000000
0!
0'
0/
#104170000000
1!
1'
1/
#104180000000
0!
1"
0'
1(
0/
10
#104190000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#104200000000
0!
1$
0'
1+
0/
#104210000000
1!
1'
1/
#104220000000
0!
0'
0/
#104230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#104240000000
0!
0'
0/
#104250000000
1!
1'
1/
#104260000000
0!
0'
0/
#104270000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#104280000000
0!
0'
0/
#104290000000
1!
1'
1/
#104300000000
0!
0'
0/
#104310000000
1!
1'
1/
#104320000000
0!
0'
0/
#104330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#104340000000
0!
0'
0/
#104350000000
1!
1'
1/
#104360000000
0!
0'
0/
#104370000000
1!
1'
1/
#104380000000
0!
0'
0/
#104390000000
1!
1'
1/
#104400000000
0!
0'
0/
#104410000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#104420000000
0!
0'
0/
#104430000000
1!
1'
1/
#104440000000
0!
0'
0/
#104450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#104460000000
0!
0'
0/
#104470000000
1!
1'
1/
#104480000000
0!
0'
0/
#104490000000
#104500000000
1!
1'
1/
#104510000000
0!
0'
0/
#104520000000
1!
1'
1/
#104530000000
0!
1"
0'
1(
0/
10
#104540000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#104550000000
0!
0'
0/
#104560000000
1!
1'
1/
#104570000000
0!
0'
0/
#104580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#104590000000
0!
0'
0/
#104600000000
1!
1'
1/
#104610000000
0!
1"
0'
1(
0/
10
#104620000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#104630000000
0!
1$
0'
1+
0/
#104640000000
1!
1'
1/
#104650000000
0!
0'
0/
#104660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#104670000000
0!
0'
0/
#104680000000
1!
1'
1/
#104690000000
0!
0'
0/
#104700000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#104710000000
0!
0'
0/
#104720000000
1!
1'
1/
#104730000000
0!
0'
0/
#104740000000
1!
1'
1/
#104750000000
0!
0'
0/
#104760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#104770000000
0!
0'
0/
#104780000000
1!
1'
1/
#104790000000
0!
0'
0/
#104800000000
1!
1'
1/
#104810000000
0!
0'
0/
#104820000000
1!
1'
1/
#104830000000
0!
0'
0/
#104840000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#104850000000
0!
0'
0/
#104860000000
1!
1'
1/
#104870000000
0!
0'
0/
#104880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#104890000000
0!
0'
0/
#104900000000
1!
1'
1/
#104910000000
0!
0'
0/
#104920000000
#104930000000
1!
1'
1/
#104940000000
0!
0'
0/
#104950000000
1!
1'
1/
#104960000000
0!
1"
0'
1(
0/
10
#104970000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#104980000000
0!
0'
0/
#104990000000
1!
1'
1/
#105000000000
0!
0'
0/
#105010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#105020000000
0!
0'
0/
#105030000000
1!
1'
1/
#105040000000
0!
1"
0'
1(
0/
10
#105050000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#105060000000
0!
1$
0'
1+
0/
#105070000000
1!
1'
1/
#105080000000
0!
0'
0/
#105090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#105100000000
0!
0'
0/
#105110000000
1!
1'
1/
#105120000000
0!
0'
0/
#105130000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#105140000000
0!
0'
0/
#105150000000
1!
1'
1/
#105160000000
0!
0'
0/
#105170000000
1!
1'
1/
#105180000000
0!
0'
0/
#105190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#105200000000
0!
0'
0/
#105210000000
1!
1'
1/
#105220000000
0!
0'
0/
#105230000000
1!
1'
1/
#105240000000
0!
0'
0/
#105250000000
1!
1'
1/
#105260000000
0!
0'
0/
#105270000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#105280000000
0!
0'
0/
#105290000000
1!
1'
1/
#105300000000
0!
0'
0/
#105310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#105320000000
0!
0'
0/
#105330000000
1!
1'
1/
#105340000000
0!
0'
0/
#105350000000
#105360000000
1!
1'
1/
#105370000000
0!
0'
0/
#105380000000
1!
1'
1/
#105390000000
0!
1"
0'
1(
0/
10
#105400000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#105410000000
0!
0'
0/
#105420000000
1!
1'
1/
#105430000000
0!
0'
0/
#105440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#105450000000
0!
0'
0/
#105460000000
1!
1'
1/
#105470000000
0!
1"
0'
1(
0/
10
#105480000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#105490000000
0!
1$
0'
1+
0/
#105500000000
1!
1'
1/
#105510000000
0!
0'
0/
#105520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#105530000000
0!
0'
0/
#105540000000
1!
1'
1/
#105550000000
0!
0'
0/
#105560000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#105570000000
0!
0'
0/
#105580000000
1!
1'
1/
#105590000000
0!
0'
0/
#105600000000
1!
1'
1/
#105610000000
0!
0'
0/
#105620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#105630000000
0!
0'
0/
#105640000000
1!
1'
1/
#105650000000
0!
0'
0/
#105660000000
1!
1'
1/
#105670000000
0!
0'
0/
#105680000000
1!
1'
1/
#105690000000
0!
0'
0/
#105700000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#105710000000
0!
0'
0/
#105720000000
1!
1'
1/
#105730000000
0!
0'
0/
#105740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#105750000000
0!
0'
0/
#105760000000
1!
1'
1/
#105770000000
0!
0'
0/
#105780000000
#105790000000
1!
1'
1/
#105800000000
0!
0'
0/
#105810000000
1!
1'
1/
#105820000000
0!
1"
0'
1(
0/
10
#105830000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#105840000000
0!
0'
0/
#105850000000
1!
1'
1/
#105860000000
0!
0'
0/
#105870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#105880000000
0!
0'
0/
#105890000000
1!
1'
1/
#105900000000
0!
1"
0'
1(
0/
10
#105910000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#105920000000
0!
1$
0'
1+
0/
#105930000000
1!
1'
1/
#105940000000
0!
0'
0/
#105950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#105960000000
0!
0'
0/
#105970000000
1!
1'
1/
#105980000000
0!
0'
0/
#105990000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#106000000000
0!
0'
0/
#106010000000
1!
1'
1/
#106020000000
0!
0'
0/
#106030000000
1!
1'
1/
#106040000000
0!
0'
0/
#106050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#106060000000
0!
0'
0/
#106070000000
1!
1'
1/
#106080000000
0!
0'
0/
#106090000000
1!
1'
1/
#106100000000
0!
0'
0/
#106110000000
1!
1'
1/
#106120000000
0!
0'
0/
#106130000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#106140000000
0!
0'
0/
#106150000000
1!
1'
1/
#106160000000
0!
0'
0/
#106170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#106180000000
0!
0'
0/
#106190000000
1!
1'
1/
#106200000000
0!
0'
0/
#106210000000
#106220000000
1!
1'
1/
#106230000000
0!
0'
0/
#106240000000
1!
1'
1/
#106250000000
0!
1"
0'
1(
0/
10
#106260000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#106270000000
0!
0'
0/
#106280000000
1!
1'
1/
#106290000000
0!
0'
0/
#106300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#106310000000
0!
0'
0/
#106320000000
1!
1'
1/
#106330000000
0!
1"
0'
1(
0/
10
#106340000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#106350000000
0!
1$
0'
1+
0/
#106360000000
1!
1'
1/
#106370000000
0!
0'
0/
#106380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#106390000000
0!
0'
0/
#106400000000
1!
1'
1/
#106410000000
0!
0'
0/
#106420000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#106430000000
0!
0'
0/
#106440000000
1!
1'
1/
#106450000000
0!
0'
0/
#106460000000
1!
1'
1/
#106470000000
0!
0'
0/
#106480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#106490000000
0!
0'
0/
#106500000000
1!
1'
1/
#106510000000
0!
0'
0/
#106520000000
1!
1'
1/
#106530000000
0!
0'
0/
#106540000000
1!
1'
1/
#106550000000
0!
0'
0/
#106560000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#106570000000
0!
0'
0/
#106580000000
1!
1'
1/
#106590000000
0!
0'
0/
#106600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#106610000000
0!
0'
0/
#106620000000
1!
1'
1/
#106630000000
0!
0'
0/
#106640000000
#106650000000
1!
1'
1/
#106660000000
0!
0'
0/
#106670000000
1!
1'
1/
#106680000000
0!
1"
0'
1(
0/
10
#106690000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#106700000000
0!
0'
0/
#106710000000
1!
1'
1/
#106720000000
0!
0'
0/
#106730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#106740000000
0!
0'
0/
#106750000000
1!
1'
1/
#106760000000
0!
1"
0'
1(
0/
10
#106770000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#106780000000
0!
1$
0'
1+
0/
#106790000000
1!
1'
1/
#106800000000
0!
0'
0/
#106810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#106820000000
0!
0'
0/
#106830000000
1!
1'
1/
#106840000000
0!
0'
0/
#106850000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#106860000000
0!
0'
0/
#106870000000
1!
1'
1/
#106880000000
0!
0'
0/
#106890000000
1!
1'
1/
#106900000000
0!
0'
0/
#106910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#106920000000
0!
0'
0/
#106930000000
1!
1'
1/
#106940000000
0!
0'
0/
#106950000000
1!
1'
1/
#106960000000
0!
0'
0/
#106970000000
1!
1'
1/
#106980000000
0!
0'
0/
#106990000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#107000000000
0!
0'
0/
#107010000000
1!
1'
1/
#107020000000
0!
0'
0/
#107030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#107040000000
0!
0'
0/
#107050000000
1!
1'
1/
#107060000000
0!
0'
0/
#107070000000
#107080000000
1!
1'
1/
#107090000000
0!
0'
0/
#107100000000
1!
1'
1/
#107110000000
0!
1"
0'
1(
0/
10
#107120000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#107130000000
0!
0'
0/
#107140000000
1!
1'
1/
#107150000000
0!
0'
0/
#107160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#107170000000
0!
0'
0/
#107180000000
1!
1'
1/
#107190000000
0!
1"
0'
1(
0/
10
#107200000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#107210000000
0!
1$
0'
1+
0/
#107220000000
1!
1'
1/
#107230000000
0!
0'
0/
#107240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#107250000000
0!
0'
0/
#107260000000
1!
1'
1/
#107270000000
0!
0'
0/
#107280000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#107290000000
0!
0'
0/
#107300000000
1!
1'
1/
#107310000000
0!
0'
0/
#107320000000
1!
1'
1/
#107330000000
0!
0'
0/
#107340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#107350000000
0!
0'
0/
#107360000000
1!
1'
1/
#107370000000
0!
0'
0/
#107380000000
1!
1'
1/
#107390000000
0!
0'
0/
#107400000000
1!
1'
1/
#107410000000
0!
0'
0/
#107420000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#107430000000
0!
0'
0/
#107440000000
1!
1'
1/
#107450000000
0!
0'
0/
#107460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#107470000000
0!
0'
0/
#107480000000
1!
1'
1/
#107490000000
0!
0'
0/
#107500000000
#107510000000
1!
1'
1/
#107520000000
0!
0'
0/
#107530000000
1!
1'
1/
#107540000000
0!
1"
0'
1(
0/
10
#107550000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#107560000000
0!
0'
0/
#107570000000
1!
1'
1/
#107580000000
0!
0'
0/
#107590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#107600000000
0!
0'
0/
#107610000000
1!
1'
1/
#107620000000
0!
1"
0'
1(
0/
10
#107630000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#107640000000
0!
1$
0'
1+
0/
#107650000000
1!
1'
1/
#107660000000
0!
0'
0/
#107670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#107680000000
0!
0'
0/
#107690000000
1!
1'
1/
#107700000000
0!
0'
0/
#107710000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#107720000000
0!
0'
0/
#107730000000
1!
1'
1/
#107740000000
0!
0'
0/
#107750000000
1!
1'
1/
#107760000000
0!
0'
0/
#107770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#107780000000
0!
0'
0/
#107790000000
1!
1'
1/
#107800000000
0!
0'
0/
#107810000000
1!
1'
1/
#107820000000
0!
0'
0/
#107830000000
1!
1'
1/
#107840000000
0!
0'
0/
#107850000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#107860000000
0!
0'
0/
#107870000000
1!
1'
1/
#107880000000
0!
0'
0/
#107890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#107900000000
0!
0'
0/
#107910000000
1!
1'
1/
#107920000000
0!
0'
0/
#107930000000
#107940000000
1!
1'
1/
#107950000000
0!
0'
0/
#107960000000
1!
1'
1/
#107970000000
0!
1"
0'
1(
0/
10
#107980000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#107990000000
0!
0'
0/
#108000000000
1!
1'
1/
#108010000000
0!
0'
0/
#108020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#108030000000
0!
0'
0/
#108040000000
1!
1'
1/
#108050000000
0!
1"
0'
1(
0/
10
#108060000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#108070000000
0!
1$
0'
1+
0/
#108080000000
1!
1'
1/
#108090000000
0!
0'
0/
#108100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#108110000000
0!
0'
0/
#108120000000
1!
1'
1/
#108130000000
0!
0'
0/
#108140000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#108150000000
0!
0'
0/
#108160000000
1!
1'
1/
#108170000000
0!
0'
0/
#108180000000
1!
1'
1/
#108190000000
0!
0'
0/
#108200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#108210000000
0!
0'
0/
#108220000000
1!
1'
1/
#108230000000
0!
0'
0/
#108240000000
1!
1'
1/
#108250000000
0!
0'
0/
#108260000000
1!
1'
1/
#108270000000
0!
0'
0/
#108280000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#108290000000
0!
0'
0/
#108300000000
1!
1'
1/
#108310000000
0!
0'
0/
#108320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#108330000000
0!
0'
0/
#108340000000
1!
1'
1/
#108350000000
0!
0'
0/
#108360000000
#108370000000
1!
1'
1/
#108380000000
0!
0'
0/
#108390000000
1!
1'
1/
#108400000000
0!
1"
0'
1(
0/
10
#108410000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#108420000000
0!
0'
0/
#108430000000
1!
1'
1/
#108440000000
0!
0'
0/
#108450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#108460000000
0!
0'
0/
#108470000000
1!
1'
1/
#108480000000
0!
1"
0'
1(
0/
10
#108490000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#108500000000
0!
1$
0'
1+
0/
#108510000000
1!
1'
1/
#108520000000
0!
0'
0/
#108530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#108540000000
0!
0'
0/
#108550000000
1!
1'
1/
#108560000000
0!
0'
0/
#108570000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#108580000000
0!
0'
0/
#108590000000
1!
1'
1/
#108600000000
0!
0'
0/
#108610000000
1!
1'
1/
#108620000000
0!
0'
0/
#108630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#108640000000
0!
0'
0/
#108650000000
1!
1'
1/
#108660000000
0!
0'
0/
#108670000000
1!
1'
1/
#108680000000
0!
0'
0/
#108690000000
1!
1'
1/
#108700000000
0!
0'
0/
#108710000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#108720000000
0!
0'
0/
#108730000000
1!
1'
1/
#108740000000
0!
0'
0/
#108750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#108760000000
0!
0'
0/
#108770000000
1!
1'
1/
#108780000000
0!
0'
0/
#108790000000
#108800000000
1!
1'
1/
#108810000000
0!
0'
0/
#108820000000
1!
1'
1/
#108830000000
0!
1"
0'
1(
0/
10
#108840000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#108850000000
0!
0'
0/
#108860000000
1!
1'
1/
#108870000000
0!
0'
0/
#108880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#108890000000
0!
0'
0/
#108900000000
1!
1'
1/
#108910000000
0!
1"
0'
1(
0/
10
#108920000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#108930000000
0!
1$
0'
1+
0/
#108940000000
1!
1'
1/
#108950000000
0!
0'
0/
#108960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#108970000000
0!
0'
0/
#108980000000
1!
1'
1/
#108990000000
0!
0'
0/
#109000000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#109010000000
0!
0'
0/
#109020000000
1!
1'
1/
#109030000000
0!
0'
0/
#109040000000
1!
1'
1/
#109050000000
0!
0'
0/
#109060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#109070000000
0!
0'
0/
#109080000000
1!
1'
1/
#109090000000
0!
0'
0/
#109100000000
1!
1'
1/
#109110000000
0!
0'
0/
#109120000000
1!
1'
1/
#109130000000
0!
0'
0/
#109140000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#109150000000
0!
0'
0/
#109160000000
1!
1'
1/
#109170000000
0!
0'
0/
#109180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#109190000000
0!
0'
0/
#109200000000
1!
1'
1/
#109210000000
0!
0'
0/
#109220000000
#109230000000
1!
1'
1/
#109240000000
0!
0'
0/
#109250000000
1!
1'
1/
#109260000000
0!
1"
0'
1(
0/
10
#109270000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#109280000000
0!
0'
0/
#109290000000
1!
1'
1/
#109300000000
0!
0'
0/
#109310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#109320000000
0!
0'
0/
#109330000000
1!
1'
1/
#109340000000
0!
1"
0'
1(
0/
10
#109350000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#109360000000
0!
1$
0'
1+
0/
#109370000000
1!
1'
1/
#109380000000
0!
0'
0/
#109390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#109400000000
0!
0'
0/
#109410000000
1!
1'
1/
#109420000000
0!
0'
0/
#109430000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#109440000000
0!
0'
0/
#109450000000
1!
1'
1/
#109460000000
0!
0'
0/
#109470000000
1!
1'
1/
#109480000000
0!
0'
0/
#109490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#109500000000
0!
0'
0/
#109510000000
1!
1'
1/
#109520000000
0!
0'
0/
#109530000000
1!
1'
1/
#109540000000
0!
0'
0/
#109550000000
1!
1'
1/
#109560000000
0!
0'
0/
#109570000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#109580000000
0!
0'
0/
#109590000000
1!
1'
1/
#109600000000
0!
0'
0/
#109610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#109620000000
0!
0'
0/
#109630000000
1!
1'
1/
#109640000000
0!
0'
0/
#109650000000
#109660000000
1!
1'
1/
#109670000000
0!
0'
0/
#109680000000
1!
1'
1/
#109690000000
0!
1"
0'
1(
0/
10
#109700000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#109710000000
0!
0'
0/
#109720000000
1!
1'
1/
#109730000000
0!
0'
0/
#109740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#109750000000
0!
0'
0/
#109760000000
1!
1'
1/
#109770000000
0!
1"
0'
1(
0/
10
#109780000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#109790000000
0!
1$
0'
1+
0/
#109800000000
1!
1'
1/
#109810000000
0!
0'
0/
#109820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#109830000000
0!
0'
0/
#109840000000
1!
1'
1/
#109850000000
0!
0'
0/
#109860000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#109870000000
0!
0'
0/
#109880000000
1!
1'
1/
#109890000000
0!
0'
0/
#109900000000
1!
1'
1/
#109910000000
0!
0'
0/
#109920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#109930000000
0!
0'
0/
#109940000000
1!
1'
1/
#109950000000
0!
0'
0/
#109960000000
1!
1'
1/
#109970000000
0!
0'
0/
#109980000000
1!
1'
1/
#109990000000
0!
0'
0/
#110000000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#110010000000
0!
0'
0/
#110020000000
1!
1'
1/
#110030000000
0!
0'
0/
#110040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#110050000000
0!
0'
0/
#110060000000
1!
1'
1/
#110070000000
0!
0'
0/
#110080000000
#110090000000
1!
1'
1/
#110100000000
0!
0'
0/
#110110000000
1!
1'
1/
#110120000000
0!
1"
0'
1(
0/
10
#110130000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#110140000000
0!
0'
0/
#110150000000
1!
1'
1/
#110160000000
0!
0'
0/
#110170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#110180000000
0!
0'
0/
#110190000000
1!
1'
1/
#110200000000
0!
1"
0'
1(
0/
10
#110210000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#110220000000
0!
1$
0'
1+
0/
#110230000000
1!
1'
1/
#110240000000
0!
0'
0/
#110250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#110260000000
0!
0'
0/
#110270000000
1!
1'
1/
#110280000000
0!
0'
0/
#110290000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#110300000000
0!
0'
0/
#110310000000
1!
1'
1/
#110320000000
0!
0'
0/
#110330000000
1!
1'
1/
#110340000000
0!
0'
0/
#110350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#110360000000
0!
0'
0/
#110370000000
1!
1'
1/
#110380000000
0!
0'
0/
#110390000000
1!
1'
1/
#110400000000
0!
0'
0/
#110410000000
1!
1'
1/
#110420000000
0!
0'
0/
#110430000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#110440000000
0!
0'
0/
#110450000000
1!
1'
1/
#110460000000
0!
0'
0/
#110470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#110480000000
0!
0'
0/
#110490000000
1!
1'
1/
#110500000000
0!
0'
0/
#110510000000
#110520000000
1!
1'
1/
#110530000000
0!
0'
0/
#110540000000
1!
1'
1/
#110550000000
0!
1"
0'
1(
0/
10
#110560000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#110570000000
0!
0'
0/
#110580000000
1!
1'
1/
#110590000000
0!
0'
0/
#110600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#110610000000
0!
0'
0/
#110620000000
1!
1'
1/
#110630000000
0!
1"
0'
1(
0/
10
#110640000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#110650000000
0!
1$
0'
1+
0/
#110660000000
1!
1'
1/
#110670000000
0!
0'
0/
#110680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#110690000000
0!
0'
0/
#110700000000
1!
1'
1/
#110710000000
0!
0'
0/
#110720000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#110730000000
0!
0'
0/
#110740000000
1!
1'
1/
#110750000000
0!
0'
0/
#110760000000
1!
1'
1/
#110770000000
0!
0'
0/
#110780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#110790000000
0!
0'
0/
#110800000000
1!
1'
1/
#110810000000
0!
0'
0/
#110820000000
1!
1'
1/
#110830000000
0!
0'
0/
#110840000000
1!
1'
1/
#110850000000
0!
0'
0/
#110860000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#110870000000
0!
0'
0/
#110880000000
1!
1'
1/
#110890000000
0!
0'
0/
#110900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#110910000000
0!
0'
0/
#110920000000
1!
1'
1/
#110930000000
0!
0'
0/
#110940000000
#110950000000
1!
1'
1/
#110960000000
0!
0'
0/
#110970000000
1!
1'
1/
#110980000000
0!
1"
0'
1(
0/
10
#110990000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#111000000000
0!
0'
0/
#111010000000
1!
1'
1/
#111020000000
0!
0'
0/
#111030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#111040000000
0!
0'
0/
#111050000000
1!
1'
1/
#111060000000
0!
1"
0'
1(
0/
10
#111070000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#111080000000
0!
1$
0'
1+
0/
#111090000000
1!
1'
1/
#111100000000
0!
0'
0/
#111110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#111120000000
0!
0'
0/
#111130000000
1!
1'
1/
#111140000000
0!
0'
0/
#111150000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#111160000000
0!
0'
0/
#111170000000
1!
1'
1/
#111180000000
0!
0'
0/
#111190000000
1!
1'
1/
#111200000000
0!
0'
0/
#111210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#111220000000
0!
0'
0/
#111230000000
1!
1'
1/
#111240000000
0!
0'
0/
#111250000000
1!
1'
1/
#111260000000
0!
0'
0/
#111270000000
1!
1'
1/
#111280000000
0!
0'
0/
#111290000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#111300000000
0!
0'
0/
#111310000000
1!
1'
1/
#111320000000
0!
0'
0/
#111330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#111340000000
0!
0'
0/
#111350000000
1!
1'
1/
#111360000000
0!
0'
0/
#111370000000
#111380000000
1!
1'
1/
#111390000000
0!
0'
0/
#111400000000
1!
1'
1/
#111410000000
0!
1"
0'
1(
0/
10
#111420000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#111430000000
0!
0'
0/
#111440000000
1!
1'
1/
#111450000000
0!
0'
0/
#111460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#111470000000
0!
0'
0/
#111480000000
1!
1'
1/
#111490000000
0!
1"
0'
1(
0/
10
#111500000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#111510000000
0!
1$
0'
1+
0/
#111520000000
1!
1'
1/
#111530000000
0!
0'
0/
#111540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#111550000000
0!
0'
0/
#111560000000
1!
1'
1/
#111570000000
0!
0'
0/
#111580000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#111590000000
0!
0'
0/
#111600000000
1!
1'
1/
#111610000000
0!
0'
0/
#111620000000
1!
1'
1/
#111630000000
0!
0'
0/
#111640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#111650000000
0!
0'
0/
#111660000000
1!
1'
1/
#111670000000
0!
0'
0/
#111680000000
1!
1'
1/
#111690000000
0!
0'
0/
#111700000000
1!
1'
1/
#111710000000
0!
0'
0/
#111720000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#111730000000
0!
0'
0/
#111740000000
1!
1'
1/
#111750000000
0!
0'
0/
#111760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#111770000000
0!
0'
0/
#111780000000
1!
1'
1/
#111790000000
0!
0'
0/
#111800000000
#111810000000
1!
1'
1/
#111820000000
0!
0'
0/
#111830000000
1!
1'
1/
#111840000000
0!
1"
0'
1(
0/
10
#111850000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#111860000000
0!
0'
0/
#111870000000
1!
1'
1/
#111880000000
0!
0'
0/
#111890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#111900000000
0!
0'
0/
#111910000000
1!
1'
1/
#111920000000
0!
1"
0'
1(
0/
10
#111930000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#111940000000
0!
1$
0'
1+
0/
#111950000000
1!
1'
1/
#111960000000
0!
0'
0/
#111970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#111980000000
0!
0'
0/
#111990000000
1!
1'
1/
#112000000000
0!
0'
0/
#112010000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#112020000000
0!
0'
0/
#112030000000
1!
1'
1/
#112040000000
0!
0'
0/
#112050000000
1!
1'
1/
#112060000000
0!
0'
0/
#112070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#112080000000
0!
0'
0/
#112090000000
1!
1'
1/
#112100000000
0!
0'
0/
#112110000000
1!
1'
1/
#112120000000
0!
0'
0/
#112130000000
1!
1'
1/
#112140000000
0!
0'
0/
#112150000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#112160000000
0!
0'
0/
#112170000000
1!
1'
1/
#112180000000
0!
0'
0/
#112190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#112200000000
0!
0'
0/
#112210000000
1!
1'
1/
#112220000000
0!
0'
0/
#112230000000
#112240000000
1!
1'
1/
#112250000000
0!
0'
0/
#112260000000
1!
1'
1/
#112270000000
0!
1"
0'
1(
0/
10
#112280000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#112290000000
0!
0'
0/
#112300000000
1!
1'
1/
#112310000000
0!
0'
0/
#112320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#112330000000
0!
0'
0/
#112340000000
1!
1'
1/
#112350000000
0!
1"
0'
1(
0/
10
#112360000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#112370000000
0!
1$
0'
1+
0/
#112380000000
1!
1'
1/
#112390000000
0!
0'
0/
#112400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#112410000000
0!
0'
0/
#112420000000
1!
1'
1/
#112430000000
0!
0'
0/
#112440000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#112450000000
0!
0'
0/
#112460000000
1!
1'
1/
#112470000000
0!
0'
0/
#112480000000
1!
1'
1/
#112490000000
0!
0'
0/
#112500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#112510000000
0!
0'
0/
#112520000000
1!
1'
1/
#112530000000
0!
0'
0/
#112540000000
1!
1'
1/
#112550000000
0!
0'
0/
#112560000000
1!
1'
1/
#112570000000
0!
0'
0/
#112580000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#112590000000
0!
0'
0/
#112600000000
1!
1'
1/
#112610000000
0!
0'
0/
#112620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#112630000000
0!
0'
0/
#112640000000
1!
1'
1/
#112650000000
0!
0'
0/
#112660000000
#112670000000
1!
1'
1/
#112680000000
0!
0'
0/
#112690000000
1!
1'
1/
#112700000000
0!
1"
0'
1(
0/
10
#112710000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#112720000000
0!
0'
0/
#112730000000
1!
1'
1/
#112740000000
0!
0'
0/
#112750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#112760000000
0!
0'
0/
#112770000000
1!
1'
1/
#112780000000
0!
1"
0'
1(
0/
10
#112790000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#112800000000
0!
1$
0'
1+
0/
#112810000000
1!
1'
1/
#112820000000
0!
0'
0/
#112830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#112840000000
0!
0'
0/
#112850000000
1!
1'
1/
#112860000000
0!
0'
0/
#112870000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#112880000000
0!
0'
0/
#112890000000
1!
1'
1/
#112900000000
0!
0'
0/
#112910000000
1!
1'
1/
#112920000000
0!
0'
0/
#112930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#112940000000
0!
0'
0/
#112950000000
1!
1'
1/
#112960000000
0!
0'
0/
#112970000000
1!
1'
1/
#112980000000
0!
0'
0/
#112990000000
1!
1'
1/
#113000000000
0!
0'
0/
#113010000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#113020000000
0!
0'
0/
#113030000000
1!
1'
1/
#113040000000
0!
0'
0/
#113050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#113060000000
0!
0'
0/
#113070000000
1!
1'
1/
#113080000000
0!
0'
0/
#113090000000
#113100000000
1!
1'
1/
#113110000000
0!
0'
0/
#113120000000
1!
1'
1/
#113130000000
0!
1"
0'
1(
0/
10
#113140000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#113150000000
0!
0'
0/
#113160000000
1!
1'
1/
#113170000000
0!
0'
0/
#113180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#113190000000
0!
0'
0/
#113200000000
1!
1'
1/
#113210000000
0!
1"
0'
1(
0/
10
#113220000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#113230000000
0!
1$
0'
1+
0/
#113240000000
1!
1'
1/
#113250000000
0!
0'
0/
#113260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#113270000000
0!
0'
0/
#113280000000
1!
1'
1/
#113290000000
0!
0'
0/
#113300000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#113310000000
0!
0'
0/
#113320000000
1!
1'
1/
#113330000000
0!
0'
0/
#113340000000
1!
1'
1/
#113350000000
0!
0'
0/
#113360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#113370000000
0!
0'
0/
#113380000000
1!
1'
1/
#113390000000
0!
0'
0/
#113400000000
1!
1'
1/
#113410000000
0!
0'
0/
#113420000000
1!
1'
1/
#113430000000
0!
0'
0/
#113440000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#113450000000
0!
0'
0/
#113460000000
1!
1'
1/
#113470000000
0!
0'
0/
#113480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#113490000000
0!
0'
0/
#113500000000
1!
1'
1/
#113510000000
0!
0'
0/
#113520000000
#113530000000
1!
1'
1/
#113540000000
0!
0'
0/
#113550000000
1!
1'
1/
#113560000000
0!
1"
0'
1(
0/
10
#113570000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#113580000000
0!
0'
0/
#113590000000
1!
1'
1/
#113600000000
0!
0'
0/
#113610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#113620000000
0!
0'
0/
#113630000000
1!
1'
1/
#113640000000
0!
1"
0'
1(
0/
10
#113650000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#113660000000
0!
1$
0'
1+
0/
#113670000000
1!
1'
1/
#113680000000
0!
0'
0/
#113690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#113700000000
0!
0'
0/
#113710000000
1!
1'
1/
#113720000000
0!
0'
0/
#113730000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#113740000000
0!
0'
0/
#113750000000
1!
1'
1/
#113760000000
0!
0'
0/
#113770000000
1!
1'
1/
#113780000000
0!
0'
0/
#113790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#113800000000
0!
0'
0/
#113810000000
1!
1'
1/
#113820000000
0!
0'
0/
#113830000000
1!
1'
1/
#113840000000
0!
0'
0/
#113850000000
1!
1'
1/
#113860000000
0!
0'
0/
#113870000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#113880000000
0!
0'
0/
#113890000000
1!
1'
1/
#113900000000
0!
0'
0/
#113910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#113920000000
0!
0'
0/
#113930000000
1!
1'
1/
#113940000000
0!
0'
0/
#113950000000
#113960000000
1!
1'
1/
#113970000000
0!
0'
0/
#113980000000
1!
1'
1/
#113990000000
0!
1"
0'
1(
0/
10
#114000000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#114010000000
0!
0'
0/
#114020000000
1!
1'
1/
#114030000000
0!
0'
0/
#114040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#114050000000
0!
0'
0/
#114060000000
1!
1'
1/
#114070000000
0!
1"
0'
1(
0/
10
#114080000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#114090000000
0!
1$
0'
1+
0/
#114100000000
1!
1'
1/
#114110000000
0!
0'
0/
#114120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#114130000000
0!
0'
0/
#114140000000
1!
1'
1/
#114150000000
0!
0'
0/
#114160000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#114170000000
0!
0'
0/
#114180000000
1!
1'
1/
#114190000000
0!
0'
0/
#114200000000
1!
1'
1/
#114210000000
0!
0'
0/
#114220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#114230000000
0!
0'
0/
#114240000000
1!
1'
1/
#114250000000
0!
0'
0/
#114260000000
1!
1'
1/
#114270000000
0!
0'
0/
#114280000000
1!
1'
1/
#114290000000
0!
0'
0/
#114300000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#114310000000
0!
0'
0/
#114320000000
1!
1'
1/
#114330000000
0!
0'
0/
#114340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#114350000000
0!
0'
0/
#114360000000
1!
1'
1/
#114370000000
0!
0'
0/
#114380000000
#114390000000
1!
1'
1/
#114400000000
0!
0'
0/
#114410000000
1!
1'
1/
#114420000000
0!
1"
0'
1(
0/
10
#114430000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#114440000000
0!
0'
0/
#114450000000
1!
1'
1/
#114460000000
0!
0'
0/
#114470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#114480000000
0!
0'
0/
#114490000000
1!
1'
1/
#114500000000
0!
1"
0'
1(
0/
10
#114510000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#114520000000
0!
1$
0'
1+
0/
#114530000000
1!
1'
1/
#114540000000
0!
0'
0/
#114550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#114560000000
0!
0'
0/
#114570000000
1!
1'
1/
#114580000000
0!
0'
0/
#114590000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#114600000000
0!
0'
0/
#114610000000
1!
1'
1/
#114620000000
0!
0'
0/
#114630000000
1!
1'
1/
#114640000000
0!
0'
0/
#114650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#114660000000
0!
0'
0/
#114670000000
1!
1'
1/
#114680000000
0!
0'
0/
#114690000000
1!
1'
1/
#114700000000
0!
0'
0/
#114710000000
1!
1'
1/
#114720000000
0!
0'
0/
#114730000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#114740000000
0!
0'
0/
#114750000000
1!
1'
1/
#114760000000
0!
0'
0/
#114770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#114780000000
0!
0'
0/
#114790000000
1!
1'
1/
#114800000000
0!
0'
0/
#114810000000
#114820000000
1!
1'
1/
#114830000000
0!
0'
0/
#114840000000
1!
1'
1/
#114850000000
0!
1"
0'
1(
0/
10
#114860000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#114870000000
0!
0'
0/
#114880000000
1!
1'
1/
#114890000000
0!
0'
0/
#114900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#114910000000
0!
0'
0/
#114920000000
1!
1'
1/
#114930000000
0!
1"
0'
1(
0/
10
#114940000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#114950000000
0!
1$
0'
1+
0/
#114960000000
1!
1'
1/
#114970000000
0!
0'
0/
#114980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#114990000000
0!
0'
0/
#115000000000
1!
1'
1/
#115010000000
0!
0'
0/
#115020000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#115030000000
0!
0'
0/
#115040000000
1!
1'
1/
#115050000000
0!
0'
0/
#115060000000
1!
1'
1/
#115070000000
0!
0'
0/
#115080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#115090000000
0!
0'
0/
#115100000000
1!
1'
1/
#115110000000
0!
0'
0/
#115120000000
1!
1'
1/
#115130000000
0!
0'
0/
#115140000000
1!
1'
1/
#115150000000
0!
0'
0/
#115160000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#115170000000
0!
0'
0/
#115180000000
1!
1'
1/
#115190000000
0!
0'
0/
#115200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#115210000000
0!
0'
0/
#115220000000
1!
1'
1/
#115230000000
0!
0'
0/
#115240000000
#115250000000
1!
1'
1/
#115260000000
0!
0'
0/
#115270000000
1!
1'
1/
#115280000000
0!
1"
0'
1(
0/
10
#115290000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#115300000000
0!
0'
0/
#115310000000
1!
1'
1/
#115320000000
0!
0'
0/
#115330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#115340000000
0!
0'
0/
#115350000000
1!
1'
1/
#115360000000
0!
1"
0'
1(
0/
10
#115370000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#115380000000
0!
1$
0'
1+
0/
#115390000000
1!
1'
1/
#115400000000
0!
0'
0/
#115410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#115420000000
0!
0'
0/
#115430000000
1!
1'
1/
#115440000000
0!
0'
0/
#115450000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#115460000000
0!
0'
0/
#115470000000
1!
1'
1/
#115480000000
0!
0'
0/
#115490000000
1!
1'
1/
#115500000000
0!
0'
0/
#115510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#115520000000
0!
0'
0/
#115530000000
1!
1'
1/
#115540000000
0!
0'
0/
#115550000000
1!
1'
1/
#115560000000
0!
0'
0/
#115570000000
1!
1'
1/
#115580000000
0!
0'
0/
#115590000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#115600000000
0!
0'
0/
#115610000000
1!
1'
1/
#115620000000
0!
0'
0/
#115630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#115640000000
0!
0'
0/
#115650000000
1!
1'
1/
#115660000000
0!
0'
0/
#115670000000
#115680000000
1!
1'
1/
#115690000000
0!
0'
0/
#115700000000
1!
1'
1/
#115710000000
0!
1"
0'
1(
0/
10
#115720000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#115730000000
0!
0'
0/
#115740000000
1!
1'
1/
#115750000000
0!
0'
0/
#115760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#115770000000
0!
0'
0/
#115780000000
1!
1'
1/
#115790000000
0!
1"
0'
1(
0/
10
#115800000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#115810000000
0!
1$
0'
1+
0/
#115820000000
1!
1'
1/
#115830000000
0!
0'
0/
#115840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#115850000000
0!
0'
0/
#115860000000
1!
1'
1/
#115870000000
0!
0'
0/
#115880000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#115890000000
0!
0'
0/
#115900000000
1!
1'
1/
#115910000000
0!
0'
0/
#115920000000
1!
1'
1/
#115930000000
0!
0'
0/
#115940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#115950000000
0!
0'
0/
#115960000000
1!
1'
1/
#115970000000
0!
0'
0/
#115980000000
1!
1'
1/
#115990000000
0!
0'
0/
#116000000000
1!
1'
1/
#116010000000
0!
0'
0/
#116020000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#116030000000
0!
0'
0/
#116040000000
1!
1'
1/
#116050000000
0!
0'
0/
#116060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#116070000000
0!
0'
0/
#116080000000
1!
1'
1/
#116090000000
0!
0'
0/
#116100000000
#116110000000
1!
1'
1/
#116120000000
0!
0'
0/
#116130000000
1!
1'
1/
#116140000000
0!
1"
0'
1(
0/
10
#116150000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#116160000000
0!
0'
0/
#116170000000
1!
1'
1/
#116180000000
0!
0'
0/
#116190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#116200000000
0!
0'
0/
#116210000000
1!
1'
1/
#116220000000
0!
1"
0'
1(
0/
10
#116230000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#116240000000
0!
1$
0'
1+
0/
#116250000000
1!
1'
1/
#116260000000
0!
0'
0/
#116270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#116280000000
0!
0'
0/
#116290000000
1!
1'
1/
#116300000000
0!
0'
0/
#116310000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#116320000000
0!
0'
0/
#116330000000
1!
1'
1/
#116340000000
0!
0'
0/
#116350000000
1!
1'
1/
#116360000000
0!
0'
0/
#116370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#116380000000
0!
0'
0/
#116390000000
1!
1'
1/
#116400000000
0!
0'
0/
#116410000000
1!
1'
1/
#116420000000
0!
0'
0/
#116430000000
1!
1'
1/
#116440000000
0!
0'
0/
#116450000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#116460000000
0!
0'
0/
#116470000000
1!
1'
1/
#116480000000
0!
0'
0/
#116490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#116500000000
0!
0'
0/
#116510000000
1!
1'
1/
#116520000000
0!
0'
0/
#116530000000
#116540000000
1!
1'
1/
#116550000000
0!
0'
0/
#116560000000
1!
1'
1/
#116570000000
0!
1"
0'
1(
0/
10
#116580000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#116590000000
0!
0'
0/
#116600000000
1!
1'
1/
#116610000000
0!
0'
0/
#116620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#116630000000
0!
0'
0/
#116640000000
1!
1'
1/
#116650000000
0!
1"
0'
1(
0/
10
#116660000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#116670000000
0!
1$
0'
1+
0/
#116680000000
1!
1'
1/
#116690000000
0!
0'
0/
#116700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#116710000000
0!
0'
0/
#116720000000
1!
1'
1/
#116730000000
0!
0'
0/
#116740000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#116750000000
0!
0'
0/
#116760000000
1!
1'
1/
#116770000000
0!
0'
0/
#116780000000
1!
1'
1/
#116790000000
0!
0'
0/
#116800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#116810000000
0!
0'
0/
#116820000000
1!
1'
1/
#116830000000
0!
0'
0/
#116840000000
1!
1'
1/
#116850000000
0!
0'
0/
#116860000000
1!
1'
1/
#116870000000
0!
0'
0/
#116880000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#116890000000
0!
0'
0/
#116900000000
1!
1'
1/
#116910000000
0!
0'
0/
#116920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#116930000000
0!
0'
0/
#116940000000
1!
1'
1/
#116950000000
0!
0'
0/
#116960000000
#116970000000
1!
1'
1/
#116980000000
0!
0'
0/
#116990000000
1!
1'
1/
#117000000000
0!
1"
0'
1(
0/
10
#117010000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#117020000000
0!
0'
0/
#117030000000
1!
1'
1/
#117040000000
0!
0'
0/
#117050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#117060000000
0!
0'
0/
#117070000000
1!
1'
1/
#117080000000
0!
1"
0'
1(
0/
10
#117090000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#117100000000
0!
1$
0'
1+
0/
#117110000000
1!
1'
1/
#117120000000
0!
0'
0/
#117130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#117140000000
0!
0'
0/
#117150000000
1!
1'
1/
#117160000000
0!
0'
0/
#117170000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#117180000000
0!
0'
0/
#117190000000
1!
1'
1/
#117200000000
0!
0'
0/
#117210000000
1!
1'
1/
#117220000000
0!
0'
0/
#117230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#117240000000
0!
0'
0/
#117250000000
1!
1'
1/
#117260000000
0!
0'
0/
#117270000000
1!
1'
1/
#117280000000
0!
0'
0/
#117290000000
1!
1'
1/
#117300000000
0!
0'
0/
#117310000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#117320000000
0!
0'
0/
#117330000000
1!
1'
1/
#117340000000
0!
0'
0/
#117350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#117360000000
0!
0'
0/
#117370000000
1!
1'
1/
#117380000000
0!
0'
0/
#117390000000
#117400000000
1!
1'
1/
#117410000000
0!
0'
0/
#117420000000
1!
1'
1/
#117430000000
0!
1"
0'
1(
0/
10
#117440000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#117450000000
0!
0'
0/
#117460000000
1!
1'
1/
#117470000000
0!
0'
0/
#117480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#117490000000
0!
0'
0/
#117500000000
1!
1'
1/
#117510000000
0!
1"
0'
1(
0/
10
#117520000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#117530000000
0!
1$
0'
1+
0/
#117540000000
1!
1'
1/
#117550000000
0!
0'
0/
#117560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#117570000000
0!
0'
0/
#117580000000
1!
1'
1/
#117590000000
0!
0'
0/
#117600000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#117610000000
0!
0'
0/
#117620000000
1!
1'
1/
#117630000000
0!
0'
0/
#117640000000
1!
1'
1/
#117650000000
0!
0'
0/
#117660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#117670000000
0!
0'
0/
#117680000000
1!
1'
1/
#117690000000
0!
0'
0/
#117700000000
1!
1'
1/
#117710000000
0!
0'
0/
#117720000000
1!
1'
1/
#117730000000
0!
0'
0/
#117740000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#117750000000
0!
0'
0/
#117760000000
1!
1'
1/
#117770000000
0!
0'
0/
#117780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#117790000000
0!
0'
0/
#117800000000
1!
1'
1/
#117810000000
0!
0'
0/
#117820000000
#117830000000
1!
1'
1/
#117840000000
0!
0'
0/
#117850000000
1!
1'
1/
#117860000000
0!
1"
0'
1(
0/
10
#117870000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#117880000000
0!
0'
0/
#117890000000
1!
1'
1/
#117900000000
0!
0'
0/
#117910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#117920000000
0!
0'
0/
#117930000000
1!
1'
1/
#117940000000
0!
1"
0'
1(
0/
10
#117950000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#117960000000
0!
1$
0'
1+
0/
#117970000000
1!
1'
1/
#117980000000
0!
0'
0/
#117990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#118000000000
0!
0'
0/
#118010000000
1!
1'
1/
#118020000000
0!
0'
0/
#118030000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#118040000000
0!
0'
0/
#118050000000
1!
1'
1/
#118060000000
0!
0'
0/
#118070000000
1!
1'
1/
#118080000000
0!
0'
0/
#118090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#118100000000
0!
0'
0/
#118110000000
1!
1'
1/
#118120000000
0!
0'
0/
#118130000000
1!
1'
1/
#118140000000
0!
0'
0/
#118150000000
1!
1'
1/
#118160000000
0!
0'
0/
#118170000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#118180000000
0!
0'
0/
#118190000000
1!
1'
1/
#118200000000
0!
0'
0/
#118210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#118220000000
0!
0'
0/
#118230000000
1!
1'
1/
#118240000000
0!
0'
0/
#118250000000
#118260000000
1!
1'
1/
#118270000000
0!
0'
0/
#118280000000
1!
1'
1/
#118290000000
0!
1"
0'
1(
0/
10
#118300000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#118310000000
0!
0'
0/
#118320000000
1!
1'
1/
#118330000000
0!
0'
0/
#118340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#118350000000
0!
0'
0/
#118360000000
1!
1'
1/
#118370000000
0!
1"
0'
1(
0/
10
#118380000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#118390000000
0!
1$
0'
1+
0/
#118400000000
1!
1'
1/
#118410000000
0!
0'
0/
#118420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#118430000000
0!
0'
0/
#118440000000
1!
1'
1/
#118450000000
0!
0'
0/
#118460000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#118470000000
0!
0'
0/
#118480000000
1!
1'
1/
#118490000000
0!
0'
0/
#118500000000
1!
1'
1/
#118510000000
0!
0'
0/
#118520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#118530000000
0!
0'
0/
#118540000000
1!
1'
1/
#118550000000
0!
0'
0/
#118560000000
1!
1'
1/
#118570000000
0!
0'
0/
#118580000000
1!
1'
1/
#118590000000
0!
0'
0/
#118600000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#118610000000
0!
0'
0/
#118620000000
1!
1'
1/
#118630000000
0!
0'
0/
#118640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#118650000000
0!
0'
0/
#118660000000
1!
1'
1/
#118670000000
0!
0'
0/
#118680000000
#118690000000
1!
1'
1/
#118700000000
0!
0'
0/
#118710000000
1!
1'
1/
#118720000000
0!
1"
0'
1(
0/
10
#118730000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#118740000000
0!
0'
0/
#118750000000
1!
1'
1/
#118760000000
0!
0'
0/
#118770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#118780000000
0!
0'
0/
#118790000000
1!
1'
1/
#118800000000
0!
1"
0'
1(
0/
10
#118810000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#118820000000
0!
1$
0'
1+
0/
#118830000000
1!
1'
1/
#118840000000
0!
0'
0/
#118850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#118860000000
0!
0'
0/
#118870000000
1!
1'
1/
#118880000000
0!
0'
0/
#118890000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#118900000000
0!
0'
0/
#118910000000
1!
1'
1/
#118920000000
0!
0'
0/
#118930000000
1!
1'
1/
#118940000000
0!
0'
0/
#118950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#118960000000
0!
0'
0/
#118970000000
1!
1'
1/
#118980000000
0!
0'
0/
#118990000000
1!
1'
1/
#119000000000
0!
0'
0/
#119010000000
1!
1'
1/
#119020000000
0!
0'
0/
#119030000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#119040000000
0!
0'
0/
#119050000000
1!
1'
1/
#119060000000
0!
0'
0/
#119070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#119080000000
0!
0'
0/
#119090000000
1!
1'
1/
#119100000000
0!
0'
0/
#119110000000
#119120000000
1!
1'
1/
#119130000000
0!
0'
0/
#119140000000
1!
1'
1/
#119150000000
0!
1"
0'
1(
0/
10
#119160000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#119170000000
0!
0'
0/
#119180000000
1!
1'
1/
#119190000000
0!
0'
0/
#119200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#119210000000
0!
0'
0/
#119220000000
1!
1'
1/
#119230000000
0!
1"
0'
1(
0/
10
#119240000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#119250000000
0!
1$
0'
1+
0/
#119260000000
1!
1'
1/
#119270000000
0!
0'
0/
#119280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#119290000000
0!
0'
0/
#119300000000
1!
1'
1/
#119310000000
0!
0'
0/
#119320000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#119330000000
0!
0'
0/
#119340000000
1!
1'
1/
#119350000000
0!
0'
0/
#119360000000
1!
1'
1/
#119370000000
0!
0'
0/
#119380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#119390000000
0!
0'
0/
#119400000000
1!
1'
1/
#119410000000
0!
0'
0/
#119420000000
1!
1'
1/
#119430000000
0!
0'
0/
#119440000000
1!
1'
1/
#119450000000
0!
0'
0/
#119460000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#119470000000
0!
0'
0/
#119480000000
1!
1'
1/
#119490000000
0!
0'
0/
#119500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#119510000000
0!
0'
0/
#119520000000
1!
1'
1/
#119530000000
0!
0'
0/
#119540000000
#119550000000
1!
1'
1/
#119560000000
0!
0'
0/
#119570000000
1!
1'
1/
#119580000000
0!
1"
0'
1(
0/
10
#119590000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#119600000000
0!
0'
0/
#119610000000
1!
1'
1/
#119620000000
0!
0'
0/
#119630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#119640000000
0!
0'
0/
#119650000000
1!
1'
1/
#119660000000
0!
1"
0'
1(
0/
10
#119670000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#119680000000
0!
1$
0'
1+
0/
#119690000000
1!
1'
1/
#119700000000
0!
0'
0/
#119710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#119720000000
0!
0'
0/
#119730000000
1!
1'
1/
#119740000000
0!
0'
0/
#119750000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#119760000000
0!
0'
0/
#119770000000
1!
1'
1/
#119780000000
0!
0'
0/
#119790000000
1!
1'
1/
#119800000000
0!
0'
0/
#119810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#119820000000
0!
0'
0/
#119830000000
1!
1'
1/
#119840000000
0!
0'
0/
#119850000000
1!
1'
1/
#119860000000
0!
0'
0/
#119870000000
1!
1'
1/
#119880000000
0!
0'
0/
#119890000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#119900000000
0!
0'
0/
#119910000000
1!
1'
1/
#119920000000
0!
0'
0/
#119930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#119940000000
0!
0'
0/
#119950000000
1!
1'
1/
#119960000000
0!
0'
0/
#119970000000
#119980000000
1!
1'
1/
#119990000000
0!
0'
0/
#120000000000
1!
1'
1/
#120010000000
0!
1"
0'
1(
0/
10
#120020000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#120030000000
0!
0'
0/
#120040000000
1!
1'
1/
#120050000000
0!
0'
0/
#120060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#120070000000
0!
0'
0/
#120080000000
1!
1'
1/
#120090000000
0!
1"
0'
1(
0/
10
#120100000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#120110000000
0!
1$
0'
1+
0/
#120120000000
1!
1'
1/
#120130000000
0!
0'
0/
#120140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#120150000000
0!
0'
0/
#120160000000
1!
1'
1/
#120170000000
0!
0'
0/
#120180000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#120190000000
0!
0'
0/
#120200000000
1!
1'
1/
#120210000000
0!
0'
0/
#120220000000
1!
1'
1/
#120230000000
0!
0'
0/
#120240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#120250000000
0!
0'
0/
#120260000000
1!
1'
1/
#120270000000
0!
0'
0/
#120280000000
1!
1'
1/
#120290000000
0!
0'
0/
#120300000000
1!
1'
1/
#120310000000
0!
0'
0/
#120320000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#120330000000
0!
0'
0/
#120340000000
1!
1'
1/
#120350000000
0!
0'
0/
#120360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#120370000000
0!
0'
0/
#120380000000
1!
1'
1/
#120390000000
0!
0'
0/
#120400000000
#120410000000
1!
1'
1/
#120420000000
0!
0'
0/
#120430000000
1!
1'
1/
#120440000000
0!
1"
0'
1(
0/
10
#120450000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#120460000000
0!
0'
0/
#120470000000
1!
1'
1/
#120480000000
0!
0'
0/
#120490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#120500000000
0!
0'
0/
#120510000000
1!
1'
1/
#120520000000
0!
1"
0'
1(
0/
10
#120530000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#120540000000
0!
1$
0'
1+
0/
#120550000000
1!
1'
1/
#120560000000
0!
0'
0/
#120570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#120580000000
0!
0'
0/
#120590000000
1!
1'
1/
#120600000000
0!
0'
0/
#120610000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#120620000000
0!
0'
0/
#120630000000
1!
1'
1/
#120640000000
0!
0'
0/
#120650000000
1!
1'
1/
#120660000000
0!
0'
0/
#120670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#120680000000
0!
0'
0/
#120690000000
1!
1'
1/
#120700000000
0!
0'
0/
#120710000000
1!
1'
1/
#120720000000
0!
0'
0/
#120730000000
1!
1'
1/
#120740000000
0!
0'
0/
#120750000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#120760000000
0!
0'
0/
#120770000000
1!
1'
1/
#120780000000
0!
0'
0/
#120790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#120800000000
0!
0'
0/
#120810000000
1!
1'
1/
#120820000000
0!
0'
0/
#120830000000
#120840000000
1!
1'
1/
#120850000000
0!
0'
0/
#120860000000
1!
1'
1/
#120870000000
0!
1"
0'
1(
0/
10
#120880000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#120890000000
0!
0'
0/
#120900000000
1!
1'
1/
#120910000000
0!
0'
0/
#120920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#120930000000
0!
0'
0/
#120940000000
1!
1'
1/
#120950000000
0!
1"
0'
1(
0/
10
#120960000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#120970000000
0!
1$
0'
1+
0/
#120980000000
1!
1'
1/
#120990000000
0!
0'
0/
#121000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#121010000000
0!
0'
0/
#121020000000
1!
1'
1/
#121030000000
0!
0'
0/
#121040000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#121050000000
0!
0'
0/
#121060000000
1!
1'
1/
#121070000000
0!
0'
0/
#121080000000
1!
1'
1/
#121090000000
0!
0'
0/
#121100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#121110000000
0!
0'
0/
#121120000000
1!
1'
1/
#121130000000
0!
0'
0/
#121140000000
1!
1'
1/
#121150000000
0!
0'
0/
#121160000000
1!
1'
1/
#121170000000
0!
0'
0/
#121180000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#121190000000
0!
0'
0/
#121200000000
1!
1'
1/
#121210000000
0!
0'
0/
#121220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#121230000000
0!
0'
0/
#121240000000
1!
1'
1/
#121250000000
0!
0'
0/
#121260000000
#121270000000
1!
1'
1/
#121280000000
0!
0'
0/
#121290000000
1!
1'
1/
#121300000000
0!
1"
0'
1(
0/
10
#121310000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#121320000000
0!
0'
0/
#121330000000
1!
1'
1/
#121340000000
0!
0'
0/
#121350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#121360000000
0!
0'
0/
#121370000000
1!
1'
1/
#121380000000
0!
1"
0'
1(
0/
10
#121390000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#121400000000
0!
1$
0'
1+
0/
#121410000000
1!
1'
1/
#121420000000
0!
0'
0/
#121430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#121440000000
0!
0'
0/
#121450000000
1!
1'
1/
#121460000000
0!
0'
0/
#121470000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#121480000000
0!
0'
0/
#121490000000
1!
1'
1/
#121500000000
0!
0'
0/
#121510000000
1!
1'
1/
#121520000000
0!
0'
0/
#121530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#121540000000
0!
0'
0/
#121550000000
1!
1'
1/
#121560000000
0!
0'
0/
#121570000000
1!
1'
1/
#121580000000
0!
0'
0/
#121590000000
1!
1'
1/
#121600000000
0!
0'
0/
#121610000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#121620000000
0!
0'
0/
#121630000000
1!
1'
1/
#121640000000
0!
0'
0/
#121650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#121660000000
0!
0'
0/
#121670000000
1!
1'
1/
#121680000000
0!
0'
0/
#121690000000
#121700000000
1!
1'
1/
#121710000000
0!
0'
0/
#121720000000
1!
1'
1/
#121730000000
0!
1"
0'
1(
0/
10
#121740000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#121750000000
0!
0'
0/
#121760000000
1!
1'
1/
#121770000000
0!
0'
0/
#121780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#121790000000
0!
0'
0/
#121800000000
1!
1'
1/
#121810000000
0!
1"
0'
1(
0/
10
#121820000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#121830000000
0!
1$
0'
1+
0/
#121840000000
1!
1'
1/
#121850000000
0!
0'
0/
#121860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#121870000000
0!
0'
0/
#121880000000
1!
1'
1/
#121890000000
0!
0'
0/
#121900000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#121910000000
0!
0'
0/
#121920000000
1!
1'
1/
#121930000000
0!
0'
0/
#121940000000
1!
1'
1/
#121950000000
0!
0'
0/
#121960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#121970000000
0!
0'
0/
#121980000000
1!
1'
1/
#121990000000
0!
0'
0/
#122000000000
1!
1'
1/
#122010000000
0!
0'
0/
#122020000000
1!
1'
1/
#122030000000
0!
0'
0/
#122040000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#122050000000
0!
0'
0/
#122060000000
1!
1'
1/
#122070000000
0!
0'
0/
#122080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#122090000000
0!
0'
0/
#122100000000
1!
1'
1/
#122110000000
0!
0'
0/
#122120000000
#122130000000
1!
1'
1/
#122140000000
0!
0'
0/
#122150000000
1!
1'
1/
#122160000000
0!
1"
0'
1(
0/
10
#122170000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#122180000000
0!
0'
0/
#122190000000
1!
1'
1/
#122200000000
0!
0'
0/
#122210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#122220000000
0!
0'
0/
#122230000000
1!
1'
1/
#122240000000
0!
1"
0'
1(
0/
10
#122250000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#122260000000
0!
1$
0'
1+
0/
#122270000000
1!
1'
1/
#122280000000
0!
0'
0/
#122290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#122300000000
0!
0'
0/
#122310000000
1!
1'
1/
#122320000000
0!
0'
0/
#122330000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#122340000000
0!
0'
0/
#122350000000
1!
1'
1/
#122360000000
0!
0'
0/
#122370000000
1!
1'
1/
#122380000000
0!
0'
0/
#122390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#122400000000
0!
0'
0/
#122410000000
1!
1'
1/
#122420000000
0!
0'
0/
#122430000000
1!
1'
1/
#122440000000
0!
0'
0/
#122450000000
1!
1'
1/
#122460000000
0!
0'
0/
#122470000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#122480000000
0!
0'
0/
#122490000000
1!
1'
1/
#122500000000
0!
0'
0/
#122510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#122520000000
0!
0'
0/
#122530000000
1!
1'
1/
#122540000000
0!
0'
0/
#122550000000
#122560000000
1!
1'
1/
#122570000000
0!
0'
0/
#122580000000
1!
1'
1/
#122590000000
0!
1"
0'
1(
0/
10
#122600000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#122610000000
0!
0'
0/
#122620000000
1!
1'
1/
#122630000000
0!
0'
0/
#122640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#122650000000
0!
0'
0/
#122660000000
1!
1'
1/
#122670000000
0!
1"
0'
1(
0/
10
#122680000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#122690000000
0!
1$
0'
1+
0/
#122700000000
1!
1'
1/
#122710000000
0!
0'
0/
#122720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#122730000000
0!
0'
0/
#122740000000
1!
1'
1/
#122750000000
0!
0'
0/
#122760000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#122770000000
0!
0'
0/
#122780000000
1!
1'
1/
#122790000000
0!
0'
0/
#122800000000
1!
1'
1/
#122810000000
0!
0'
0/
#122820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#122830000000
0!
0'
0/
#122840000000
1!
1'
1/
#122850000000
0!
0'
0/
#122860000000
1!
1'
1/
#122870000000
0!
0'
0/
#122880000000
1!
1'
1/
#122890000000
0!
0'
0/
#122900000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#122910000000
0!
0'
0/
#122920000000
1!
1'
1/
#122930000000
0!
0'
0/
#122940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#122950000000
0!
0'
0/
#122960000000
1!
1'
1/
#122970000000
0!
0'
0/
#122980000000
#122990000000
1!
1'
1/
#123000000000
0!
0'
0/
#123010000000
1!
1'
1/
#123020000000
0!
1"
0'
1(
0/
10
#123030000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#123040000000
0!
0'
0/
#123050000000
1!
1'
1/
#123060000000
0!
0'
0/
#123070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#123080000000
0!
0'
0/
#123090000000
1!
1'
1/
#123100000000
0!
1"
0'
1(
0/
10
#123110000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#123120000000
0!
1$
0'
1+
0/
#123130000000
1!
1'
1/
#123140000000
0!
0'
0/
#123150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#123160000000
0!
0'
0/
#123170000000
1!
1'
1/
#123180000000
0!
0'
0/
#123190000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#123200000000
0!
0'
0/
#123210000000
1!
1'
1/
#123220000000
0!
0'
0/
#123230000000
1!
1'
1/
#123240000000
0!
0'
0/
#123250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#123260000000
0!
0'
0/
#123270000000
1!
1'
1/
#123280000000
0!
0'
0/
#123290000000
1!
1'
1/
#123300000000
0!
0'
0/
#123310000000
1!
1'
1/
#123320000000
0!
0'
0/
#123330000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#123340000000
0!
0'
0/
#123350000000
1!
1'
1/
#123360000000
0!
0'
0/
#123370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#123380000000
0!
0'
0/
#123390000000
1!
1'
1/
#123400000000
0!
0'
0/
#123410000000
#123420000000
1!
1'
1/
#123430000000
0!
0'
0/
#123440000000
1!
1'
1/
#123450000000
0!
1"
0'
1(
0/
10
#123460000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#123470000000
0!
0'
0/
#123480000000
1!
1'
1/
#123490000000
0!
0'
0/
#123500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#123510000000
0!
0'
0/
#123520000000
1!
1'
1/
#123530000000
0!
1"
0'
1(
0/
10
#123540000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#123550000000
0!
1$
0'
1+
0/
#123560000000
1!
1'
1/
#123570000000
0!
0'
0/
#123580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#123590000000
0!
0'
0/
#123600000000
1!
1'
1/
#123610000000
0!
0'
0/
#123620000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#123630000000
0!
0'
0/
#123640000000
1!
1'
1/
#123650000000
0!
0'
0/
#123660000000
1!
1'
1/
#123670000000
0!
0'
0/
#123680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#123690000000
0!
0'
0/
#123700000000
1!
1'
1/
#123710000000
0!
0'
0/
#123720000000
1!
1'
1/
#123730000000
0!
0'
0/
#123740000000
1!
1'
1/
#123750000000
0!
0'
0/
#123760000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#123770000000
0!
0'
0/
#123780000000
1!
1'
1/
#123790000000
0!
0'
0/
#123800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#123810000000
0!
0'
0/
#123820000000
1!
1'
1/
#123830000000
0!
0'
0/
#123840000000
#123850000000
1!
1'
1/
#123860000000
0!
0'
0/
#123870000000
1!
1'
1/
#123880000000
0!
1"
0'
1(
0/
10
#123890000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#123900000000
0!
0'
0/
#123910000000
1!
1'
1/
#123920000000
0!
0'
0/
#123930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#123940000000
0!
0'
0/
#123950000000
1!
1'
1/
#123960000000
0!
1"
0'
1(
0/
10
#123970000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#123980000000
0!
1$
0'
1+
0/
#123990000000
1!
1'
1/
#124000000000
0!
0'
0/
#124010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#124020000000
0!
0'
0/
#124030000000
1!
1'
1/
#124040000000
0!
0'
0/
#124050000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#124060000000
0!
0'
0/
#124070000000
1!
1'
1/
#124080000000
0!
0'
0/
#124090000000
1!
1'
1/
#124100000000
0!
0'
0/
#124110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#124120000000
0!
0'
0/
#124130000000
1!
1'
1/
#124140000000
0!
0'
0/
#124150000000
1!
1'
1/
#124160000000
0!
0'
0/
#124170000000
1!
1'
1/
#124180000000
0!
0'
0/
#124190000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#124200000000
0!
0'
0/
#124210000000
1!
1'
1/
#124220000000
0!
0'
0/
#124230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#124240000000
0!
0'
0/
#124250000000
1!
1'
1/
#124260000000
0!
0'
0/
#124270000000
#124280000000
1!
1'
1/
#124290000000
0!
0'
0/
#124300000000
1!
1'
1/
#124310000000
0!
1"
0'
1(
0/
10
#124320000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#124330000000
0!
0'
0/
#124340000000
1!
1'
1/
#124350000000
0!
0'
0/
#124360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#124370000000
0!
0'
0/
#124380000000
1!
1'
1/
#124390000000
0!
1"
0'
1(
0/
10
#124400000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#124410000000
0!
1$
0'
1+
0/
#124420000000
1!
1'
1/
#124430000000
0!
0'
0/
#124440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#124450000000
0!
0'
0/
#124460000000
1!
1'
1/
#124470000000
0!
0'
0/
#124480000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#124490000000
0!
0'
0/
#124500000000
1!
1'
1/
#124510000000
0!
0'
0/
#124520000000
1!
1'
1/
#124530000000
0!
0'
0/
#124540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#124550000000
0!
0'
0/
#124560000000
1!
1'
1/
#124570000000
0!
0'
0/
#124580000000
1!
1'
1/
#124590000000
0!
0'
0/
#124600000000
1!
1'
1/
#124610000000
0!
0'
0/
#124620000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#124630000000
0!
0'
0/
#124640000000
1!
1'
1/
#124650000000
0!
0'
0/
#124660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#124670000000
0!
0'
0/
#124680000000
1!
1'
1/
#124690000000
0!
0'
0/
#124700000000
#124710000000
1!
1'
1/
#124720000000
0!
0'
0/
#124730000000
1!
1'
1/
#124740000000
0!
1"
0'
1(
0/
10
#124750000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#124760000000
0!
0'
0/
#124770000000
1!
1'
1/
#124780000000
0!
0'
0/
#124790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#124800000000
0!
0'
0/
#124810000000
1!
1'
1/
#124820000000
0!
1"
0'
1(
0/
10
#124830000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#124840000000
0!
1$
0'
1+
0/
#124850000000
1!
1'
1/
#124860000000
0!
0'
0/
#124870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#124880000000
0!
0'
0/
#124890000000
1!
1'
1/
#124900000000
0!
0'
0/
#124910000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#124920000000
0!
0'
0/
#124930000000
1!
1'
1/
#124940000000
0!
0'
0/
#124950000000
1!
1'
1/
#124960000000
0!
0'
0/
#124970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#124980000000
0!
0'
0/
#124990000000
1!
1'
1/
#125000000000
0!
0'
0/
#125010000000
1!
1'
1/
#125020000000
0!
0'
0/
#125030000000
1!
1'
1/
#125040000000
0!
0'
0/
#125050000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#125060000000
0!
0'
0/
#125070000000
1!
1'
1/
#125080000000
0!
0'
0/
#125090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#125100000000
0!
0'
0/
#125110000000
1!
1'
1/
#125120000000
0!
0'
0/
#125130000000
#125140000000
1!
1'
1/
#125150000000
0!
0'
0/
#125160000000
1!
1'
1/
#125170000000
0!
1"
0'
1(
0/
10
#125180000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#125190000000
0!
0'
0/
#125200000000
1!
1'
1/
#125210000000
0!
0'
0/
#125220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#125230000000
0!
0'
0/
#125240000000
1!
1'
1/
#125250000000
0!
1"
0'
1(
0/
10
#125260000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#125270000000
0!
1$
0'
1+
0/
#125280000000
1!
1'
1/
#125290000000
0!
0'
0/
#125300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#125310000000
0!
0'
0/
#125320000000
1!
1'
1/
#125330000000
0!
0'
0/
#125340000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#125350000000
0!
0'
0/
#125360000000
1!
1'
1/
#125370000000
0!
0'
0/
#125380000000
1!
1'
1/
#125390000000
0!
0'
0/
#125400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#125410000000
0!
0'
0/
#125420000000
1!
1'
1/
#125430000000
0!
0'
0/
#125440000000
1!
1'
1/
#125450000000
0!
0'
0/
#125460000000
1!
1'
1/
#125470000000
0!
0'
0/
#125480000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#125490000000
0!
0'
0/
#125500000000
1!
1'
1/
#125510000000
0!
0'
0/
#125520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#125530000000
0!
0'
0/
#125540000000
1!
1'
1/
#125550000000
0!
0'
0/
#125560000000
#125570000000
1!
1'
1/
#125580000000
0!
0'
0/
#125590000000
1!
1'
1/
#125600000000
0!
1"
0'
1(
0/
10
#125610000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#125620000000
0!
0'
0/
#125630000000
1!
1'
1/
#125640000000
0!
0'
0/
#125650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#125660000000
0!
0'
0/
#125670000000
1!
1'
1/
#125680000000
0!
1"
0'
1(
0/
10
#125690000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#125700000000
0!
1$
0'
1+
0/
#125710000000
1!
1'
1/
#125720000000
0!
0'
0/
#125730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#125740000000
0!
0'
0/
#125750000000
1!
1'
1/
#125760000000
0!
0'
0/
#125770000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#125780000000
0!
0'
0/
#125790000000
1!
1'
1/
#125800000000
0!
0'
0/
#125810000000
1!
1'
1/
#125820000000
0!
0'
0/
#125830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#125840000000
0!
0'
0/
#125850000000
1!
1'
1/
#125860000000
0!
0'
0/
#125870000000
1!
1'
1/
#125880000000
0!
0'
0/
#125890000000
1!
1'
1/
#125900000000
0!
0'
0/
#125910000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#125920000000
0!
0'
0/
#125930000000
1!
1'
1/
#125940000000
0!
0'
0/
#125950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#125960000000
0!
0'
0/
#125970000000
1!
1'
1/
#125980000000
0!
0'
0/
#125990000000
#126000000000
1!
1'
1/
#126010000000
0!
0'
0/
#126020000000
1!
1'
1/
#126030000000
0!
1"
0'
1(
0/
10
#126040000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#126050000000
0!
0'
0/
#126060000000
1!
1'
1/
#126070000000
0!
0'
0/
#126080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#126090000000
0!
0'
0/
#126100000000
1!
1'
1/
#126110000000
0!
1"
0'
1(
0/
10
#126120000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#126130000000
0!
1$
0'
1+
0/
#126140000000
1!
1'
1/
#126150000000
0!
0'
0/
#126160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#126170000000
0!
0'
0/
#126180000000
1!
1'
1/
#126190000000
0!
0'
0/
#126200000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#126210000000
0!
0'
0/
#126220000000
1!
1'
1/
#126230000000
0!
0'
0/
#126240000000
1!
1'
1/
#126250000000
0!
0'
0/
#126260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#126270000000
0!
0'
0/
#126280000000
1!
1'
1/
#126290000000
0!
0'
0/
#126300000000
1!
1'
1/
#126310000000
0!
0'
0/
#126320000000
1!
1'
1/
#126330000000
0!
0'
0/
#126340000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#126350000000
0!
0'
0/
#126360000000
1!
1'
1/
#126370000000
0!
0'
0/
#126380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#126390000000
0!
0'
0/
#126400000000
1!
1'
1/
#126410000000
0!
0'
0/
#126420000000
#126430000000
1!
1'
1/
#126440000000
0!
0'
0/
#126450000000
1!
1'
1/
#126460000000
0!
1"
0'
1(
0/
10
#126470000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#126480000000
0!
0'
0/
#126490000000
1!
1'
1/
#126500000000
0!
0'
0/
#126510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#126520000000
0!
0'
0/
#126530000000
1!
1'
1/
#126540000000
0!
1"
0'
1(
0/
10
#126550000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#126560000000
0!
1$
0'
1+
0/
#126570000000
1!
1'
1/
#126580000000
0!
0'
0/
#126590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#126600000000
0!
0'
0/
#126610000000
1!
1'
1/
#126620000000
0!
0'
0/
#126630000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#126640000000
0!
0'
0/
#126650000000
1!
1'
1/
#126660000000
0!
0'
0/
#126670000000
1!
1'
1/
#126680000000
0!
0'
0/
#126690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#126700000000
0!
0'
0/
#126710000000
1!
1'
1/
#126720000000
0!
0'
0/
#126730000000
1!
1'
1/
#126740000000
0!
0'
0/
#126750000000
1!
1'
1/
#126760000000
0!
0'
0/
#126770000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#126780000000
0!
0'
0/
#126790000000
1!
1'
1/
#126800000000
0!
0'
0/
#126810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#126820000000
0!
0'
0/
#126830000000
1!
1'
1/
#126840000000
0!
0'
0/
#126850000000
#126860000000
1!
1'
1/
#126870000000
0!
0'
0/
#126880000000
1!
1'
1/
#126890000000
0!
1"
0'
1(
0/
10
#126900000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#126910000000
0!
0'
0/
#126920000000
1!
1'
1/
#126930000000
0!
0'
0/
#126940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#126950000000
0!
0'
0/
#126960000000
1!
1'
1/
#126970000000
0!
1"
0'
1(
0/
10
#126980000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#126990000000
0!
1$
0'
1+
0/
#127000000000
1!
1'
1/
#127010000000
0!
0'
0/
#127020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#127030000000
0!
0'
0/
#127040000000
1!
1'
1/
#127050000000
0!
0'
0/
#127060000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#127070000000
0!
0'
0/
#127080000000
1!
1'
1/
#127090000000
0!
0'
0/
#127100000000
1!
1'
1/
#127110000000
0!
0'
0/
#127120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#127130000000
0!
0'
0/
#127140000000
1!
1'
1/
#127150000000
0!
0'
0/
#127160000000
1!
1'
1/
#127170000000
0!
0'
0/
#127180000000
1!
1'
1/
#127190000000
0!
0'
0/
#127200000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#127210000000
0!
0'
0/
#127220000000
1!
1'
1/
#127230000000
0!
0'
0/
#127240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#127250000000
0!
0'
0/
#127260000000
1!
1'
1/
#127270000000
0!
0'
0/
#127280000000
#127290000000
1!
1'
1/
#127300000000
0!
0'
0/
#127310000000
1!
1'
1/
#127320000000
0!
1"
0'
1(
0/
10
#127330000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#127340000000
0!
0'
0/
#127350000000
1!
1'
1/
#127360000000
0!
0'
0/
#127370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#127380000000
0!
0'
0/
#127390000000
1!
1'
1/
#127400000000
0!
1"
0'
1(
0/
10
#127410000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#127420000000
0!
1$
0'
1+
0/
#127430000000
1!
1'
1/
#127440000000
0!
0'
0/
#127450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#127460000000
0!
0'
0/
#127470000000
1!
1'
1/
#127480000000
0!
0'
0/
#127490000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#127500000000
0!
0'
0/
#127510000000
1!
1'
1/
#127520000000
0!
0'
0/
#127530000000
1!
1'
1/
#127540000000
0!
0'
0/
#127550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#127560000000
0!
0'
0/
#127570000000
1!
1'
1/
#127580000000
0!
0'
0/
#127590000000
1!
1'
1/
#127600000000
0!
0'
0/
#127610000000
1!
1'
1/
#127620000000
0!
0'
0/
#127630000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#127640000000
0!
0'
0/
#127650000000
1!
1'
1/
#127660000000
0!
0'
0/
#127670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#127680000000
0!
0'
0/
#127690000000
1!
1'
1/
#127700000000
0!
0'
0/
#127710000000
#127720000000
1!
1'
1/
#127730000000
0!
0'
0/
#127740000000
1!
1'
1/
#127750000000
0!
1"
0'
1(
0/
10
#127760000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#127770000000
0!
0'
0/
#127780000000
1!
1'
1/
#127790000000
0!
0'
0/
#127800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#127810000000
0!
0'
0/
#127820000000
1!
1'
1/
#127830000000
0!
1"
0'
1(
0/
10
#127840000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#127850000000
0!
1$
0'
1+
0/
#127860000000
1!
1'
1/
#127870000000
0!
0'
0/
#127880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#127890000000
0!
0'
0/
#127900000000
1!
1'
1/
#127910000000
0!
0'
0/
#127920000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#127930000000
0!
0'
0/
#127940000000
1!
1'
1/
#127950000000
0!
0'
0/
#127960000000
1!
1'
1/
#127970000000
0!
0'
0/
#127980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#127990000000
0!
0'
0/
#128000000000
1!
1'
1/
#128010000000
0!
0'
0/
#128020000000
1!
1'
1/
#128030000000
0!
0'
0/
#128040000000
1!
1'
1/
#128050000000
0!
0'
0/
#128060000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#128070000000
0!
0'
0/
#128080000000
1!
1'
1/
#128090000000
0!
0'
0/
#128100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#128110000000
0!
0'
0/
#128120000000
1!
1'
1/
#128130000000
0!
0'
0/
#128140000000
#128150000000
1!
1'
1/
#128160000000
0!
0'
0/
#128170000000
1!
1'
1/
#128180000000
0!
1"
0'
1(
0/
10
#128190000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#128200000000
0!
0'
0/
#128210000000
1!
1'
1/
#128220000000
0!
0'
0/
#128230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#128240000000
0!
0'
0/
#128250000000
1!
1'
1/
#128260000000
0!
1"
0'
1(
0/
10
#128270000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#128280000000
0!
1$
0'
1+
0/
#128290000000
1!
1'
1/
#128300000000
0!
0'
0/
#128310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#128320000000
0!
0'
0/
#128330000000
1!
1'
1/
#128340000000
0!
0'
0/
#128350000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#128360000000
0!
0'
0/
#128370000000
1!
1'
1/
#128380000000
0!
0'
0/
#128390000000
1!
1'
1/
#128400000000
0!
0'
0/
#128410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#128420000000
0!
0'
0/
#128430000000
1!
1'
1/
#128440000000
0!
0'
0/
#128450000000
1!
1'
1/
#128460000000
0!
0'
0/
#128470000000
1!
1'
1/
#128480000000
0!
0'
0/
#128490000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#128500000000
0!
0'
0/
#128510000000
1!
1'
1/
#128520000000
0!
0'
0/
#128530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#128540000000
0!
0'
0/
#128550000000
1!
1'
1/
#128560000000
0!
0'
0/
#128570000000
#128580000000
1!
1'
1/
#128590000000
0!
0'
0/
#128600000000
1!
1'
1/
#128610000000
0!
1"
0'
1(
0/
10
#128620000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#128630000000
0!
0'
0/
#128640000000
1!
1'
1/
#128650000000
0!
0'
0/
#128660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#128670000000
0!
0'
0/
#128680000000
1!
1'
1/
#128690000000
0!
1"
0'
1(
0/
10
#128700000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#128710000000
0!
1$
0'
1+
0/
#128720000000
1!
1'
1/
#128730000000
0!
0'
0/
#128740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#128750000000
0!
0'
0/
#128760000000
1!
1'
1/
#128770000000
0!
0'
0/
#128780000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#128790000000
0!
0'
0/
#128800000000
1!
1'
1/
#128810000000
0!
0'
0/
#128820000000
1!
1'
1/
#128830000000
0!
0'
0/
#128840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#128850000000
0!
0'
0/
#128860000000
1!
1'
1/
#128870000000
0!
0'
0/
#128880000000
1!
1'
1/
#128890000000
0!
0'
0/
#128900000000
1!
1'
1/
#128910000000
0!
0'
0/
#128920000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#128930000000
0!
0'
0/
#128940000000
1!
1'
1/
#128950000000
0!
0'
0/
#128960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#128970000000
0!
0'
0/
#128980000000
1!
1'
1/
#128990000000
0!
0'
0/
#129000000000
#129010000000
1!
1'
1/
#129020000000
0!
0'
0/
#129030000000
1!
1'
1/
#129040000000
0!
1"
0'
1(
0/
10
#129050000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#129060000000
0!
0'
0/
#129070000000
1!
1'
1/
#129080000000
0!
0'
0/
#129090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#129100000000
0!
0'
0/
#129110000000
1!
1'
1/
#129120000000
0!
1"
0'
1(
0/
10
#129130000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#129140000000
0!
1$
0'
1+
0/
#129150000000
1!
1'
1/
#129160000000
0!
0'
0/
#129170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#129180000000
0!
0'
0/
#129190000000
1!
1'
1/
#129200000000
0!
0'
0/
#129210000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#129220000000
0!
0'
0/
#129230000000
1!
1'
1/
#129240000000
0!
0'
0/
#129250000000
1!
1'
1/
#129260000000
0!
0'
0/
#129270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#129280000000
0!
0'
0/
#129290000000
1!
1'
1/
#129300000000
0!
0'
0/
#129310000000
1!
1'
1/
#129320000000
0!
0'
0/
#129330000000
1!
1'
1/
#129340000000
0!
0'
0/
#129350000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#129360000000
0!
0'
0/
#129370000000
1!
1'
1/
#129380000000
0!
0'
0/
#129390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#129400000000
0!
0'
0/
#129410000000
1!
1'
1/
#129420000000
0!
0'
0/
#129430000000
#129440000000
1!
1'
1/
#129450000000
0!
0'
0/
#129460000000
1!
1'
1/
#129470000000
0!
1"
0'
1(
0/
10
#129480000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#129490000000
0!
0'
0/
#129500000000
1!
1'
1/
#129510000000
0!
0'
0/
#129520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#129530000000
0!
0'
0/
#129540000000
1!
1'
1/
#129550000000
0!
1"
0'
1(
0/
10
#129560000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#129570000000
0!
1$
0'
1+
0/
#129580000000
1!
1'
1/
#129590000000
0!
0'
0/
#129600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#129610000000
0!
0'
0/
#129620000000
1!
1'
1/
#129630000000
0!
0'
0/
#129640000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#129650000000
0!
0'
0/
#129660000000
1!
1'
1/
#129670000000
0!
0'
0/
#129680000000
1!
1'
1/
#129690000000
0!
0'
0/
#129700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#129710000000
0!
0'
0/
#129720000000
1!
1'
1/
#129730000000
0!
0'
0/
#129740000000
1!
1'
1/
#129750000000
0!
0'
0/
#129760000000
1!
1'
1/
#129770000000
0!
0'
0/
#129780000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#129790000000
0!
0'
0/
#129800000000
1!
1'
1/
#129810000000
0!
0'
0/
#129820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#129830000000
0!
0'
0/
#129840000000
1!
1'
1/
#129850000000
0!
0'
0/
#129860000000
#129870000000
1!
1'
1/
#129880000000
0!
0'
0/
#129890000000
1!
1'
1/
#129900000000
0!
1"
0'
1(
0/
10
#129910000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#129920000000
0!
0'
0/
#129930000000
1!
1'
1/
#129940000000
0!
0'
0/
#129950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#129960000000
0!
0'
0/
#129970000000
1!
1'
1/
#129980000000
0!
1"
0'
1(
0/
10
#129990000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#130000000000
0!
1$
0'
1+
0/
#130010000000
1!
1'
1/
#130020000000
0!
0'
0/
#130030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#130040000000
0!
0'
0/
#130050000000
1!
1'
1/
#130060000000
0!
0'
0/
#130070000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#130080000000
0!
0'
0/
#130090000000
1!
1'
1/
#130100000000
0!
0'
0/
#130110000000
1!
1'
1/
#130120000000
0!
0'
0/
#130130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#130140000000
0!
0'
0/
#130150000000
1!
1'
1/
#130160000000
0!
0'
0/
#130170000000
1!
1'
1/
#130180000000
0!
0'
0/
#130190000000
1!
1'
1/
#130200000000
0!
0'
0/
#130210000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#130220000000
0!
0'
0/
#130230000000
1!
1'
1/
#130240000000
0!
0'
0/
#130250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#130260000000
0!
0'
0/
#130270000000
1!
1'
1/
#130280000000
0!
0'
0/
#130290000000
#130300000000
1!
1'
1/
#130310000000
0!
0'
0/
#130320000000
1!
1'
1/
#130330000000
0!
1"
0'
1(
0/
10
#130340000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#130350000000
0!
0'
0/
#130360000000
1!
1'
1/
#130370000000
0!
0'
0/
#130380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#130390000000
0!
0'
0/
#130400000000
1!
1'
1/
#130410000000
0!
1"
0'
1(
0/
10
#130420000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#130430000000
0!
1$
0'
1+
0/
#130440000000
1!
1'
1/
#130450000000
0!
0'
0/
#130460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#130470000000
0!
0'
0/
#130480000000
1!
1'
1/
#130490000000
0!
0'
0/
#130500000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#130510000000
0!
0'
0/
#130520000000
1!
1'
1/
#130530000000
0!
0'
0/
#130540000000
1!
1'
1/
#130550000000
0!
0'
0/
#130560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#130570000000
0!
0'
0/
#130580000000
1!
1'
1/
#130590000000
0!
0'
0/
#130600000000
1!
1'
1/
#130610000000
0!
0'
0/
#130620000000
1!
1'
1/
#130630000000
0!
0'
0/
#130640000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#130650000000
0!
0'
0/
#130660000000
1!
1'
1/
#130670000000
0!
0'
0/
#130680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#130690000000
0!
0'
0/
#130700000000
1!
1'
1/
#130710000000
0!
0'
0/
#130720000000
#130730000000
1!
1'
1/
#130740000000
0!
0'
0/
#130750000000
1!
1'
1/
#130760000000
0!
1"
0'
1(
0/
10
#130770000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#130780000000
0!
0'
0/
#130790000000
1!
1'
1/
#130800000000
0!
0'
0/
#130810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#130820000000
0!
0'
0/
#130830000000
1!
1'
1/
#130840000000
0!
1"
0'
1(
0/
10
#130850000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#130860000000
0!
1$
0'
1+
0/
#130870000000
1!
1'
1/
#130880000000
0!
0'
0/
#130890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#130900000000
0!
0'
0/
#130910000000
1!
1'
1/
#130920000000
0!
0'
0/
#130930000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#130940000000
0!
0'
0/
#130950000000
1!
1'
1/
#130960000000
0!
0'
0/
#130970000000
1!
1'
1/
#130980000000
0!
0'
0/
#130990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#131000000000
0!
0'
0/
#131010000000
1!
1'
1/
#131020000000
0!
0'
0/
#131030000000
1!
1'
1/
#131040000000
0!
0'
0/
#131050000000
1!
1'
1/
#131060000000
0!
0'
0/
#131070000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#131080000000
0!
0'
0/
#131090000000
1!
1'
1/
#131100000000
0!
0'
0/
#131110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#131120000000
0!
0'
0/
#131130000000
1!
1'
1/
#131140000000
0!
0'
0/
#131150000000
#131160000000
1!
1'
1/
#131170000000
0!
0'
0/
#131180000000
1!
1'
1/
#131190000000
0!
1"
0'
1(
0/
10
#131200000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#131210000000
0!
0'
0/
#131220000000
1!
1'
1/
#131230000000
0!
0'
0/
#131240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#131250000000
0!
0'
0/
#131260000000
1!
1'
1/
#131270000000
0!
1"
0'
1(
0/
10
#131280000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#131290000000
0!
1$
0'
1+
0/
#131300000000
1!
1'
1/
#131310000000
0!
0'
0/
#131320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#131330000000
0!
0'
0/
#131340000000
1!
1'
1/
#131350000000
0!
0'
0/
#131360000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#131370000000
0!
0'
0/
#131380000000
1!
1'
1/
#131390000000
0!
0'
0/
#131400000000
1!
1'
1/
#131410000000
0!
0'
0/
#131420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#131430000000
0!
0'
0/
#131440000000
1!
1'
1/
#131450000000
0!
0'
0/
#131460000000
1!
1'
1/
#131470000000
0!
0'
0/
#131480000000
1!
1'
1/
#131490000000
0!
0'
0/
#131500000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#131510000000
0!
0'
0/
#131520000000
1!
1'
1/
#131530000000
0!
0'
0/
#131540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#131550000000
0!
0'
0/
#131560000000
1!
1'
1/
#131570000000
0!
0'
0/
#131580000000
#131590000000
1!
1'
1/
#131600000000
0!
0'
0/
#131610000000
1!
1'
1/
#131620000000
0!
1"
0'
1(
0/
10
#131630000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#131640000000
0!
0'
0/
#131650000000
1!
1'
1/
#131660000000
0!
0'
0/
#131670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#131680000000
0!
0'
0/
#131690000000
1!
1'
1/
#131700000000
0!
1"
0'
1(
0/
10
#131710000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#131720000000
0!
1$
0'
1+
0/
#131730000000
1!
1'
1/
#131740000000
0!
0'
0/
#131750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#131760000000
0!
0'
0/
#131770000000
1!
1'
1/
#131780000000
0!
0'
0/
#131790000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#131800000000
0!
0'
0/
#131810000000
1!
1'
1/
#131820000000
0!
0'
0/
#131830000000
1!
1'
1/
#131840000000
0!
0'
0/
#131850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#131860000000
0!
0'
0/
#131870000000
1!
1'
1/
#131880000000
0!
0'
0/
#131890000000
1!
1'
1/
#131900000000
0!
0'
0/
#131910000000
1!
1'
1/
#131920000000
0!
0'
0/
#131930000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#131940000000
0!
0'
0/
#131950000000
1!
1'
1/
#131960000000
0!
0'
0/
#131970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#131980000000
0!
0'
0/
#131990000000
1!
1'
1/
#132000000000
0!
0'
0/
#132010000000
#132020000000
1!
1'
1/
#132030000000
0!
0'
0/
#132040000000
1!
1'
1/
#132050000000
0!
1"
0'
1(
0/
10
#132060000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#132070000000
0!
0'
0/
#132080000000
1!
1'
1/
#132090000000
0!
0'
0/
#132100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#132110000000
0!
0'
0/
#132120000000
1!
1'
1/
#132130000000
0!
1"
0'
1(
0/
10
#132140000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#132150000000
0!
1$
0'
1+
0/
#132160000000
1!
1'
1/
#132170000000
0!
0'
0/
#132180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#132190000000
0!
0'
0/
#132200000000
1!
1'
1/
#132210000000
0!
0'
0/
#132220000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#132230000000
0!
0'
0/
#132240000000
1!
1'
1/
#132250000000
0!
0'
0/
#132260000000
1!
1'
1/
#132270000000
0!
0'
0/
#132280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#132290000000
0!
0'
0/
#132300000000
1!
1'
1/
#132310000000
0!
0'
0/
#132320000000
1!
1'
1/
#132330000000
0!
0'
0/
#132340000000
1!
1'
1/
#132350000000
0!
0'
0/
#132360000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#132370000000
0!
0'
0/
#132380000000
1!
1'
1/
#132390000000
0!
0'
0/
#132400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#132410000000
0!
0'
0/
#132420000000
1!
1'
1/
#132430000000
0!
0'
0/
#132440000000
#132450000000
1!
1'
1/
#132460000000
0!
0'
0/
#132470000000
1!
1'
1/
#132480000000
0!
1"
0'
1(
0/
10
#132490000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#132500000000
0!
0'
0/
#132510000000
1!
1'
1/
#132520000000
0!
0'
0/
#132530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#132540000000
0!
0'
0/
#132550000000
1!
1'
1/
#132560000000
0!
1"
0'
1(
0/
10
#132570000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#132580000000
0!
1$
0'
1+
0/
#132590000000
1!
1'
1/
#132600000000
0!
0'
0/
#132610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#132620000000
0!
0'
0/
#132630000000
1!
1'
1/
#132640000000
0!
0'
0/
#132650000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#132660000000
0!
0'
0/
#132670000000
1!
1'
1/
#132680000000
0!
0'
0/
#132690000000
1!
1'
1/
#132700000000
0!
0'
0/
#132710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#132720000000
0!
0'
0/
#132730000000
1!
1'
1/
#132740000000
0!
0'
0/
#132750000000
1!
1'
1/
#132760000000
0!
0'
0/
#132770000000
1!
1'
1/
#132780000000
0!
0'
0/
#132790000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#132800000000
0!
0'
0/
#132810000000
1!
1'
1/
#132820000000
0!
0'
0/
#132830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#132840000000
0!
0'
0/
#132850000000
1!
1'
1/
#132860000000
0!
0'
0/
#132870000000
#132880000000
1!
1'
1/
#132890000000
0!
0'
0/
#132900000000
1!
1'
1/
#132910000000
0!
1"
0'
1(
0/
10
#132920000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#132930000000
0!
0'
0/
#132940000000
1!
1'
1/
#132950000000
0!
0'
0/
#132960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#132970000000
0!
0'
0/
#132980000000
1!
1'
1/
#132990000000
0!
1"
0'
1(
0/
10
#133000000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#133010000000
0!
1$
0'
1+
0/
#133020000000
1!
1'
1/
#133030000000
0!
0'
0/
#133040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#133050000000
0!
0'
0/
#133060000000
1!
1'
1/
#133070000000
0!
0'
0/
#133080000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#133090000000
0!
0'
0/
#133100000000
1!
1'
1/
#133110000000
0!
0'
0/
#133120000000
1!
1'
1/
#133130000000
0!
0'
0/
#133140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#133150000000
0!
0'
0/
#133160000000
1!
1'
1/
#133170000000
0!
0'
0/
#133180000000
1!
1'
1/
#133190000000
0!
0'
0/
#133200000000
1!
1'
1/
#133210000000
0!
0'
0/
#133220000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#133230000000
0!
0'
0/
#133240000000
1!
1'
1/
#133250000000
0!
0'
0/
#133260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#133270000000
0!
0'
0/
#133280000000
1!
1'
1/
#133290000000
0!
0'
0/
#133300000000
#133310000000
1!
1'
1/
#133320000000
0!
0'
0/
#133330000000
1!
1'
1/
#133340000000
0!
1"
0'
1(
0/
10
#133350000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#133360000000
0!
0'
0/
#133370000000
1!
1'
1/
#133380000000
0!
0'
0/
#133390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#133400000000
0!
0'
0/
#133410000000
1!
1'
1/
#133420000000
0!
1"
0'
1(
0/
10
#133430000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#133440000000
0!
1$
0'
1+
0/
#133450000000
1!
1'
1/
#133460000000
0!
0'
0/
#133470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#133480000000
0!
0'
0/
#133490000000
1!
1'
1/
#133500000000
0!
0'
0/
#133510000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#133520000000
0!
0'
0/
#133530000000
1!
1'
1/
#133540000000
0!
0'
0/
#133550000000
1!
1'
1/
#133560000000
0!
0'
0/
#133570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#133580000000
0!
0'
0/
#133590000000
1!
1'
1/
#133600000000
0!
0'
0/
#133610000000
1!
1'
1/
#133620000000
0!
0'
0/
#133630000000
1!
1'
1/
#133640000000
0!
0'
0/
#133650000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#133660000000
0!
0'
0/
#133670000000
1!
1'
1/
#133680000000
0!
0'
0/
#133690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#133700000000
0!
0'
0/
#133710000000
1!
1'
1/
#133720000000
0!
0'
0/
#133730000000
#133740000000
1!
1'
1/
#133750000000
0!
0'
0/
#133760000000
1!
1'
1/
#133770000000
0!
1"
0'
1(
0/
10
#133780000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#133790000000
0!
0'
0/
#133800000000
1!
1'
1/
#133810000000
0!
0'
0/
#133820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#133830000000
0!
0'
0/
#133840000000
1!
1'
1/
#133850000000
0!
1"
0'
1(
0/
10
#133860000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#133870000000
0!
1$
0'
1+
0/
#133880000000
1!
1'
1/
#133890000000
0!
0'
0/
#133900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#133910000000
0!
0'
0/
#133920000000
1!
1'
1/
#133930000000
0!
0'
0/
#133940000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#133950000000
0!
0'
0/
#133960000000
1!
1'
1/
#133970000000
0!
0'
0/
#133980000000
1!
1'
1/
#133990000000
0!
0'
0/
#134000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#134010000000
0!
0'
0/
#134020000000
1!
1'
1/
#134030000000
0!
0'
0/
#134040000000
1!
1'
1/
#134050000000
0!
0'
0/
#134060000000
1!
1'
1/
#134070000000
0!
0'
0/
#134080000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#134090000000
0!
0'
0/
#134100000000
1!
1'
1/
#134110000000
0!
0'
0/
#134120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#134130000000
0!
0'
0/
#134140000000
1!
1'
1/
#134150000000
0!
0'
0/
#134160000000
#134170000000
1!
1'
1/
#134180000000
0!
0'
0/
#134190000000
1!
1'
1/
#134200000000
0!
1"
0'
1(
0/
10
#134210000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#134220000000
0!
0'
0/
#134230000000
1!
1'
1/
#134240000000
0!
0'
0/
#134250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#134260000000
0!
0'
0/
#134270000000
1!
1'
1/
#134280000000
0!
1"
0'
1(
0/
10
#134290000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#134300000000
0!
1$
0'
1+
0/
#134310000000
1!
1'
1/
#134320000000
0!
0'
0/
#134330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#134340000000
0!
0'
0/
#134350000000
1!
1'
1/
#134360000000
0!
0'
0/
#134370000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#134380000000
0!
0'
0/
#134390000000
1!
1'
1/
#134400000000
0!
0'
0/
#134410000000
1!
1'
1/
#134420000000
0!
0'
0/
#134430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#134440000000
0!
0'
0/
#134450000000
1!
1'
1/
#134460000000
0!
0'
0/
#134470000000
1!
1'
1/
#134480000000
0!
0'
0/
#134490000000
1!
1'
1/
#134500000000
0!
0'
0/
#134510000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#134520000000
0!
0'
0/
#134530000000
1!
1'
1/
#134540000000
0!
0'
0/
#134550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#134560000000
0!
0'
0/
#134570000000
1!
1'
1/
#134580000000
0!
0'
0/
#134590000000
#134600000000
1!
1'
1/
#134610000000
0!
0'
0/
#134620000000
1!
1'
1/
#134630000000
0!
1"
0'
1(
0/
10
#134640000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#134650000000
0!
0'
0/
#134660000000
1!
1'
1/
#134670000000
0!
0'
0/
#134680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#134690000000
0!
0'
0/
#134700000000
1!
1'
1/
#134710000000
0!
1"
0'
1(
0/
10
#134720000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#134730000000
0!
1$
0'
1+
0/
#134740000000
1!
1'
1/
#134750000000
0!
0'
0/
#134760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#134770000000
0!
0'
0/
#134780000000
1!
1'
1/
#134790000000
0!
0'
0/
#134800000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#134810000000
0!
0'
0/
#134820000000
1!
1'
1/
#134830000000
0!
0'
0/
#134840000000
1!
1'
1/
#134850000000
0!
0'
0/
#134860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#134870000000
0!
0'
0/
#134880000000
1!
1'
1/
#134890000000
0!
0'
0/
#134900000000
1!
1'
1/
#134910000000
0!
0'
0/
#134920000000
1!
1'
1/
#134930000000
0!
0'
0/
#134940000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#134950000000
0!
0'
0/
#134960000000
1!
1'
1/
#134970000000
0!
0'
0/
#134980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#134990000000
0!
0'
0/
#135000000000
1!
1'
1/
#135010000000
0!
0'
0/
#135020000000
#135030000000
1!
1'
1/
#135040000000
0!
0'
0/
#135050000000
1!
1'
1/
#135060000000
0!
1"
0'
1(
0/
10
#135070000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#135080000000
0!
0'
0/
#135090000000
1!
1'
1/
#135100000000
0!
0'
0/
#135110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#135120000000
0!
0'
0/
#135130000000
1!
1'
1/
#135140000000
0!
1"
0'
1(
0/
10
#135150000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#135160000000
0!
1$
0'
1+
0/
#135170000000
1!
1'
1/
#135180000000
0!
0'
0/
#135190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#135200000000
0!
0'
0/
#135210000000
1!
1'
1/
#135220000000
0!
0'
0/
#135230000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#135240000000
0!
0'
0/
#135250000000
1!
1'
1/
#135260000000
0!
0'
0/
#135270000000
1!
1'
1/
#135280000000
0!
0'
0/
#135290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#135300000000
0!
0'
0/
#135310000000
1!
1'
1/
#135320000000
0!
0'
0/
#135330000000
1!
1'
1/
#135340000000
0!
0'
0/
#135350000000
1!
1'
1/
#135360000000
0!
0'
0/
#135370000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#135380000000
0!
0'
0/
#135390000000
1!
1'
1/
#135400000000
0!
0'
0/
#135410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#135420000000
0!
0'
0/
#135430000000
1!
1'
1/
#135440000000
0!
0'
0/
#135450000000
#135460000000
1!
1'
1/
#135470000000
0!
0'
0/
#135480000000
1!
1'
1/
#135490000000
0!
1"
0'
1(
0/
10
#135500000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#135510000000
0!
0'
0/
#135520000000
1!
1'
1/
#135530000000
0!
0'
0/
#135540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#135550000000
0!
0'
0/
#135560000000
1!
1'
1/
#135570000000
0!
1"
0'
1(
0/
10
#135580000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#135590000000
0!
1$
0'
1+
0/
#135600000000
1!
1'
1/
#135610000000
0!
0'
0/
#135620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#135630000000
0!
0'
0/
#135640000000
1!
1'
1/
#135650000000
0!
0'
0/
#135660000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#135670000000
0!
0'
0/
#135680000000
1!
1'
1/
#135690000000
0!
0'
0/
#135700000000
1!
1'
1/
#135710000000
0!
0'
0/
#135720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#135730000000
0!
0'
0/
#135740000000
1!
1'
1/
#135750000000
0!
0'
0/
#135760000000
1!
1'
1/
#135770000000
0!
0'
0/
#135780000000
1!
1'
1/
#135790000000
0!
0'
0/
#135800000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#135810000000
0!
0'
0/
#135820000000
1!
1'
1/
#135830000000
0!
0'
0/
#135840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#135850000000
0!
0'
0/
#135860000000
1!
1'
1/
#135870000000
0!
0'
0/
#135880000000
#135890000000
1!
1'
1/
#135900000000
0!
0'
0/
#135910000000
1!
1'
1/
#135920000000
0!
1"
0'
1(
0/
10
#135930000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#135940000000
0!
0'
0/
#135950000000
1!
1'
1/
#135960000000
0!
0'
0/
#135970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#135980000000
0!
0'
0/
#135990000000
1!
1'
1/
#136000000000
0!
1"
0'
1(
0/
10
#136010000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#136020000000
0!
1$
0'
1+
0/
#136030000000
1!
1'
1/
#136040000000
0!
0'
0/
#136050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#136060000000
0!
0'
0/
#136070000000
1!
1'
1/
#136080000000
0!
0'
0/
#136090000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#136100000000
0!
0'
0/
#136110000000
1!
1'
1/
#136120000000
0!
0'
0/
#136130000000
1!
1'
1/
#136140000000
0!
0'
0/
#136150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#136160000000
0!
0'
0/
#136170000000
1!
1'
1/
#136180000000
0!
0'
0/
#136190000000
1!
1'
1/
#136200000000
0!
0'
0/
#136210000000
1!
1'
1/
#136220000000
0!
0'
0/
#136230000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#136240000000
0!
0'
0/
#136250000000
1!
1'
1/
#136260000000
0!
0'
0/
#136270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#136280000000
0!
0'
0/
#136290000000
1!
1'
1/
#136300000000
0!
0'
0/
#136310000000
#136320000000
1!
1'
1/
#136330000000
0!
0'
0/
#136340000000
1!
1'
1/
#136350000000
0!
1"
0'
1(
0/
10
#136360000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#136370000000
0!
0'
0/
#136380000000
1!
1'
1/
#136390000000
0!
0'
0/
#136400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#136410000000
0!
0'
0/
#136420000000
1!
1'
1/
#136430000000
0!
1"
0'
1(
0/
10
#136440000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#136450000000
0!
1$
0'
1+
0/
#136460000000
1!
1'
1/
#136470000000
0!
0'
0/
#136480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#136490000000
0!
0'
0/
#136500000000
1!
1'
1/
#136510000000
0!
0'
0/
#136520000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#136530000000
0!
0'
0/
#136540000000
1!
1'
1/
#136550000000
0!
0'
0/
#136560000000
1!
1'
1/
#136570000000
0!
0'
0/
#136580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#136590000000
0!
0'
0/
#136600000000
1!
1'
1/
#136610000000
0!
0'
0/
#136620000000
1!
1'
1/
#136630000000
0!
0'
0/
#136640000000
1!
1'
1/
#136650000000
0!
0'
0/
#136660000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#136670000000
0!
0'
0/
#136680000000
1!
1'
1/
#136690000000
0!
0'
0/
#136700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#136710000000
0!
0'
0/
#136720000000
1!
1'
1/
#136730000000
0!
0'
0/
#136740000000
#136750000000
1!
1'
1/
#136760000000
0!
0'
0/
#136770000000
1!
1'
1/
#136780000000
0!
1"
0'
1(
0/
10
#136790000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#136800000000
0!
0'
0/
#136810000000
1!
1'
1/
#136820000000
0!
0'
0/
#136830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#136840000000
0!
0'
0/
#136850000000
1!
1'
1/
#136860000000
0!
1"
0'
1(
0/
10
#136870000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#136880000000
0!
1$
0'
1+
0/
#136890000000
1!
1'
1/
#136900000000
0!
0'
0/
#136910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#136920000000
0!
0'
0/
#136930000000
1!
1'
1/
#136940000000
0!
0'
0/
#136950000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#136960000000
0!
0'
0/
#136970000000
1!
1'
1/
#136980000000
0!
0'
0/
#136990000000
1!
1'
1/
#137000000000
0!
0'
0/
#137010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#137020000000
0!
0'
0/
#137030000000
1!
1'
1/
#137040000000
0!
0'
0/
#137050000000
1!
1'
1/
#137060000000
0!
0'
0/
#137070000000
1!
1'
1/
#137080000000
0!
0'
0/
#137090000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#137100000000
0!
0'
0/
#137110000000
1!
1'
1/
#137120000000
0!
0'
0/
#137130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#137140000000
0!
0'
0/
#137150000000
1!
1'
1/
#137160000000
0!
0'
0/
#137170000000
#137180000000
1!
1'
1/
#137190000000
0!
0'
0/
#137200000000
1!
1'
1/
#137210000000
0!
1"
0'
1(
0/
10
#137220000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#137230000000
0!
0'
0/
#137240000000
1!
1'
1/
#137250000000
0!
0'
0/
#137260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#137270000000
0!
0'
0/
#137280000000
1!
1'
1/
#137290000000
0!
1"
0'
1(
0/
10
#137300000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#137310000000
0!
1$
0'
1+
0/
#137320000000
1!
1'
1/
#137330000000
0!
0'
0/
#137340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#137350000000
0!
0'
0/
#137360000000
1!
1'
1/
#137370000000
0!
0'
0/
#137380000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#137390000000
0!
0'
0/
#137400000000
1!
1'
1/
#137410000000
0!
0'
0/
#137420000000
1!
1'
1/
#137430000000
0!
0'
0/
#137440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#137450000000
0!
0'
0/
#137460000000
1!
1'
1/
#137470000000
0!
0'
0/
#137480000000
1!
1'
1/
#137490000000
0!
0'
0/
#137500000000
1!
1'
1/
#137510000000
0!
0'
0/
#137520000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#137530000000
0!
0'
0/
#137540000000
1!
1'
1/
#137550000000
0!
0'
0/
#137560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#137570000000
0!
0'
0/
#137580000000
1!
1'
1/
#137590000000
0!
0'
0/
#137600000000
#137610000000
1!
1'
1/
#137620000000
0!
0'
0/
#137630000000
1!
1'
1/
#137640000000
0!
1"
0'
1(
0/
10
#137650000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#137660000000
0!
0'
0/
#137670000000
1!
1'
1/
#137680000000
0!
0'
0/
#137690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#137700000000
0!
0'
0/
#137710000000
1!
1'
1/
#137720000000
0!
1"
0'
1(
0/
10
#137730000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#137740000000
0!
1$
0'
1+
0/
#137750000000
1!
1'
1/
#137760000000
0!
0'
0/
#137770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#137780000000
0!
0'
0/
#137790000000
1!
1'
1/
#137800000000
0!
0'
0/
#137810000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#137820000000
0!
0'
0/
#137830000000
1!
1'
1/
#137840000000
0!
0'
0/
#137850000000
1!
1'
1/
#137860000000
0!
0'
0/
#137870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#137880000000
0!
0'
0/
#137890000000
1!
1'
1/
#137900000000
0!
0'
0/
#137910000000
1!
1'
1/
#137920000000
0!
0'
0/
#137930000000
1!
1'
1/
#137940000000
0!
0'
0/
#137950000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#137960000000
0!
0'
0/
#137970000000
1!
1'
1/
#137980000000
0!
0'
0/
#137990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#138000000000
0!
0'
0/
#138010000000
1!
1'
1/
#138020000000
0!
0'
0/
#138030000000
#138040000000
1!
1'
1/
#138050000000
0!
0'
0/
#138060000000
1!
1'
1/
#138070000000
0!
1"
0'
1(
0/
10
#138080000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#138090000000
0!
0'
0/
#138100000000
1!
1'
1/
#138110000000
0!
0'
0/
#138120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#138130000000
0!
0'
0/
#138140000000
1!
1'
1/
#138150000000
0!
1"
0'
1(
0/
10
#138160000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#138170000000
0!
1$
0'
1+
0/
#138180000000
1!
1'
1/
#138190000000
0!
0'
0/
#138200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#138210000000
0!
0'
0/
#138220000000
1!
1'
1/
#138230000000
0!
0'
0/
#138240000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#138250000000
0!
0'
0/
#138260000000
1!
1'
1/
#138270000000
0!
0'
0/
#138280000000
1!
1'
1/
#138290000000
0!
0'
0/
#138300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#138310000000
0!
0'
0/
#138320000000
1!
1'
1/
#138330000000
0!
0'
0/
#138340000000
1!
1'
1/
#138350000000
0!
0'
0/
#138360000000
1!
1'
1/
#138370000000
0!
0'
0/
#138380000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#138390000000
0!
0'
0/
#138400000000
1!
1'
1/
#138410000000
0!
0'
0/
#138420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#138430000000
0!
0'
0/
#138440000000
1!
1'
1/
#138450000000
0!
0'
0/
#138460000000
#138470000000
1!
1'
1/
#138480000000
0!
0'
0/
#138490000000
1!
1'
1/
#138500000000
0!
1"
0'
1(
0/
10
#138510000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#138520000000
0!
0'
0/
#138530000000
1!
1'
1/
#138540000000
0!
0'
0/
#138550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#138560000000
0!
0'
0/
#138570000000
1!
1'
1/
#138580000000
0!
1"
0'
1(
0/
10
#138590000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#138600000000
0!
1$
0'
1+
0/
#138610000000
1!
1'
1/
#138620000000
0!
0'
0/
#138630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#138640000000
0!
0'
0/
#138650000000
1!
1'
1/
#138660000000
0!
0'
0/
#138670000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#138680000000
0!
0'
0/
#138690000000
1!
1'
1/
#138700000000
0!
0'
0/
#138710000000
1!
1'
1/
#138720000000
0!
0'
0/
#138730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#138740000000
0!
0'
0/
#138750000000
1!
1'
1/
#138760000000
0!
0'
0/
#138770000000
1!
1'
1/
#138780000000
0!
0'
0/
#138790000000
1!
1'
1/
#138800000000
0!
0'
0/
#138810000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#138820000000
0!
0'
0/
#138830000000
1!
1'
1/
#138840000000
0!
0'
0/
#138850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#138860000000
0!
0'
0/
#138870000000
1!
1'
1/
#138880000000
0!
0'
0/
#138890000000
#138900000000
1!
1'
1/
#138910000000
0!
0'
0/
#138920000000
1!
1'
1/
#138930000000
0!
1"
0'
1(
0/
10
#138940000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#138950000000
0!
0'
0/
#138960000000
1!
1'
1/
#138970000000
0!
0'
0/
#138980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#138990000000
0!
0'
0/
#139000000000
1!
1'
1/
#139010000000
0!
1"
0'
1(
0/
10
#139020000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#139030000000
0!
1$
0'
1+
0/
#139040000000
1!
1'
1/
#139050000000
0!
0'
0/
#139060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#139070000000
0!
0'
0/
#139080000000
1!
1'
1/
#139090000000
0!
0'
0/
#139100000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#139110000000
0!
0'
0/
#139120000000
1!
1'
1/
#139130000000
0!
0'
0/
#139140000000
1!
1'
1/
#139150000000
0!
0'
0/
#139160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#139170000000
0!
0'
0/
#139180000000
1!
1'
1/
#139190000000
0!
0'
0/
#139200000000
1!
1'
1/
#139210000000
0!
0'
0/
#139220000000
1!
1'
1/
#139230000000
0!
0'
0/
#139240000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#139250000000
0!
0'
0/
#139260000000
1!
1'
1/
#139270000000
0!
0'
0/
#139280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#139290000000
0!
0'
0/
#139300000000
1!
1'
1/
#139310000000
0!
0'
0/
#139320000000
#139330000000
1!
1'
1/
#139340000000
0!
0'
0/
#139350000000
1!
1'
1/
#139360000000
0!
1"
0'
1(
0/
10
#139370000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#139380000000
0!
0'
0/
#139390000000
1!
1'
1/
#139400000000
0!
0'
0/
#139410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#139420000000
0!
0'
0/
#139430000000
1!
1'
1/
#139440000000
0!
1"
0'
1(
0/
10
#139450000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#139460000000
0!
1$
0'
1+
0/
#139470000000
1!
1'
1/
#139480000000
0!
0'
0/
#139490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#139500000000
0!
0'
0/
#139510000000
1!
1'
1/
#139520000000
0!
0'
0/
#139530000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#139540000000
0!
0'
0/
#139550000000
1!
1'
1/
#139560000000
0!
0'
0/
#139570000000
1!
1'
1/
#139580000000
0!
0'
0/
#139590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#139600000000
0!
0'
0/
#139610000000
1!
1'
1/
#139620000000
0!
0'
0/
#139630000000
1!
1'
1/
#139640000000
0!
0'
0/
#139650000000
1!
1'
1/
#139660000000
0!
0'
0/
#139670000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#139680000000
0!
0'
0/
#139690000000
1!
1'
1/
#139700000000
0!
0'
0/
#139710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#139720000000
0!
0'
0/
#139730000000
1!
1'
1/
#139740000000
0!
0'
0/
#139750000000
#139760000000
1!
1'
1/
#139770000000
0!
0'
0/
#139780000000
1!
1'
1/
#139790000000
0!
1"
0'
1(
0/
10
#139800000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#139810000000
0!
0'
0/
#139820000000
1!
1'
1/
#139830000000
0!
0'
0/
#139840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#139850000000
0!
0'
0/
#139860000000
1!
1'
1/
#139870000000
0!
1"
0'
1(
0/
10
#139880000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#139890000000
0!
1$
0'
1+
0/
#139900000000
1!
1'
1/
#139910000000
0!
0'
0/
#139920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#139930000000
0!
0'
0/
#139940000000
1!
1'
1/
#139950000000
0!
0'
0/
#139960000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#139970000000
0!
0'
0/
#139980000000
1!
1'
1/
#139990000000
0!
0'
0/
#140000000000
1!
1'
1/
#140010000000
0!
0'
0/
#140020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#140030000000
0!
0'
0/
#140040000000
1!
1'
1/
#140050000000
0!
0'
0/
#140060000000
1!
1'
1/
#140070000000
0!
0'
0/
#140080000000
1!
1'
1/
#140090000000
0!
0'
0/
#140100000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#140110000000
0!
0'
0/
#140120000000
1!
1'
1/
#140130000000
0!
0'
0/
#140140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#140150000000
0!
0'
0/
#140160000000
1!
1'
1/
#140170000000
0!
0'
0/
#140180000000
#140190000000
1!
1'
1/
#140200000000
0!
0'
0/
#140210000000
1!
1'
1/
#140220000000
0!
1"
0'
1(
0/
10
#140230000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#140240000000
0!
0'
0/
#140250000000
1!
1'
1/
#140260000000
0!
0'
0/
#140270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#140280000000
0!
0'
0/
#140290000000
1!
1'
1/
#140300000000
0!
1"
0'
1(
0/
10
#140310000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#140320000000
0!
1$
0'
1+
0/
#140330000000
1!
1'
1/
#140340000000
0!
0'
0/
#140350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#140360000000
0!
0'
0/
#140370000000
1!
1'
1/
#140380000000
0!
0'
0/
#140390000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#140400000000
0!
0'
0/
#140410000000
1!
1'
1/
#140420000000
0!
0'
0/
#140430000000
1!
1'
1/
#140440000000
0!
0'
0/
#140450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#140460000000
0!
0'
0/
#140470000000
1!
1'
1/
#140480000000
0!
0'
0/
#140490000000
1!
1'
1/
#140500000000
0!
0'
0/
#140510000000
1!
1'
1/
#140520000000
0!
0'
0/
#140530000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#140540000000
0!
0'
0/
#140550000000
1!
1'
1/
#140560000000
0!
0'
0/
#140570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#140580000000
0!
0'
0/
#140590000000
1!
1'
1/
#140600000000
0!
0'
0/
#140610000000
#140620000000
1!
1'
1/
#140630000000
0!
0'
0/
#140640000000
1!
1'
1/
#140650000000
0!
1"
0'
1(
0/
10
#140660000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#140670000000
0!
0'
0/
#140680000000
1!
1'
1/
#140690000000
0!
0'
0/
#140700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#140710000000
0!
0'
0/
#140720000000
1!
1'
1/
#140730000000
0!
1"
0'
1(
0/
10
#140740000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#140750000000
0!
1$
0'
1+
0/
#140760000000
1!
1'
1/
#140770000000
0!
0'
0/
#140780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#140790000000
0!
0'
0/
#140800000000
1!
1'
1/
#140810000000
0!
0'
0/
#140820000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#140830000000
0!
0'
0/
#140840000000
1!
1'
1/
#140850000000
0!
0'
0/
#140860000000
1!
1'
1/
#140870000000
0!
0'
0/
#140880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#140890000000
0!
0'
0/
#140900000000
1!
1'
1/
#140910000000
0!
0'
0/
#140920000000
1!
1'
1/
#140930000000
0!
0'
0/
#140940000000
1!
1'
1/
#140950000000
0!
0'
0/
#140960000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#140970000000
0!
0'
0/
#140980000000
1!
1'
1/
#140990000000
0!
0'
0/
#141000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#141010000000
0!
0'
0/
#141020000000
1!
1'
1/
#141030000000
0!
0'
0/
#141040000000
#141050000000
1!
1'
1/
#141060000000
0!
0'
0/
#141070000000
1!
1'
1/
#141080000000
0!
1"
0'
1(
0/
10
#141090000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#141100000000
0!
0'
0/
#141110000000
1!
1'
1/
#141120000000
0!
0'
0/
#141130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#141140000000
0!
0'
0/
#141150000000
1!
1'
1/
#141160000000
0!
1"
0'
1(
0/
10
#141170000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#141180000000
0!
1$
0'
1+
0/
#141190000000
1!
1'
1/
#141200000000
0!
0'
0/
#141210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#141220000000
0!
0'
0/
#141230000000
1!
1'
1/
#141240000000
0!
0'
0/
#141250000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#141260000000
0!
0'
0/
#141270000000
1!
1'
1/
#141280000000
0!
0'
0/
#141290000000
1!
1'
1/
#141300000000
0!
0'
0/
#141310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#141320000000
0!
0'
0/
#141330000000
1!
1'
1/
#141340000000
0!
0'
0/
#141350000000
1!
1'
1/
#141360000000
0!
0'
0/
#141370000000
1!
1'
1/
#141380000000
0!
0'
0/
#141390000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#141400000000
0!
0'
0/
#141410000000
1!
1'
1/
#141420000000
0!
0'
0/
#141430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#141440000000
0!
0'
0/
#141450000000
1!
1'
1/
#141460000000
0!
0'
0/
#141470000000
#141480000000
1!
1'
1/
#141490000000
0!
0'
0/
#141500000000
1!
1'
1/
#141510000000
0!
1"
0'
1(
0/
10
#141520000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#141530000000
0!
0'
0/
#141540000000
1!
1'
1/
#141550000000
0!
0'
0/
#141560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#141570000000
0!
0'
0/
#141580000000
1!
1'
1/
#141590000000
0!
1"
0'
1(
0/
10
#141600000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#141610000000
0!
1$
0'
1+
0/
#141620000000
1!
1'
1/
#141630000000
0!
0'
0/
#141640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#141650000000
0!
0'
0/
#141660000000
1!
1'
1/
#141670000000
0!
0'
0/
#141680000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#141690000000
0!
0'
0/
#141700000000
1!
1'
1/
#141710000000
0!
0'
0/
#141720000000
1!
1'
1/
#141730000000
0!
0'
0/
#141740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#141750000000
0!
0'
0/
#141760000000
1!
1'
1/
#141770000000
0!
0'
0/
#141780000000
1!
1'
1/
#141790000000
0!
0'
0/
#141800000000
1!
1'
1/
#141810000000
0!
0'
0/
#141820000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#141830000000
0!
0'
0/
#141840000000
1!
1'
1/
#141850000000
0!
0'
0/
#141860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#141870000000
0!
0'
0/
#141880000000
1!
1'
1/
#141890000000
0!
0'
0/
#141900000000
#141910000000
1!
1'
1/
#141920000000
0!
0'
0/
#141930000000
1!
1'
1/
#141940000000
0!
1"
0'
1(
0/
10
#141950000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#141960000000
0!
0'
0/
#141970000000
1!
1'
1/
#141980000000
0!
0'
0/
#141990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#142000000000
0!
0'
0/
#142010000000
1!
1'
1/
#142020000000
0!
1"
0'
1(
0/
10
#142030000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#142040000000
0!
1$
0'
1+
0/
#142050000000
1!
1'
1/
#142060000000
0!
0'
0/
#142070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#142080000000
0!
0'
0/
#142090000000
1!
1'
1/
#142100000000
0!
0'
0/
#142110000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#142120000000
0!
0'
0/
#142130000000
1!
1'
1/
#142140000000
0!
0'
0/
#142150000000
1!
1'
1/
#142160000000
0!
0'
0/
#142170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#142180000000
0!
0'
0/
#142190000000
1!
1'
1/
#142200000000
0!
0'
0/
#142210000000
1!
1'
1/
#142220000000
0!
0'
0/
#142230000000
1!
1'
1/
#142240000000
0!
0'
0/
#142250000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#142260000000
0!
0'
0/
#142270000000
1!
1'
1/
#142280000000
0!
0'
0/
#142290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#142300000000
0!
0'
0/
#142310000000
1!
1'
1/
#142320000000
0!
0'
0/
#142330000000
#142340000000
1!
1'
1/
#142350000000
0!
0'
0/
#142360000000
1!
1'
1/
#142370000000
0!
1"
0'
1(
0/
10
#142380000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#142390000000
0!
0'
0/
#142400000000
1!
1'
1/
#142410000000
0!
0'
0/
#142420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#142430000000
0!
0'
0/
#142440000000
1!
1'
1/
#142450000000
0!
1"
0'
1(
0/
10
#142460000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#142470000000
0!
1$
0'
1+
0/
#142480000000
1!
1'
1/
#142490000000
0!
0'
0/
#142500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#142510000000
0!
0'
0/
#142520000000
1!
1'
1/
#142530000000
0!
0'
0/
#142540000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#142550000000
0!
0'
0/
#142560000000
1!
1'
1/
#142570000000
0!
0'
0/
#142580000000
1!
1'
1/
#142590000000
0!
0'
0/
#142600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#142610000000
0!
0'
0/
#142620000000
1!
1'
1/
#142630000000
0!
0'
0/
#142640000000
1!
1'
1/
#142650000000
0!
0'
0/
#142660000000
1!
1'
1/
#142670000000
0!
0'
0/
#142680000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#142690000000
0!
0'
0/
#142700000000
1!
1'
1/
#142710000000
0!
0'
0/
#142720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#142730000000
0!
0'
0/
#142740000000
1!
1'
1/
#142750000000
0!
0'
0/
#142760000000
#142770000000
1!
1'
1/
#142780000000
0!
0'
0/
#142790000000
1!
1'
1/
#142800000000
0!
1"
0'
1(
0/
10
#142810000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#142820000000
0!
0'
0/
#142830000000
1!
1'
1/
#142840000000
0!
0'
0/
#142850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#142860000000
0!
0'
0/
#142870000000
1!
1'
1/
#142880000000
0!
1"
0'
1(
0/
10
#142890000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#142900000000
0!
1$
0'
1+
0/
#142910000000
1!
1'
1/
#142920000000
0!
0'
0/
#142930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#142940000000
0!
0'
0/
#142950000000
1!
1'
1/
#142960000000
0!
0'
0/
#142970000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#142980000000
0!
0'
0/
#142990000000
1!
1'
1/
#143000000000
0!
0'
0/
#143010000000
1!
1'
1/
#143020000000
0!
0'
0/
#143030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#143040000000
0!
0'
0/
#143050000000
1!
1'
1/
#143060000000
0!
0'
0/
#143070000000
1!
1'
1/
#143080000000
0!
0'
0/
#143090000000
1!
1'
1/
#143100000000
0!
0'
0/
#143110000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#143120000000
0!
0'
0/
#143130000000
1!
1'
1/
#143140000000
0!
0'
0/
#143150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#143160000000
0!
0'
0/
#143170000000
1!
1'
1/
#143180000000
0!
0'
0/
#143190000000
#143200000000
1!
1'
1/
#143210000000
0!
0'
0/
#143220000000
1!
1'
1/
#143230000000
0!
1"
0'
1(
0/
10
#143240000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#143250000000
0!
0'
0/
#143260000000
1!
1'
1/
#143270000000
0!
0'
0/
#143280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#143290000000
0!
0'
0/
#143300000000
1!
1'
1/
#143310000000
0!
1"
0'
1(
0/
10
#143320000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#143330000000
0!
1$
0'
1+
0/
#143340000000
1!
1'
1/
#143350000000
0!
0'
0/
#143360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#143370000000
0!
0'
0/
#143380000000
1!
1'
1/
#143390000000
0!
0'
0/
#143400000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#143410000000
0!
0'
0/
#143420000000
1!
1'
1/
#143430000000
0!
0'
0/
#143440000000
1!
1'
1/
#143450000000
0!
0'
0/
#143460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#143470000000
0!
0'
0/
#143480000000
1!
1'
1/
#143490000000
0!
0'
0/
#143500000000
1!
1'
1/
#143510000000
0!
0'
0/
#143520000000
1!
1'
1/
#143530000000
0!
0'
0/
#143540000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#143550000000
0!
0'
0/
#143560000000
1!
1'
1/
#143570000000
0!
0'
0/
#143580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#143590000000
0!
0'
0/
#143600000000
1!
1'
1/
#143610000000
0!
0'
0/
#143620000000
#143630000000
1!
1'
1/
#143640000000
0!
0'
0/
#143650000000
1!
1'
1/
#143660000000
0!
1"
0'
1(
0/
10
#143670000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#143680000000
0!
0'
0/
#143690000000
1!
1'
1/
#143700000000
0!
0'
0/
#143710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#143720000000
0!
0'
0/
#143730000000
1!
1'
1/
#143740000000
0!
1"
0'
1(
0/
10
#143750000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#143760000000
0!
1$
0'
1+
0/
#143770000000
1!
1'
1/
#143780000000
0!
0'
0/
#143790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#143800000000
0!
0'
0/
#143810000000
1!
1'
1/
#143820000000
0!
0'
0/
#143830000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#143840000000
0!
0'
0/
#143850000000
1!
1'
1/
#143860000000
0!
0'
0/
#143870000000
1!
1'
1/
#143880000000
0!
0'
0/
#143890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#143900000000
0!
0'
0/
#143910000000
1!
1'
1/
#143920000000
0!
0'
0/
#143930000000
1!
1'
1/
#143940000000
0!
0'
0/
#143950000000
1!
1'
1/
#143960000000
0!
0'
0/
#143970000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#143980000000
0!
0'
0/
#143990000000
1!
1'
1/
#144000000000
0!
0'
0/
#144010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#144020000000
0!
0'
0/
#144030000000
1!
1'
1/
#144040000000
0!
0'
0/
#144050000000
#144060000000
1!
1'
1/
#144070000000
0!
0'
0/
#144080000000
1!
1'
1/
#144090000000
0!
1"
0'
1(
0/
10
#144100000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#144110000000
0!
0'
0/
#144120000000
1!
1'
1/
#144130000000
0!
0'
0/
#144140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#144150000000
0!
0'
0/
#144160000000
1!
1'
1/
#144170000000
0!
1"
0'
1(
0/
10
#144180000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#144190000000
0!
1$
0'
1+
0/
#144200000000
1!
1'
1/
#144210000000
0!
0'
0/
#144220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#144230000000
0!
0'
0/
#144240000000
1!
1'
1/
#144250000000
0!
0'
0/
#144260000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#144270000000
0!
0'
0/
#144280000000
1!
1'
1/
#144290000000
0!
0'
0/
#144300000000
1!
1'
1/
#144310000000
0!
0'
0/
#144320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#144330000000
0!
0'
0/
#144340000000
1!
1'
1/
#144350000000
0!
0'
0/
#144360000000
1!
1'
1/
#144370000000
0!
0'
0/
#144380000000
1!
1'
1/
#144390000000
0!
0'
0/
#144400000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#144410000000
0!
0'
0/
#144420000000
1!
1'
1/
#144430000000
0!
0'
0/
#144440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#144450000000
0!
0'
0/
#144460000000
1!
1'
1/
#144470000000
0!
0'
0/
#144480000000
#144490000000
1!
1'
1/
#144500000000
0!
0'
0/
#144510000000
1!
1'
1/
#144520000000
0!
1"
0'
1(
0/
10
#144530000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#144540000000
0!
0'
0/
#144550000000
1!
1'
1/
#144560000000
0!
0'
0/
#144570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#144580000000
0!
0'
0/
#144590000000
1!
1'
1/
#144600000000
0!
1"
0'
1(
0/
10
#144610000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#144620000000
0!
1$
0'
1+
0/
#144630000000
1!
1'
1/
#144640000000
0!
0'
0/
#144650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#144660000000
0!
0'
0/
#144670000000
1!
1'
1/
#144680000000
0!
0'
0/
#144690000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#144700000000
0!
0'
0/
#144710000000
1!
1'
1/
#144720000000
0!
0'
0/
#144730000000
1!
1'
1/
#144740000000
0!
0'
0/
#144750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#144760000000
0!
0'
0/
#144770000000
1!
1'
1/
#144780000000
0!
0'
0/
#144790000000
1!
1'
1/
#144800000000
0!
0'
0/
#144810000000
1!
1'
1/
#144820000000
0!
0'
0/
#144830000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#144840000000
0!
0'
0/
#144850000000
1!
1'
1/
#144860000000
0!
0'
0/
#144870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#144880000000
0!
0'
0/
#144890000000
1!
1'
1/
#144900000000
0!
0'
0/
#144910000000
#144920000000
1!
1'
1/
#144930000000
0!
0'
0/
#144940000000
1!
1'
1/
#144950000000
0!
1"
0'
1(
0/
10
#144960000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#144970000000
0!
0'
0/
#144980000000
1!
1'
1/
#144990000000
0!
0'
0/
#145000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#145010000000
0!
0'
0/
#145020000000
1!
1'
1/
#145030000000
0!
1"
0'
1(
0/
10
#145040000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#145050000000
0!
1$
0'
1+
0/
#145060000000
1!
1'
1/
#145070000000
0!
0'
0/
#145080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#145090000000
0!
0'
0/
#145100000000
1!
1'
1/
#145110000000
0!
0'
0/
#145120000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#145130000000
0!
0'
0/
#145140000000
1!
1'
1/
#145150000000
0!
0'
0/
#145160000000
1!
1'
1/
#145170000000
0!
0'
0/
#145180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#145190000000
0!
0'
0/
#145200000000
1!
1'
1/
#145210000000
0!
0'
0/
#145220000000
1!
1'
1/
#145230000000
0!
0'
0/
#145240000000
1!
1'
1/
#145250000000
0!
0'
0/
#145260000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#145270000000
0!
0'
0/
#145280000000
1!
1'
1/
#145290000000
0!
0'
0/
#145300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#145310000000
0!
0'
0/
#145320000000
1!
1'
1/
#145330000000
0!
0'
0/
#145340000000
#145350000000
1!
1'
1/
#145360000000
0!
0'
0/
#145370000000
1!
1'
1/
#145380000000
0!
1"
0'
1(
0/
10
#145390000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#145400000000
0!
0'
0/
#145410000000
1!
1'
1/
#145420000000
0!
0'
0/
#145430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#145440000000
0!
0'
0/
#145450000000
1!
1'
1/
#145460000000
0!
1"
0'
1(
0/
10
#145470000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#145480000000
0!
1$
0'
1+
0/
#145490000000
1!
1'
1/
#145500000000
0!
0'
0/
#145510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#145520000000
0!
0'
0/
#145530000000
1!
1'
1/
#145540000000
0!
0'
0/
#145550000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#145560000000
0!
0'
0/
#145570000000
1!
1'
1/
#145580000000
0!
0'
0/
#145590000000
1!
1'
1/
#145600000000
0!
0'
0/
#145610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#145620000000
0!
0'
0/
#145630000000
1!
1'
1/
#145640000000
0!
0'
0/
#145650000000
1!
1'
1/
#145660000000
0!
0'
0/
#145670000000
1!
1'
1/
#145680000000
0!
0'
0/
#145690000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#145700000000
0!
0'
0/
#145710000000
1!
1'
1/
#145720000000
0!
0'
0/
#145730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#145740000000
0!
0'
0/
#145750000000
1!
1'
1/
#145760000000
0!
0'
0/
#145770000000
#145780000000
1!
1'
1/
#145790000000
0!
0'
0/
#145800000000
1!
1'
1/
#145810000000
0!
1"
0'
1(
0/
10
#145820000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#145830000000
0!
0'
0/
#145840000000
1!
1'
1/
#145850000000
0!
0'
0/
#145860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#145870000000
0!
0'
0/
#145880000000
1!
1'
1/
#145890000000
0!
1"
0'
1(
0/
10
#145900000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#145910000000
0!
1$
0'
1+
0/
#145920000000
1!
1'
1/
#145930000000
0!
0'
0/
#145940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#145950000000
0!
0'
0/
#145960000000
1!
1'
1/
#145970000000
0!
0'
0/
#145980000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#145990000000
0!
0'
0/
#146000000000
1!
1'
1/
#146010000000
0!
0'
0/
#146020000000
1!
1'
1/
#146030000000
0!
0'
0/
#146040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#146050000000
0!
0'
0/
#146060000000
1!
1'
1/
#146070000000
0!
0'
0/
#146080000000
1!
1'
1/
#146090000000
0!
0'
0/
#146100000000
1!
1'
1/
#146110000000
0!
0'
0/
#146120000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#146130000000
0!
0'
0/
#146140000000
1!
1'
1/
#146150000000
0!
0'
0/
#146160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#146170000000
0!
0'
0/
#146180000000
1!
1'
1/
#146190000000
0!
0'
0/
#146200000000
#146210000000
1!
1'
1/
#146220000000
0!
0'
0/
#146230000000
1!
1'
1/
#146240000000
0!
1"
0'
1(
0/
10
#146250000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#146260000000
0!
0'
0/
#146270000000
1!
1'
1/
#146280000000
0!
0'
0/
#146290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#146300000000
0!
0'
0/
#146310000000
1!
1'
1/
#146320000000
0!
1"
0'
1(
0/
10
#146330000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#146340000000
0!
1$
0'
1+
0/
#146350000000
1!
1'
1/
#146360000000
0!
0'
0/
#146370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#146380000000
0!
0'
0/
#146390000000
1!
1'
1/
#146400000000
0!
0'
0/
#146410000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#146420000000
0!
0'
0/
#146430000000
1!
1'
1/
#146440000000
0!
0'
0/
#146450000000
1!
1'
1/
#146460000000
0!
0'
0/
#146470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#146480000000
0!
0'
0/
#146490000000
1!
1'
1/
#146500000000
0!
0'
0/
#146510000000
1!
1'
1/
#146520000000
0!
0'
0/
#146530000000
1!
1'
1/
#146540000000
0!
0'
0/
#146550000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#146560000000
0!
0'
0/
#146570000000
1!
1'
1/
#146580000000
0!
0'
0/
#146590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#146600000000
0!
0'
0/
#146610000000
1!
1'
1/
#146620000000
0!
0'
0/
#146630000000
#146640000000
1!
1'
1/
#146650000000
0!
0'
0/
#146660000000
1!
1'
1/
#146670000000
0!
1"
0'
1(
0/
10
#146680000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#146690000000
0!
0'
0/
#146700000000
1!
1'
1/
#146710000000
0!
0'
0/
#146720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#146730000000
0!
0'
0/
#146740000000
1!
1'
1/
#146750000000
0!
1"
0'
1(
0/
10
#146760000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#146770000000
0!
1$
0'
1+
0/
#146780000000
1!
1'
1/
#146790000000
0!
0'
0/
#146800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#146810000000
0!
0'
0/
#146820000000
1!
1'
1/
#146830000000
0!
0'
0/
#146840000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#146850000000
0!
0'
0/
#146860000000
1!
1'
1/
#146870000000
0!
0'
0/
#146880000000
1!
1'
1/
#146890000000
0!
0'
0/
#146900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#146910000000
0!
0'
0/
#146920000000
1!
1'
1/
#146930000000
0!
0'
0/
#146940000000
1!
1'
1/
#146950000000
0!
0'
0/
#146960000000
1!
1'
1/
#146970000000
0!
0'
0/
#146980000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#146990000000
0!
0'
0/
#147000000000
1!
1'
1/
#147010000000
0!
0'
0/
#147020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#147030000000
0!
0'
0/
#147040000000
1!
1'
1/
#147050000000
0!
0'
0/
#147060000000
#147070000000
1!
1'
1/
#147080000000
0!
0'
0/
#147090000000
1!
1'
1/
#147100000000
0!
1"
0'
1(
0/
10
#147110000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#147120000000
0!
0'
0/
#147130000000
1!
1'
1/
#147140000000
0!
0'
0/
#147150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#147160000000
0!
0'
0/
#147170000000
1!
1'
1/
#147180000000
0!
1"
0'
1(
0/
10
#147190000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#147200000000
0!
1$
0'
1+
0/
#147210000000
1!
1'
1/
#147220000000
0!
0'
0/
#147230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#147240000000
0!
0'
0/
#147250000000
1!
1'
1/
#147260000000
0!
0'
0/
#147270000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#147280000000
0!
0'
0/
#147290000000
1!
1'
1/
#147300000000
0!
0'
0/
#147310000000
1!
1'
1/
#147320000000
0!
0'
0/
#147330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#147340000000
0!
0'
0/
#147350000000
1!
1'
1/
#147360000000
0!
0'
0/
#147370000000
1!
1'
1/
#147380000000
0!
0'
0/
#147390000000
1!
1'
1/
#147400000000
0!
0'
0/
#147410000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#147420000000
0!
0'
0/
#147430000000
1!
1'
1/
#147440000000
0!
0'
0/
#147450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#147460000000
0!
0'
0/
#147470000000
1!
1'
1/
#147480000000
0!
0'
0/
#147490000000
#147500000000
1!
1'
1/
#147510000000
0!
0'
0/
#147520000000
1!
1'
1/
#147530000000
0!
1"
0'
1(
0/
10
#147540000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#147550000000
0!
0'
0/
#147560000000
1!
1'
1/
#147570000000
0!
0'
0/
#147580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#147590000000
0!
0'
0/
#147600000000
1!
1'
1/
#147610000000
0!
1"
0'
1(
0/
10
#147620000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#147630000000
0!
1$
0'
1+
0/
#147640000000
1!
1'
1/
#147650000000
0!
0'
0/
#147660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#147670000000
0!
0'
0/
#147680000000
1!
1'
1/
#147690000000
0!
0'
0/
#147700000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#147710000000
0!
0'
0/
#147720000000
1!
1'
1/
#147730000000
0!
0'
0/
#147740000000
1!
1'
1/
#147750000000
0!
0'
0/
#147760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#147770000000
0!
0'
0/
#147780000000
1!
1'
1/
#147790000000
0!
0'
0/
#147800000000
1!
1'
1/
#147810000000
0!
0'
0/
#147820000000
1!
1'
1/
#147830000000
0!
0'
0/
#147840000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#147850000000
0!
0'
0/
#147860000000
1!
1'
1/
#147870000000
0!
0'
0/
#147880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#147890000000
0!
0'
0/
#147900000000
1!
1'
1/
#147910000000
0!
0'
0/
#147920000000
#147930000000
1!
1'
1/
#147940000000
0!
0'
0/
#147950000000
1!
1'
1/
#147960000000
0!
1"
0'
1(
0/
10
#147970000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#147980000000
0!
0'
0/
#147990000000
1!
1'
1/
#148000000000
0!
0'
0/
#148010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#148020000000
0!
0'
0/
#148030000000
1!
1'
1/
#148040000000
0!
1"
0'
1(
0/
10
#148050000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#148060000000
0!
1$
0'
1+
0/
#148070000000
1!
1'
1/
#148080000000
0!
0'
0/
#148090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#148100000000
0!
0'
0/
#148110000000
1!
1'
1/
#148120000000
0!
0'
0/
#148130000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#148140000000
0!
0'
0/
#148150000000
1!
1'
1/
#148160000000
0!
0'
0/
#148170000000
1!
1'
1/
#148180000000
0!
0'
0/
#148190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#148200000000
0!
0'
0/
#148210000000
1!
1'
1/
#148220000000
0!
0'
0/
#148230000000
1!
1'
1/
#148240000000
0!
0'
0/
#148250000000
1!
1'
1/
#148260000000
0!
0'
0/
#148270000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#148280000000
0!
0'
0/
#148290000000
1!
1'
1/
#148300000000
0!
0'
0/
#148310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#148320000000
0!
0'
0/
#148330000000
1!
1'
1/
#148340000000
0!
0'
0/
#148350000000
#148360000000
1!
1'
1/
#148370000000
0!
0'
0/
#148380000000
1!
1'
1/
#148390000000
0!
1"
0'
1(
0/
10
#148400000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#148410000000
0!
0'
0/
#148420000000
1!
1'
1/
#148430000000
0!
0'
0/
#148440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#148450000000
0!
0'
0/
#148460000000
1!
1'
1/
#148470000000
0!
1"
0'
1(
0/
10
#148480000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#148490000000
0!
1$
0'
1+
0/
#148500000000
1!
1'
1/
#148510000000
0!
0'
0/
#148520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#148530000000
0!
0'
0/
#148540000000
1!
1'
1/
#148550000000
0!
0'
0/
#148560000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#148570000000
0!
0'
0/
#148580000000
1!
1'
1/
#148590000000
0!
0'
0/
#148600000000
1!
1'
1/
#148610000000
0!
0'
0/
#148620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#148630000000
0!
0'
0/
#148640000000
1!
1'
1/
#148650000000
0!
0'
0/
#148660000000
1!
1'
1/
#148670000000
0!
0'
0/
#148680000000
1!
1'
1/
#148690000000
0!
0'
0/
#148700000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#148710000000
0!
0'
0/
#148720000000
1!
1'
1/
#148730000000
0!
0'
0/
#148740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#148750000000
0!
0'
0/
#148760000000
1!
1'
1/
#148770000000
0!
0'
0/
#148780000000
#148790000000
1!
1'
1/
#148800000000
0!
0'
0/
#148810000000
1!
1'
1/
#148820000000
0!
1"
0'
1(
0/
10
#148830000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#148840000000
0!
0'
0/
#148850000000
1!
1'
1/
#148860000000
0!
0'
0/
#148870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#148880000000
0!
0'
0/
#148890000000
1!
1'
1/
#148900000000
0!
1"
0'
1(
0/
10
#148910000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#148920000000
0!
1$
0'
1+
0/
#148930000000
1!
1'
1/
#148940000000
0!
0'
0/
#148950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#148960000000
0!
0'
0/
#148970000000
1!
1'
1/
#148980000000
0!
0'
0/
#148990000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#149000000000
0!
0'
0/
#149010000000
1!
1'
1/
#149020000000
0!
0'
0/
#149030000000
1!
1'
1/
#149040000000
0!
0'
0/
#149050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#149060000000
0!
0'
0/
#149070000000
1!
1'
1/
#149080000000
0!
0'
0/
#149090000000
1!
1'
1/
#149100000000
0!
0'
0/
#149110000000
1!
1'
1/
#149120000000
0!
0'
0/
#149130000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#149140000000
0!
0'
0/
#149150000000
1!
1'
1/
#149160000000
0!
0'
0/
#149170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#149180000000
0!
0'
0/
#149190000000
1!
1'
1/
#149200000000
0!
0'
0/
#149210000000
#149220000000
1!
1'
1/
#149230000000
0!
0'
0/
#149240000000
1!
1'
1/
#149250000000
0!
1"
0'
1(
0/
10
#149260000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#149270000000
0!
0'
0/
#149280000000
1!
1'
1/
#149290000000
0!
0'
0/
#149300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#149310000000
0!
0'
0/
#149320000000
1!
1'
1/
#149330000000
0!
1"
0'
1(
0/
10
#149340000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#149350000000
0!
1$
0'
1+
0/
#149360000000
1!
1'
1/
#149370000000
0!
0'
0/
#149380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#149390000000
0!
0'
0/
#149400000000
1!
1'
1/
#149410000000
0!
0'
0/
#149420000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#149430000000
0!
0'
0/
#149440000000
1!
1'
1/
#149450000000
0!
0'
0/
#149460000000
1!
1'
1/
#149470000000
0!
0'
0/
#149480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#149490000000
0!
0'
0/
#149500000000
1!
1'
1/
#149510000000
0!
0'
0/
#149520000000
1!
1'
1/
#149530000000
0!
0'
0/
#149540000000
1!
1'
1/
#149550000000
0!
0'
0/
#149560000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#149570000000
0!
0'
0/
#149580000000
1!
1'
1/
#149590000000
0!
0'
0/
#149600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#149610000000
0!
0'
0/
#149620000000
1!
1'
1/
#149630000000
0!
0'
0/
#149640000000
#149650000000
1!
1'
1/
#149660000000
0!
0'
0/
#149670000000
1!
1'
1/
#149680000000
0!
1"
0'
1(
0/
10
#149690000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#149700000000
0!
0'
0/
#149710000000
1!
1'
1/
#149720000000
0!
0'
0/
#149730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#149740000000
0!
0'
0/
#149750000000
1!
1'
1/
#149760000000
0!
1"
0'
1(
0/
10
#149770000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#149780000000
0!
1$
0'
1+
0/
#149790000000
1!
1'
1/
#149800000000
0!
0'
0/
#149810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#149820000000
0!
0'
0/
#149830000000
1!
1'
1/
#149840000000
0!
0'
0/
#149850000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#149860000000
0!
0'
0/
#149870000000
1!
1'
1/
#149880000000
0!
0'
0/
#149890000000
1!
1'
1/
#149900000000
0!
0'
0/
#149910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#149920000000
0!
0'
0/
#149930000000
1!
1'
1/
#149940000000
0!
0'
0/
#149950000000
1!
1'
1/
#149960000000
0!
0'
0/
#149970000000
1!
1'
1/
#149980000000
0!
0'
0/
#149990000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#150000000000
0!
0'
0/
#150010000000
1!
1'
1/
#150020000000
0!
0'
0/
#150030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#150040000000
0!
0'
0/
#150050000000
1!
1'
1/
#150060000000
0!
0'
0/
#150070000000
#150080000000
1!
1'
1/
#150090000000
0!
0'
0/
#150100000000
1!
1'
1/
#150110000000
0!
1"
0'
1(
0/
10
#150120000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#150130000000
0!
0'
0/
#150140000000
1!
1'
1/
#150150000000
0!
0'
0/
#150160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#150170000000
0!
0'
0/
#150180000000
1!
1'
1/
#150190000000
0!
1"
0'
1(
0/
10
#150200000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#150210000000
0!
1$
0'
1+
0/
#150220000000
1!
1'
1/
#150230000000
0!
0'
0/
#150240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#150250000000
0!
0'
0/
#150260000000
1!
1'
1/
#150270000000
0!
0'
0/
#150280000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#150290000000
0!
0'
0/
#150300000000
1!
1'
1/
#150310000000
0!
0'
0/
#150320000000
1!
1'
1/
#150330000000
0!
0'
0/
#150340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#150350000000
0!
0'
0/
#150360000000
1!
1'
1/
#150370000000
0!
0'
0/
#150380000000
1!
1'
1/
#150390000000
0!
0'
0/
#150400000000
1!
1'
1/
#150410000000
0!
0'
0/
#150420000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#150430000000
0!
0'
0/
#150440000000
1!
1'
1/
#150450000000
0!
0'
0/
#150460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#150470000000
0!
0'
0/
#150480000000
1!
1'
1/
#150490000000
0!
0'
0/
#150500000000
#150510000000
1!
1'
1/
#150520000000
0!
0'
0/
#150530000000
1!
1'
1/
#150540000000
0!
1"
0'
1(
0/
10
#150550000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#150560000000
0!
0'
0/
#150570000000
1!
1'
1/
#150580000000
0!
0'
0/
#150590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#150600000000
0!
0'
0/
#150610000000
1!
1'
1/
#150620000000
0!
1"
0'
1(
0/
10
#150630000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#150640000000
0!
1$
0'
1+
0/
#150650000000
1!
1'
1/
#150660000000
0!
0'
0/
#150670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#150680000000
0!
0'
0/
#150690000000
1!
1'
1/
#150700000000
0!
0'
0/
#150710000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#150720000000
0!
0'
0/
#150730000000
1!
1'
1/
#150740000000
0!
0'
0/
#150750000000
1!
1'
1/
#150760000000
0!
0'
0/
#150770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#150780000000
0!
0'
0/
#150790000000
1!
1'
1/
#150800000000
0!
0'
0/
#150810000000
1!
1'
1/
#150820000000
0!
0'
0/
#150830000000
1!
1'
1/
#150840000000
0!
0'
0/
#150850000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#150860000000
0!
0'
0/
#150870000000
1!
1'
1/
#150880000000
0!
0'
0/
#150890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#150900000000
0!
0'
0/
#150910000000
1!
1'
1/
#150920000000
0!
0'
0/
#150930000000
#150940000000
1!
1'
1/
#150950000000
0!
0'
0/
#150960000000
1!
1'
1/
#150970000000
0!
1"
0'
1(
0/
10
#150980000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#150990000000
0!
0'
0/
#151000000000
1!
1'
1/
#151010000000
0!
0'
0/
#151020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#151030000000
0!
0'
0/
#151040000000
1!
1'
1/
#151050000000
0!
1"
0'
1(
0/
10
#151060000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#151070000000
0!
1$
0'
1+
0/
#151080000000
1!
1'
1/
#151090000000
0!
0'
0/
#151100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#151110000000
0!
0'
0/
#151120000000
1!
1'
1/
#151130000000
0!
0'
0/
#151140000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#151150000000
0!
0'
0/
#151160000000
1!
1'
1/
#151170000000
0!
0'
0/
#151180000000
1!
1'
1/
#151190000000
0!
0'
0/
#151200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#151210000000
0!
0'
0/
#151220000000
1!
1'
1/
#151230000000
0!
0'
0/
#151240000000
1!
1'
1/
#151250000000
0!
0'
0/
#151260000000
1!
1'
1/
#151270000000
0!
0'
0/
#151280000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#151290000000
0!
0'
0/
#151300000000
1!
1'
1/
#151310000000
0!
0'
0/
#151320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#151330000000
0!
0'
0/
#151340000000
1!
1'
1/
#151350000000
0!
0'
0/
#151360000000
#151370000000
1!
1'
1/
#151380000000
0!
0'
0/
#151390000000
1!
1'
1/
#151400000000
0!
1"
0'
1(
0/
10
#151410000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#151420000000
0!
0'
0/
#151430000000
1!
1'
1/
#151440000000
0!
0'
0/
#151450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#151460000000
0!
0'
0/
#151470000000
1!
1'
1/
#151480000000
0!
1"
0'
1(
0/
10
#151490000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#151500000000
0!
1$
0'
1+
0/
#151510000000
1!
1'
1/
#151520000000
0!
0'
0/
#151530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#151540000000
0!
0'
0/
#151550000000
1!
1'
1/
#151560000000
0!
0'
0/
#151570000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#151580000000
0!
0'
0/
#151590000000
1!
1'
1/
#151600000000
0!
0'
0/
#151610000000
1!
1'
1/
#151620000000
0!
0'
0/
#151630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#151640000000
0!
0'
0/
#151650000000
1!
1'
1/
#151660000000
0!
0'
0/
#151670000000
1!
1'
1/
#151680000000
0!
0'
0/
#151690000000
1!
1'
1/
#151700000000
0!
0'
0/
#151710000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#151720000000
0!
0'
0/
#151730000000
1!
1'
1/
#151740000000
0!
0'
0/
#151750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#151760000000
0!
0'
0/
#151770000000
1!
1'
1/
#151780000000
0!
0'
0/
#151790000000
#151800000000
1!
1'
1/
#151810000000
0!
0'
0/
#151820000000
1!
1'
1/
#151830000000
0!
1"
0'
1(
0/
10
#151840000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#151850000000
0!
0'
0/
#151860000000
1!
1'
1/
#151870000000
0!
0'
0/
#151880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#151890000000
0!
0'
0/
#151900000000
1!
1'
1/
#151910000000
0!
1"
0'
1(
0/
10
#151920000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#151930000000
0!
1$
0'
1+
0/
#151940000000
1!
1'
1/
#151950000000
0!
0'
0/
#151960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#151970000000
0!
0'
0/
#151980000000
1!
1'
1/
#151990000000
0!
0'
0/
#152000000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#152010000000
0!
0'
0/
#152020000000
1!
1'
1/
#152030000000
0!
0'
0/
#152040000000
1!
1'
1/
#152050000000
0!
0'
0/
#152060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#152070000000
0!
0'
0/
#152080000000
1!
1'
1/
#152090000000
0!
0'
0/
#152100000000
1!
1'
1/
#152110000000
0!
0'
0/
#152120000000
1!
1'
1/
#152130000000
0!
0'
0/
#152140000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#152150000000
0!
0'
0/
#152160000000
1!
1'
1/
#152170000000
0!
0'
0/
#152180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#152190000000
0!
0'
0/
#152200000000
1!
1'
1/
#152210000000
0!
0'
0/
#152220000000
#152230000000
1!
1'
1/
#152240000000
0!
0'
0/
#152250000000
1!
1'
1/
#152260000000
0!
1"
0'
1(
0/
10
#152270000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#152280000000
0!
0'
0/
#152290000000
1!
1'
1/
#152300000000
0!
0'
0/
#152310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#152320000000
0!
0'
0/
#152330000000
1!
1'
1/
#152340000000
0!
1"
0'
1(
0/
10
#152350000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#152360000000
0!
1$
0'
1+
0/
#152370000000
1!
1'
1/
#152380000000
0!
0'
0/
#152390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#152400000000
0!
0'
0/
#152410000000
1!
1'
1/
#152420000000
0!
0'
0/
#152430000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#152440000000
0!
0'
0/
#152450000000
1!
1'
1/
#152460000000
0!
0'
0/
#152470000000
1!
1'
1/
#152480000000
0!
0'
0/
#152490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#152500000000
0!
0'
0/
#152510000000
1!
1'
1/
#152520000000
0!
0'
0/
#152530000000
1!
1'
1/
#152540000000
0!
0'
0/
#152550000000
1!
1'
1/
#152560000000
0!
0'
0/
#152570000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#152580000000
0!
0'
0/
#152590000000
1!
1'
1/
#152600000000
0!
0'
0/
#152610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#152620000000
0!
0'
0/
#152630000000
1!
1'
1/
#152640000000
0!
0'
0/
#152650000000
#152660000000
1!
1'
1/
#152670000000
0!
0'
0/
#152680000000
1!
1'
1/
#152690000000
0!
1"
0'
1(
0/
10
#152700000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#152710000000
0!
0'
0/
#152720000000
1!
1'
1/
#152730000000
0!
0'
0/
#152740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#152750000000
0!
0'
0/
#152760000000
1!
1'
1/
#152770000000
0!
1"
0'
1(
0/
10
#152780000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#152790000000
0!
1$
0'
1+
0/
#152800000000
1!
1'
1/
#152810000000
0!
0'
0/
#152820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#152830000000
0!
0'
0/
#152840000000
1!
1'
1/
#152850000000
0!
0'
0/
#152860000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#152870000000
0!
0'
0/
#152880000000
1!
1'
1/
#152890000000
0!
0'
0/
#152900000000
1!
1'
1/
#152910000000
0!
0'
0/
#152920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#152930000000
0!
0'
0/
#152940000000
1!
1'
1/
#152950000000
0!
0'
0/
#152960000000
1!
1'
1/
#152970000000
0!
0'
0/
#152980000000
1!
1'
1/
#152990000000
0!
0'
0/
#153000000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#153010000000
0!
0'
0/
#153020000000
1!
1'
1/
#153030000000
0!
0'
0/
#153040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#153050000000
0!
0'
0/
#153060000000
1!
1'
1/
#153070000000
0!
0'
0/
#153080000000
#153090000000
1!
1'
1/
#153100000000
0!
0'
0/
#153110000000
1!
1'
1/
#153120000000
0!
1"
0'
1(
0/
10
#153130000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#153140000000
0!
0'
0/
#153150000000
1!
1'
1/
#153160000000
0!
0'
0/
#153170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#153180000000
0!
0'
0/
#153190000000
1!
1'
1/
#153200000000
0!
1"
0'
1(
0/
10
#153210000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#153220000000
0!
1$
0'
1+
0/
#153230000000
1!
1'
1/
#153240000000
0!
0'
0/
#153250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#153260000000
0!
0'
0/
#153270000000
1!
1'
1/
#153280000000
0!
0'
0/
#153290000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#153300000000
0!
0'
0/
#153310000000
1!
1'
1/
#153320000000
0!
0'
0/
#153330000000
1!
1'
1/
#153340000000
0!
0'
0/
#153350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#153360000000
0!
0'
0/
#153370000000
1!
1'
1/
#153380000000
0!
0'
0/
#153390000000
1!
1'
1/
#153400000000
0!
0'
0/
#153410000000
1!
1'
1/
#153420000000
0!
0'
0/
#153430000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#153440000000
0!
0'
0/
#153450000000
1!
1'
1/
#153460000000
0!
0'
0/
#153470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#153480000000
0!
0'
0/
#153490000000
1!
1'
1/
#153500000000
0!
0'
0/
#153510000000
#153520000000
1!
1'
1/
#153530000000
0!
0'
0/
#153540000000
1!
1'
1/
#153550000000
0!
1"
0'
1(
0/
10
#153560000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#153570000000
0!
0'
0/
#153580000000
1!
1'
1/
#153590000000
0!
0'
0/
#153600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#153610000000
0!
0'
0/
#153620000000
1!
1'
1/
#153630000000
0!
1"
0'
1(
0/
10
#153640000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#153650000000
0!
1$
0'
1+
0/
#153660000000
1!
1'
1/
#153670000000
0!
0'
0/
#153680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#153690000000
0!
0'
0/
#153700000000
1!
1'
1/
#153710000000
0!
0'
0/
#153720000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#153730000000
0!
0'
0/
#153740000000
1!
1'
1/
#153750000000
0!
0'
0/
#153760000000
1!
1'
1/
#153770000000
0!
0'
0/
#153780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#153790000000
0!
0'
0/
#153800000000
1!
1'
1/
#153810000000
0!
0'
0/
#153820000000
1!
1'
1/
#153830000000
0!
0'
0/
#153840000000
1!
1'
1/
#153850000000
0!
0'
0/
#153860000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#153870000000
0!
0'
0/
#153880000000
1!
1'
1/
#153890000000
0!
0'
0/
#153900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#153910000000
0!
0'
0/
#153920000000
1!
1'
1/
#153930000000
0!
0'
0/
#153940000000
#153950000000
1!
1'
1/
#153960000000
0!
0'
0/
#153970000000
1!
1'
1/
#153980000000
0!
1"
0'
1(
0/
10
#153990000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#154000000000
0!
0'
0/
#154010000000
1!
1'
1/
#154020000000
0!
0'
0/
#154030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#154040000000
0!
0'
0/
#154050000000
1!
1'
1/
#154060000000
0!
1"
0'
1(
0/
10
#154070000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#154080000000
0!
1$
0'
1+
0/
#154090000000
1!
1'
1/
#154100000000
0!
0'
0/
#154110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#154120000000
0!
0'
0/
#154130000000
1!
1'
1/
#154140000000
0!
0'
0/
#154150000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#154160000000
0!
0'
0/
#154170000000
1!
1'
1/
#154180000000
0!
0'
0/
#154190000000
1!
1'
1/
#154200000000
0!
0'
0/
#154210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#154220000000
0!
0'
0/
#154230000000
1!
1'
1/
#154240000000
0!
0'
0/
#154250000000
1!
1'
1/
#154260000000
0!
0'
0/
#154270000000
1!
1'
1/
#154280000000
0!
0'
0/
#154290000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#154300000000
0!
0'
0/
#154310000000
1!
1'
1/
#154320000000
0!
0'
0/
#154330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#154340000000
0!
0'
0/
#154350000000
1!
1'
1/
#154360000000
0!
0'
0/
#154370000000
#154380000000
1!
1'
1/
#154390000000
0!
0'
0/
#154400000000
1!
1'
1/
#154410000000
0!
1"
0'
1(
0/
10
#154420000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#154430000000
0!
0'
0/
#154440000000
1!
1'
1/
#154450000000
0!
0'
0/
#154460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#154470000000
0!
0'
0/
#154480000000
1!
1'
1/
#154490000000
0!
1"
0'
1(
0/
10
#154500000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#154510000000
0!
1$
0'
1+
0/
#154520000000
1!
1'
1/
#154530000000
0!
0'
0/
#154540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#154550000000
0!
0'
0/
#154560000000
1!
1'
1/
#154570000000
0!
0'
0/
#154580000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#154590000000
0!
0'
0/
#154600000000
1!
1'
1/
#154610000000
0!
0'
0/
#154620000000
1!
1'
1/
#154630000000
0!
0'
0/
#154640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#154650000000
0!
0'
0/
#154660000000
1!
1'
1/
#154670000000
0!
0'
0/
#154680000000
1!
1'
1/
#154690000000
0!
0'
0/
#154700000000
1!
1'
1/
#154710000000
0!
0'
0/
#154720000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#154730000000
0!
0'
0/
#154740000000
1!
1'
1/
#154750000000
0!
0'
0/
#154760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#154770000000
0!
0'
0/
#154780000000
1!
1'
1/
#154790000000
0!
0'
0/
#154800000000
#154810000000
1!
1'
1/
#154820000000
0!
0'
0/
#154830000000
1!
1'
1/
#154840000000
0!
1"
0'
1(
0/
10
#154850000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#154860000000
0!
0'
0/
#154870000000
1!
1'
1/
#154880000000
0!
0'
0/
#154890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#154900000000
0!
0'
0/
#154910000000
1!
1'
1/
#154920000000
0!
1"
0'
1(
0/
10
#154930000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#154940000000
0!
1$
0'
1+
0/
#154950000000
1!
1'
1/
#154960000000
0!
0'
0/
#154970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#154980000000
0!
0'
0/
#154990000000
1!
1'
1/
#155000000000
0!
0'
0/
#155010000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#155020000000
0!
0'
0/
#155030000000
1!
1'
1/
#155040000000
0!
0'
0/
#155050000000
1!
1'
1/
#155060000000
0!
0'
0/
#155070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#155080000000
0!
0'
0/
#155090000000
1!
1'
1/
#155100000000
0!
0'
0/
#155110000000
1!
1'
1/
#155120000000
0!
0'
0/
#155130000000
1!
1'
1/
#155140000000
0!
0'
0/
#155150000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#155160000000
0!
0'
0/
#155170000000
1!
1'
1/
#155180000000
0!
0'
0/
#155190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#155200000000
0!
0'
0/
#155210000000
1!
1'
1/
#155220000000
0!
0'
0/
#155230000000
#155240000000
1!
1'
1/
#155250000000
0!
0'
0/
#155260000000
1!
1'
1/
#155270000000
0!
1"
0'
1(
0/
10
#155280000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#155290000000
0!
0'
0/
#155300000000
1!
1'
1/
#155310000000
0!
0'
0/
#155320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#155330000000
0!
0'
0/
#155340000000
1!
1'
1/
#155350000000
0!
1"
0'
1(
0/
10
#155360000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#155370000000
0!
1$
0'
1+
0/
#155380000000
1!
1'
1/
#155390000000
0!
0'
0/
#155400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#155410000000
0!
0'
0/
#155420000000
1!
1'
1/
#155430000000
0!
0'
0/
#155440000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#155450000000
0!
0'
0/
#155460000000
1!
1'
1/
#155470000000
0!
0'
0/
#155480000000
1!
1'
1/
#155490000000
0!
0'
0/
#155500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#155510000000
0!
0'
0/
#155520000000
1!
1'
1/
#155530000000
0!
0'
0/
#155540000000
1!
1'
1/
#155550000000
0!
0'
0/
#155560000000
1!
1'
1/
#155570000000
0!
0'
0/
#155580000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#155590000000
0!
0'
0/
#155600000000
1!
1'
1/
#155610000000
0!
0'
0/
#155620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#155630000000
0!
0'
0/
#155640000000
1!
1'
1/
#155650000000
0!
0'
0/
#155660000000
#155670000000
1!
1'
1/
#155680000000
0!
0'
0/
#155690000000
1!
1'
1/
#155700000000
0!
1"
0'
1(
0/
10
#155710000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#155720000000
0!
0'
0/
#155730000000
1!
1'
1/
#155740000000
0!
0'
0/
#155750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#155760000000
0!
0'
0/
#155770000000
1!
1'
1/
#155780000000
0!
1"
0'
1(
0/
10
#155790000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#155800000000
0!
1$
0'
1+
0/
#155810000000
1!
1'
1/
#155820000000
0!
0'
0/
#155830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#155840000000
0!
0'
0/
#155850000000
1!
1'
1/
#155860000000
0!
0'
0/
#155870000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#155880000000
0!
0'
0/
#155890000000
1!
1'
1/
#155900000000
0!
0'
0/
#155910000000
1!
1'
1/
#155920000000
0!
0'
0/
#155930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#155940000000
0!
0'
0/
#155950000000
1!
1'
1/
#155960000000
0!
0'
0/
#155970000000
1!
1'
1/
#155980000000
0!
0'
0/
#155990000000
1!
1'
1/
#156000000000
0!
0'
0/
#156010000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#156020000000
0!
0'
0/
#156030000000
1!
1'
1/
#156040000000
0!
0'
0/
#156050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#156060000000
0!
0'
0/
#156070000000
1!
1'
1/
#156080000000
0!
0'
0/
#156090000000
#156100000000
1!
1'
1/
#156110000000
0!
0'
0/
#156120000000
1!
1'
1/
#156130000000
0!
1"
0'
1(
0/
10
#156140000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#156150000000
0!
0'
0/
#156160000000
1!
1'
1/
#156170000000
0!
0'
0/
#156180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#156190000000
0!
0'
0/
#156200000000
1!
1'
1/
#156210000000
0!
1"
0'
1(
0/
10
#156220000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#156230000000
0!
1$
0'
1+
0/
#156240000000
1!
1'
1/
#156250000000
0!
0'
0/
#156260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#156270000000
0!
0'
0/
#156280000000
1!
1'
1/
#156290000000
0!
0'
0/
#156300000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#156310000000
0!
0'
0/
#156320000000
1!
1'
1/
#156330000000
0!
0'
0/
#156340000000
1!
1'
1/
#156350000000
0!
0'
0/
#156360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#156370000000
0!
0'
0/
#156380000000
1!
1'
1/
#156390000000
0!
0'
0/
#156400000000
1!
1'
1/
#156410000000
0!
0'
0/
#156420000000
1!
1'
1/
#156430000000
0!
0'
0/
#156440000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#156450000000
0!
0'
0/
#156460000000
1!
1'
1/
#156470000000
0!
0'
0/
#156480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#156490000000
0!
0'
0/
#156500000000
1!
1'
1/
#156510000000
0!
0'
0/
#156520000000
#156530000000
1!
1'
1/
#156540000000
0!
0'
0/
#156550000000
1!
1'
1/
#156560000000
0!
1"
0'
1(
0/
10
#156570000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#156580000000
0!
0'
0/
#156590000000
1!
1'
1/
#156600000000
0!
0'
0/
#156610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#156620000000
0!
0'
0/
#156630000000
1!
1'
1/
#156640000000
0!
1"
0'
1(
0/
10
#156650000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#156660000000
0!
1$
0'
1+
0/
#156670000000
1!
1'
1/
#156680000000
0!
0'
0/
#156690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#156700000000
0!
0'
0/
#156710000000
1!
1'
1/
#156720000000
0!
0'
0/
#156730000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#156740000000
0!
0'
0/
#156750000000
1!
1'
1/
#156760000000
0!
0'
0/
#156770000000
1!
1'
1/
#156780000000
0!
0'
0/
#156790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#156800000000
0!
0'
0/
#156810000000
1!
1'
1/
#156820000000
0!
0'
0/
#156830000000
1!
1'
1/
#156840000000
0!
0'
0/
#156850000000
1!
1'
1/
#156860000000
0!
0'
0/
#156870000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#156880000000
0!
0'
0/
#156890000000
1!
1'
1/
#156900000000
0!
0'
0/
#156910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#156920000000
0!
0'
0/
#156930000000
1!
1'
1/
#156940000000
0!
0'
0/
#156950000000
#156960000000
1!
1'
1/
#156970000000
0!
0'
0/
#156980000000
1!
1'
1/
#156990000000
0!
1"
0'
1(
0/
10
#157000000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#157010000000
0!
0'
0/
#157020000000
1!
1'
1/
#157030000000
0!
0'
0/
#157040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#157050000000
0!
0'
0/
#157060000000
1!
1'
1/
#157070000000
0!
1"
0'
1(
0/
10
#157080000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#157090000000
0!
1$
0'
1+
0/
#157100000000
1!
1'
1/
#157110000000
0!
0'
0/
#157120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#157130000000
0!
0'
0/
#157140000000
1!
1'
1/
#157150000000
0!
0'
0/
#157160000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#157170000000
0!
0'
0/
#157180000000
1!
1'
1/
#157190000000
0!
0'
0/
#157200000000
1!
1'
1/
#157210000000
0!
0'
0/
#157220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#157230000000
0!
0'
0/
#157240000000
1!
1'
1/
#157250000000
0!
0'
0/
#157260000000
1!
1'
1/
#157270000000
0!
0'
0/
#157280000000
1!
1'
1/
#157290000000
0!
0'
0/
#157300000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#157310000000
0!
0'
0/
#157320000000
1!
1'
1/
#157330000000
0!
0'
0/
#157340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#157350000000
0!
0'
0/
#157360000000
1!
1'
1/
#157370000000
0!
0'
0/
#157380000000
#157390000000
1!
1'
1/
#157400000000
0!
0'
0/
#157410000000
1!
1'
1/
#157420000000
0!
1"
0'
1(
0/
10
#157430000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#157440000000
0!
0'
0/
#157450000000
1!
1'
1/
#157460000000
0!
0'
0/
#157470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#157480000000
0!
0'
0/
#157490000000
1!
1'
1/
#157500000000
0!
1"
0'
1(
0/
10
#157510000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#157520000000
0!
1$
0'
1+
0/
#157530000000
1!
1'
1/
#157540000000
0!
0'
0/
#157550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#157560000000
0!
0'
0/
#157570000000
1!
1'
1/
#157580000000
0!
0'
0/
#157590000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#157600000000
0!
0'
0/
#157610000000
1!
1'
1/
#157620000000
0!
0'
0/
#157630000000
1!
1'
1/
#157640000000
0!
0'
0/
#157650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#157660000000
0!
0'
0/
#157670000000
1!
1'
1/
#157680000000
0!
0'
0/
#157690000000
1!
1'
1/
#157700000000
0!
0'
0/
#157710000000
1!
1'
1/
#157720000000
0!
0'
0/
#157730000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#157740000000
0!
0'
0/
#157750000000
1!
1'
1/
#157760000000
0!
0'
0/
#157770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#157780000000
0!
0'
0/
#157790000000
1!
1'
1/
#157800000000
0!
0'
0/
#157810000000
#157820000000
1!
1'
1/
#157830000000
0!
0'
0/
#157840000000
1!
1'
1/
#157850000000
0!
1"
0'
1(
0/
10
#157860000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#157870000000
0!
0'
0/
#157880000000
1!
1'
1/
#157890000000
0!
0'
0/
#157900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#157910000000
0!
0'
0/
#157920000000
1!
1'
1/
#157930000000
0!
1"
0'
1(
0/
10
#157940000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#157950000000
0!
1$
0'
1+
0/
#157960000000
1!
1'
1/
#157970000000
0!
0'
0/
#157980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#157990000000
0!
0'
0/
#158000000000
1!
1'
1/
#158010000000
0!
0'
0/
#158020000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#158030000000
0!
0'
0/
#158040000000
1!
1'
1/
#158050000000
0!
0'
0/
#158060000000
1!
1'
1/
#158070000000
0!
0'
0/
#158080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#158090000000
0!
0'
0/
#158100000000
1!
1'
1/
#158110000000
0!
0'
0/
#158120000000
1!
1'
1/
#158130000000
0!
0'
0/
#158140000000
1!
1'
1/
#158150000000
0!
0'
0/
#158160000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#158170000000
0!
0'
0/
#158180000000
1!
1'
1/
#158190000000
0!
0'
0/
#158200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#158210000000
0!
0'
0/
#158220000000
1!
1'
1/
#158230000000
0!
0'
0/
#158240000000
#158250000000
1!
1'
1/
#158260000000
0!
0'
0/
#158270000000
1!
1'
1/
#158280000000
0!
1"
0'
1(
0/
10
#158290000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#158300000000
0!
0'
0/
#158310000000
1!
1'
1/
#158320000000
0!
0'
0/
#158330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#158340000000
0!
0'
0/
#158350000000
1!
1'
1/
#158360000000
0!
1"
0'
1(
0/
10
#158370000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#158380000000
0!
1$
0'
1+
0/
#158390000000
1!
1'
1/
#158400000000
0!
0'
0/
#158410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#158420000000
0!
0'
0/
#158430000000
1!
1'
1/
#158440000000
0!
0'
0/
#158450000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#158460000000
0!
0'
0/
#158470000000
1!
1'
1/
#158480000000
0!
0'
0/
#158490000000
1!
1'
1/
#158500000000
0!
0'
0/
#158510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#158520000000
0!
0'
0/
#158530000000
1!
1'
1/
#158540000000
0!
0'
0/
#158550000000
1!
1'
1/
#158560000000
0!
0'
0/
#158570000000
1!
1'
1/
#158580000000
0!
0'
0/
#158590000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#158600000000
0!
0'
0/
#158610000000
1!
1'
1/
#158620000000
0!
0'
0/
#158630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#158640000000
0!
0'
0/
#158650000000
1!
1'
1/
#158660000000
0!
0'
0/
#158670000000
#158680000000
1!
1'
1/
#158690000000
0!
0'
0/
#158700000000
1!
1'
1/
#158710000000
0!
1"
0'
1(
0/
10
#158720000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#158730000000
0!
0'
0/
#158740000000
1!
1'
1/
#158750000000
0!
0'
0/
#158760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#158770000000
0!
0'
0/
#158780000000
1!
1'
1/
#158790000000
0!
1"
0'
1(
0/
10
#158800000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#158810000000
0!
1$
0'
1+
0/
#158820000000
1!
1'
1/
#158830000000
0!
0'
0/
#158840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#158850000000
0!
0'
0/
#158860000000
1!
1'
1/
#158870000000
0!
0'
0/
#158880000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#158890000000
0!
0'
0/
#158900000000
1!
1'
1/
#158910000000
0!
0'
0/
#158920000000
1!
1'
1/
#158930000000
0!
0'
0/
#158940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#158950000000
0!
0'
0/
#158960000000
1!
1'
1/
#158970000000
0!
0'
0/
#158980000000
1!
1'
1/
#158990000000
0!
0'
0/
#159000000000
1!
1'
1/
#159010000000
0!
0'
0/
#159020000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#159030000000
0!
0'
0/
#159040000000
1!
1'
1/
#159050000000
0!
0'
0/
#159060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#159070000000
0!
0'
0/
#159080000000
1!
1'
1/
#159090000000
0!
0'
0/
#159100000000
#159110000000
1!
1'
1/
#159120000000
0!
0'
0/
#159130000000
1!
1'
1/
#159140000000
0!
1"
0'
1(
0/
10
#159150000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#159160000000
0!
0'
0/
#159170000000
1!
1'
1/
#159180000000
0!
0'
0/
#159190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#159200000000
0!
0'
0/
#159210000000
1!
1'
1/
#159220000000
0!
1"
0'
1(
0/
10
#159230000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#159240000000
0!
1$
0'
1+
0/
#159250000000
1!
1'
1/
#159260000000
0!
0'
0/
#159270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#159280000000
0!
0'
0/
#159290000000
1!
1'
1/
#159300000000
0!
0'
0/
#159310000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#159320000000
0!
0'
0/
#159330000000
1!
1'
1/
#159340000000
0!
0'
0/
#159350000000
1!
1'
1/
#159360000000
0!
0'
0/
#159370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#159380000000
0!
0'
0/
#159390000000
1!
1'
1/
#159400000000
0!
0'
0/
#159410000000
1!
1'
1/
#159420000000
0!
0'
0/
#159430000000
1!
1'
1/
#159440000000
0!
0'
0/
#159450000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#159460000000
0!
0'
0/
#159470000000
1!
1'
1/
#159480000000
0!
0'
0/
#159490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#159500000000
0!
0'
0/
#159510000000
1!
1'
1/
#159520000000
0!
0'
0/
#159530000000
#159540000000
1!
1'
1/
#159550000000
0!
0'
0/
#159560000000
1!
1'
1/
#159570000000
0!
1"
0'
1(
0/
10
#159580000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#159590000000
0!
0'
0/
#159600000000
1!
1'
1/
#159610000000
0!
0'
0/
#159620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#159630000000
0!
0'
0/
#159640000000
1!
1'
1/
#159650000000
0!
1"
0'
1(
0/
10
#159660000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#159670000000
0!
1$
0'
1+
0/
#159680000000
1!
1'
1/
#159690000000
0!
0'
0/
#159700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#159710000000
0!
0'
0/
#159720000000
1!
1'
1/
#159730000000
0!
0'
0/
#159740000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#159750000000
0!
0'
0/
#159760000000
1!
1'
1/
#159770000000
0!
0'
0/
#159780000000
1!
1'
1/
#159790000000
0!
0'
0/
#159800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#159810000000
0!
0'
0/
#159820000000
1!
1'
1/
#159830000000
0!
0'
0/
#159840000000
1!
1'
1/
#159850000000
0!
0'
0/
#159860000000
1!
1'
1/
#159870000000
0!
0'
0/
#159880000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#159890000000
0!
0'
0/
#159900000000
1!
1'
1/
#159910000000
0!
0'
0/
#159920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#159930000000
0!
0'
0/
#159940000000
1!
1'
1/
#159950000000
0!
0'
0/
#159960000000
#159970000000
1!
1'
1/
#159980000000
0!
0'
0/
#159990000000
1!
1'
1/
#160000000000
0!
1"
0'
1(
0/
10
#160010000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#160020000000
0!
0'
0/
#160030000000
1!
1'
1/
#160040000000
0!
0'
0/
#160050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#160060000000
0!
0'
0/
#160070000000
1!
1'
1/
#160080000000
0!
1"
0'
1(
0/
10
#160090000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#160100000000
0!
1$
0'
1+
0/
#160110000000
1!
1'
1/
#160120000000
0!
0'
0/
#160130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#160140000000
0!
0'
0/
#160150000000
1!
1'
1/
#160160000000
0!
0'
0/
#160170000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#160180000000
0!
0'
0/
#160190000000
1!
1'
1/
#160200000000
0!
0'
0/
#160210000000
1!
1'
1/
#160220000000
0!
0'
0/
#160230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#160240000000
0!
0'
0/
#160250000000
1!
1'
1/
#160260000000
0!
0'
0/
#160270000000
1!
1'
1/
#160280000000
0!
0'
0/
#160290000000
1!
1'
1/
#160300000000
0!
0'
0/
#160310000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#160320000000
0!
0'
0/
#160330000000
1!
1'
1/
#160340000000
0!
0'
0/
#160350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#160360000000
0!
0'
0/
#160370000000
1!
1'
1/
#160380000000
0!
0'
0/
#160390000000
#160400000000
1!
1'
1/
#160410000000
0!
0'
0/
#160420000000
1!
1'
1/
#160430000000
0!
1"
0'
1(
0/
10
#160440000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#160450000000
0!
0'
0/
#160460000000
1!
1'
1/
#160470000000
0!
0'
0/
#160480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#160490000000
0!
0'
0/
#160500000000
1!
1'
1/
#160510000000
0!
1"
0'
1(
0/
10
#160520000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#160530000000
0!
1$
0'
1+
0/
#160540000000
1!
1'
1/
#160550000000
0!
0'
0/
#160560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#160570000000
0!
0'
0/
#160580000000
1!
1'
1/
#160590000000
0!
0'
0/
#160600000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#160610000000
0!
0'
0/
#160620000000
1!
1'
1/
#160630000000
0!
0'
0/
#160640000000
1!
1'
1/
#160650000000
0!
0'
0/
#160660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#160670000000
0!
0'
0/
#160680000000
1!
1'
1/
#160690000000
0!
0'
0/
#160700000000
1!
1'
1/
#160710000000
0!
0'
0/
#160720000000
1!
1'
1/
#160730000000
0!
0'
0/
#160740000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#160750000000
0!
0'
0/
#160760000000
1!
1'
1/
#160770000000
0!
0'
0/
#160780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#160790000000
0!
0'
0/
#160800000000
1!
1'
1/
#160810000000
0!
0'
0/
#160820000000
#160830000000
1!
1'
1/
#160840000000
0!
0'
0/
#160850000000
1!
1'
1/
#160860000000
0!
1"
0'
1(
0/
10
#160870000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#160880000000
0!
0'
0/
#160890000000
1!
1'
1/
#160900000000
0!
0'
0/
#160910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#160920000000
0!
0'
0/
#160930000000
1!
1'
1/
#160940000000
0!
1"
0'
1(
0/
10
#160950000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#160960000000
0!
1$
0'
1+
0/
#160970000000
1!
1'
1/
#160980000000
0!
0'
0/
#160990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#161000000000
0!
0'
0/
#161010000000
1!
1'
1/
#161020000000
0!
0'
0/
#161030000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#161040000000
0!
0'
0/
#161050000000
1!
1'
1/
#161060000000
0!
0'
0/
#161070000000
1!
1'
1/
#161080000000
0!
0'
0/
#161090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#161100000000
0!
0'
0/
#161110000000
1!
1'
1/
#161120000000
0!
0'
0/
#161130000000
1!
1'
1/
#161140000000
0!
0'
0/
#161150000000
1!
1'
1/
#161160000000
0!
0'
0/
#161170000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#161180000000
0!
0'
0/
#161190000000
1!
1'
1/
#161200000000
0!
0'
0/
#161210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#161220000000
0!
0'
0/
#161230000000
1!
1'
1/
#161240000000
0!
0'
0/
#161250000000
#161260000000
1!
1'
1/
#161270000000
0!
0'
0/
#161280000000
1!
1'
1/
#161290000000
0!
1"
0'
1(
0/
10
#161300000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#161310000000
0!
0'
0/
#161320000000
1!
1'
1/
#161330000000
0!
0'
0/
#161340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#161350000000
0!
0'
0/
#161360000000
1!
1'
1/
#161370000000
0!
1"
0'
1(
0/
10
#161380000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#161390000000
0!
1$
0'
1+
0/
#161400000000
1!
1'
1/
#161410000000
0!
0'
0/
#161420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#161430000000
0!
0'
0/
#161440000000
1!
1'
1/
#161450000000
0!
0'
0/
#161460000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#161470000000
0!
0'
0/
#161480000000
1!
1'
1/
#161490000000
0!
0'
0/
#161500000000
1!
1'
1/
#161510000000
0!
0'
0/
#161520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#161530000000
0!
0'
0/
#161540000000
1!
1'
1/
#161550000000
0!
0'
0/
#161560000000
1!
1'
1/
#161570000000
0!
0'
0/
#161580000000
1!
1'
1/
#161590000000
0!
0'
0/
#161600000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#161610000000
0!
0'
0/
#161620000000
1!
1'
1/
#161630000000
0!
0'
0/
#161640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#161650000000
0!
0'
0/
#161660000000
1!
1'
1/
#161670000000
0!
0'
0/
#161680000000
#161690000000
1!
1'
1/
#161700000000
0!
0'
0/
#161710000000
1!
1'
1/
#161720000000
0!
1"
0'
1(
0/
10
#161730000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#161740000000
0!
0'
0/
#161750000000
1!
1'
1/
#161760000000
0!
0'
0/
#161770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#161780000000
0!
0'
0/
#161790000000
1!
1'
1/
#161800000000
0!
1"
0'
1(
0/
10
#161810000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#161820000000
0!
1$
0'
1+
0/
#161830000000
1!
1'
1/
#161840000000
0!
0'
0/
#161850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#161860000000
0!
0'
0/
#161870000000
1!
1'
1/
#161880000000
0!
0'
0/
#161890000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#161900000000
0!
0'
0/
#161910000000
1!
1'
1/
#161920000000
0!
0'
0/
#161930000000
1!
1'
1/
#161940000000
0!
0'
0/
#161950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#161960000000
0!
0'
0/
#161970000000
1!
1'
1/
#161980000000
0!
0'
0/
#161990000000
1!
1'
1/
#162000000000
0!
0'
0/
#162010000000
1!
1'
1/
#162020000000
0!
0'
0/
#162030000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#162040000000
0!
0'
0/
#162050000000
1!
1'
1/
#162060000000
0!
0'
0/
#162070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#162080000000
0!
0'
0/
#162090000000
1!
1'
1/
#162100000000
0!
0'
0/
#162110000000
#162120000000
1!
1'
1/
#162130000000
0!
0'
0/
#162140000000
1!
1'
1/
#162150000000
0!
1"
0'
1(
0/
10
#162160000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#162170000000
0!
0'
0/
#162180000000
1!
1'
1/
#162190000000
0!
0'
0/
#162200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#162210000000
0!
0'
0/
#162220000000
1!
1'
1/
#162230000000
0!
1"
0'
1(
0/
10
#162240000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#162250000000
0!
1$
0'
1+
0/
#162260000000
1!
1'
1/
#162270000000
0!
0'
0/
#162280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#162290000000
0!
0'
0/
#162300000000
1!
1'
1/
#162310000000
0!
0'
0/
#162320000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#162330000000
0!
0'
0/
#162340000000
1!
1'
1/
#162350000000
0!
0'
0/
#162360000000
1!
1'
1/
#162370000000
0!
0'
0/
#162380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#162390000000
0!
0'
0/
#162400000000
1!
1'
1/
#162410000000
0!
0'
0/
#162420000000
1!
1'
1/
#162430000000
0!
0'
0/
#162440000000
1!
1'
1/
#162450000000
0!
0'
0/
#162460000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#162470000000
0!
0'
0/
#162480000000
1!
1'
1/
#162490000000
0!
0'
0/
#162500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#162510000000
0!
0'
0/
#162520000000
1!
1'
1/
#162530000000
0!
0'
0/
#162540000000
#162550000000
1!
1'
1/
#162560000000
0!
0'
0/
#162570000000
1!
1'
1/
#162580000000
0!
1"
0'
1(
0/
10
#162590000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#162600000000
0!
0'
0/
#162610000000
1!
1'
1/
#162620000000
0!
0'
0/
#162630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#162640000000
0!
0'
0/
#162650000000
1!
1'
1/
#162660000000
0!
1"
0'
1(
0/
10
#162670000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#162680000000
0!
1$
0'
1+
0/
#162690000000
1!
1'
1/
#162700000000
0!
0'
0/
#162710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#162720000000
0!
0'
0/
#162730000000
1!
1'
1/
#162740000000
0!
0'
0/
#162750000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#162760000000
0!
0'
0/
#162770000000
1!
1'
1/
#162780000000
0!
0'
0/
#162790000000
1!
1'
1/
#162800000000
0!
0'
0/
#162810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#162820000000
0!
0'
0/
#162830000000
1!
1'
1/
#162840000000
0!
0'
0/
#162850000000
1!
1'
1/
#162860000000
0!
0'
0/
#162870000000
1!
1'
1/
#162880000000
0!
0'
0/
#162890000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#162900000000
0!
0'
0/
#162910000000
1!
1'
1/
#162920000000
0!
0'
0/
#162930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#162940000000
0!
0'
0/
#162950000000
1!
1'
1/
#162960000000
0!
0'
0/
#162970000000
#162980000000
1!
1'
1/
#162990000000
0!
0'
0/
#163000000000
1!
1'
1/
#163010000000
0!
1"
0'
1(
0/
10
#163020000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#163030000000
0!
0'
0/
#163040000000
1!
1'
1/
#163050000000
0!
0'
0/
#163060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#163070000000
0!
0'
0/
#163080000000
1!
1'
1/
#163090000000
0!
1"
0'
1(
0/
10
#163100000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#163110000000
0!
1$
0'
1+
0/
#163120000000
1!
1'
1/
#163130000000
0!
0'
0/
#163140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#163150000000
0!
0'
0/
#163160000000
1!
1'
1/
#163170000000
0!
0'
0/
#163180000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#163190000000
0!
0'
0/
#163200000000
1!
1'
1/
#163210000000
0!
0'
0/
#163220000000
1!
1'
1/
#163230000000
0!
0'
0/
#163240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#163250000000
0!
0'
0/
#163260000000
1!
1'
1/
#163270000000
0!
0'
0/
#163280000000
1!
1'
1/
#163290000000
0!
0'
0/
#163300000000
1!
1'
1/
#163310000000
0!
0'
0/
#163320000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#163330000000
0!
0'
0/
#163340000000
1!
1'
1/
#163350000000
0!
0'
0/
#163360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#163370000000
0!
0'
0/
#163380000000
1!
1'
1/
#163390000000
0!
0'
0/
#163400000000
#163410000000
1!
1'
1/
#163420000000
0!
0'
0/
#163430000000
1!
1'
1/
#163440000000
0!
1"
0'
1(
0/
10
#163450000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#163460000000
0!
0'
0/
#163470000000
1!
1'
1/
#163480000000
0!
0'
0/
#163490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#163500000000
0!
0'
0/
#163510000000
1!
1'
1/
#163520000000
0!
1"
0'
1(
0/
10
#163530000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#163540000000
0!
1$
0'
1+
0/
#163550000000
1!
1'
1/
#163560000000
0!
0'
0/
#163570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#163580000000
0!
0'
0/
#163590000000
1!
1'
1/
#163600000000
0!
0'
0/
#163610000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#163620000000
0!
0'
0/
#163630000000
1!
1'
1/
#163640000000
0!
0'
0/
#163650000000
1!
1'
1/
#163660000000
0!
0'
0/
#163670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#163680000000
0!
0'
0/
#163690000000
1!
1'
1/
#163700000000
0!
0'
0/
#163710000000
1!
1'
1/
#163720000000
0!
0'
0/
#163730000000
1!
1'
1/
#163740000000
0!
0'
0/
#163750000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#163760000000
0!
0'
0/
#163770000000
1!
1'
1/
#163780000000
0!
0'
0/
#163790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#163800000000
0!
0'
0/
#163810000000
1!
1'
1/
#163820000000
0!
0'
0/
#163830000000
#163840000000
1!
1'
1/
#163850000000
0!
0'
0/
#163860000000
1!
1'
1/
#163870000000
0!
1"
0'
1(
0/
10
#163880000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#163890000000
0!
0'
0/
#163900000000
1!
1'
1/
#163910000000
0!
0'
0/
#163920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#163930000000
0!
0'
0/
#163940000000
1!
1'
1/
#163950000000
0!
1"
0'
1(
0/
10
#163960000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#163970000000
0!
1$
0'
1+
0/
#163980000000
1!
1'
1/
#163990000000
0!
0'
0/
#164000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#164010000000
0!
0'
0/
#164020000000
1!
1'
1/
#164030000000
0!
0'
0/
#164040000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#164050000000
0!
0'
0/
#164060000000
1!
1'
1/
#164070000000
0!
0'
0/
#164080000000
1!
1'
1/
#164090000000
0!
0'
0/
#164100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#164110000000
0!
0'
0/
#164120000000
1!
1'
1/
#164130000000
0!
0'
0/
#164140000000
1!
1'
1/
#164150000000
0!
0'
0/
#164160000000
1!
1'
1/
#164170000000
0!
0'
0/
#164180000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#164190000000
0!
0'
0/
#164200000000
1!
1'
1/
#164210000000
0!
0'
0/
#164220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#164230000000
0!
0'
0/
#164240000000
1!
1'
1/
#164250000000
0!
0'
0/
#164260000000
#164270000000
1!
1'
1/
#164280000000
0!
0'
0/
#164290000000
1!
1'
1/
#164300000000
0!
1"
0'
1(
0/
10
#164310000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#164320000000
0!
0'
0/
#164330000000
1!
1'
1/
#164340000000
0!
0'
0/
#164350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#164360000000
0!
0'
0/
#164370000000
1!
1'
1/
#164380000000
0!
1"
0'
1(
0/
10
#164390000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#164400000000
0!
1$
0'
1+
0/
#164410000000
1!
1'
1/
#164420000000
0!
0'
0/
#164430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#164440000000
0!
0'
0/
#164450000000
1!
1'
1/
#164460000000
0!
0'
0/
#164470000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#164480000000
0!
0'
0/
#164490000000
1!
1'
1/
#164500000000
0!
0'
0/
#164510000000
1!
1'
1/
#164520000000
0!
0'
0/
#164530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#164540000000
0!
0'
0/
#164550000000
1!
1'
1/
#164560000000
0!
0'
0/
#164570000000
1!
1'
1/
#164580000000
0!
0'
0/
#164590000000
1!
1'
1/
#164600000000
0!
0'
0/
#164610000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#164620000000
0!
0'
0/
#164630000000
1!
1'
1/
#164640000000
0!
0'
0/
#164650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#164660000000
0!
0'
0/
#164670000000
1!
1'
1/
#164680000000
0!
0'
0/
#164690000000
#164700000000
1!
1'
1/
#164710000000
0!
0'
0/
#164720000000
1!
1'
1/
#164730000000
0!
1"
0'
1(
0/
10
#164740000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#164750000000
0!
0'
0/
#164760000000
1!
1'
1/
#164770000000
0!
0'
0/
#164780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#164790000000
0!
0'
0/
#164800000000
1!
1'
1/
#164810000000
0!
1"
0'
1(
0/
10
#164820000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#164830000000
0!
1$
0'
1+
0/
#164840000000
1!
1'
1/
#164850000000
0!
0'
0/
#164860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#164870000000
0!
0'
0/
#164880000000
1!
1'
1/
#164890000000
0!
0'
0/
#164900000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#164910000000
0!
0'
0/
#164920000000
1!
1'
1/
#164930000000
0!
0'
0/
#164940000000
1!
1'
1/
#164950000000
0!
0'
0/
#164960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#164970000000
0!
0'
0/
#164980000000
1!
1'
1/
#164990000000
0!
0'
0/
#165000000000
1!
1'
1/
#165010000000
0!
0'
0/
#165020000000
1!
1'
1/
#165030000000
0!
0'
0/
#165040000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#165050000000
0!
0'
0/
#165060000000
1!
1'
1/
#165070000000
0!
0'
0/
#165080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#165090000000
0!
0'
0/
#165100000000
1!
1'
1/
#165110000000
0!
0'
0/
#165120000000
#165130000000
1!
1'
1/
#165140000000
0!
0'
0/
#165150000000
1!
1'
1/
#165160000000
0!
1"
0'
1(
0/
10
#165170000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#165180000000
0!
0'
0/
#165190000000
1!
1'
1/
#165200000000
0!
0'
0/
#165210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#165220000000
0!
0'
0/
#165230000000
1!
1'
1/
#165240000000
0!
1"
0'
1(
0/
10
#165250000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#165260000000
0!
1$
0'
1+
0/
#165270000000
1!
1'
1/
#165280000000
0!
0'
0/
#165290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#165300000000
0!
0'
0/
#165310000000
1!
1'
1/
#165320000000
0!
0'
0/
#165330000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#165340000000
0!
0'
0/
#165350000000
1!
1'
1/
#165360000000
0!
0'
0/
#165370000000
1!
1'
1/
#165380000000
0!
0'
0/
#165390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#165400000000
0!
0'
0/
#165410000000
1!
1'
1/
#165420000000
0!
0'
0/
#165430000000
1!
1'
1/
#165440000000
0!
0'
0/
#165450000000
1!
1'
1/
#165460000000
0!
0'
0/
#165470000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#165480000000
0!
0'
0/
#165490000000
1!
1'
1/
#165500000000
0!
0'
0/
#165510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#165520000000
0!
0'
0/
#165530000000
1!
1'
1/
#165540000000
0!
0'
0/
#165550000000
#165560000000
1!
1'
1/
#165570000000
0!
0'
0/
#165580000000
1!
1'
1/
#165590000000
0!
1"
0'
1(
0/
10
#165600000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#165610000000
0!
0'
0/
#165620000000
1!
1'
1/
#165630000000
0!
0'
0/
#165640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#165650000000
0!
0'
0/
#165660000000
1!
1'
1/
#165670000000
0!
1"
0'
1(
0/
10
#165680000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#165690000000
0!
1$
0'
1+
0/
#165700000000
1!
1'
1/
#165710000000
0!
0'
0/
#165720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#165730000000
0!
0'
0/
#165740000000
1!
1'
1/
#165750000000
0!
0'
0/
#165760000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#165770000000
0!
0'
0/
#165780000000
1!
1'
1/
#165790000000
0!
0'
0/
#165800000000
1!
1'
1/
#165810000000
0!
0'
0/
#165820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#165830000000
0!
0'
0/
#165840000000
1!
1'
1/
#165850000000
0!
0'
0/
#165860000000
1!
1'
1/
#165870000000
0!
0'
0/
#165880000000
1!
1'
1/
#165890000000
0!
0'
0/
#165900000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#165910000000
0!
0'
0/
#165920000000
1!
1'
1/
#165930000000
0!
0'
0/
#165940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#165950000000
0!
0'
0/
#165960000000
1!
1'
1/
#165970000000
0!
0'
0/
#165980000000
#165990000000
1!
1'
1/
#166000000000
0!
0'
0/
#166010000000
1!
1'
1/
#166020000000
0!
1"
0'
1(
0/
10
#166030000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#166040000000
0!
0'
0/
#166050000000
1!
1'
1/
#166060000000
0!
0'
0/
#166070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#166080000000
0!
0'
0/
#166090000000
1!
1'
1/
#166100000000
0!
1"
0'
1(
0/
10
#166110000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#166120000000
0!
1$
0'
1+
0/
#166130000000
1!
1'
1/
#166140000000
0!
0'
0/
#166150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#166160000000
0!
0'
0/
#166170000000
1!
1'
1/
#166180000000
0!
0'
0/
#166190000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#166200000000
0!
0'
0/
#166210000000
1!
1'
1/
#166220000000
0!
0'
0/
#166230000000
1!
1'
1/
#166240000000
0!
0'
0/
#166250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#166260000000
0!
0'
0/
#166270000000
1!
1'
1/
#166280000000
0!
0'
0/
#166290000000
1!
1'
1/
#166300000000
0!
0'
0/
#166310000000
1!
1'
1/
#166320000000
0!
0'
0/
#166330000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#166340000000
0!
0'
0/
#166350000000
1!
1'
1/
#166360000000
0!
0'
0/
#166370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#166380000000
0!
0'
0/
#166390000000
1!
1'
1/
#166400000000
0!
0'
0/
#166410000000
#166420000000
1!
1'
1/
#166430000000
0!
0'
0/
#166440000000
1!
1'
1/
#166450000000
0!
1"
0'
1(
0/
10
#166460000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#166470000000
0!
0'
0/
#166480000000
1!
1'
1/
#166490000000
0!
0'
0/
#166500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#166510000000
0!
0'
0/
#166520000000
1!
1'
1/
#166530000000
0!
1"
0'
1(
0/
10
#166540000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#166550000000
0!
1$
0'
1+
0/
#166560000000
1!
1'
1/
#166570000000
0!
0'
0/
#166580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#166590000000
0!
0'
0/
#166600000000
1!
1'
1/
#166610000000
0!
0'
0/
#166620000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#166630000000
0!
0'
0/
#166640000000
1!
1'
1/
#166650000000
0!
0'
0/
#166660000000
1!
1'
1/
#166670000000
0!
0'
0/
#166680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#166690000000
0!
0'
0/
#166700000000
1!
1'
1/
#166710000000
0!
0'
0/
#166720000000
1!
1'
1/
#166730000000
0!
0'
0/
#166740000000
1!
1'
1/
#166750000000
0!
0'
0/
#166760000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#166770000000
0!
0'
0/
#166780000000
1!
1'
1/
#166790000000
0!
0'
0/
#166800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#166810000000
0!
0'
0/
#166820000000
1!
1'
1/
#166830000000
0!
0'
0/
#166840000000
#166850000000
1!
1'
1/
#166860000000
0!
0'
0/
#166870000000
1!
1'
1/
#166880000000
0!
1"
0'
1(
0/
10
#166890000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#166900000000
0!
0'
0/
#166910000000
1!
1'
1/
#166920000000
0!
0'
0/
#166930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#166940000000
0!
0'
0/
#166950000000
1!
1'
1/
#166960000000
0!
1"
0'
1(
0/
10
#166970000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#166980000000
0!
1$
0'
1+
0/
#166990000000
1!
1'
1/
#167000000000
0!
0'
0/
#167010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#167020000000
0!
0'
0/
#167030000000
1!
1'
1/
#167040000000
0!
0'
0/
#167050000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#167060000000
0!
0'
0/
#167070000000
1!
1'
1/
#167080000000
0!
0'
0/
#167090000000
1!
1'
1/
#167100000000
0!
0'
0/
#167110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#167120000000
0!
0'
0/
#167130000000
1!
1'
1/
#167140000000
0!
0'
0/
#167150000000
1!
1'
1/
#167160000000
0!
0'
0/
#167170000000
1!
1'
1/
#167180000000
0!
0'
0/
#167190000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#167200000000
0!
0'
0/
#167210000000
1!
1'
1/
#167220000000
0!
0'
0/
#167230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#167240000000
0!
0'
0/
#167250000000
1!
1'
1/
#167260000000
0!
0'
0/
#167270000000
#167280000000
1!
1'
1/
#167290000000
0!
0'
0/
#167300000000
1!
1'
1/
#167310000000
0!
1"
0'
1(
0/
10
#167320000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#167330000000
0!
0'
0/
#167340000000
1!
1'
1/
#167350000000
0!
0'
0/
#167360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#167370000000
0!
0'
0/
#167380000000
1!
1'
1/
#167390000000
0!
1"
0'
1(
0/
10
#167400000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#167410000000
0!
1$
0'
1+
0/
#167420000000
1!
1'
1/
#167430000000
0!
0'
0/
#167440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#167450000000
0!
0'
0/
#167460000000
1!
1'
1/
#167470000000
0!
0'
0/
#167480000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#167490000000
0!
0'
0/
#167500000000
1!
1'
1/
#167510000000
0!
0'
0/
#167520000000
1!
1'
1/
#167530000000
0!
0'
0/
#167540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#167550000000
0!
0'
0/
#167560000000
1!
1'
1/
#167570000000
0!
0'
0/
#167580000000
1!
1'
1/
#167590000000
0!
0'
0/
#167600000000
1!
1'
1/
#167610000000
0!
0'
0/
#167620000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#167630000000
0!
0'
0/
#167640000000
1!
1'
1/
#167650000000
0!
0'
0/
#167660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#167670000000
0!
0'
0/
#167680000000
1!
1'
1/
#167690000000
0!
0'
0/
#167700000000
#167710000000
1!
1'
1/
#167720000000
0!
0'
0/
#167730000000
1!
1'
1/
#167740000000
0!
1"
0'
1(
0/
10
#167750000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#167760000000
0!
0'
0/
#167770000000
1!
1'
1/
#167780000000
0!
0'
0/
#167790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#167800000000
0!
0'
0/
#167810000000
1!
1'
1/
#167820000000
0!
1"
0'
1(
0/
10
#167830000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#167840000000
0!
1$
0'
1+
0/
#167850000000
1!
1'
1/
#167860000000
0!
0'
0/
#167870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#167880000000
0!
0'
0/
#167890000000
1!
1'
1/
#167900000000
0!
0'
0/
#167910000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#167920000000
0!
0'
0/
#167930000000
1!
1'
1/
#167940000000
0!
0'
0/
#167950000000
1!
1'
1/
#167960000000
0!
0'
0/
#167970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#167980000000
0!
0'
0/
#167990000000
1!
1'
1/
#168000000000
0!
0'
0/
#168010000000
1!
1'
1/
#168020000000
0!
0'
0/
#168030000000
1!
1'
1/
#168040000000
0!
0'
0/
#168050000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#168060000000
0!
0'
0/
#168070000000
1!
1'
1/
#168080000000
0!
0'
0/
#168090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#168100000000
0!
0'
0/
#168110000000
1!
1'
1/
#168120000000
0!
0'
0/
#168130000000
#168140000000
1!
1'
1/
#168150000000
0!
0'
0/
#168160000000
1!
1'
1/
#168170000000
0!
1"
0'
1(
0/
10
#168180000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#168190000000
0!
0'
0/
#168200000000
1!
1'
1/
#168210000000
0!
0'
0/
#168220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#168230000000
0!
0'
0/
#168240000000
1!
1'
1/
#168250000000
0!
1"
0'
1(
0/
10
#168260000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#168270000000
0!
1$
0'
1+
0/
#168280000000
1!
1'
1/
#168290000000
0!
0'
0/
#168300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#168310000000
0!
0'
0/
#168320000000
1!
1'
1/
#168330000000
0!
0'
0/
#168340000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#168350000000
0!
0'
0/
#168360000000
1!
1'
1/
#168370000000
0!
0'
0/
#168380000000
1!
1'
1/
#168390000000
0!
0'
0/
#168400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#168410000000
0!
0'
0/
#168420000000
1!
1'
1/
#168430000000
0!
0'
0/
#168440000000
1!
1'
1/
#168450000000
0!
0'
0/
#168460000000
1!
1'
1/
#168470000000
0!
0'
0/
#168480000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#168490000000
0!
0'
0/
#168500000000
1!
1'
1/
#168510000000
0!
0'
0/
#168520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#168530000000
0!
0'
0/
#168540000000
1!
1'
1/
#168550000000
0!
0'
0/
#168560000000
#168570000000
1!
1'
1/
#168580000000
0!
0'
0/
#168590000000
1!
1'
1/
#168600000000
0!
1"
0'
1(
0/
10
#168610000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#168620000000
0!
0'
0/
#168630000000
1!
1'
1/
#168640000000
0!
0'
0/
#168650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#168660000000
0!
0'
0/
#168670000000
1!
1'
1/
#168680000000
0!
1"
0'
1(
0/
10
#168690000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#168700000000
0!
1$
0'
1+
0/
#168710000000
1!
1'
1/
#168720000000
0!
0'
0/
#168730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#168740000000
0!
0'
0/
#168750000000
1!
1'
1/
#168760000000
0!
0'
0/
#168770000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#168780000000
0!
0'
0/
#168790000000
1!
1'
1/
#168800000000
0!
0'
0/
#168810000000
1!
1'
1/
#168820000000
0!
0'
0/
#168830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#168840000000
0!
0'
0/
#168850000000
1!
1'
1/
#168860000000
0!
0'
0/
#168870000000
1!
1'
1/
#168880000000
0!
0'
0/
#168890000000
1!
1'
1/
#168900000000
0!
0'
0/
#168910000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#168920000000
0!
0'
0/
#168930000000
1!
1'
1/
#168940000000
0!
0'
0/
#168950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#168960000000
0!
0'
0/
#168970000000
1!
1'
1/
#168980000000
0!
0'
0/
#168990000000
#169000000000
1!
1'
1/
#169010000000
0!
0'
0/
#169020000000
1!
1'
1/
#169030000000
0!
1"
0'
1(
0/
10
#169040000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#169050000000
0!
0'
0/
#169060000000
1!
1'
1/
#169070000000
0!
0'
0/
#169080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#169090000000
0!
0'
0/
#169100000000
1!
1'
1/
#169110000000
0!
1"
0'
1(
0/
10
#169120000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#169130000000
0!
1$
0'
1+
0/
#169140000000
1!
1'
1/
#169150000000
0!
0'
0/
#169160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#169170000000
0!
0'
0/
#169180000000
1!
1'
1/
#169190000000
0!
0'
0/
#169200000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#169210000000
0!
0'
0/
#169220000000
1!
1'
1/
#169230000000
0!
0'
0/
#169240000000
1!
1'
1/
#169250000000
0!
0'
0/
#169260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#169270000000
0!
0'
0/
#169280000000
1!
1'
1/
#169290000000
0!
0'
0/
#169300000000
1!
1'
1/
#169310000000
0!
0'
0/
#169320000000
1!
1'
1/
#169330000000
0!
0'
0/
#169340000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#169350000000
0!
0'
0/
#169360000000
1!
1'
1/
#169370000000
0!
0'
0/
#169380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#169390000000
0!
0'
0/
#169400000000
1!
1'
1/
#169410000000
0!
0'
0/
#169420000000
#169430000000
1!
1'
1/
#169440000000
0!
0'
0/
#169450000000
1!
1'
1/
#169460000000
0!
1"
0'
1(
0/
10
#169470000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#169480000000
0!
0'
0/
#169490000000
1!
1'
1/
#169500000000
0!
0'
0/
#169510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#169520000000
0!
0'
0/
#169530000000
1!
1'
1/
#169540000000
0!
1"
0'
1(
0/
10
#169550000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#169560000000
0!
1$
0'
1+
0/
#169570000000
1!
1'
1/
#169580000000
0!
0'
0/
#169590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#169600000000
0!
0'
0/
#169610000000
1!
1'
1/
#169620000000
0!
0'
0/
#169630000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#169640000000
0!
0'
0/
#169650000000
1!
1'
1/
#169660000000
0!
0'
0/
#169670000000
1!
1'
1/
#169680000000
0!
0'
0/
#169690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#169700000000
0!
0'
0/
#169710000000
1!
1'
1/
#169720000000
0!
0'
0/
#169730000000
1!
1'
1/
#169740000000
0!
0'
0/
#169750000000
1!
1'
1/
#169760000000
0!
0'
0/
#169770000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#169780000000
0!
0'
0/
#169790000000
1!
1'
1/
#169800000000
0!
0'
0/
#169810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#169820000000
0!
0'
0/
#169830000000
1!
1'
1/
#169840000000
0!
0'
0/
#169850000000
#169860000000
1!
1'
1/
#169870000000
0!
0'
0/
#169880000000
1!
1'
1/
#169890000000
0!
1"
0'
1(
0/
10
#169900000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#169910000000
0!
0'
0/
#169920000000
1!
1'
1/
#169930000000
0!
0'
0/
#169940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#169950000000
0!
0'
0/
#169960000000
1!
1'
1/
#169970000000
0!
1"
0'
1(
0/
10
#169980000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#169990000000
0!
1$
0'
1+
0/
#170000000000
1!
1'
1/
#170010000000
0!
0'
0/
#170020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#170030000000
0!
0'
0/
#170040000000
1!
1'
1/
#170050000000
0!
0'
0/
#170060000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#170070000000
0!
0'
0/
#170080000000
1!
1'
1/
#170090000000
0!
0'
0/
#170100000000
1!
1'
1/
#170110000000
0!
0'
0/
#170120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#170130000000
0!
0'
0/
#170140000000
1!
1'
1/
#170150000000
0!
0'
0/
#170160000000
1!
1'
1/
#170170000000
0!
0'
0/
#170180000000
1!
1'
1/
#170190000000
0!
0'
0/
#170200000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#170210000000
0!
0'
0/
#170220000000
1!
1'
1/
#170230000000
0!
0'
0/
#170240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#170250000000
0!
0'
0/
#170260000000
1!
1'
1/
#170270000000
0!
0'
0/
#170280000000
#170290000000
1!
1'
1/
#170300000000
0!
0'
0/
#170310000000
1!
1'
1/
#170320000000
0!
1"
0'
1(
0/
10
#170330000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#170340000000
0!
0'
0/
#170350000000
1!
1'
1/
#170360000000
0!
0'
0/
#170370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#170380000000
0!
0'
0/
#170390000000
1!
1'
1/
#170400000000
0!
1"
0'
1(
0/
10
#170410000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#170420000000
0!
1$
0'
1+
0/
#170430000000
1!
1'
1/
#170440000000
0!
0'
0/
#170450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#170460000000
0!
0'
0/
#170470000000
1!
1'
1/
#170480000000
0!
0'
0/
#170490000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#170500000000
0!
0'
0/
#170510000000
1!
1'
1/
#170520000000
0!
0'
0/
#170530000000
1!
1'
1/
#170540000000
0!
0'
0/
#170550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#170560000000
0!
0'
0/
#170570000000
1!
1'
1/
#170580000000
0!
0'
0/
#170590000000
1!
1'
1/
#170600000000
0!
0'
0/
#170610000000
1!
1'
1/
#170620000000
0!
0'
0/
#170630000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#170640000000
0!
0'
0/
#170650000000
1!
1'
1/
#170660000000
0!
0'
0/
#170670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#170680000000
0!
0'
0/
#170690000000
1!
1'
1/
#170700000000
0!
0'
0/
#170710000000
#170720000000
1!
1'
1/
#170730000000
0!
0'
0/
#170740000000
1!
1'
1/
#170750000000
0!
1"
0'
1(
0/
10
#170760000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#170770000000
0!
0'
0/
#170780000000
1!
1'
1/
#170790000000
0!
0'
0/
#170800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#170810000000
0!
0'
0/
#170820000000
1!
1'
1/
#170830000000
0!
1"
0'
1(
0/
10
#170840000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#170850000000
0!
1$
0'
1+
0/
#170860000000
1!
1'
1/
#170870000000
0!
0'
0/
#170880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#170890000000
0!
0'
0/
#170900000000
1!
1'
1/
#170910000000
0!
0'
0/
#170920000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#170930000000
0!
0'
0/
#170940000000
1!
1'
1/
#170950000000
0!
0'
0/
#170960000000
1!
1'
1/
#170970000000
0!
0'
0/
#170980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#170990000000
0!
0'
0/
#171000000000
1!
1'
1/
#171010000000
0!
0'
0/
#171020000000
1!
1'
1/
#171030000000
0!
0'
0/
#171040000000
1!
1'
1/
#171050000000
0!
0'
0/
#171060000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#171070000000
0!
0'
0/
#171080000000
1!
1'
1/
#171090000000
0!
0'
0/
#171100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#171110000000
0!
0'
0/
#171120000000
1!
1'
1/
#171130000000
0!
0'
0/
#171140000000
#171150000000
1!
1'
1/
#171160000000
0!
0'
0/
#171170000000
1!
1'
1/
#171180000000
0!
1"
0'
1(
0/
10
#171190000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#171200000000
0!
0'
0/
#171210000000
1!
1'
1/
#171220000000
0!
0'
0/
#171230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#171240000000
0!
0'
0/
#171250000000
1!
1'
1/
#171260000000
0!
1"
0'
1(
0/
10
#171270000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#171280000000
0!
1$
0'
1+
0/
#171290000000
1!
1'
1/
#171300000000
0!
0'
0/
#171310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#171320000000
0!
0'
0/
#171330000000
1!
1'
1/
#171340000000
0!
0'
0/
#171350000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#171360000000
0!
0'
0/
#171370000000
1!
1'
1/
#171380000000
0!
0'
0/
#171390000000
1!
1'
1/
#171400000000
0!
0'
0/
#171410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#171420000000
0!
0'
0/
#171430000000
1!
1'
1/
#171440000000
0!
0'
0/
#171450000000
1!
1'
1/
#171460000000
0!
0'
0/
#171470000000
1!
1'
1/
#171480000000
0!
0'
0/
#171490000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#171500000000
0!
0'
0/
#171510000000
1!
1'
1/
#171520000000
0!
0'
0/
#171530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#171540000000
0!
0'
0/
#171550000000
1!
1'
1/
#171560000000
0!
0'
0/
#171570000000
#171580000000
1!
1'
1/
#171590000000
0!
0'
0/
#171600000000
1!
1'
1/
#171610000000
0!
1"
0'
1(
0/
10
#171620000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#171630000000
0!
0'
0/
#171640000000
1!
1'
1/
#171650000000
0!
0'
0/
#171660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#171670000000
0!
0'
0/
#171680000000
1!
1'
1/
#171690000000
0!
1"
0'
1(
0/
10
#171700000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#171710000000
0!
1$
0'
1+
0/
#171720000000
1!
1'
1/
#171730000000
0!
0'
0/
#171740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#171750000000
0!
0'
0/
#171760000000
1!
1'
1/
#171770000000
0!
0'
0/
#171780000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#171790000000
0!
0'
0/
#171800000000
1!
1'
1/
#171810000000
0!
0'
0/
#171820000000
1!
1'
1/
#171830000000
0!
0'
0/
#171840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#171850000000
0!
0'
0/
#171860000000
1!
1'
1/
#171870000000
0!
0'
0/
#171880000000
1!
1'
1/
#171890000000
0!
0'
0/
#171900000000
1!
1'
1/
#171910000000
0!
0'
0/
#171920000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#171930000000
0!
0'
0/
#171940000000
1!
1'
1/
#171950000000
0!
0'
0/
#171960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#171970000000
0!
0'
0/
#171980000000
1!
1'
1/
#171990000000
0!
0'
0/
#172000000000
#172010000000
1!
1'
1/
#172020000000
0!
0'
0/
#172030000000
1!
1'
1/
#172040000000
0!
1"
0'
1(
0/
10
#172050000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#172060000000
0!
0'
0/
#172070000000
1!
1'
1/
#172080000000
0!
0'
0/
#172090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#172100000000
0!
0'
0/
#172110000000
1!
1'
1/
#172120000000
0!
1"
0'
1(
0/
10
#172130000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#172140000000
0!
1$
0'
1+
0/
#172150000000
1!
1'
1/
#172160000000
0!
0'
0/
#172170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#172180000000
0!
0'
0/
#172190000000
1!
1'
1/
#172200000000
0!
0'
0/
#172210000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#172220000000
0!
0'
0/
#172230000000
1!
1'
1/
#172240000000
0!
0'
0/
#172250000000
1!
1'
1/
#172260000000
0!
0'
0/
#172270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#172280000000
0!
0'
0/
#172290000000
1!
1'
1/
#172300000000
0!
0'
0/
#172310000000
1!
1'
1/
#172320000000
0!
0'
0/
#172330000000
1!
1'
1/
#172340000000
0!
0'
0/
#172350000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#172360000000
0!
0'
0/
#172370000000
1!
1'
1/
#172380000000
0!
0'
0/
#172390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#172400000000
0!
0'
0/
#172410000000
1!
1'
1/
#172420000000
0!
0'
0/
#172430000000
#172440000000
1!
1'
1/
#172450000000
0!
0'
0/
#172460000000
1!
1'
1/
#172470000000
0!
1"
0'
1(
0/
10
#172480000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#172490000000
0!
0'
0/
#172500000000
1!
1'
1/
#172510000000
0!
0'
0/
#172520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#172530000000
0!
0'
0/
#172540000000
1!
1'
1/
#172550000000
0!
1"
0'
1(
0/
10
#172560000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#172570000000
0!
1$
0'
1+
0/
#172580000000
1!
1'
1/
#172590000000
0!
0'
0/
#172600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#172610000000
0!
0'
0/
#172620000000
1!
1'
1/
#172630000000
0!
0'
0/
#172640000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#172650000000
0!
0'
0/
#172660000000
1!
1'
1/
#172670000000
0!
0'
0/
#172680000000
1!
1'
1/
#172690000000
0!
0'
0/
#172700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#172710000000
0!
0'
0/
#172720000000
1!
1'
1/
#172730000000
0!
0'
0/
#172740000000
1!
1'
1/
#172750000000
0!
0'
0/
#172760000000
1!
1'
1/
#172770000000
0!
0'
0/
#172780000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#172790000000
0!
0'
0/
#172800000000
1!
1'
1/
#172810000000
0!
0'
0/
#172820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#172830000000
0!
0'
0/
#172840000000
1!
1'
1/
#172850000000
0!
0'
0/
#172860000000
#172870000000
1!
1'
1/
#172880000000
0!
0'
0/
#172890000000
1!
1'
1/
#172900000000
0!
1"
0'
1(
0/
10
#172910000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#172920000000
0!
0'
0/
#172930000000
1!
1'
1/
#172940000000
0!
0'
0/
#172950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#172960000000
0!
0'
0/
#172970000000
1!
1'
1/
#172980000000
0!
1"
0'
1(
0/
10
#172990000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#173000000000
0!
1$
0'
1+
0/
#173010000000
1!
1'
1/
#173020000000
0!
0'
0/
#173030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#173040000000
0!
0'
0/
#173050000000
1!
1'
1/
#173060000000
0!
0'
0/
#173070000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#173080000000
0!
0'
0/
#173090000000
1!
1'
1/
#173100000000
0!
0'
0/
#173110000000
1!
1'
1/
#173120000000
0!
0'
0/
#173130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#173140000000
0!
0'
0/
#173150000000
1!
1'
1/
#173160000000
0!
0'
0/
#173170000000
1!
1'
1/
#173180000000
0!
0'
0/
#173190000000
1!
1'
1/
#173200000000
0!
0'
0/
#173210000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#173220000000
0!
0'
0/
#173230000000
1!
1'
1/
#173240000000
0!
0'
0/
#173250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#173260000000
0!
0'
0/
#173270000000
1!
1'
1/
#173280000000
0!
0'
0/
#173290000000
#173300000000
1!
1'
1/
#173310000000
0!
0'
0/
#173320000000
1!
1'
1/
#173330000000
0!
1"
0'
1(
0/
10
#173340000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#173350000000
0!
0'
0/
#173360000000
1!
1'
1/
#173370000000
0!
0'
0/
#173380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#173390000000
0!
0'
0/
#173400000000
1!
1'
1/
#173410000000
0!
1"
0'
1(
0/
10
#173420000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#173430000000
0!
1$
0'
1+
0/
#173440000000
1!
1'
1/
#173450000000
0!
0'
0/
#173460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#173470000000
0!
0'
0/
#173480000000
1!
1'
1/
#173490000000
0!
0'
0/
#173500000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#173510000000
0!
0'
0/
#173520000000
1!
1'
1/
#173530000000
0!
0'
0/
#173540000000
1!
1'
1/
#173550000000
0!
0'
0/
#173560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#173570000000
0!
0'
0/
#173580000000
1!
1'
1/
#173590000000
0!
0'
0/
#173600000000
1!
1'
1/
#173610000000
0!
0'
0/
#173620000000
1!
1'
1/
#173630000000
0!
0'
0/
#173640000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#173650000000
0!
0'
0/
#173660000000
1!
1'
1/
#173670000000
0!
0'
0/
#173680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#173690000000
0!
0'
0/
#173700000000
1!
1'
1/
#173710000000
0!
0'
0/
#173720000000
#173730000000
1!
1'
1/
#173740000000
0!
0'
0/
#173750000000
1!
1'
1/
#173760000000
0!
1"
0'
1(
0/
10
#173770000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#173780000000
0!
0'
0/
#173790000000
1!
1'
1/
#173800000000
0!
0'
0/
#173810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#173820000000
0!
0'
0/
#173830000000
1!
1'
1/
#173840000000
0!
1"
0'
1(
0/
10
#173850000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#173860000000
0!
1$
0'
1+
0/
#173870000000
1!
1'
1/
#173880000000
0!
0'
0/
#173890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#173900000000
0!
0'
0/
#173910000000
1!
1'
1/
#173920000000
0!
0'
0/
#173930000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#173940000000
0!
0'
0/
#173950000000
1!
1'
1/
#173960000000
0!
0'
0/
#173970000000
1!
1'
1/
#173980000000
0!
0'
0/
#173990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#174000000000
0!
0'
0/
#174010000000
1!
1'
1/
#174020000000
0!
0'
0/
#174030000000
1!
1'
1/
#174040000000
0!
0'
0/
#174050000000
1!
1'
1/
#174060000000
0!
0'
0/
#174070000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#174080000000
0!
0'
0/
#174090000000
1!
1'
1/
#174100000000
0!
0'
0/
#174110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#174120000000
0!
0'
0/
#174130000000
1!
1'
1/
#174140000000
0!
0'
0/
#174150000000
#174160000000
1!
1'
1/
#174170000000
0!
0'
0/
#174180000000
1!
1'
1/
#174190000000
0!
1"
0'
1(
0/
10
#174200000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#174210000000
0!
0'
0/
#174220000000
1!
1'
1/
#174230000000
0!
0'
0/
#174240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#174250000000
0!
0'
0/
#174260000000
1!
1'
1/
#174270000000
0!
1"
0'
1(
0/
10
#174280000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#174290000000
0!
1$
0'
1+
0/
#174300000000
1!
1'
1/
#174310000000
0!
0'
0/
#174320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#174330000000
0!
0'
0/
#174340000000
1!
1'
1/
#174350000000
0!
0'
0/
#174360000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#174370000000
0!
0'
0/
#174380000000
1!
1'
1/
#174390000000
0!
0'
0/
#174400000000
1!
1'
1/
#174410000000
0!
0'
0/
#174420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#174430000000
0!
0'
0/
#174440000000
1!
1'
1/
#174450000000
0!
0'
0/
#174460000000
1!
1'
1/
#174470000000
0!
0'
0/
#174480000000
1!
1'
1/
#174490000000
0!
0'
0/
#174500000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#174510000000
0!
0'
0/
#174520000000
1!
1'
1/
#174530000000
0!
0'
0/
#174540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#174550000000
0!
0'
0/
#174560000000
1!
1'
1/
#174570000000
0!
0'
0/
#174580000000
#174590000000
1!
1'
1/
#174600000000
0!
0'
0/
#174610000000
1!
1'
1/
#174620000000
0!
1"
0'
1(
0/
10
#174630000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#174640000000
0!
0'
0/
#174650000000
1!
1'
1/
#174660000000
0!
0'
0/
#174670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#174680000000
0!
0'
0/
#174690000000
1!
1'
1/
#174700000000
0!
1"
0'
1(
0/
10
#174710000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#174720000000
0!
1$
0'
1+
0/
#174730000000
1!
1'
1/
#174740000000
0!
0'
0/
#174750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#174760000000
0!
0'
0/
#174770000000
1!
1'
1/
#174780000000
0!
0'
0/
#174790000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#174800000000
0!
0'
0/
#174810000000
1!
1'
1/
#174820000000
0!
0'
0/
#174830000000
1!
1'
1/
#174840000000
0!
0'
0/
#174850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#174860000000
0!
0'
0/
#174870000000
1!
1'
1/
#174880000000
0!
0'
0/
#174890000000
1!
1'
1/
#174900000000
0!
0'
0/
#174910000000
1!
1'
1/
#174920000000
0!
0'
0/
#174930000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#174940000000
0!
0'
0/
#174950000000
1!
1'
1/
#174960000000
0!
0'
0/
#174970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#174980000000
0!
0'
0/
#174990000000
1!
1'
1/
#175000000000
0!
0'
0/
#175010000000
#175020000000
1!
1'
1/
#175030000000
0!
0'
0/
#175040000000
1!
1'
1/
#175050000000
0!
1"
0'
1(
0/
10
#175060000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#175070000000
0!
0'
0/
#175080000000
1!
1'
1/
#175090000000
0!
0'
0/
#175100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#175110000000
0!
0'
0/
#175120000000
1!
1'
1/
#175130000000
0!
1"
0'
1(
0/
10
#175140000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#175150000000
0!
1$
0'
1+
0/
#175160000000
1!
1'
1/
#175170000000
0!
0'
0/
#175180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#175190000000
0!
0'
0/
#175200000000
1!
1'
1/
#175210000000
0!
0'
0/
#175220000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#175230000000
0!
0'
0/
#175240000000
1!
1'
1/
#175250000000
0!
0'
0/
#175260000000
1!
1'
1/
#175270000000
0!
0'
0/
#175280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#175290000000
0!
0'
0/
#175300000000
1!
1'
1/
#175310000000
0!
0'
0/
#175320000000
1!
1'
1/
#175330000000
0!
0'
0/
#175340000000
1!
1'
1/
#175350000000
0!
0'
0/
#175360000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#175370000000
0!
0'
0/
#175380000000
1!
1'
1/
#175390000000
0!
0'
0/
#175400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#175410000000
0!
0'
0/
#175420000000
1!
1'
1/
#175430000000
0!
0'
0/
#175440000000
#175450000000
1!
1'
1/
#175460000000
0!
0'
0/
#175470000000
1!
1'
1/
#175480000000
0!
1"
0'
1(
0/
10
#175490000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#175500000000
0!
0'
0/
#175510000000
1!
1'
1/
#175520000000
0!
0'
0/
#175530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#175540000000
0!
0'
0/
#175550000000
1!
1'
1/
#175560000000
0!
1"
0'
1(
0/
10
#175570000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#175580000000
0!
1$
0'
1+
0/
#175590000000
1!
1'
1/
#175600000000
0!
0'
0/
#175610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#175620000000
0!
0'
0/
#175630000000
1!
1'
1/
#175640000000
0!
0'
0/
#175650000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#175660000000
0!
0'
0/
#175670000000
1!
1'
1/
#175680000000
0!
0'
0/
#175690000000
1!
1'
1/
#175700000000
0!
0'
0/
#175710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#175720000000
0!
0'
0/
#175730000000
1!
1'
1/
#175740000000
0!
0'
0/
#175750000000
1!
1'
1/
#175760000000
0!
0'
0/
#175770000000
1!
1'
1/
#175780000000
0!
0'
0/
#175790000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#175800000000
0!
0'
0/
#175810000000
1!
1'
1/
#175820000000
0!
0'
0/
#175830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#175840000000
0!
0'
0/
#175850000000
1!
1'
1/
#175860000000
0!
0'
0/
#175870000000
#175880000000
1!
1'
1/
#175890000000
0!
0'
0/
#175900000000
1!
1'
1/
#175910000000
0!
1"
0'
1(
0/
10
#175920000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#175930000000
0!
0'
0/
#175940000000
1!
1'
1/
#175950000000
0!
0'
0/
#175960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#175970000000
0!
0'
0/
#175980000000
1!
1'
1/
#175990000000
0!
1"
0'
1(
0/
10
#176000000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#176010000000
0!
1$
0'
1+
0/
#176020000000
1!
1'
1/
#176030000000
0!
0'
0/
#176040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#176050000000
0!
0'
0/
#176060000000
1!
1'
1/
#176070000000
0!
0'
0/
#176080000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#176090000000
0!
0'
0/
#176100000000
1!
1'
1/
#176110000000
0!
0'
0/
#176120000000
1!
1'
1/
#176130000000
0!
0'
0/
#176140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#176150000000
0!
0'
0/
#176160000000
1!
1'
1/
#176170000000
0!
0'
0/
#176180000000
1!
1'
1/
#176190000000
0!
0'
0/
#176200000000
1!
1'
1/
#176210000000
0!
0'
0/
#176220000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#176230000000
0!
0'
0/
#176240000000
1!
1'
1/
#176250000000
0!
0'
0/
#176260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#176270000000
0!
0'
0/
#176280000000
1!
1'
1/
#176290000000
0!
0'
0/
#176300000000
#176310000000
1!
1'
1/
#176320000000
0!
0'
0/
#176330000000
1!
1'
1/
#176340000000
0!
1"
0'
1(
0/
10
#176350000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#176360000000
0!
0'
0/
#176370000000
1!
1'
1/
#176380000000
0!
0'
0/
#176390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#176400000000
0!
0'
0/
#176410000000
1!
1'
1/
#176420000000
0!
1"
0'
1(
0/
10
#176430000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#176440000000
0!
1$
0'
1+
0/
#176450000000
1!
1'
1/
#176460000000
0!
0'
0/
#176470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#176480000000
0!
0'
0/
#176490000000
1!
1'
1/
#176500000000
0!
0'
0/
#176510000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#176520000000
0!
0'
0/
#176530000000
1!
1'
1/
#176540000000
0!
0'
0/
#176550000000
1!
1'
1/
#176560000000
0!
0'
0/
#176570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#176580000000
0!
0'
0/
#176590000000
1!
1'
1/
#176600000000
0!
0'
0/
#176610000000
1!
1'
1/
#176620000000
0!
0'
0/
#176630000000
1!
1'
1/
#176640000000
0!
0'
0/
#176650000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#176660000000
0!
0'
0/
#176670000000
1!
1'
1/
#176680000000
0!
0'
0/
#176690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#176700000000
0!
0'
0/
#176710000000
1!
1'
1/
#176720000000
0!
0'
0/
#176730000000
#176740000000
1!
1'
1/
#176750000000
0!
0'
0/
#176760000000
1!
1'
1/
#176770000000
0!
1"
0'
1(
0/
10
#176780000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#176790000000
0!
0'
0/
#176800000000
1!
1'
1/
#176810000000
0!
0'
0/
#176820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#176830000000
0!
0'
0/
#176840000000
1!
1'
1/
#176850000000
0!
1"
0'
1(
0/
10
#176860000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#176870000000
0!
1$
0'
1+
0/
#176880000000
1!
1'
1/
#176890000000
0!
0'
0/
#176900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#176910000000
0!
0'
0/
#176920000000
1!
1'
1/
#176930000000
0!
0'
0/
#176940000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#176950000000
0!
0'
0/
#176960000000
1!
1'
1/
#176970000000
0!
0'
0/
#176980000000
1!
1'
1/
#176990000000
0!
0'
0/
#177000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#177010000000
0!
0'
0/
#177020000000
1!
1'
1/
#177030000000
0!
0'
0/
#177040000000
1!
1'
1/
#177050000000
0!
0'
0/
#177060000000
1!
1'
1/
#177070000000
0!
0'
0/
#177080000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#177090000000
0!
0'
0/
#177100000000
1!
1'
1/
#177110000000
0!
0'
0/
#177120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#177130000000
0!
0'
0/
#177140000000
1!
1'
1/
#177150000000
0!
0'
0/
#177160000000
#177170000000
1!
1'
1/
#177180000000
0!
0'
0/
#177190000000
1!
1'
1/
#177200000000
0!
1"
0'
1(
0/
10
#177210000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#177220000000
0!
0'
0/
#177230000000
1!
1'
1/
#177240000000
0!
0'
0/
#177250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#177260000000
0!
0'
0/
#177270000000
1!
1'
1/
#177280000000
0!
1"
0'
1(
0/
10
#177290000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#177300000000
0!
1$
0'
1+
0/
#177310000000
1!
1'
1/
#177320000000
0!
0'
0/
#177330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#177340000000
0!
0'
0/
#177350000000
1!
1'
1/
#177360000000
0!
0'
0/
#177370000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#177380000000
0!
0'
0/
#177390000000
1!
1'
1/
#177400000000
0!
0'
0/
#177410000000
1!
1'
1/
#177420000000
0!
0'
0/
#177430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#177440000000
0!
0'
0/
#177450000000
1!
1'
1/
#177460000000
0!
0'
0/
#177470000000
1!
1'
1/
#177480000000
0!
0'
0/
#177490000000
1!
1'
1/
#177500000000
0!
0'
0/
#177510000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#177520000000
0!
0'
0/
#177530000000
1!
1'
1/
#177540000000
0!
0'
0/
#177550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#177560000000
0!
0'
0/
#177570000000
1!
1'
1/
#177580000000
0!
0'
0/
#177590000000
#177600000000
1!
1'
1/
#177610000000
0!
0'
0/
#177620000000
1!
1'
1/
#177630000000
0!
1"
0'
1(
0/
10
#177640000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#177650000000
0!
0'
0/
#177660000000
1!
1'
1/
#177670000000
0!
0'
0/
#177680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#177690000000
0!
0'
0/
#177700000000
1!
1'
1/
#177710000000
0!
1"
0'
1(
0/
10
#177720000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#177730000000
0!
1$
0'
1+
0/
#177740000000
1!
1'
1/
#177750000000
0!
0'
0/
#177760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#177770000000
0!
0'
0/
#177780000000
1!
1'
1/
#177790000000
0!
0'
0/
#177800000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#177810000000
0!
0'
0/
#177820000000
1!
1'
1/
#177830000000
0!
0'
0/
#177840000000
1!
1'
1/
#177850000000
0!
0'
0/
#177860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#177870000000
0!
0'
0/
#177880000000
1!
1'
1/
#177890000000
0!
0'
0/
#177900000000
1!
1'
1/
#177910000000
0!
0'
0/
#177920000000
1!
1'
1/
#177930000000
0!
0'
0/
#177940000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#177950000000
0!
0'
0/
#177960000000
1!
1'
1/
#177970000000
0!
0'
0/
#177980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#177990000000
0!
0'
0/
#178000000000
1!
1'
1/
#178010000000
0!
0'
0/
#178020000000
#178030000000
1!
1'
1/
#178040000000
0!
0'
0/
#178050000000
1!
1'
1/
#178060000000
0!
1"
0'
1(
0/
10
#178070000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#178080000000
0!
0'
0/
#178090000000
1!
1'
1/
#178100000000
0!
0'
0/
#178110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#178120000000
0!
0'
0/
#178130000000
1!
1'
1/
#178140000000
0!
1"
0'
1(
0/
10
#178150000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#178160000000
0!
1$
0'
1+
0/
#178170000000
1!
1'
1/
#178180000000
0!
0'
0/
#178190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#178200000000
0!
0'
0/
#178210000000
1!
1'
1/
#178220000000
0!
0'
0/
#178230000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#178240000000
0!
0'
0/
#178250000000
1!
1'
1/
#178260000000
0!
0'
0/
#178270000000
1!
1'
1/
#178280000000
0!
0'
0/
#178290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#178300000000
0!
0'
0/
#178310000000
1!
1'
1/
#178320000000
0!
0'
0/
#178330000000
1!
1'
1/
#178340000000
0!
0'
0/
#178350000000
1!
1'
1/
#178360000000
0!
0'
0/
#178370000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#178380000000
0!
0'
0/
#178390000000
1!
1'
1/
#178400000000
0!
0'
0/
#178410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#178420000000
0!
0'
0/
#178430000000
1!
1'
1/
#178440000000
0!
0'
0/
#178450000000
#178460000000
1!
1'
1/
#178470000000
0!
0'
0/
#178480000000
1!
1'
1/
#178490000000
0!
1"
0'
1(
0/
10
#178500000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#178510000000
0!
0'
0/
#178520000000
1!
1'
1/
#178530000000
0!
0'
0/
#178540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#178550000000
0!
0'
0/
#178560000000
1!
1'
1/
#178570000000
0!
1"
0'
1(
0/
10
#178580000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#178590000000
0!
1$
0'
1+
0/
#178600000000
1!
1'
1/
#178610000000
0!
0'
0/
#178620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#178630000000
0!
0'
0/
#178640000000
1!
1'
1/
#178650000000
0!
0'
0/
#178660000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#178670000000
0!
0'
0/
#178680000000
1!
1'
1/
#178690000000
0!
0'
0/
#178700000000
1!
1'
1/
#178710000000
0!
0'
0/
#178720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#178730000000
0!
0'
0/
#178740000000
1!
1'
1/
#178750000000
0!
0'
0/
#178760000000
1!
1'
1/
#178770000000
0!
0'
0/
#178780000000
1!
1'
1/
#178790000000
0!
0'
0/
#178800000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#178810000000
0!
0'
0/
#178820000000
1!
1'
1/
#178830000000
0!
0'
0/
#178840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#178850000000
0!
0'
0/
#178860000000
1!
1'
1/
#178870000000
0!
0'
0/
#178880000000
#178890000000
1!
1'
1/
#178900000000
0!
0'
0/
#178910000000
1!
1'
1/
#178920000000
0!
1"
0'
1(
0/
10
#178930000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#178940000000
0!
0'
0/
#178950000000
1!
1'
1/
#178960000000
0!
0'
0/
#178970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#178980000000
0!
0'
0/
#178990000000
1!
1'
1/
#179000000000
0!
1"
0'
1(
0/
10
#179010000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#179020000000
0!
1$
0'
1+
0/
#179030000000
1!
1'
1/
#179040000000
0!
0'
0/
#179050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#179060000000
0!
0'
0/
#179070000000
1!
1'
1/
#179080000000
0!
0'
0/
#179090000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#179100000000
0!
0'
0/
#179110000000
1!
1'
1/
#179120000000
0!
0'
0/
#179130000000
1!
1'
1/
#179140000000
0!
0'
0/
#179150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#179160000000
0!
0'
0/
#179170000000
1!
1'
1/
#179180000000
0!
0'
0/
#179190000000
1!
1'
1/
#179200000000
0!
0'
0/
#179210000000
1!
1'
1/
#179220000000
0!
0'
0/
#179230000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#179240000000
0!
0'
0/
#179250000000
1!
1'
1/
#179260000000
0!
0'
0/
#179270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#179280000000
0!
0'
0/
#179290000000
1!
1'
1/
#179300000000
0!
0'
0/
#179310000000
#179320000000
1!
1'
1/
#179330000000
0!
0'
0/
#179340000000
1!
1'
1/
#179350000000
0!
1"
0'
1(
0/
10
#179360000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#179370000000
0!
0'
0/
#179380000000
1!
1'
1/
#179390000000
0!
0'
0/
#179400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#179410000000
0!
0'
0/
#179420000000
1!
1'
1/
#179430000000
0!
1"
0'
1(
0/
10
#179440000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#179450000000
0!
1$
0'
1+
0/
#179460000000
1!
1'
1/
#179470000000
0!
0'
0/
#179480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#179490000000
0!
0'
0/
#179500000000
1!
1'
1/
#179510000000
0!
0'
0/
#179520000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#179530000000
0!
0'
0/
#179540000000
1!
1'
1/
#179550000000
0!
0'
0/
#179560000000
1!
1'
1/
#179570000000
0!
0'
0/
#179580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#179590000000
0!
0'
0/
#179600000000
1!
1'
1/
#179610000000
0!
0'
0/
#179620000000
1!
1'
1/
#179630000000
0!
0'
0/
#179640000000
1!
1'
1/
#179650000000
0!
0'
0/
#179660000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#179670000000
0!
0'
0/
#179680000000
1!
1'
1/
#179690000000
0!
0'
0/
#179700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#179710000000
0!
0'
0/
#179720000000
1!
1'
1/
#179730000000
0!
0'
0/
#179740000000
#179750000000
1!
1'
1/
#179760000000
0!
0'
0/
#179770000000
1!
1'
1/
#179780000000
0!
1"
0'
1(
0/
10
#179790000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#179800000000
0!
0'
0/
#179810000000
1!
1'
1/
#179820000000
0!
0'
0/
#179830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#179840000000
0!
0'
0/
#179850000000
1!
1'
1/
#179860000000
0!
1"
0'
1(
0/
10
#179870000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#179880000000
0!
1$
0'
1+
0/
#179890000000
1!
1'
1/
#179900000000
0!
0'
0/
#179910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#179920000000
0!
0'
0/
#179930000000
1!
1'
1/
#179940000000
0!
0'
0/
#179950000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#179960000000
0!
0'
0/
#179970000000
1!
1'
1/
#179980000000
0!
0'
0/
#179990000000
1!
1'
1/
#180000000000
0!
0'
0/
#180010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#180020000000
0!
0'
0/
#180030000000
1!
1'
1/
#180040000000
0!
0'
0/
#180050000000
1!
1'
1/
#180060000000
0!
0'
0/
#180070000000
1!
1'
1/
#180080000000
0!
0'
0/
#180090000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#180100000000
0!
0'
0/
#180110000000
1!
1'
1/
#180120000000
0!
0'
0/
#180130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#180140000000
0!
0'
0/
#180150000000
1!
1'
1/
#180160000000
0!
0'
0/
#180170000000
#180180000000
1!
1'
1/
#180190000000
0!
0'
0/
#180200000000
1!
1'
1/
#180210000000
0!
1"
0'
1(
0/
10
#180220000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#180230000000
0!
0'
0/
#180240000000
1!
1'
1/
#180250000000
0!
0'
0/
#180260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#180270000000
0!
0'
0/
#180280000000
1!
1'
1/
#180290000000
0!
1"
0'
1(
0/
10
#180300000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#180310000000
0!
1$
0'
1+
0/
#180320000000
1!
1'
1/
#180330000000
0!
0'
0/
#180340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#180350000000
0!
0'
0/
#180360000000
1!
1'
1/
#180370000000
0!
0'
0/
#180380000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#180390000000
0!
0'
0/
#180400000000
1!
1'
1/
#180410000000
0!
0'
0/
#180420000000
1!
1'
1/
#180430000000
0!
0'
0/
#180440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#180450000000
0!
0'
0/
#180460000000
1!
1'
1/
#180470000000
0!
0'
0/
#180480000000
1!
1'
1/
#180490000000
0!
0'
0/
#180500000000
1!
1'
1/
#180510000000
0!
0'
0/
#180520000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#180530000000
0!
0'
0/
#180540000000
1!
1'
1/
#180550000000
0!
0'
0/
#180560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#180570000000
0!
0'
0/
#180580000000
1!
1'
1/
#180590000000
0!
0'
0/
#180600000000
#180610000000
1!
1'
1/
#180620000000
0!
0'
0/
#180630000000
1!
1'
1/
#180640000000
0!
1"
0'
1(
0/
10
#180650000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#180660000000
0!
0'
0/
#180670000000
1!
1'
1/
#180680000000
0!
0'
0/
#180690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#180700000000
0!
0'
0/
#180710000000
1!
1'
1/
#180720000000
0!
1"
0'
1(
0/
10
#180730000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#180740000000
0!
1$
0'
1+
0/
#180750000000
1!
1'
1/
#180760000000
0!
0'
0/
#180770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#180780000000
0!
0'
0/
#180790000000
1!
1'
1/
#180800000000
0!
0'
0/
#180810000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#180820000000
0!
0'
0/
#180830000000
1!
1'
1/
#180840000000
0!
0'
0/
#180850000000
1!
1'
1/
#180860000000
0!
0'
0/
#180870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#180880000000
0!
0'
0/
#180890000000
1!
1'
1/
#180900000000
0!
0'
0/
#180910000000
1!
1'
1/
#180920000000
0!
0'
0/
#180930000000
1!
1'
1/
#180940000000
0!
0'
0/
#180950000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#180960000000
0!
0'
0/
#180970000000
1!
1'
1/
#180980000000
0!
0'
0/
#180990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#181000000000
0!
0'
0/
#181010000000
1!
1'
1/
#181020000000
0!
0'
0/
#181030000000
#181040000000
1!
1'
1/
#181050000000
0!
0'
0/
#181060000000
1!
1'
1/
#181070000000
0!
1"
0'
1(
0/
10
#181080000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#181090000000
0!
0'
0/
#181100000000
1!
1'
1/
#181110000000
0!
0'
0/
#181120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#181130000000
0!
0'
0/
#181140000000
1!
1'
1/
#181150000000
0!
1"
0'
1(
0/
10
#181160000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#181170000000
0!
1$
0'
1+
0/
#181180000000
1!
1'
1/
#181190000000
0!
0'
0/
#181200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#181210000000
0!
0'
0/
#181220000000
1!
1'
1/
#181230000000
0!
0'
0/
#181240000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#181250000000
0!
0'
0/
#181260000000
1!
1'
1/
#181270000000
0!
0'
0/
#181280000000
1!
1'
1/
#181290000000
0!
0'
0/
#181300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#181310000000
0!
0'
0/
#181320000000
1!
1'
1/
#181330000000
0!
0'
0/
#181340000000
1!
1'
1/
#181350000000
0!
0'
0/
#181360000000
1!
1'
1/
#181370000000
0!
0'
0/
#181380000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#181390000000
0!
0'
0/
#181400000000
1!
1'
1/
#181410000000
0!
0'
0/
#181420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#181430000000
0!
0'
0/
#181440000000
1!
1'
1/
#181450000000
0!
0'
0/
#181460000000
#181470000000
1!
1'
1/
#181480000000
0!
0'
0/
#181490000000
1!
1'
1/
#181500000000
0!
1"
0'
1(
0/
10
#181510000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#181520000000
0!
0'
0/
#181530000000
1!
1'
1/
#181540000000
0!
0'
0/
#181550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#181560000000
0!
0'
0/
#181570000000
1!
1'
1/
#181580000000
0!
1"
0'
1(
0/
10
#181590000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#181600000000
0!
1$
0'
1+
0/
#181610000000
1!
1'
1/
#181620000000
0!
0'
0/
#181630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#181640000000
0!
0'
0/
#181650000000
1!
1'
1/
#181660000000
0!
0'
0/
#181670000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#181680000000
0!
0'
0/
#181690000000
1!
1'
1/
#181700000000
0!
0'
0/
#181710000000
1!
1'
1/
#181720000000
0!
0'
0/
#181730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#181740000000
0!
0'
0/
#181750000000
1!
1'
1/
#181760000000
0!
0'
0/
#181770000000
1!
1'
1/
#181780000000
0!
0'
0/
#181790000000
1!
1'
1/
#181800000000
0!
0'
0/
#181810000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#181820000000
0!
0'
0/
#181830000000
1!
1'
1/
#181840000000
0!
0'
0/
#181850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#181860000000
0!
0'
0/
#181870000000
1!
1'
1/
#181880000000
0!
0'
0/
#181890000000
#181900000000
1!
1'
1/
#181910000000
0!
0'
0/
#181920000000
1!
1'
1/
#181930000000
0!
1"
0'
1(
0/
10
#181940000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#181950000000
0!
0'
0/
#181960000000
1!
1'
1/
#181970000000
0!
0'
0/
#181980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#181990000000
0!
0'
0/
#182000000000
1!
1'
1/
#182010000000
0!
1"
0'
1(
0/
10
#182020000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#182030000000
0!
1$
0'
1+
0/
#182040000000
1!
1'
1/
#182050000000
0!
0'
0/
#182060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#182070000000
0!
0'
0/
#182080000000
1!
1'
1/
#182090000000
0!
0'
0/
#182100000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#182110000000
0!
0'
0/
#182120000000
1!
1'
1/
#182130000000
0!
0'
0/
#182140000000
1!
1'
1/
#182150000000
0!
0'
0/
#182160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#182170000000
0!
0'
0/
#182180000000
1!
1'
1/
#182190000000
0!
0'
0/
#182200000000
1!
1'
1/
#182210000000
0!
0'
0/
#182220000000
1!
1'
1/
#182230000000
0!
0'
0/
#182240000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#182250000000
0!
0'
0/
#182260000000
1!
1'
1/
#182270000000
0!
0'
0/
#182280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#182290000000
0!
0'
0/
#182300000000
1!
1'
1/
#182310000000
0!
0'
0/
#182320000000
#182330000000
1!
1'
1/
#182340000000
0!
0'
0/
#182350000000
1!
1'
1/
#182360000000
0!
1"
0'
1(
0/
10
#182370000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#182380000000
0!
0'
0/
#182390000000
1!
1'
1/
#182400000000
0!
0'
0/
#182410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#182420000000
0!
0'
0/
#182430000000
1!
1'
1/
#182440000000
0!
1"
0'
1(
0/
10
#182450000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#182460000000
0!
1$
0'
1+
0/
#182470000000
1!
1'
1/
#182480000000
0!
0'
0/
#182490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#182500000000
0!
0'
0/
#182510000000
1!
1'
1/
#182520000000
0!
0'
0/
#182530000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#182540000000
0!
0'
0/
#182550000000
1!
1'
1/
#182560000000
0!
0'
0/
#182570000000
1!
1'
1/
#182580000000
0!
0'
0/
#182590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#182600000000
0!
0'
0/
#182610000000
1!
1'
1/
#182620000000
0!
0'
0/
#182630000000
1!
1'
1/
#182640000000
0!
0'
0/
#182650000000
1!
1'
1/
#182660000000
0!
0'
0/
#182670000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#182680000000
0!
0'
0/
#182690000000
1!
1'
1/
#182700000000
0!
0'
0/
#182710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#182720000000
0!
0'
0/
#182730000000
1!
1'
1/
#182740000000
0!
0'
0/
#182750000000
#182760000000
1!
1'
1/
#182770000000
0!
0'
0/
#182780000000
1!
1'
1/
#182790000000
0!
1"
0'
1(
0/
10
#182800000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#182810000000
0!
0'
0/
#182820000000
1!
1'
1/
#182830000000
0!
0'
0/
#182840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#182850000000
0!
0'
0/
#182860000000
1!
1'
1/
#182870000000
0!
1"
0'
1(
0/
10
#182880000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#182890000000
0!
1$
0'
1+
0/
#182900000000
1!
1'
1/
#182910000000
0!
0'
0/
#182920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#182930000000
0!
0'
0/
#182940000000
1!
1'
1/
#182950000000
0!
0'
0/
#182960000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#182970000000
0!
0'
0/
#182980000000
1!
1'
1/
#182990000000
0!
0'
0/
#183000000000
1!
1'
1/
#183010000000
0!
0'
0/
#183020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#183030000000
0!
0'
0/
#183040000000
1!
1'
1/
#183050000000
0!
0'
0/
#183060000000
1!
1'
1/
#183070000000
0!
0'
0/
#183080000000
1!
1'
1/
#183090000000
0!
0'
0/
#183100000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#183110000000
0!
0'
0/
#183120000000
1!
1'
1/
#183130000000
0!
0'
0/
#183140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#183150000000
0!
0'
0/
#183160000000
1!
1'
1/
#183170000000
0!
0'
0/
#183180000000
#183190000000
1!
1'
1/
#183200000000
0!
0'
0/
#183210000000
1!
1'
1/
#183220000000
0!
1"
0'
1(
0/
10
#183230000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#183240000000
0!
0'
0/
#183250000000
1!
1'
1/
#183260000000
0!
0'
0/
#183270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#183280000000
0!
0'
0/
#183290000000
1!
1'
1/
#183300000000
0!
1"
0'
1(
0/
10
#183310000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#183320000000
0!
1$
0'
1+
0/
#183330000000
1!
1'
1/
#183340000000
0!
0'
0/
#183350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#183360000000
0!
0'
0/
#183370000000
1!
1'
1/
#183380000000
0!
0'
0/
#183390000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#183400000000
0!
0'
0/
#183410000000
1!
1'
1/
#183420000000
0!
0'
0/
#183430000000
1!
1'
1/
#183440000000
0!
0'
0/
#183450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#183460000000
0!
0'
0/
#183470000000
1!
1'
1/
#183480000000
0!
0'
0/
#183490000000
1!
1'
1/
#183500000000
0!
0'
0/
#183510000000
1!
1'
1/
#183520000000
0!
0'
0/
#183530000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#183540000000
0!
0'
0/
#183550000000
1!
1'
1/
#183560000000
0!
0'
0/
#183570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#183580000000
0!
0'
0/
#183590000000
1!
1'
1/
#183600000000
0!
0'
0/
#183610000000
#183620000000
1!
1'
1/
#183630000000
0!
0'
0/
#183640000000
1!
1'
1/
#183650000000
0!
1"
0'
1(
0/
10
#183660000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#183670000000
0!
0'
0/
#183680000000
1!
1'
1/
#183690000000
0!
0'
0/
#183700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#183710000000
0!
0'
0/
#183720000000
1!
1'
1/
#183730000000
0!
1"
0'
1(
0/
10
#183740000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#183750000000
0!
1$
0'
1+
0/
#183760000000
1!
1'
1/
#183770000000
0!
0'
0/
#183780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#183790000000
0!
0'
0/
#183800000000
1!
1'
1/
#183810000000
0!
0'
0/
#183820000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#183830000000
0!
0'
0/
#183840000000
1!
1'
1/
#183850000000
0!
0'
0/
#183860000000
1!
1'
1/
#183870000000
0!
0'
0/
#183880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#183890000000
0!
0'
0/
#183900000000
1!
1'
1/
#183910000000
0!
0'
0/
#183920000000
1!
1'
1/
#183930000000
0!
0'
0/
#183940000000
1!
1'
1/
#183950000000
0!
0'
0/
#183960000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#183970000000
0!
0'
0/
#183980000000
1!
1'
1/
#183990000000
0!
0'
0/
#184000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#184010000000
0!
0'
0/
#184020000000
1!
1'
1/
#184030000000
0!
0'
0/
#184040000000
#184050000000
1!
1'
1/
#184060000000
0!
0'
0/
#184070000000
1!
1'
1/
#184080000000
0!
1"
0'
1(
0/
10
#184090000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#184100000000
0!
0'
0/
#184110000000
1!
1'
1/
#184120000000
0!
0'
0/
#184130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#184140000000
0!
0'
0/
#184150000000
1!
1'
1/
#184160000000
0!
1"
0'
1(
0/
10
#184170000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#184180000000
0!
1$
0'
1+
0/
#184190000000
1!
1'
1/
#184200000000
0!
0'
0/
#184210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#184220000000
0!
0'
0/
#184230000000
1!
1'
1/
#184240000000
0!
0'
0/
#184250000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#184260000000
0!
0'
0/
#184270000000
1!
1'
1/
#184280000000
0!
0'
0/
#184290000000
1!
1'
1/
#184300000000
0!
0'
0/
#184310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#184320000000
0!
0'
0/
#184330000000
1!
1'
1/
#184340000000
0!
0'
0/
#184350000000
1!
1'
1/
#184360000000
0!
0'
0/
#184370000000
1!
1'
1/
#184380000000
0!
0'
0/
#184390000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#184400000000
0!
0'
0/
#184410000000
1!
1'
1/
#184420000000
0!
0'
0/
#184430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#184440000000
0!
0'
0/
#184450000000
1!
1'
1/
#184460000000
0!
0'
0/
#184470000000
#184480000000
1!
1'
1/
#184490000000
0!
0'
0/
#184500000000
1!
1'
1/
#184510000000
0!
1"
0'
1(
0/
10
#184520000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#184530000000
0!
0'
0/
#184540000000
1!
1'
1/
#184550000000
0!
0'
0/
#184560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#184570000000
0!
0'
0/
#184580000000
1!
1'
1/
#184590000000
0!
1"
0'
1(
0/
10
#184600000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#184610000000
0!
1$
0'
1+
0/
#184620000000
1!
1'
1/
#184630000000
0!
0'
0/
#184640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#184650000000
0!
0'
0/
#184660000000
1!
1'
1/
#184670000000
0!
0'
0/
#184680000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#184690000000
0!
0'
0/
#184700000000
1!
1'
1/
#184710000000
0!
0'
0/
#184720000000
1!
1'
1/
#184730000000
0!
0'
0/
#184740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#184750000000
0!
0'
0/
#184760000000
1!
1'
1/
#184770000000
0!
0'
0/
#184780000000
1!
1'
1/
#184790000000
0!
0'
0/
#184800000000
1!
1'
1/
#184810000000
0!
0'
0/
#184820000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#184830000000
0!
0'
0/
#184840000000
1!
1'
1/
#184850000000
0!
0'
0/
#184860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#184870000000
0!
0'
0/
#184880000000
1!
1'
1/
#184890000000
0!
0'
0/
#184900000000
#184910000000
1!
1'
1/
#184920000000
0!
0'
0/
#184930000000
1!
1'
1/
#184940000000
0!
1"
0'
1(
0/
10
#184950000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#184960000000
0!
0'
0/
#184970000000
1!
1'
1/
#184980000000
0!
0'
0/
#184990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#185000000000
0!
0'
0/
#185010000000
1!
1'
1/
#185020000000
0!
1"
0'
1(
0/
10
#185030000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#185040000000
0!
1$
0'
1+
0/
#185050000000
1!
1'
1/
#185060000000
0!
0'
0/
#185070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#185080000000
0!
0'
0/
#185090000000
1!
1'
1/
#185100000000
0!
0'
0/
#185110000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#185120000000
0!
0'
0/
#185130000000
1!
1'
1/
#185140000000
0!
0'
0/
#185150000000
1!
1'
1/
#185160000000
0!
0'
0/
#185170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#185180000000
0!
0'
0/
#185190000000
1!
1'
1/
#185200000000
0!
0'
0/
#185210000000
1!
1'
1/
#185220000000
0!
0'
0/
#185230000000
1!
1'
1/
#185240000000
0!
0'
0/
#185250000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#185260000000
0!
0'
0/
#185270000000
1!
1'
1/
#185280000000
0!
0'
0/
#185290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#185300000000
0!
0'
0/
#185310000000
1!
1'
1/
#185320000000
0!
0'
0/
#185330000000
#185340000000
1!
1'
1/
#185350000000
0!
0'
0/
#185360000000
1!
1'
1/
#185370000000
0!
1"
0'
1(
0/
10
#185380000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#185390000000
0!
0'
0/
#185400000000
1!
1'
1/
#185410000000
0!
0'
0/
#185420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#185430000000
0!
0'
0/
#185440000000
1!
1'
1/
#185450000000
0!
1"
0'
1(
0/
10
#185460000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#185470000000
0!
1$
0'
1+
0/
#185480000000
1!
1'
1/
#185490000000
0!
0'
0/
#185500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#185510000000
0!
0'
0/
#185520000000
1!
1'
1/
#185530000000
0!
0'
0/
#185540000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#185550000000
0!
0'
0/
#185560000000
1!
1'
1/
#185570000000
0!
0'
0/
#185580000000
1!
1'
1/
#185590000000
0!
0'
0/
#185600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#185610000000
0!
0'
0/
#185620000000
1!
1'
1/
#185630000000
0!
0'
0/
#185640000000
1!
1'
1/
#185650000000
0!
0'
0/
#185660000000
1!
1'
1/
#185670000000
0!
0'
0/
#185680000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#185690000000
0!
0'
0/
#185700000000
1!
1'
1/
#185710000000
0!
0'
0/
#185720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#185730000000
0!
0'
0/
#185740000000
1!
1'
1/
#185750000000
0!
0'
0/
#185760000000
#185770000000
1!
1'
1/
#185780000000
0!
0'
0/
#185790000000
1!
1'
1/
#185800000000
0!
1"
0'
1(
0/
10
#185810000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#185820000000
0!
0'
0/
#185830000000
1!
1'
1/
#185840000000
0!
0'
0/
#185850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#185860000000
0!
0'
0/
#185870000000
1!
1'
1/
#185880000000
0!
1"
0'
1(
0/
10
#185890000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#185900000000
0!
1$
0'
1+
0/
#185910000000
1!
1'
1/
#185920000000
0!
0'
0/
#185930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#185940000000
0!
0'
0/
#185950000000
1!
1'
1/
#185960000000
0!
0'
0/
#185970000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#185980000000
0!
0'
0/
#185990000000
1!
1'
1/
#186000000000
0!
0'
0/
#186010000000
1!
1'
1/
#186020000000
0!
0'
0/
#186030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#186040000000
0!
0'
0/
#186050000000
1!
1'
1/
#186060000000
0!
0'
0/
#186070000000
1!
1'
1/
#186080000000
0!
0'
0/
#186090000000
1!
1'
1/
#186100000000
0!
0'
0/
#186110000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#186120000000
0!
0'
0/
#186130000000
1!
1'
1/
#186140000000
0!
0'
0/
#186150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#186160000000
0!
0'
0/
#186170000000
1!
1'
1/
#186180000000
0!
0'
0/
#186190000000
#186200000000
1!
1'
1/
#186210000000
0!
0'
0/
#186220000000
1!
1'
1/
#186230000000
0!
1"
0'
1(
0/
10
#186240000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#186250000000
0!
0'
0/
#186260000000
1!
1'
1/
#186270000000
0!
0'
0/
#186280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#186290000000
0!
0'
0/
#186300000000
1!
1'
1/
#186310000000
0!
1"
0'
1(
0/
10
#186320000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#186330000000
0!
1$
0'
1+
0/
#186340000000
1!
1'
1/
#186350000000
0!
0'
0/
#186360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#186370000000
0!
0'
0/
#186380000000
1!
1'
1/
#186390000000
0!
0'
0/
#186400000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#186410000000
0!
0'
0/
#186420000000
1!
1'
1/
#186430000000
0!
0'
0/
#186440000000
1!
1'
1/
#186450000000
0!
0'
0/
#186460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#186470000000
0!
0'
0/
#186480000000
1!
1'
1/
#186490000000
0!
0'
0/
#186500000000
1!
1'
1/
#186510000000
0!
0'
0/
#186520000000
1!
1'
1/
#186530000000
0!
0'
0/
#186540000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#186550000000
0!
0'
0/
#186560000000
1!
1'
1/
#186570000000
0!
0'
0/
#186580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#186590000000
0!
0'
0/
#186600000000
1!
1'
1/
#186610000000
0!
0'
0/
#186620000000
#186630000000
1!
1'
1/
#186640000000
0!
0'
0/
#186650000000
1!
1'
1/
#186660000000
0!
1"
0'
1(
0/
10
#186670000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#186680000000
0!
0'
0/
#186690000000
1!
1'
1/
#186700000000
0!
0'
0/
#186710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#186720000000
0!
0'
0/
#186730000000
1!
1'
1/
#186740000000
0!
1"
0'
1(
0/
10
#186750000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#186760000000
0!
1$
0'
1+
0/
#186770000000
1!
1'
1/
#186780000000
0!
0'
0/
#186790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#186800000000
0!
0'
0/
#186810000000
1!
1'
1/
#186820000000
0!
0'
0/
#186830000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#186840000000
0!
0'
0/
#186850000000
1!
1'
1/
#186860000000
0!
0'
0/
#186870000000
1!
1'
1/
#186880000000
0!
0'
0/
#186890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#186900000000
0!
0'
0/
#186910000000
1!
1'
1/
#186920000000
0!
0'
0/
#186930000000
1!
1'
1/
#186940000000
0!
0'
0/
#186950000000
1!
1'
1/
#186960000000
0!
0'
0/
#186970000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#186980000000
0!
0'
0/
#186990000000
1!
1'
1/
#187000000000
0!
0'
0/
#187010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#187020000000
0!
0'
0/
#187030000000
1!
1'
1/
#187040000000
0!
0'
0/
#187050000000
#187060000000
1!
1'
1/
#187070000000
0!
0'
0/
#187080000000
1!
1'
1/
#187090000000
0!
1"
0'
1(
0/
10
#187100000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#187110000000
0!
0'
0/
#187120000000
1!
1'
1/
#187130000000
0!
0'
0/
#187140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#187150000000
0!
0'
0/
#187160000000
1!
1'
1/
#187170000000
0!
1"
0'
1(
0/
10
#187180000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#187190000000
0!
1$
0'
1+
0/
#187200000000
1!
1'
1/
#187210000000
0!
0'
0/
#187220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#187230000000
0!
0'
0/
#187240000000
1!
1'
1/
#187250000000
0!
0'
0/
#187260000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#187270000000
0!
0'
0/
#187280000000
1!
1'
1/
#187290000000
0!
0'
0/
#187300000000
1!
1'
1/
#187310000000
0!
0'
0/
#187320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#187330000000
0!
0'
0/
#187340000000
1!
1'
1/
#187350000000
0!
0'
0/
#187360000000
1!
1'
1/
#187370000000
0!
0'
0/
#187380000000
1!
1'
1/
#187390000000
0!
0'
0/
#187400000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#187410000000
0!
0'
0/
#187420000000
1!
1'
1/
#187430000000
0!
0'
0/
#187440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#187450000000
0!
0'
0/
#187460000000
1!
1'
1/
#187470000000
0!
0'
0/
#187480000000
#187490000000
1!
1'
1/
#187500000000
0!
0'
0/
#187510000000
1!
1'
1/
#187520000000
0!
1"
0'
1(
0/
10
#187530000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#187540000000
0!
0'
0/
#187550000000
1!
1'
1/
#187560000000
0!
0'
0/
#187570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#187580000000
0!
0'
0/
#187590000000
1!
1'
1/
#187600000000
0!
1"
0'
1(
0/
10
#187610000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#187620000000
0!
1$
0'
1+
0/
#187630000000
1!
1'
1/
#187640000000
0!
0'
0/
#187650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#187660000000
0!
0'
0/
#187670000000
1!
1'
1/
#187680000000
0!
0'
0/
#187690000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#187700000000
0!
0'
0/
#187710000000
1!
1'
1/
#187720000000
0!
0'
0/
#187730000000
1!
1'
1/
#187740000000
0!
0'
0/
#187750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#187760000000
0!
0'
0/
#187770000000
1!
1'
1/
#187780000000
0!
0'
0/
#187790000000
1!
1'
1/
#187800000000
0!
0'
0/
#187810000000
1!
1'
1/
#187820000000
0!
0'
0/
#187830000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#187840000000
0!
0'
0/
#187850000000
1!
1'
1/
#187860000000
0!
0'
0/
#187870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#187880000000
0!
0'
0/
#187890000000
1!
1'
1/
#187900000000
0!
0'
0/
#187910000000
#187920000000
1!
1'
1/
#187930000000
0!
0'
0/
#187940000000
1!
1'
1/
#187950000000
0!
1"
0'
1(
0/
10
#187960000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#187970000000
0!
0'
0/
#187980000000
1!
1'
1/
#187990000000
0!
0'
0/
#188000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#188010000000
0!
0'
0/
#188020000000
1!
1'
1/
#188030000000
0!
1"
0'
1(
0/
10
#188040000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#188050000000
0!
1$
0'
1+
0/
#188060000000
1!
1'
1/
#188070000000
0!
0'
0/
#188080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#188090000000
0!
0'
0/
#188100000000
1!
1'
1/
#188110000000
0!
0'
0/
#188120000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#188130000000
0!
0'
0/
#188140000000
1!
1'
1/
#188150000000
0!
0'
0/
#188160000000
1!
1'
1/
#188170000000
0!
0'
0/
#188180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#188190000000
0!
0'
0/
#188200000000
1!
1'
1/
#188210000000
0!
0'
0/
#188220000000
1!
1'
1/
#188230000000
0!
0'
0/
#188240000000
1!
1'
1/
#188250000000
0!
0'
0/
#188260000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#188270000000
0!
0'
0/
#188280000000
1!
1'
1/
#188290000000
0!
0'
0/
#188300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#188310000000
0!
0'
0/
#188320000000
1!
1'
1/
#188330000000
0!
0'
0/
#188340000000
#188350000000
1!
1'
1/
#188360000000
0!
0'
0/
#188370000000
1!
1'
1/
#188380000000
0!
1"
0'
1(
0/
10
#188390000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#188400000000
0!
0'
0/
#188410000000
1!
1'
1/
#188420000000
0!
0'
0/
#188430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#188440000000
0!
0'
0/
#188450000000
1!
1'
1/
#188460000000
0!
1"
0'
1(
0/
10
#188470000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#188480000000
0!
1$
0'
1+
0/
#188490000000
1!
1'
1/
#188500000000
0!
0'
0/
#188510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#188520000000
0!
0'
0/
#188530000000
1!
1'
1/
#188540000000
0!
0'
0/
#188550000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#188560000000
0!
0'
0/
#188570000000
1!
1'
1/
#188580000000
0!
0'
0/
#188590000000
1!
1'
1/
#188600000000
0!
0'
0/
#188610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#188620000000
0!
0'
0/
#188630000000
1!
1'
1/
#188640000000
0!
0'
0/
#188650000000
1!
1'
1/
#188660000000
0!
0'
0/
#188670000000
1!
1'
1/
#188680000000
0!
0'
0/
#188690000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#188700000000
0!
0'
0/
#188710000000
1!
1'
1/
#188720000000
0!
0'
0/
#188730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#188740000000
0!
0'
0/
#188750000000
1!
1'
1/
#188760000000
0!
0'
0/
#188770000000
#188780000000
1!
1'
1/
#188790000000
0!
0'
0/
#188800000000
1!
1'
1/
#188810000000
0!
1"
0'
1(
0/
10
#188820000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#188830000000
0!
0'
0/
#188840000000
1!
1'
1/
#188850000000
0!
0'
0/
#188860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#188870000000
0!
0'
0/
#188880000000
1!
1'
1/
#188890000000
0!
1"
0'
1(
0/
10
#188900000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#188910000000
0!
1$
0'
1+
0/
#188920000000
1!
1'
1/
#188930000000
0!
0'
0/
#188940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#188950000000
0!
0'
0/
#188960000000
1!
1'
1/
#188970000000
0!
0'
0/
#188980000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#188990000000
0!
0'
0/
#189000000000
1!
1'
1/
#189010000000
0!
0'
0/
#189020000000
1!
1'
1/
#189030000000
0!
0'
0/
#189040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#189050000000
0!
0'
0/
#189060000000
1!
1'
1/
#189070000000
0!
0'
0/
#189080000000
1!
1'
1/
#189090000000
0!
0'
0/
#189100000000
1!
1'
1/
#189110000000
0!
0'
0/
#189120000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#189130000000
0!
0'
0/
#189140000000
1!
1'
1/
#189150000000
0!
0'
0/
#189160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#189170000000
0!
0'
0/
#189180000000
1!
1'
1/
#189190000000
0!
0'
0/
#189200000000
#189210000000
1!
1'
1/
#189220000000
0!
0'
0/
#189230000000
1!
1'
1/
#189240000000
0!
1"
0'
1(
0/
10
#189250000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#189260000000
0!
0'
0/
#189270000000
1!
1'
1/
#189280000000
0!
0'
0/
#189290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#189300000000
0!
0'
0/
#189310000000
1!
1'
1/
#189320000000
0!
1"
0'
1(
0/
10
#189330000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#189340000000
0!
1$
0'
1+
0/
#189350000000
1!
1'
1/
#189360000000
0!
0'
0/
#189370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#189380000000
0!
0'
0/
#189390000000
1!
1'
1/
#189400000000
0!
0'
0/
#189410000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#189420000000
0!
0'
0/
#189430000000
1!
1'
1/
#189440000000
0!
0'
0/
#189450000000
1!
1'
1/
#189460000000
0!
0'
0/
#189470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#189480000000
0!
0'
0/
#189490000000
1!
1'
1/
#189500000000
0!
0'
0/
#189510000000
1!
1'
1/
#189520000000
0!
0'
0/
#189530000000
1!
1'
1/
#189540000000
0!
0'
0/
#189550000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#189560000000
0!
0'
0/
#189570000000
1!
1'
1/
#189580000000
0!
0'
0/
#189590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#189600000000
0!
0'
0/
#189610000000
1!
1'
1/
#189620000000
0!
0'
0/
#189630000000
#189640000000
1!
1'
1/
#189650000000
0!
0'
0/
#189660000000
1!
1'
1/
#189670000000
0!
1"
0'
1(
0/
10
#189680000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#189690000000
0!
0'
0/
#189700000000
1!
1'
1/
#189710000000
0!
0'
0/
#189720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#189730000000
0!
0'
0/
#189740000000
1!
1'
1/
#189750000000
0!
1"
0'
1(
0/
10
#189760000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#189770000000
0!
1$
0'
1+
0/
#189780000000
1!
1'
1/
#189790000000
0!
0'
0/
#189800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#189810000000
0!
0'
0/
#189820000000
1!
1'
1/
#189830000000
0!
0'
0/
#189840000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#189850000000
0!
0'
0/
#189860000000
1!
1'
1/
#189870000000
0!
0'
0/
#189880000000
1!
1'
1/
#189890000000
0!
0'
0/
#189900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#189910000000
0!
0'
0/
#189920000000
1!
1'
1/
#189930000000
0!
0'
0/
#189940000000
1!
1'
1/
#189950000000
0!
0'
0/
#189960000000
1!
1'
1/
#189970000000
0!
0'
0/
#189980000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#189990000000
0!
0'
0/
#190000000000
1!
1'
1/
#190010000000
0!
0'
0/
#190020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#190030000000
0!
0'
0/
#190040000000
1!
1'
1/
#190050000000
0!
0'
0/
#190060000000
#190070000000
1!
1'
1/
#190080000000
0!
0'
0/
#190090000000
1!
1'
1/
#190100000000
0!
1"
0'
1(
0/
10
#190110000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#190120000000
0!
0'
0/
#190130000000
1!
1'
1/
#190140000000
0!
0'
0/
#190150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#190160000000
0!
0'
0/
#190170000000
1!
1'
1/
#190180000000
0!
1"
0'
1(
0/
10
#190190000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#190200000000
0!
1$
0'
1+
0/
#190210000000
1!
1'
1/
#190220000000
0!
0'
0/
#190230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#190240000000
0!
0'
0/
#190250000000
1!
1'
1/
#190260000000
0!
0'
0/
#190270000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#190280000000
0!
0'
0/
#190290000000
1!
1'
1/
#190300000000
0!
0'
0/
#190310000000
1!
1'
1/
#190320000000
0!
0'
0/
#190330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#190340000000
0!
0'
0/
#190350000000
1!
1'
1/
#190360000000
0!
0'
0/
#190370000000
1!
1'
1/
#190380000000
0!
0'
0/
#190390000000
1!
1'
1/
#190400000000
0!
0'
0/
#190410000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#190420000000
0!
0'
0/
#190430000000
1!
1'
1/
#190440000000
0!
0'
0/
#190450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#190460000000
0!
0'
0/
#190470000000
1!
1'
1/
#190480000000
0!
0'
0/
#190490000000
#190500000000
1!
1'
1/
#190510000000
0!
0'
0/
#190520000000
1!
1'
1/
#190530000000
0!
1"
0'
1(
0/
10
#190540000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#190550000000
0!
0'
0/
#190560000000
1!
1'
1/
#190570000000
0!
0'
0/
#190580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#190590000000
0!
0'
0/
#190600000000
1!
1'
1/
#190610000000
0!
1"
0'
1(
0/
10
#190620000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#190630000000
0!
1$
0'
1+
0/
#190640000000
1!
1'
1/
#190650000000
0!
0'
0/
#190660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#190670000000
0!
0'
0/
#190680000000
1!
1'
1/
#190690000000
0!
0'
0/
#190700000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#190710000000
0!
0'
0/
#190720000000
1!
1'
1/
#190730000000
0!
0'
0/
#190740000000
1!
1'
1/
#190750000000
0!
0'
0/
#190760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#190770000000
0!
0'
0/
#190780000000
1!
1'
1/
#190790000000
0!
0'
0/
#190800000000
1!
1'
1/
#190810000000
0!
0'
0/
#190820000000
1!
1'
1/
#190830000000
0!
0'
0/
#190840000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#190850000000
0!
0'
0/
#190860000000
1!
1'
1/
#190870000000
0!
0'
0/
#190880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#190890000000
0!
0'
0/
#190900000000
1!
1'
1/
#190910000000
0!
0'
0/
#190920000000
#190930000000
1!
1'
1/
#190940000000
0!
0'
0/
#190950000000
1!
1'
1/
#190960000000
0!
1"
0'
1(
0/
10
#190970000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#190980000000
0!
0'
0/
#190990000000
1!
1'
1/
#191000000000
0!
0'
0/
#191010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#191020000000
0!
0'
0/
#191030000000
1!
1'
1/
#191040000000
0!
1"
0'
1(
0/
10
#191050000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#191060000000
0!
1$
0'
1+
0/
#191070000000
1!
1'
1/
#191080000000
0!
0'
0/
#191090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#191100000000
0!
0'
0/
#191110000000
1!
1'
1/
#191120000000
0!
0'
0/
#191130000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#191140000000
0!
0'
0/
#191150000000
1!
1'
1/
#191160000000
0!
0'
0/
#191170000000
1!
1'
1/
#191180000000
0!
0'
0/
#191190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#191200000000
0!
0'
0/
#191210000000
1!
1'
1/
#191220000000
0!
0'
0/
#191230000000
1!
1'
1/
#191240000000
0!
0'
0/
#191250000000
1!
1'
1/
#191260000000
0!
0'
0/
#191270000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#191280000000
0!
0'
0/
#191290000000
1!
1'
1/
#191300000000
0!
0'
0/
#191310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#191320000000
0!
0'
0/
#191330000000
1!
1'
1/
#191340000000
0!
0'
0/
#191350000000
#191360000000
1!
1'
1/
#191370000000
0!
0'
0/
#191380000000
1!
1'
1/
#191390000000
0!
1"
0'
1(
0/
10
#191400000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#191410000000
0!
0'
0/
#191420000000
1!
1'
1/
#191430000000
0!
0'
0/
#191440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#191450000000
0!
0'
0/
#191460000000
1!
1'
1/
#191470000000
0!
1"
0'
1(
0/
10
#191480000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#191490000000
0!
1$
0'
1+
0/
#191500000000
1!
1'
1/
#191510000000
0!
0'
0/
#191520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#191530000000
0!
0'
0/
#191540000000
1!
1'
1/
#191550000000
0!
0'
0/
#191560000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#191570000000
0!
0'
0/
#191580000000
1!
1'
1/
#191590000000
0!
0'
0/
#191600000000
1!
1'
1/
#191610000000
0!
0'
0/
#191620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#191630000000
0!
0'
0/
#191640000000
1!
1'
1/
#191650000000
0!
0'
0/
#191660000000
1!
1'
1/
#191670000000
0!
0'
0/
#191680000000
1!
1'
1/
#191690000000
0!
0'
0/
#191700000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#191710000000
0!
0'
0/
#191720000000
1!
1'
1/
#191730000000
0!
0'
0/
#191740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#191750000000
0!
0'
0/
#191760000000
1!
1'
1/
#191770000000
0!
0'
0/
#191780000000
#191790000000
1!
1'
1/
#191800000000
0!
0'
0/
#191810000000
1!
1'
1/
#191820000000
0!
1"
0'
1(
0/
10
#191830000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#191840000000
0!
0'
0/
#191850000000
1!
1'
1/
#191860000000
0!
0'
0/
#191870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#191880000000
0!
0'
0/
#191890000000
1!
1'
1/
#191900000000
0!
1"
0'
1(
0/
10
#191910000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#191920000000
0!
1$
0'
1+
0/
#191930000000
1!
1'
1/
#191940000000
0!
0'
0/
#191950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#191960000000
0!
0'
0/
#191970000000
1!
1'
1/
#191980000000
0!
0'
0/
#191990000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#192000000000
0!
0'
0/
#192010000000
1!
1'
1/
#192020000000
0!
0'
0/
#192030000000
1!
1'
1/
#192040000000
0!
0'
0/
#192050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#192060000000
0!
0'
0/
#192070000000
1!
1'
1/
#192080000000
0!
0'
0/
#192090000000
1!
1'
1/
#192100000000
0!
0'
0/
#192110000000
1!
1'
1/
#192120000000
0!
0'
0/
#192130000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#192140000000
0!
0'
0/
#192150000000
1!
1'
1/
#192160000000
0!
0'
0/
#192170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#192180000000
0!
0'
0/
#192190000000
1!
1'
1/
#192200000000
0!
0'
0/
#192210000000
#192220000000
1!
1'
1/
#192230000000
0!
0'
0/
#192240000000
1!
1'
1/
#192250000000
0!
1"
0'
1(
0/
10
#192260000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#192270000000
0!
0'
0/
#192280000000
1!
1'
1/
#192290000000
0!
0'
0/
#192300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#192310000000
0!
0'
0/
#192320000000
1!
1'
1/
#192330000000
0!
1"
0'
1(
0/
10
#192340000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#192350000000
0!
1$
0'
1+
0/
#192360000000
1!
1'
1/
#192370000000
0!
0'
0/
#192380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#192390000000
0!
0'
0/
#192400000000
1!
1'
1/
#192410000000
0!
0'
0/
#192420000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#192430000000
0!
0'
0/
#192440000000
1!
1'
1/
#192450000000
0!
0'
0/
#192460000000
1!
1'
1/
#192470000000
0!
0'
0/
#192480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#192490000000
0!
0'
0/
#192500000000
1!
1'
1/
#192510000000
0!
0'
0/
#192520000000
1!
1'
1/
#192530000000
0!
0'
0/
#192540000000
1!
1'
1/
#192550000000
0!
0'
0/
#192560000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#192570000000
0!
0'
0/
#192580000000
1!
1'
1/
#192590000000
0!
0'
0/
#192600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#192610000000
0!
0'
0/
#192620000000
1!
1'
1/
#192630000000
0!
0'
0/
#192640000000
#192650000000
1!
1'
1/
#192660000000
0!
0'
0/
#192670000000
1!
1'
1/
#192680000000
0!
1"
0'
1(
0/
10
#192690000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#192700000000
0!
0'
0/
#192710000000
1!
1'
1/
#192720000000
0!
0'
0/
#192730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#192740000000
0!
0'
0/
#192750000000
1!
1'
1/
#192760000000
0!
1"
0'
1(
0/
10
#192770000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#192780000000
0!
1$
0'
1+
0/
#192790000000
1!
1'
1/
#192800000000
0!
0'
0/
#192810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#192820000000
0!
0'
0/
#192830000000
1!
1'
1/
#192840000000
0!
0'
0/
#192850000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#192860000000
0!
0'
0/
#192870000000
1!
1'
1/
#192880000000
0!
0'
0/
#192890000000
1!
1'
1/
#192900000000
0!
0'
0/
#192910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#192920000000
0!
0'
0/
#192930000000
1!
1'
1/
#192940000000
0!
0'
0/
#192950000000
1!
1'
1/
#192960000000
0!
0'
0/
#192970000000
1!
1'
1/
#192980000000
0!
0'
0/
#192990000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#193000000000
0!
0'
0/
#193010000000
1!
1'
1/
#193020000000
0!
0'
0/
#193030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#193040000000
0!
0'
0/
#193050000000
1!
1'
1/
#193060000000
0!
0'
0/
#193070000000
#193080000000
1!
1'
1/
#193090000000
0!
0'
0/
#193100000000
1!
1'
1/
#193110000000
0!
1"
0'
1(
0/
10
#193120000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#193130000000
0!
0'
0/
#193140000000
1!
1'
1/
#193150000000
0!
0'
0/
#193160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#193170000000
0!
0'
0/
#193180000000
1!
1'
1/
#193190000000
0!
1"
0'
1(
0/
10
#193200000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#193210000000
0!
1$
0'
1+
0/
#193220000000
1!
1'
1/
#193230000000
0!
0'
0/
#193240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#193250000000
0!
0'
0/
#193260000000
1!
1'
1/
#193270000000
0!
0'
0/
#193280000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#193290000000
0!
0'
0/
#193300000000
1!
1'
1/
#193310000000
0!
0'
0/
#193320000000
1!
1'
1/
#193330000000
0!
0'
0/
#193340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#193350000000
0!
0'
0/
#193360000000
1!
1'
1/
#193370000000
0!
0'
0/
#193380000000
1!
1'
1/
#193390000000
0!
0'
0/
#193400000000
1!
1'
1/
#193410000000
0!
0'
0/
#193420000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#193430000000
0!
0'
0/
#193440000000
1!
1'
1/
#193450000000
0!
0'
0/
#193460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#193470000000
0!
0'
0/
#193480000000
1!
1'
1/
#193490000000
0!
0'
0/
#193500000000
#193510000000
1!
1'
1/
#193520000000
0!
0'
0/
#193530000000
1!
1'
1/
#193540000000
0!
1"
0'
1(
0/
10
#193550000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#193560000000
0!
0'
0/
#193570000000
1!
1'
1/
#193580000000
0!
0'
0/
#193590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#193600000000
0!
0'
0/
#193610000000
1!
1'
1/
#193620000000
0!
1"
0'
1(
0/
10
#193630000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#193640000000
0!
1$
0'
1+
0/
#193650000000
1!
1'
1/
#193660000000
0!
0'
0/
#193670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#193680000000
0!
0'
0/
#193690000000
1!
1'
1/
#193700000000
0!
0'
0/
#193710000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#193720000000
0!
0'
0/
#193730000000
1!
1'
1/
#193740000000
0!
0'
0/
#193750000000
1!
1'
1/
#193760000000
0!
0'
0/
#193770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#193780000000
0!
0'
0/
#193790000000
1!
1'
1/
#193800000000
0!
0'
0/
#193810000000
1!
1'
1/
#193820000000
0!
0'
0/
#193830000000
1!
1'
1/
#193840000000
0!
0'
0/
#193850000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#193860000000
0!
0'
0/
#193870000000
1!
1'
1/
#193880000000
0!
0'
0/
#193890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#193900000000
0!
0'
0/
#193910000000
1!
1'
1/
#193920000000
0!
0'
0/
#193930000000
#193940000000
1!
1'
1/
#193950000000
0!
0'
0/
#193960000000
1!
1'
1/
#193970000000
0!
1"
0'
1(
0/
10
#193980000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#193990000000
0!
0'
0/
#194000000000
1!
1'
1/
#194010000000
0!
0'
0/
#194020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#194030000000
0!
0'
0/
#194040000000
1!
1'
1/
#194050000000
0!
1"
0'
1(
0/
10
#194060000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#194070000000
0!
1$
0'
1+
0/
#194080000000
1!
1'
1/
#194090000000
0!
0'
0/
#194100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#194110000000
0!
0'
0/
#194120000000
1!
1'
1/
#194130000000
0!
0'
0/
#194140000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#194150000000
0!
0'
0/
#194160000000
1!
1'
1/
#194170000000
0!
0'
0/
#194180000000
1!
1'
1/
#194190000000
0!
0'
0/
#194200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#194210000000
0!
0'
0/
#194220000000
1!
1'
1/
#194230000000
0!
0'
0/
#194240000000
1!
1'
1/
#194250000000
0!
0'
0/
#194260000000
1!
1'
1/
#194270000000
0!
0'
0/
#194280000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#194290000000
0!
0'
0/
#194300000000
1!
1'
1/
#194310000000
0!
0'
0/
#194320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#194330000000
0!
0'
0/
#194340000000
1!
1'
1/
#194350000000
0!
0'
0/
#194360000000
#194370000000
1!
1'
1/
#194380000000
0!
0'
0/
#194390000000
1!
1'
1/
#194400000000
0!
1"
0'
1(
0/
10
#194410000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#194420000000
0!
0'
0/
#194430000000
1!
1'
1/
#194440000000
0!
0'
0/
#194450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#194460000000
0!
0'
0/
#194470000000
1!
1'
1/
#194480000000
0!
1"
0'
1(
0/
10
#194490000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#194500000000
0!
1$
0'
1+
0/
#194510000000
1!
1'
1/
#194520000000
0!
0'
0/
#194530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#194540000000
0!
0'
0/
#194550000000
1!
1'
1/
#194560000000
0!
0'
0/
#194570000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#194580000000
0!
0'
0/
#194590000000
1!
1'
1/
#194600000000
0!
0'
0/
#194610000000
1!
1'
1/
#194620000000
0!
0'
0/
#194630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#194640000000
0!
0'
0/
#194650000000
1!
1'
1/
#194660000000
0!
0'
0/
#194670000000
1!
1'
1/
#194680000000
0!
0'
0/
#194690000000
1!
1'
1/
#194700000000
0!
0'
0/
#194710000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#194720000000
0!
0'
0/
#194730000000
1!
1'
1/
#194740000000
0!
0'
0/
#194750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#194760000000
0!
0'
0/
#194770000000
1!
1'
1/
#194780000000
0!
0'
0/
#194790000000
#194800000000
1!
1'
1/
#194810000000
0!
0'
0/
#194820000000
1!
1'
1/
#194830000000
0!
1"
0'
1(
0/
10
#194840000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#194850000000
0!
0'
0/
#194860000000
1!
1'
1/
#194870000000
0!
0'
0/
#194880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#194890000000
0!
0'
0/
#194900000000
1!
1'
1/
#194910000000
0!
1"
0'
1(
0/
10
#194920000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#194930000000
0!
1$
0'
1+
0/
#194940000000
1!
1'
1/
#194950000000
0!
0'
0/
#194960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#194970000000
0!
0'
0/
#194980000000
1!
1'
1/
#194990000000
0!
0'
0/
#195000000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#195010000000
0!
0'
0/
#195020000000
1!
1'
1/
#195030000000
0!
0'
0/
#195040000000
1!
1'
1/
#195050000000
0!
0'
0/
#195060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#195070000000
0!
0'
0/
#195080000000
1!
1'
1/
#195090000000
0!
0'
0/
#195100000000
1!
1'
1/
#195110000000
0!
0'
0/
#195120000000
1!
1'
1/
#195130000000
0!
0'
0/
#195140000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#195150000000
0!
0'
0/
#195160000000
1!
1'
1/
#195170000000
0!
0'
0/
#195180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#195190000000
0!
0'
0/
#195200000000
1!
1'
1/
#195210000000
0!
0'
0/
#195220000000
#195230000000
1!
1'
1/
#195240000000
0!
0'
0/
#195250000000
1!
1'
1/
#195260000000
0!
1"
0'
1(
0/
10
#195270000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#195280000000
0!
0'
0/
#195290000000
1!
1'
1/
#195300000000
0!
0'
0/
#195310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#195320000000
0!
0'
0/
#195330000000
1!
1'
1/
#195340000000
0!
1"
0'
1(
0/
10
#195350000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#195360000000
0!
1$
0'
1+
0/
#195370000000
1!
1'
1/
#195380000000
0!
0'
0/
#195390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#195400000000
0!
0'
0/
#195410000000
1!
1'
1/
#195420000000
0!
0'
0/
#195430000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#195440000000
0!
0'
0/
#195450000000
1!
1'
1/
#195460000000
0!
0'
0/
#195470000000
1!
1'
1/
#195480000000
0!
0'
0/
#195490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#195500000000
0!
0'
0/
#195510000000
1!
1'
1/
#195520000000
0!
0'
0/
#195530000000
1!
1'
1/
#195540000000
0!
0'
0/
#195550000000
1!
1'
1/
#195560000000
0!
0'
0/
#195570000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#195580000000
0!
0'
0/
#195590000000
1!
1'
1/
#195600000000
0!
0'
0/
#195610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#195620000000
0!
0'
0/
#195630000000
1!
1'
1/
#195640000000
0!
0'
0/
#195650000000
#195660000000
1!
1'
1/
#195670000000
0!
0'
0/
#195680000000
1!
1'
1/
#195690000000
0!
1"
0'
1(
0/
10
#195700000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#195710000000
0!
0'
0/
#195720000000
1!
1'
1/
#195730000000
0!
0'
0/
#195740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#195750000000
0!
0'
0/
#195760000000
1!
1'
1/
#195770000000
0!
1"
0'
1(
0/
10
#195780000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#195790000000
0!
1$
0'
1+
0/
#195800000000
1!
1'
1/
#195810000000
0!
0'
0/
#195820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#195830000000
0!
0'
0/
#195840000000
1!
1'
1/
#195850000000
0!
0'
0/
#195860000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#195870000000
0!
0'
0/
#195880000000
1!
1'
1/
#195890000000
0!
0'
0/
#195900000000
1!
1'
1/
#195910000000
0!
0'
0/
#195920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#195930000000
0!
0'
0/
#195940000000
1!
1'
1/
#195950000000
0!
0'
0/
#195960000000
1!
1'
1/
#195970000000
0!
0'
0/
#195980000000
1!
1'
1/
#195990000000
0!
0'
0/
#196000000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#196010000000
0!
0'
0/
#196020000000
1!
1'
1/
#196030000000
0!
0'
0/
#196040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#196050000000
0!
0'
0/
#196060000000
1!
1'
1/
#196070000000
0!
0'
0/
#196080000000
#196090000000
1!
1'
1/
#196100000000
0!
0'
0/
#196110000000
1!
1'
1/
#196120000000
0!
1"
0'
1(
0/
10
#196130000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#196140000000
0!
0'
0/
#196150000000
1!
1'
1/
#196160000000
0!
0'
0/
#196170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#196180000000
0!
0'
0/
#196190000000
1!
1'
1/
#196200000000
0!
1"
0'
1(
0/
10
#196210000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#196220000000
0!
1$
0'
1+
0/
#196230000000
1!
1'
1/
#196240000000
0!
0'
0/
#196250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#196260000000
0!
0'
0/
#196270000000
1!
1'
1/
#196280000000
0!
0'
0/
#196290000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#196300000000
0!
0'
0/
#196310000000
1!
1'
1/
#196320000000
0!
0'
0/
#196330000000
1!
1'
1/
#196340000000
0!
0'
0/
#196350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#196360000000
0!
0'
0/
#196370000000
1!
1'
1/
#196380000000
0!
0'
0/
#196390000000
1!
1'
1/
#196400000000
0!
0'
0/
#196410000000
1!
1'
1/
#196420000000
0!
0'
0/
#196430000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#196440000000
0!
0'
0/
#196450000000
1!
1'
1/
#196460000000
0!
0'
0/
#196470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#196480000000
0!
0'
0/
#196490000000
1!
1'
1/
#196500000000
0!
0'
0/
#196510000000
#196520000000
1!
1'
1/
#196530000000
0!
0'
0/
#196540000000
1!
1'
1/
#196550000000
0!
1"
0'
1(
0/
10
#196560000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#196570000000
0!
0'
0/
#196580000000
1!
1'
1/
#196590000000
0!
0'
0/
#196600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#196610000000
0!
0'
0/
#196620000000
1!
1'
1/
#196630000000
0!
1"
0'
1(
0/
10
#196640000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#196650000000
0!
1$
0'
1+
0/
#196660000000
1!
1'
1/
#196670000000
0!
0'
0/
#196680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#196690000000
0!
0'
0/
#196700000000
1!
1'
1/
#196710000000
0!
0'
0/
#196720000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#196730000000
0!
0'
0/
#196740000000
1!
1'
1/
#196750000000
0!
0'
0/
#196760000000
1!
1'
1/
#196770000000
0!
0'
0/
#196780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#196790000000
0!
0'
0/
#196800000000
1!
1'
1/
#196810000000
0!
0'
0/
#196820000000
1!
1'
1/
#196830000000
0!
0'
0/
#196840000000
1!
1'
1/
#196850000000
0!
0'
0/
#196860000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#196870000000
0!
0'
0/
#196880000000
1!
1'
1/
#196890000000
0!
0'
0/
#196900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#196910000000
0!
0'
0/
#196920000000
1!
1'
1/
#196930000000
0!
0'
0/
#196940000000
#196950000000
1!
1'
1/
#196960000000
0!
0'
0/
#196970000000
1!
1'
1/
#196980000000
0!
1"
0'
1(
0/
10
#196990000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#197000000000
0!
0'
0/
#197010000000
1!
1'
1/
#197020000000
0!
0'
0/
#197030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#197040000000
0!
0'
0/
#197050000000
1!
1'
1/
#197060000000
0!
1"
0'
1(
0/
10
#197070000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#197080000000
0!
1$
0'
1+
0/
#197090000000
1!
1'
1/
#197100000000
0!
0'
0/
#197110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#197120000000
0!
0'
0/
#197130000000
1!
1'
1/
#197140000000
0!
0'
0/
#197150000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#197160000000
0!
0'
0/
#197170000000
1!
1'
1/
#197180000000
0!
0'
0/
#197190000000
1!
1'
1/
#197200000000
0!
0'
0/
#197210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#197220000000
0!
0'
0/
#197230000000
1!
1'
1/
#197240000000
0!
0'
0/
#197250000000
1!
1'
1/
#197260000000
0!
0'
0/
#197270000000
1!
1'
1/
#197280000000
0!
0'
0/
#197290000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#197300000000
0!
0'
0/
#197310000000
1!
1'
1/
#197320000000
0!
0'
0/
#197330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#197340000000
0!
0'
0/
#197350000000
1!
1'
1/
#197360000000
0!
0'
0/
#197370000000
#197380000000
1!
1'
1/
#197390000000
0!
0'
0/
#197400000000
1!
1'
1/
#197410000000
0!
1"
0'
1(
0/
10
#197420000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#197430000000
0!
0'
0/
#197440000000
1!
1'
1/
#197450000000
0!
0'
0/
#197460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#197470000000
0!
0'
0/
#197480000000
1!
1'
1/
#197490000000
0!
1"
0'
1(
0/
10
#197500000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#197510000000
0!
1$
0'
1+
0/
#197520000000
1!
1'
1/
#197530000000
0!
0'
0/
#197540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#197550000000
0!
0'
0/
#197560000000
1!
1'
1/
#197570000000
0!
0'
0/
#197580000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#197590000000
0!
0'
0/
#197600000000
1!
1'
1/
#197610000000
0!
0'
0/
#197620000000
1!
1'
1/
#197630000000
0!
0'
0/
#197640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#197650000000
0!
0'
0/
#197660000000
1!
1'
1/
#197670000000
0!
0'
0/
#197680000000
1!
1'
1/
#197690000000
0!
0'
0/
#197700000000
1!
1'
1/
#197710000000
0!
0'
0/
#197720000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#197730000000
0!
0'
0/
#197740000000
1!
1'
1/
#197750000000
0!
0'
0/
#197760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#197770000000
0!
0'
0/
#197780000000
1!
1'
1/
#197790000000
0!
0'
0/
#197800000000
#197810000000
1!
1'
1/
#197820000000
0!
0'
0/
#197830000000
1!
1'
1/
#197840000000
0!
1"
0'
1(
0/
10
#197850000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#197860000000
0!
0'
0/
#197870000000
1!
1'
1/
#197880000000
0!
0'
0/
#197890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#197900000000
0!
0'
0/
#197910000000
1!
1'
1/
#197920000000
0!
1"
0'
1(
0/
10
#197930000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#197940000000
0!
1$
0'
1+
0/
#197950000000
1!
1'
1/
#197960000000
0!
0'
0/
#197970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#197980000000
0!
0'
0/
#197990000000
1!
1'
1/
#198000000000
0!
0'
0/
#198010000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#198020000000
0!
0'
0/
#198030000000
1!
1'
1/
#198040000000
0!
0'
0/
#198050000000
1!
1'
1/
#198060000000
0!
0'
0/
#198070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#198080000000
0!
0'
0/
#198090000000
1!
1'
1/
#198100000000
0!
0'
0/
#198110000000
1!
1'
1/
#198120000000
0!
0'
0/
#198130000000
1!
1'
1/
#198140000000
0!
0'
0/
#198150000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#198160000000
0!
0'
0/
#198170000000
1!
1'
1/
#198180000000
0!
0'
0/
#198190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#198200000000
0!
0'
0/
#198210000000
1!
1'
1/
#198220000000
0!
0'
0/
#198230000000
#198240000000
1!
1'
1/
#198250000000
0!
0'
0/
#198260000000
1!
1'
1/
#198270000000
0!
1"
0'
1(
0/
10
#198280000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#198290000000
0!
0'
0/
#198300000000
1!
1'
1/
#198310000000
0!
0'
0/
#198320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#198330000000
0!
0'
0/
#198340000000
1!
1'
1/
#198350000000
0!
1"
0'
1(
0/
10
#198360000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#198370000000
0!
1$
0'
1+
0/
#198380000000
1!
1'
1/
#198390000000
0!
0'
0/
#198400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#198410000000
0!
0'
0/
#198420000000
1!
1'
1/
#198430000000
0!
0'
0/
#198440000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#198450000000
0!
0'
0/
#198460000000
1!
1'
1/
#198470000000
0!
0'
0/
#198480000000
1!
1'
1/
#198490000000
0!
0'
0/
#198500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#198510000000
0!
0'
0/
#198520000000
1!
1'
1/
#198530000000
0!
0'
0/
#198540000000
1!
1'
1/
#198550000000
0!
0'
0/
#198560000000
1!
1'
1/
#198570000000
0!
0'
0/
#198580000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#198590000000
0!
0'
0/
#198600000000
1!
1'
1/
#198610000000
0!
0'
0/
#198620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#198630000000
0!
0'
0/
#198640000000
1!
1'
1/
#198650000000
0!
0'
0/
#198660000000
#198670000000
1!
1'
1/
#198680000000
0!
0'
0/
#198690000000
1!
1'
1/
#198700000000
0!
1"
0'
1(
0/
10
#198710000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#198720000000
0!
0'
0/
#198730000000
1!
1'
1/
#198740000000
0!
0'
0/
#198750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#198760000000
0!
0'
0/
#198770000000
1!
1'
1/
#198780000000
0!
1"
0'
1(
0/
10
#198790000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#198800000000
0!
1$
0'
1+
0/
#198810000000
1!
1'
1/
#198820000000
0!
0'
0/
#198830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#198840000000
0!
0'
0/
#198850000000
1!
1'
1/
#198860000000
0!
0'
0/
#198870000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#198880000000
0!
0'
0/
#198890000000
1!
1'
1/
#198900000000
0!
0'
0/
#198910000000
1!
1'
1/
#198920000000
0!
0'
0/
#198930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#198940000000
0!
0'
0/
#198950000000
1!
1'
1/
#198960000000
0!
0'
0/
#198970000000
1!
1'
1/
#198980000000
0!
0'
0/
#198990000000
1!
1'
1/
#199000000000
0!
0'
0/
#199010000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#199020000000
0!
0'
0/
#199030000000
1!
1'
1/
#199040000000
0!
0'
0/
#199050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#199060000000
0!
0'
0/
#199070000000
1!
1'
1/
#199080000000
0!
0'
0/
#199090000000
#199100000000
1!
1'
1/
#199110000000
0!
0'
0/
#199120000000
1!
1'
1/
#199130000000
0!
1"
0'
1(
0/
10
#199140000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#199150000000
0!
0'
0/
#199160000000
1!
1'
1/
#199170000000
0!
0'
0/
#199180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#199190000000
0!
0'
0/
#199200000000
1!
1'
1/
#199210000000
0!
1"
0'
1(
0/
10
#199220000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#199230000000
0!
1$
0'
1+
0/
#199240000000
1!
1'
1/
#199250000000
0!
0'
0/
#199260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#199270000000
0!
0'
0/
#199280000000
1!
1'
1/
#199290000000
0!
0'
0/
#199300000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#199310000000
0!
0'
0/
#199320000000
1!
1'
1/
#199330000000
0!
0'
0/
#199340000000
1!
1'
1/
#199350000000
0!
0'
0/
#199360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#199370000000
0!
0'
0/
#199380000000
1!
1'
1/
#199390000000
0!
0'
0/
#199400000000
1!
1'
1/
#199410000000
0!
0'
0/
#199420000000
1!
1'
1/
#199430000000
0!
0'
0/
#199440000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#199450000000
0!
0'
0/
#199460000000
1!
1'
1/
#199470000000
0!
0'
0/
#199480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#199490000000
0!
0'
0/
#199500000000
1!
1'
1/
#199510000000
0!
0'
0/
#199520000000
#199530000000
1!
1'
1/
#199540000000
0!
0'
0/
#199550000000
1!
1'
1/
#199560000000
0!
1"
0'
1(
0/
10
#199570000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#199580000000
0!
0'
0/
#199590000000
1!
1'
1/
#199600000000
0!
0'
0/
#199610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#199620000000
0!
0'
0/
#199630000000
1!
1'
1/
#199640000000
0!
1"
0'
1(
0/
10
#199650000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#199660000000
0!
1$
0'
1+
0/
#199670000000
1!
1'
1/
#199680000000
0!
0'
0/
#199690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#199700000000
0!
0'
0/
#199710000000
1!
1'
1/
#199720000000
0!
0'
0/
#199730000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#199740000000
0!
0'
0/
#199750000000
1!
1'
1/
#199760000000
0!
0'
0/
#199770000000
1!
1'
1/
#199780000000
0!
0'
0/
#199790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#199800000000
0!
0'
0/
#199810000000
1!
1'
1/
#199820000000
0!
0'
0/
#199830000000
1!
1'
1/
#199840000000
0!
0'
0/
#199850000000
1!
1'
1/
#199860000000
0!
0'
0/
#199870000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#199880000000
0!
0'
0/
#199890000000
1!
1'
1/
#199900000000
0!
0'
0/
#199910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#199920000000
0!
0'
0/
#199930000000
1!
1'
1/
#199940000000
0!
0'
0/
#199950000000
#199960000000
1!
1'
1/
#199970000000
0!
0'
0/
#199980000000
1!
1'
1/
#199990000000
0!
1"
0'
1(
0/
10
#200000000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#200010000000
0!
0'
0/
#200020000000
1!
1'
1/
#200030000000
0!
0'
0/
#200040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#200050000000
0!
0'
0/
#200060000000
1!
1'
1/
#200070000000
0!
1"
0'
1(
0/
10
#200080000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#200090000000
0!
1$
0'
1+
0/
#200100000000
1!
1'
1/
#200110000000
0!
0'
0/
#200120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#200130000000
0!
0'
0/
#200140000000
1!
1'
1/
#200150000000
0!
0'
0/
#200160000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#200170000000
0!
0'
0/
#200180000000
1!
1'
1/
#200190000000
0!
0'
0/
#200200000000
1!
1'
1/
#200210000000
0!
0'
0/
#200220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#200230000000
0!
0'
0/
#200240000000
1!
1'
1/
#200250000000
0!
0'
0/
#200260000000
1!
1'
1/
#200270000000
0!
0'
0/
#200280000000
1!
1'
1/
#200290000000
0!
0'
0/
#200300000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#200310000000
0!
0'
0/
#200320000000
1!
1'
1/
#200330000000
0!
0'
0/
#200340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#200350000000
0!
0'
0/
#200360000000
1!
1'
1/
#200370000000
0!
0'
0/
#200380000000
#200390000000
1!
1'
1/
#200400000000
0!
0'
0/
#200410000000
1!
1'
1/
#200420000000
0!
1"
0'
1(
0/
10
#200430000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#200440000000
0!
0'
0/
#200450000000
1!
1'
1/
#200460000000
0!
0'
0/
#200470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#200480000000
0!
0'
0/
#200490000000
1!
1'
1/
#200500000000
0!
1"
0'
1(
0/
10
#200510000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#200520000000
0!
1$
0'
1+
0/
#200530000000
1!
1'
1/
#200540000000
0!
0'
0/
#200550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#200560000000
0!
0'
0/
#200570000000
1!
1'
1/
#200580000000
0!
0'
0/
#200590000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#200600000000
0!
0'
0/
#200610000000
1!
1'
1/
#200620000000
0!
0'
0/
#200630000000
1!
1'
1/
#200640000000
0!
0'
0/
#200650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#200660000000
0!
0'
0/
#200670000000
1!
1'
1/
#200680000000
0!
0'
0/
#200690000000
1!
1'
1/
#200700000000
0!
0'
0/
#200710000000
1!
1'
1/
#200720000000
0!
0'
0/
#200730000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#200740000000
0!
0'
0/
#200750000000
1!
1'
1/
#200760000000
0!
0'
0/
#200770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#200780000000
0!
0'
0/
#200790000000
1!
1'
1/
#200800000000
0!
0'
0/
#200810000000
#200820000000
1!
1'
1/
#200830000000
0!
0'
0/
#200840000000
1!
1'
1/
#200850000000
0!
1"
0'
1(
0/
10
#200860000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#200870000000
0!
0'
0/
#200880000000
1!
1'
1/
#200890000000
0!
0'
0/
#200900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#200910000000
0!
0'
0/
#200920000000
1!
1'
1/
#200930000000
0!
1"
0'
1(
0/
10
#200940000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#200950000000
0!
1$
0'
1+
0/
#200960000000
1!
1'
1/
#200970000000
0!
0'
0/
#200980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#200990000000
0!
0'
0/
#201000000000
1!
1'
1/
#201010000000
0!
0'
0/
#201020000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#201030000000
0!
0'
0/
#201040000000
1!
1'
1/
#201050000000
0!
0'
0/
#201060000000
1!
1'
1/
#201070000000
0!
0'
0/
#201080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#201090000000
0!
0'
0/
#201100000000
1!
1'
1/
#201110000000
0!
0'
0/
#201120000000
1!
1'
1/
#201130000000
0!
0'
0/
#201140000000
1!
1'
1/
#201150000000
0!
0'
0/
#201160000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#201170000000
0!
0'
0/
#201180000000
1!
1'
1/
#201190000000
0!
0'
0/
#201200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#201210000000
0!
0'
0/
#201220000000
1!
1'
1/
#201230000000
0!
0'
0/
#201240000000
#201250000000
1!
1'
1/
#201260000000
0!
0'
0/
#201270000000
1!
1'
1/
#201280000000
0!
1"
0'
1(
0/
10
#201290000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#201300000000
0!
0'
0/
#201310000000
1!
1'
1/
#201320000000
0!
0'
0/
#201330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#201340000000
0!
0'
0/
#201350000000
1!
1'
1/
#201360000000
0!
1"
0'
1(
0/
10
#201370000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#201380000000
0!
1$
0'
1+
0/
#201390000000
1!
1'
1/
#201400000000
0!
0'
0/
#201410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#201420000000
0!
0'
0/
#201430000000
1!
1'
1/
#201440000000
0!
0'
0/
#201450000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#201460000000
0!
0'
0/
#201470000000
1!
1'
1/
#201480000000
0!
0'
0/
#201490000000
1!
1'
1/
#201500000000
0!
0'
0/
#201510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#201520000000
0!
0'
0/
#201530000000
1!
1'
1/
#201540000000
0!
0'
0/
#201550000000
1!
1'
1/
#201560000000
0!
0'
0/
#201570000000
1!
1'
1/
#201580000000
0!
0'
0/
#201590000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#201600000000
0!
0'
0/
#201610000000
1!
1'
1/
#201620000000
0!
0'
0/
#201630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#201640000000
0!
0'
0/
#201650000000
1!
1'
1/
#201660000000
0!
0'
0/
#201670000000
#201680000000
1!
1'
1/
#201690000000
0!
0'
0/
#201700000000
1!
1'
1/
#201710000000
0!
1"
0'
1(
0/
10
#201720000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#201730000000
0!
0'
0/
#201740000000
1!
1'
1/
#201750000000
0!
0'
0/
#201760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#201770000000
0!
0'
0/
#201780000000
1!
1'
1/
#201790000000
0!
1"
0'
1(
0/
10
#201800000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#201810000000
0!
1$
0'
1+
0/
#201820000000
1!
1'
1/
#201830000000
0!
0'
0/
#201840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#201850000000
0!
0'
0/
#201860000000
1!
1'
1/
#201870000000
0!
0'
0/
#201880000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#201890000000
0!
0'
0/
#201900000000
1!
1'
1/
#201910000000
0!
0'
0/
#201920000000
1!
1'
1/
#201930000000
0!
0'
0/
#201940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#201950000000
0!
0'
0/
#201960000000
1!
1'
1/
#201970000000
0!
0'
0/
#201980000000
1!
1'
1/
#201990000000
0!
0'
0/
#202000000000
1!
1'
1/
#202010000000
0!
0'
0/
#202020000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#202030000000
0!
0'
0/
#202040000000
1!
1'
1/
#202050000000
0!
0'
0/
#202060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#202070000000
0!
0'
0/
#202080000000
1!
1'
1/
#202090000000
0!
0'
0/
#202100000000
#202110000000
1!
1'
1/
#202120000000
0!
0'
0/
#202130000000
1!
1'
1/
#202140000000
0!
1"
0'
1(
0/
10
#202150000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#202160000000
0!
0'
0/
#202170000000
1!
1'
1/
#202180000000
0!
0'
0/
#202190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#202200000000
0!
0'
0/
#202210000000
1!
1'
1/
#202220000000
0!
1"
0'
1(
0/
10
#202230000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#202240000000
0!
1$
0'
1+
0/
#202250000000
1!
1'
1/
#202260000000
0!
0'
0/
#202270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#202280000000
0!
0'
0/
#202290000000
1!
1'
1/
#202300000000
0!
0'
0/
#202310000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#202320000000
0!
0'
0/
#202330000000
1!
1'
1/
#202340000000
0!
0'
0/
#202350000000
1!
1'
1/
#202360000000
0!
0'
0/
#202370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#202380000000
0!
0'
0/
#202390000000
1!
1'
1/
#202400000000
0!
0'
0/
#202410000000
1!
1'
1/
#202420000000
0!
0'
0/
#202430000000
1!
1'
1/
#202440000000
0!
0'
0/
#202450000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#202460000000
0!
0'
0/
#202470000000
1!
1'
1/
#202480000000
0!
0'
0/
#202490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#202500000000
0!
0'
0/
#202510000000
1!
1'
1/
#202520000000
0!
0'
0/
#202530000000
#202540000000
1!
1'
1/
#202550000000
0!
0'
0/
#202560000000
1!
1'
1/
#202570000000
0!
1"
0'
1(
0/
10
#202580000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#202590000000
0!
0'
0/
#202600000000
1!
1'
1/
#202610000000
0!
0'
0/
#202620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#202630000000
0!
0'
0/
#202640000000
1!
1'
1/
#202650000000
0!
1"
0'
1(
0/
10
#202660000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#202670000000
0!
1$
0'
1+
0/
#202680000000
1!
1'
1/
#202690000000
0!
0'
0/
#202700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#202710000000
0!
0'
0/
#202720000000
1!
1'
1/
#202730000000
0!
0'
0/
#202740000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#202750000000
0!
0'
0/
#202760000000
1!
1'
1/
#202770000000
0!
0'
0/
#202780000000
1!
1'
1/
#202790000000
0!
0'
0/
#202800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#202810000000
0!
0'
0/
#202820000000
1!
1'
1/
#202830000000
0!
0'
0/
#202840000000
1!
1'
1/
#202850000000
0!
0'
0/
#202860000000
1!
1'
1/
#202870000000
0!
0'
0/
#202880000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#202890000000
0!
0'
0/
#202900000000
1!
1'
1/
#202910000000
0!
0'
0/
#202920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#202930000000
0!
0'
0/
#202940000000
1!
1'
1/
#202950000000
0!
0'
0/
#202960000000
#202970000000
1!
1'
1/
#202980000000
0!
0'
0/
#202990000000
1!
1'
1/
#203000000000
0!
1"
0'
1(
0/
10
#203010000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#203020000000
0!
0'
0/
#203030000000
1!
1'
1/
#203040000000
0!
0'
0/
#203050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#203060000000
0!
0'
0/
#203070000000
1!
1'
1/
#203080000000
0!
1"
0'
1(
0/
10
#203090000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#203100000000
0!
1$
0'
1+
0/
#203110000000
1!
1'
1/
#203120000000
0!
0'
0/
#203130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#203140000000
0!
0'
0/
#203150000000
1!
1'
1/
#203160000000
0!
0'
0/
#203170000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#203180000000
0!
0'
0/
#203190000000
1!
1'
1/
#203200000000
0!
0'
0/
#203210000000
1!
1'
1/
#203220000000
0!
0'
0/
#203230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#203240000000
0!
0'
0/
#203250000000
1!
1'
1/
#203260000000
0!
0'
0/
#203270000000
1!
1'
1/
#203280000000
0!
0'
0/
#203290000000
1!
1'
1/
#203300000000
0!
0'
0/
#203310000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#203320000000
0!
0'
0/
#203330000000
1!
1'
1/
#203340000000
0!
0'
0/
#203350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#203360000000
0!
0'
0/
#203370000000
1!
1'
1/
#203380000000
0!
0'
0/
#203390000000
#203400000000
1!
1'
1/
#203410000000
0!
0'
0/
#203420000000
1!
1'
1/
#203430000000
0!
1"
0'
1(
0/
10
#203440000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#203450000000
0!
0'
0/
#203460000000
1!
1'
1/
#203470000000
0!
0'
0/
#203480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#203490000000
0!
0'
0/
#203500000000
1!
1'
1/
#203510000000
0!
1"
0'
1(
0/
10
#203520000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#203530000000
0!
1$
0'
1+
0/
#203540000000
1!
1'
1/
#203550000000
0!
0'
0/
#203560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#203570000000
0!
0'
0/
#203580000000
1!
1'
1/
#203590000000
0!
0'
0/
#203600000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#203610000000
0!
0'
0/
#203620000000
1!
1'
1/
#203630000000
0!
0'
0/
#203640000000
1!
1'
1/
#203650000000
0!
0'
0/
#203660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#203670000000
0!
0'
0/
#203680000000
1!
1'
1/
#203690000000
0!
0'
0/
#203700000000
1!
1'
1/
#203710000000
0!
0'
0/
#203720000000
1!
1'
1/
#203730000000
0!
0'
0/
#203740000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#203750000000
0!
0'
0/
#203760000000
1!
1'
1/
#203770000000
0!
0'
0/
#203780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#203790000000
0!
0'
0/
#203800000000
1!
1'
1/
#203810000000
0!
0'
0/
#203820000000
#203830000000
1!
1'
1/
#203840000000
0!
0'
0/
#203850000000
1!
1'
1/
#203860000000
0!
1"
0'
1(
0/
10
#203870000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#203880000000
0!
0'
0/
#203890000000
1!
1'
1/
#203900000000
0!
0'
0/
#203910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#203920000000
0!
0'
0/
#203930000000
1!
1'
1/
#203940000000
0!
1"
0'
1(
0/
10
#203950000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#203960000000
0!
1$
0'
1+
0/
#203970000000
1!
1'
1/
#203980000000
0!
0'
0/
#203990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#204000000000
0!
0'
0/
#204010000000
1!
1'
1/
#204020000000
0!
0'
0/
#204030000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#204040000000
0!
0'
0/
#204050000000
1!
1'
1/
#204060000000
0!
0'
0/
#204070000000
1!
1'
1/
#204080000000
0!
0'
0/
#204090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#204100000000
0!
0'
0/
#204110000000
1!
1'
1/
#204120000000
0!
0'
0/
#204130000000
1!
1'
1/
#204140000000
0!
0'
0/
#204150000000
1!
1'
1/
#204160000000
0!
0'
0/
#204170000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#204180000000
0!
0'
0/
#204190000000
1!
1'
1/
#204200000000
0!
0'
0/
#204210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#204220000000
0!
0'
0/
#204230000000
1!
1'
1/
#204240000000
0!
0'
0/
#204250000000
#204260000000
1!
1'
1/
#204270000000
0!
0'
0/
#204280000000
1!
1'
1/
#204290000000
0!
1"
0'
1(
0/
10
#204300000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#204310000000
0!
0'
0/
#204320000000
1!
1'
1/
#204330000000
0!
0'
0/
#204340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#204350000000
0!
0'
0/
#204360000000
1!
1'
1/
#204370000000
0!
1"
0'
1(
0/
10
#204380000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#204390000000
0!
1$
0'
1+
0/
#204400000000
1!
1'
1/
#204410000000
0!
0'
0/
#204420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#204430000000
0!
0'
0/
#204440000000
1!
1'
1/
#204450000000
0!
0'
0/
#204460000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#204470000000
0!
0'
0/
#204480000000
1!
1'
1/
#204490000000
0!
0'
0/
#204500000000
1!
1'
1/
#204510000000
0!
0'
0/
#204520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#204530000000
0!
0'
0/
#204540000000
1!
1'
1/
#204550000000
0!
0'
0/
#204560000000
1!
1'
1/
#204570000000
0!
0'
0/
#204580000000
1!
1'
1/
#204590000000
0!
0'
0/
#204600000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#204610000000
0!
0'
0/
#204620000000
1!
1'
1/
#204630000000
0!
0'
0/
#204640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#204650000000
0!
0'
0/
#204660000000
1!
1'
1/
#204670000000
0!
0'
0/
#204680000000
#204690000000
1!
1'
1/
#204700000000
0!
0'
0/
#204710000000
1!
1'
1/
#204720000000
0!
1"
0'
1(
0/
10
#204730000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#204740000000
0!
0'
0/
#204750000000
1!
1'
1/
#204760000000
0!
0'
0/
#204770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#204780000000
0!
0'
0/
#204790000000
1!
1'
1/
#204800000000
0!
1"
0'
1(
0/
10
#204810000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#204820000000
0!
1$
0'
1+
0/
#204830000000
1!
1'
1/
#204840000000
0!
0'
0/
#204850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#204860000000
0!
0'
0/
#204870000000
1!
1'
1/
#204880000000
0!
0'
0/
#204890000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#204900000000
0!
0'
0/
#204910000000
1!
1'
1/
#204920000000
0!
0'
0/
#204930000000
1!
1'
1/
#204940000000
0!
0'
0/
#204950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#204960000000
0!
0'
0/
#204970000000
1!
1'
1/
#204980000000
0!
0'
0/
#204990000000
1!
1'
1/
#205000000000
0!
0'
0/
#205010000000
1!
1'
1/
#205020000000
0!
0'
0/
#205030000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#205040000000
0!
0'
0/
#205050000000
1!
1'
1/
#205060000000
0!
0'
0/
#205070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#205080000000
0!
0'
0/
#205090000000
1!
1'
1/
#205100000000
0!
0'
0/
#205110000000
#205120000000
1!
1'
1/
#205130000000
0!
0'
0/
#205140000000
1!
1'
1/
#205150000000
0!
1"
0'
1(
0/
10
#205160000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#205170000000
0!
0'
0/
#205180000000
1!
1'
1/
#205190000000
0!
0'
0/
#205200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#205210000000
0!
0'
0/
#205220000000
1!
1'
1/
#205230000000
0!
1"
0'
1(
0/
10
#205240000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#205250000000
0!
1$
0'
1+
0/
#205260000000
1!
1'
1/
#205270000000
0!
0'
0/
#205280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#205290000000
0!
0'
0/
#205300000000
1!
1'
1/
#205310000000
0!
0'
0/
#205320000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#205330000000
0!
0'
0/
#205340000000
1!
1'
1/
#205350000000
0!
0'
0/
#205360000000
1!
1'
1/
#205370000000
0!
0'
0/
#205380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#205390000000
0!
0'
0/
#205400000000
1!
1'
1/
#205410000000
0!
0'
0/
#205420000000
1!
1'
1/
#205430000000
0!
0'
0/
#205440000000
1!
1'
1/
#205450000000
0!
0'
0/
#205460000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#205470000000
0!
0'
0/
#205480000000
1!
1'
1/
#205490000000
0!
0'
0/
#205500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#205510000000
0!
0'
0/
#205520000000
1!
1'
1/
#205530000000
0!
0'
0/
#205540000000
#205550000000
1!
1'
1/
#205560000000
0!
0'
0/
#205570000000
1!
1'
1/
#205580000000
0!
1"
0'
1(
0/
10
#205590000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#205600000000
0!
0'
0/
#205610000000
1!
1'
1/
#205620000000
0!
0'
0/
#205630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#205640000000
0!
0'
0/
#205650000000
1!
1'
1/
#205660000000
0!
1"
0'
1(
0/
10
#205670000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#205680000000
0!
1$
0'
1+
0/
#205690000000
1!
1'
1/
#205700000000
0!
0'
0/
#205710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#205720000000
0!
0'
0/
#205730000000
1!
1'
1/
#205740000000
0!
0'
0/
#205750000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#205760000000
0!
0'
0/
#205770000000
1!
1'
1/
#205780000000
0!
0'
0/
#205790000000
1!
1'
1/
#205800000000
0!
0'
0/
#205810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#205820000000
0!
0'
0/
#205830000000
1!
1'
1/
#205840000000
0!
0'
0/
#205850000000
1!
1'
1/
#205860000000
0!
0'
0/
#205870000000
1!
1'
1/
#205880000000
0!
0'
0/
#205890000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#205900000000
0!
0'
0/
#205910000000
1!
1'
1/
#205920000000
0!
0'
0/
#205930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#205940000000
0!
0'
0/
#205950000000
1!
1'
1/
#205960000000
0!
0'
0/
#205970000000
#205980000000
1!
1'
1/
#205990000000
0!
0'
0/
#206000000000
1!
1'
1/
#206010000000
0!
1"
0'
1(
0/
10
#206020000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#206030000000
0!
0'
0/
#206040000000
1!
1'
1/
#206050000000
0!
0'
0/
#206060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#206070000000
0!
0'
0/
#206080000000
1!
1'
1/
#206090000000
0!
1"
0'
1(
0/
10
#206100000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#206110000000
0!
1$
0'
1+
0/
#206120000000
1!
1'
1/
#206130000000
0!
0'
0/
#206140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#206150000000
0!
0'
0/
#206160000000
1!
1'
1/
#206170000000
0!
0'
0/
#206180000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#206190000000
0!
0'
0/
#206200000000
1!
1'
1/
#206210000000
0!
0'
0/
#206220000000
1!
1'
1/
#206230000000
0!
0'
0/
#206240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#206250000000
0!
0'
0/
#206260000000
1!
1'
1/
#206270000000
0!
0'
0/
#206280000000
1!
1'
1/
#206290000000
0!
0'
0/
#206300000000
1!
1'
1/
#206310000000
0!
0'
0/
#206320000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#206330000000
0!
0'
0/
#206340000000
1!
1'
1/
#206350000000
0!
0'
0/
#206360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#206370000000
0!
0'
0/
#206380000000
1!
1'
1/
#206390000000
0!
0'
0/
#206400000000
#206410000000
1!
1'
1/
#206420000000
0!
0'
0/
#206430000000
1!
1'
1/
#206440000000
0!
1"
0'
1(
0/
10
#206450000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#206460000000
0!
0'
0/
#206470000000
1!
1'
1/
#206480000000
0!
0'
0/
#206490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#206500000000
0!
0'
0/
#206510000000
1!
1'
1/
#206520000000
0!
1"
0'
1(
0/
10
#206530000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#206540000000
0!
1$
0'
1+
0/
#206550000000
1!
1'
1/
#206560000000
0!
0'
0/
#206570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#206580000000
0!
0'
0/
#206590000000
1!
1'
1/
#206600000000
0!
0'
0/
#206610000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#206620000000
0!
0'
0/
#206630000000
1!
1'
1/
#206640000000
0!
0'
0/
#206650000000
1!
1'
1/
#206660000000
0!
0'
0/
#206670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#206680000000
0!
0'
0/
#206690000000
1!
1'
1/
#206700000000
0!
0'
0/
#206710000000
1!
1'
1/
#206720000000
0!
0'
0/
#206730000000
1!
1'
1/
#206740000000
0!
0'
0/
#206750000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#206760000000
0!
0'
0/
#206770000000
1!
1'
1/
#206780000000
0!
0'
0/
#206790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#206800000000
0!
0'
0/
#206810000000
1!
1'
1/
#206820000000
0!
0'
0/
#206830000000
#206840000000
1!
1'
1/
#206850000000
0!
0'
0/
#206860000000
1!
1'
1/
#206870000000
0!
1"
0'
1(
0/
10
#206880000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#206890000000
0!
0'
0/
#206900000000
1!
1'
1/
#206910000000
0!
0'
0/
#206920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#206930000000
0!
0'
0/
#206940000000
1!
1'
1/
#206950000000
0!
1"
0'
1(
0/
10
#206960000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#206970000000
0!
1$
0'
1+
0/
#206980000000
1!
1'
1/
#206990000000
0!
0'
0/
#207000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#207010000000
0!
0'
0/
#207020000000
1!
1'
1/
#207030000000
0!
0'
0/
#207040000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#207050000000
0!
0'
0/
#207060000000
1!
1'
1/
#207070000000
0!
0'
0/
#207080000000
1!
1'
1/
#207090000000
0!
0'
0/
#207100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#207110000000
0!
0'
0/
#207120000000
1!
1'
1/
#207130000000
0!
0'
0/
#207140000000
1!
1'
1/
#207150000000
0!
0'
0/
#207160000000
1!
1'
1/
#207170000000
0!
0'
0/
#207180000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#207190000000
0!
0'
0/
#207200000000
1!
1'
1/
#207210000000
0!
0'
0/
#207220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#207230000000
0!
0'
0/
#207240000000
1!
1'
1/
#207250000000
0!
0'
0/
#207260000000
#207270000000
1!
1'
1/
#207280000000
0!
0'
0/
#207290000000
1!
1'
1/
#207300000000
0!
1"
0'
1(
0/
10
#207310000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#207320000000
0!
0'
0/
#207330000000
1!
1'
1/
#207340000000
0!
0'
0/
#207350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#207360000000
0!
0'
0/
#207370000000
1!
1'
1/
#207380000000
0!
1"
0'
1(
0/
10
#207390000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#207400000000
0!
1$
0'
1+
0/
#207410000000
1!
1'
1/
#207420000000
0!
0'
0/
#207430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#207440000000
0!
0'
0/
#207450000000
1!
1'
1/
#207460000000
0!
0'
0/
#207470000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#207480000000
0!
0'
0/
#207490000000
1!
1'
1/
#207500000000
0!
0'
0/
#207510000000
1!
1'
1/
#207520000000
0!
0'
0/
#207530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#207540000000
0!
0'
0/
#207550000000
1!
1'
1/
#207560000000
0!
0'
0/
#207570000000
1!
1'
1/
#207580000000
0!
0'
0/
#207590000000
1!
1'
1/
#207600000000
0!
0'
0/
#207610000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#207620000000
0!
0'
0/
#207630000000
1!
1'
1/
#207640000000
0!
0'
0/
#207650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#207660000000
0!
0'
0/
#207670000000
1!
1'
1/
#207680000000
0!
0'
0/
#207690000000
#207700000000
1!
1'
1/
#207710000000
0!
0'
0/
#207720000000
1!
1'
1/
#207730000000
0!
1"
0'
1(
0/
10
#207740000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#207750000000
0!
0'
0/
#207760000000
1!
1'
1/
#207770000000
0!
0'
0/
#207780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#207790000000
0!
0'
0/
#207800000000
1!
1'
1/
#207810000000
0!
1"
0'
1(
0/
10
#207820000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#207830000000
0!
1$
0'
1+
0/
#207840000000
1!
1'
1/
#207850000000
0!
0'
0/
#207860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#207870000000
0!
0'
0/
#207880000000
1!
1'
1/
#207890000000
0!
0'
0/
#207900000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#207910000000
0!
0'
0/
#207920000000
1!
1'
1/
#207930000000
0!
0'
0/
#207940000000
1!
1'
1/
#207950000000
0!
0'
0/
#207960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#207970000000
0!
0'
0/
#207980000000
1!
1'
1/
#207990000000
0!
0'
0/
#208000000000
1!
1'
1/
#208010000000
0!
0'
0/
#208020000000
1!
1'
1/
#208030000000
0!
0'
0/
#208040000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#208050000000
0!
0'
0/
#208060000000
1!
1'
1/
#208070000000
0!
0'
0/
#208080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#208090000000
0!
0'
0/
#208100000000
1!
1'
1/
#208110000000
0!
0'
0/
#208120000000
#208130000000
1!
1'
1/
#208140000000
0!
0'
0/
#208150000000
1!
1'
1/
#208160000000
0!
1"
0'
1(
0/
10
#208170000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#208180000000
0!
0'
0/
#208190000000
1!
1'
1/
#208200000000
0!
0'
0/
#208210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#208220000000
0!
0'
0/
#208230000000
1!
1'
1/
#208240000000
0!
1"
0'
1(
0/
10
#208250000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#208260000000
0!
1$
0'
1+
0/
#208270000000
1!
1'
1/
#208280000000
0!
0'
0/
#208290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#208300000000
0!
0'
0/
#208310000000
1!
1'
1/
#208320000000
0!
0'
0/
#208330000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#208340000000
0!
0'
0/
#208350000000
1!
1'
1/
#208360000000
0!
0'
0/
#208370000000
1!
1'
1/
#208380000000
0!
0'
0/
#208390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#208400000000
0!
0'
0/
#208410000000
1!
1'
1/
#208420000000
0!
0'
0/
#208430000000
1!
1'
1/
#208440000000
0!
0'
0/
#208450000000
1!
1'
1/
#208460000000
0!
0'
0/
#208470000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#208480000000
0!
0'
0/
#208490000000
1!
1'
1/
#208500000000
0!
0'
0/
#208510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#208520000000
0!
0'
0/
#208530000000
1!
1'
1/
#208540000000
0!
0'
0/
#208550000000
#208560000000
1!
1'
1/
#208570000000
0!
0'
0/
#208580000000
1!
1'
1/
#208590000000
0!
1"
0'
1(
0/
10
#208600000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#208610000000
0!
0'
0/
#208620000000
1!
1'
1/
#208630000000
0!
0'
0/
#208640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#208650000000
0!
0'
0/
#208660000000
1!
1'
1/
#208670000000
0!
1"
0'
1(
0/
10
#208680000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#208690000000
0!
1$
0'
1+
0/
#208700000000
1!
1'
1/
#208710000000
0!
0'
0/
#208720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#208730000000
0!
0'
0/
#208740000000
1!
1'
1/
#208750000000
0!
0'
0/
#208760000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#208770000000
0!
0'
0/
#208780000000
1!
1'
1/
#208790000000
0!
0'
0/
#208800000000
1!
1'
1/
#208810000000
0!
0'
0/
#208820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#208830000000
0!
0'
0/
#208840000000
1!
1'
1/
#208850000000
0!
0'
0/
#208860000000
1!
1'
1/
#208870000000
0!
0'
0/
#208880000000
1!
1'
1/
#208890000000
0!
0'
0/
#208900000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#208910000000
0!
0'
0/
#208920000000
1!
1'
1/
#208930000000
0!
0'
0/
#208940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#208950000000
0!
0'
0/
#208960000000
1!
1'
1/
#208970000000
0!
0'
0/
#208980000000
#208990000000
1!
1'
1/
#209000000000
0!
0'
0/
#209010000000
1!
1'
1/
#209020000000
0!
1"
0'
1(
0/
10
#209030000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#209040000000
0!
0'
0/
#209050000000
1!
1'
1/
#209060000000
0!
0'
0/
#209070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#209080000000
0!
0'
0/
#209090000000
1!
1'
1/
#209100000000
0!
1"
0'
1(
0/
10
#209110000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#209120000000
0!
1$
0'
1+
0/
#209130000000
1!
1'
1/
#209140000000
0!
0'
0/
#209150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#209160000000
0!
0'
0/
#209170000000
1!
1'
1/
#209180000000
0!
0'
0/
#209190000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#209200000000
0!
0'
0/
#209210000000
1!
1'
1/
#209220000000
0!
0'
0/
#209230000000
1!
1'
1/
#209240000000
0!
0'
0/
#209250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#209260000000
0!
0'
0/
#209270000000
1!
1'
1/
#209280000000
0!
0'
0/
#209290000000
1!
1'
1/
#209300000000
0!
0'
0/
#209310000000
1!
1'
1/
#209320000000
0!
0'
0/
#209330000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#209340000000
0!
0'
0/
#209350000000
1!
1'
1/
#209360000000
0!
0'
0/
#209370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#209380000000
0!
0'
0/
#209390000000
1!
1'
1/
#209400000000
0!
0'
0/
#209410000000
#209420000000
1!
1'
1/
#209430000000
0!
0'
0/
#209440000000
1!
1'
1/
#209450000000
0!
1"
0'
1(
0/
10
#209460000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#209470000000
0!
0'
0/
#209480000000
1!
1'
1/
#209490000000
0!
0'
0/
#209500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#209510000000
0!
0'
0/
#209520000000
1!
1'
1/
#209530000000
0!
1"
0'
1(
0/
10
#209540000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#209550000000
0!
1$
0'
1+
0/
#209560000000
1!
1'
1/
#209570000000
0!
0'
0/
#209580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#209590000000
0!
0'
0/
#209600000000
1!
1'
1/
#209610000000
0!
0'
0/
#209620000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#209630000000
0!
0'
0/
#209640000000
1!
1'
1/
#209650000000
0!
0'
0/
#209660000000
1!
1'
1/
#209670000000
0!
0'
0/
#209680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#209690000000
0!
0'
0/
#209700000000
1!
1'
1/
#209710000000
0!
0'
0/
#209720000000
1!
1'
1/
#209730000000
0!
0'
0/
#209740000000
1!
1'
1/
#209750000000
0!
0'
0/
#209760000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#209770000000
0!
0'
0/
#209780000000
1!
1'
1/
#209790000000
0!
0'
0/
#209800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#209810000000
0!
0'
0/
#209820000000
1!
1'
1/
#209830000000
0!
0'
0/
#209840000000
#209850000000
1!
1'
1/
#209860000000
0!
0'
0/
#209870000000
1!
1'
1/
#209880000000
0!
1"
0'
1(
0/
10
#209890000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#209900000000
0!
0'
0/
#209910000000
1!
1'
1/
#209920000000
0!
0'
0/
#209930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#209940000000
0!
0'
0/
#209950000000
1!
1'
1/
#209960000000
0!
1"
0'
1(
0/
10
#209970000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#209980000000
0!
1$
0'
1+
0/
#209990000000
1!
1'
1/
#210000000000
0!
0'
0/
#210010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#210020000000
0!
0'
0/
#210030000000
1!
1'
1/
#210040000000
0!
0'
0/
#210050000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#210060000000
0!
0'
0/
#210070000000
1!
1'
1/
#210080000000
0!
0'
0/
#210090000000
1!
1'
1/
#210100000000
0!
0'
0/
#210110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#210120000000
0!
0'
0/
#210130000000
1!
1'
1/
#210140000000
0!
0'
0/
#210150000000
1!
1'
1/
#210160000000
0!
0'
0/
#210170000000
1!
1'
1/
#210180000000
0!
0'
0/
#210190000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#210200000000
0!
0'
0/
#210210000000
1!
1'
1/
#210220000000
0!
0'
0/
#210230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#210240000000
0!
0'
0/
#210250000000
1!
1'
1/
#210260000000
0!
0'
0/
#210270000000
#210280000000
1!
1'
1/
#210290000000
0!
0'
0/
#210300000000
1!
1'
1/
#210310000000
0!
1"
0'
1(
0/
10
#210320000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#210330000000
0!
0'
0/
#210340000000
1!
1'
1/
#210350000000
0!
0'
0/
#210360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#210370000000
0!
0'
0/
#210380000000
1!
1'
1/
#210390000000
0!
1"
0'
1(
0/
10
#210400000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#210410000000
0!
1$
0'
1+
0/
#210420000000
1!
1'
1/
#210430000000
0!
0'
0/
#210440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#210450000000
0!
0'
0/
#210460000000
1!
1'
1/
#210470000000
0!
0'
0/
#210480000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#210490000000
0!
0'
0/
#210500000000
1!
1'
1/
#210510000000
0!
0'
0/
#210520000000
1!
1'
1/
#210530000000
0!
0'
0/
#210540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#210550000000
0!
0'
0/
#210560000000
1!
1'
1/
#210570000000
0!
0'
0/
#210580000000
1!
1'
1/
#210590000000
0!
0'
0/
#210600000000
1!
1'
1/
#210610000000
0!
0'
0/
#210620000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#210630000000
0!
0'
0/
#210640000000
1!
1'
1/
#210650000000
0!
0'
0/
#210660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#210670000000
0!
0'
0/
#210680000000
1!
1'
1/
#210690000000
0!
0'
0/
#210700000000
#210710000000
1!
1'
1/
#210720000000
0!
0'
0/
#210730000000
1!
1'
1/
#210740000000
0!
1"
0'
1(
0/
10
#210750000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#210760000000
0!
0'
0/
#210770000000
1!
1'
1/
#210780000000
0!
0'
0/
#210790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#210800000000
0!
0'
0/
#210810000000
1!
1'
1/
#210820000000
0!
1"
0'
1(
0/
10
#210830000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#210840000000
0!
1$
0'
1+
0/
#210850000000
1!
1'
1/
#210860000000
0!
0'
0/
#210870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#210880000000
0!
0'
0/
#210890000000
1!
1'
1/
#210900000000
0!
0'
0/
#210910000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#210920000000
0!
0'
0/
#210930000000
1!
1'
1/
#210940000000
0!
0'
0/
#210950000000
1!
1'
1/
#210960000000
0!
0'
0/
#210970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#210980000000
0!
0'
0/
#210990000000
1!
1'
1/
#211000000000
0!
0'
0/
#211010000000
1!
1'
1/
#211020000000
0!
0'
0/
#211030000000
1!
1'
1/
#211040000000
0!
0'
0/
#211050000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#211060000000
0!
0'
0/
#211070000000
1!
1'
1/
#211080000000
0!
0'
0/
#211090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#211100000000
0!
0'
0/
#211110000000
1!
1'
1/
#211120000000
0!
0'
0/
#211130000000
#211140000000
1!
1'
1/
#211150000000
0!
0'
0/
#211160000000
1!
1'
1/
#211170000000
0!
1"
0'
1(
0/
10
#211180000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#211190000000
0!
0'
0/
#211200000000
1!
1'
1/
#211210000000
0!
0'
0/
#211220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#211230000000
0!
0'
0/
#211240000000
1!
1'
1/
#211250000000
0!
1"
0'
1(
0/
10
#211260000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#211270000000
0!
1$
0'
1+
0/
#211280000000
1!
1'
1/
#211290000000
0!
0'
0/
#211300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#211310000000
0!
0'
0/
#211320000000
1!
1'
1/
#211330000000
0!
0'
0/
#211340000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#211350000000
0!
0'
0/
#211360000000
1!
1'
1/
#211370000000
0!
0'
0/
#211380000000
1!
1'
1/
#211390000000
0!
0'
0/
#211400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#211410000000
0!
0'
0/
#211420000000
1!
1'
1/
#211430000000
0!
0'
0/
#211440000000
1!
1'
1/
#211450000000
0!
0'
0/
#211460000000
1!
1'
1/
#211470000000
0!
0'
0/
#211480000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#211490000000
0!
0'
0/
#211500000000
1!
1'
1/
#211510000000
0!
0'
0/
#211520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#211530000000
0!
0'
0/
#211540000000
1!
1'
1/
#211550000000
0!
0'
0/
#211560000000
#211570000000
1!
1'
1/
#211580000000
0!
0'
0/
#211590000000
1!
1'
1/
#211600000000
0!
1"
0'
1(
0/
10
#211610000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#211620000000
0!
0'
0/
#211630000000
1!
1'
1/
#211640000000
0!
0'
0/
#211650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#211660000000
0!
0'
0/
#211670000000
1!
1'
1/
#211680000000
0!
1"
0'
1(
0/
10
#211690000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#211700000000
0!
1$
0'
1+
0/
#211710000000
1!
1'
1/
#211720000000
0!
0'
0/
#211730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#211740000000
0!
0'
0/
#211750000000
1!
1'
1/
#211760000000
0!
0'
0/
#211770000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#211780000000
0!
0'
0/
#211790000000
1!
1'
1/
#211800000000
0!
0'
0/
#211810000000
1!
1'
1/
#211820000000
0!
0'
0/
#211830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#211840000000
0!
0'
0/
#211850000000
1!
1'
1/
#211860000000
0!
0'
0/
#211870000000
1!
1'
1/
#211880000000
0!
0'
0/
#211890000000
1!
1'
1/
#211900000000
0!
0'
0/
#211910000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#211920000000
0!
0'
0/
#211930000000
1!
1'
1/
#211940000000
0!
0'
0/
#211950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#211960000000
0!
0'
0/
#211970000000
1!
1'
1/
#211980000000
0!
0'
0/
#211990000000
#212000000000
1!
1'
1/
#212010000000
0!
0'
0/
#212020000000
1!
1'
1/
#212030000000
0!
1"
0'
1(
0/
10
#212040000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#212050000000
0!
0'
0/
#212060000000
1!
1'
1/
#212070000000
0!
0'
0/
#212080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#212090000000
0!
0'
0/
#212100000000
1!
1'
1/
#212110000000
0!
1"
0'
1(
0/
10
#212120000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#212130000000
0!
1$
0'
1+
0/
#212140000000
1!
1'
1/
#212150000000
0!
0'
0/
#212160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#212170000000
0!
0'
0/
#212180000000
1!
1'
1/
#212190000000
0!
0'
0/
#212200000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#212210000000
0!
0'
0/
#212220000000
1!
1'
1/
#212230000000
0!
0'
0/
#212240000000
1!
1'
1/
#212250000000
0!
0'
0/
#212260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#212270000000
0!
0'
0/
#212280000000
1!
1'
1/
#212290000000
0!
0'
0/
#212300000000
1!
1'
1/
#212310000000
0!
0'
0/
#212320000000
1!
1'
1/
#212330000000
0!
0'
0/
#212340000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#212350000000
0!
0'
0/
#212360000000
1!
1'
1/
#212370000000
0!
0'
0/
#212380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#212390000000
0!
0'
0/
#212400000000
1!
1'
1/
#212410000000
0!
0'
0/
#212420000000
#212430000000
1!
1'
1/
#212440000000
0!
0'
0/
#212450000000
1!
1'
1/
#212460000000
0!
1"
0'
1(
0/
10
#212470000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#212480000000
0!
0'
0/
#212490000000
1!
1'
1/
#212500000000
0!
0'
0/
#212510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#212520000000
0!
0'
0/
#212530000000
1!
1'
1/
#212540000000
0!
1"
0'
1(
0/
10
#212550000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#212560000000
0!
1$
0'
1+
0/
#212570000000
1!
1'
1/
#212580000000
0!
0'
0/
#212590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#212600000000
0!
0'
0/
#212610000000
1!
1'
1/
#212620000000
0!
0'
0/
#212630000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#212640000000
0!
0'
0/
#212650000000
1!
1'
1/
#212660000000
0!
0'
0/
#212670000000
1!
1'
1/
#212680000000
0!
0'
0/
#212690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#212700000000
0!
0'
0/
#212710000000
1!
1'
1/
#212720000000
0!
0'
0/
#212730000000
1!
1'
1/
#212740000000
0!
0'
0/
#212750000000
1!
1'
1/
#212760000000
0!
0'
0/
#212770000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#212780000000
0!
0'
0/
#212790000000
1!
1'
1/
#212800000000
0!
0'
0/
#212810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#212820000000
0!
0'
0/
#212830000000
1!
1'
1/
#212840000000
0!
0'
0/
#212850000000
#212860000000
1!
1'
1/
#212870000000
0!
0'
0/
#212880000000
1!
1'
1/
#212890000000
0!
1"
0'
1(
0/
10
#212900000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#212910000000
0!
0'
0/
#212920000000
1!
1'
1/
#212930000000
0!
0'
0/
#212940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#212950000000
0!
0'
0/
#212960000000
1!
1'
1/
#212970000000
0!
1"
0'
1(
0/
10
#212980000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#212990000000
0!
1$
0'
1+
0/
#213000000000
1!
1'
1/
#213010000000
0!
0'
0/
#213020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#213030000000
0!
0'
0/
#213040000000
1!
1'
1/
#213050000000
0!
0'
0/
#213060000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#213070000000
0!
0'
0/
#213080000000
1!
1'
1/
#213090000000
0!
0'
0/
#213100000000
1!
1'
1/
#213110000000
0!
0'
0/
#213120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#213130000000
0!
0'
0/
#213140000000
1!
1'
1/
#213150000000
0!
0'
0/
#213160000000
1!
1'
1/
#213170000000
0!
0'
0/
#213180000000
1!
1'
1/
#213190000000
0!
0'
0/
#213200000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#213210000000
0!
0'
0/
#213220000000
1!
1'
1/
#213230000000
0!
0'
0/
#213240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#213250000000
0!
0'
0/
#213260000000
1!
1'
1/
#213270000000
0!
0'
0/
#213280000000
#213290000000
1!
1'
1/
#213300000000
0!
0'
0/
#213310000000
1!
1'
1/
#213320000000
0!
1"
0'
1(
0/
10
#213330000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#213340000000
0!
0'
0/
#213350000000
1!
1'
1/
#213360000000
0!
0'
0/
#213370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#213380000000
0!
0'
0/
#213390000000
1!
1'
1/
#213400000000
0!
1"
0'
1(
0/
10
#213410000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#213420000000
0!
1$
0'
1+
0/
#213430000000
1!
1'
1/
#213440000000
0!
0'
0/
#213450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#213460000000
0!
0'
0/
#213470000000
1!
1'
1/
#213480000000
0!
0'
0/
#213490000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#213500000000
0!
0'
0/
#213510000000
1!
1'
1/
#213520000000
0!
0'
0/
#213530000000
1!
1'
1/
#213540000000
0!
0'
0/
#213550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#213560000000
0!
0'
0/
#213570000000
1!
1'
1/
#213580000000
0!
0'
0/
#213590000000
1!
1'
1/
#213600000000
0!
0'
0/
#213610000000
1!
1'
1/
#213620000000
0!
0'
0/
#213630000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#213640000000
0!
0'
0/
#213650000000
1!
1'
1/
#213660000000
0!
0'
0/
#213670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#213680000000
0!
0'
0/
#213690000000
1!
1'
1/
#213700000000
0!
0'
0/
#213710000000
#213720000000
1!
1'
1/
#213730000000
0!
0'
0/
#213740000000
1!
1'
1/
#213750000000
0!
1"
0'
1(
0/
10
#213760000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#213770000000
0!
0'
0/
#213780000000
1!
1'
1/
#213790000000
0!
0'
0/
#213800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#213810000000
0!
0'
0/
#213820000000
1!
1'
1/
#213830000000
0!
1"
0'
1(
0/
10
#213840000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#213850000000
0!
1$
0'
1+
0/
#213860000000
1!
1'
1/
#213870000000
0!
0'
0/
#213880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#213890000000
0!
0'
0/
#213900000000
1!
1'
1/
#213910000000
0!
0'
0/
#213920000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#213930000000
0!
0'
0/
#213940000000
1!
1'
1/
#213950000000
0!
0'
0/
#213960000000
1!
1'
1/
#213970000000
0!
0'
0/
#213980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#213990000000
0!
0'
0/
#214000000000
1!
1'
1/
#214010000000
0!
0'
0/
#214020000000
1!
1'
1/
#214030000000
0!
0'
0/
#214040000000
1!
1'
1/
#214050000000
0!
0'
0/
#214060000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#214070000000
0!
0'
0/
#214080000000
1!
1'
1/
#214090000000
0!
0'
0/
#214100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#214110000000
0!
0'
0/
#214120000000
1!
1'
1/
#214130000000
0!
0'
0/
#214140000000
#214150000000
1!
1'
1/
#214160000000
0!
0'
0/
#214170000000
1!
1'
1/
#214180000000
0!
1"
0'
1(
0/
10
#214190000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#214200000000
0!
0'
0/
#214210000000
1!
1'
1/
#214220000000
0!
0'
0/
#214230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#214240000000
0!
0'
0/
#214250000000
1!
1'
1/
#214260000000
0!
1"
0'
1(
0/
10
#214270000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#214280000000
0!
1$
0'
1+
0/
#214290000000
1!
1'
1/
#214300000000
0!
0'
0/
#214310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#214320000000
0!
0'
0/
#214330000000
1!
1'
1/
#214340000000
0!
0'
0/
#214350000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#214360000000
0!
0'
0/
#214370000000
1!
1'
1/
#214380000000
0!
0'
0/
#214390000000
1!
1'
1/
#214400000000
0!
0'
0/
#214410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#214420000000
0!
0'
0/
#214430000000
1!
1'
1/
#214440000000
0!
0'
0/
#214450000000
1!
1'
1/
#214460000000
0!
0'
0/
#214470000000
1!
1'
1/
#214480000000
0!
0'
0/
#214490000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#214500000000
0!
0'
0/
#214510000000
1!
1'
1/
#214520000000
0!
0'
0/
#214530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#214540000000
0!
0'
0/
#214550000000
1!
1'
1/
#214560000000
0!
0'
0/
#214570000000
#214580000000
1!
1'
1/
#214590000000
0!
0'
0/
#214600000000
1!
1'
1/
#214610000000
0!
1"
0'
1(
0/
10
#214620000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#214630000000
0!
0'
0/
#214640000000
1!
1'
1/
#214650000000
0!
0'
0/
#214660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#214670000000
0!
0'
0/
#214680000000
1!
1'
1/
#214690000000
0!
1"
0'
1(
0/
10
#214700000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#214710000000
0!
1$
0'
1+
0/
#214720000000
1!
1'
1/
#214730000000
0!
0'
0/
#214740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#214750000000
0!
0'
0/
#214760000000
1!
1'
1/
#214770000000
0!
0'
0/
#214780000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#214790000000
0!
0'
0/
#214800000000
1!
1'
1/
#214810000000
0!
0'
0/
#214820000000
1!
1'
1/
#214830000000
0!
0'
0/
#214840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#214850000000
0!
0'
0/
#214860000000
1!
1'
1/
#214870000000
0!
0'
0/
#214880000000
1!
1'
1/
#214890000000
0!
0'
0/
#214900000000
1!
1'
1/
#214910000000
0!
0'
0/
#214920000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#214930000000
0!
0'
0/
#214940000000
1!
1'
1/
#214950000000
0!
0'
0/
#214960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#214970000000
0!
0'
0/
#214980000000
1!
1'
1/
#214990000000
0!
0'
0/
#215000000000
#215010000000
1!
1'
1/
#215020000000
0!
0'
0/
#215030000000
1!
1'
1/
#215040000000
0!
1"
0'
1(
0/
10
#215050000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#215060000000
0!
0'
0/
#215070000000
1!
1'
1/
#215080000000
0!
0'
0/
#215090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#215100000000
0!
0'
0/
#215110000000
1!
1'
1/
#215120000000
0!
1"
0'
1(
0/
10
#215130000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#215140000000
0!
1$
0'
1+
0/
#215150000000
1!
1'
1/
#215160000000
0!
0'
0/
#215170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#215180000000
0!
0'
0/
#215190000000
1!
1'
1/
#215200000000
0!
0'
0/
#215210000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#215220000000
0!
0'
0/
#215230000000
1!
1'
1/
#215240000000
0!
0'
0/
#215250000000
1!
1'
1/
#215260000000
0!
0'
0/
#215270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#215280000000
0!
0'
0/
#215290000000
1!
1'
1/
#215300000000
0!
0'
0/
#215310000000
1!
1'
1/
#215320000000
0!
0'
0/
#215330000000
1!
1'
1/
#215340000000
0!
0'
0/
#215350000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#215360000000
0!
0'
0/
#215370000000
1!
1'
1/
#215380000000
0!
0'
0/
#215390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#215400000000
0!
0'
0/
#215410000000
1!
1'
1/
#215420000000
0!
0'
0/
#215430000000
#215440000000
1!
1'
1/
#215450000000
0!
0'
0/
#215460000000
1!
1'
1/
#215470000000
0!
1"
0'
1(
0/
10
#215480000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#215490000000
0!
0'
0/
#215500000000
1!
1'
1/
#215510000000
0!
0'
0/
#215520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#215530000000
0!
0'
0/
#215540000000
1!
1'
1/
#215550000000
0!
1"
0'
1(
0/
10
#215560000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#215570000000
0!
1$
0'
1+
0/
#215580000000
1!
1'
1/
#215590000000
0!
0'
0/
#215600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#215610000000
0!
0'
0/
#215620000000
1!
1'
1/
#215630000000
0!
0'
0/
#215640000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#215650000000
0!
0'
0/
#215660000000
1!
1'
1/
#215670000000
0!
0'
0/
#215680000000
1!
1'
1/
#215690000000
0!
0'
0/
#215700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#215710000000
0!
0'
0/
#215720000000
1!
1'
1/
#215730000000
0!
0'
0/
#215740000000
1!
1'
1/
#215750000000
0!
0'
0/
#215760000000
1!
1'
1/
#215770000000
0!
0'
0/
#215780000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#215790000000
0!
0'
0/
#215800000000
1!
1'
1/
#215810000000
0!
0'
0/
#215820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#215830000000
0!
0'
0/
#215840000000
1!
1'
1/
#215850000000
0!
0'
0/
#215860000000
#215870000000
1!
1'
1/
#215880000000
0!
0'
0/
#215890000000
1!
1'
1/
#215900000000
0!
1"
0'
1(
0/
10
#215910000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#215920000000
0!
0'
0/
#215930000000
1!
1'
1/
#215940000000
0!
0'
0/
#215950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#215960000000
0!
0'
0/
#215970000000
1!
1'
1/
#215980000000
0!
1"
0'
1(
0/
10
#215990000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#216000000000
0!
1$
0'
1+
0/
#216010000000
1!
1'
1/
#216020000000
0!
0'
0/
#216030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#216040000000
0!
0'
0/
#216050000000
1!
1'
1/
#216060000000
0!
0'
0/
#216070000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#216080000000
0!
0'
0/
#216090000000
1!
1'
1/
#216100000000
0!
0'
0/
#216110000000
1!
1'
1/
#216120000000
0!
0'
0/
#216130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#216140000000
0!
0'
0/
#216150000000
1!
1'
1/
#216160000000
0!
0'
0/
#216170000000
1!
1'
1/
#216180000000
0!
0'
0/
#216190000000
1!
1'
1/
#216200000000
0!
0'
0/
#216210000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#216220000000
0!
0'
0/
#216230000000
1!
1'
1/
#216240000000
0!
0'
0/
#216250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#216260000000
0!
0'
0/
#216270000000
1!
1'
1/
#216280000000
0!
0'
0/
#216290000000
#216300000000
1!
1'
1/
#216310000000
0!
0'
0/
#216320000000
1!
1'
1/
#216330000000
0!
1"
0'
1(
0/
10
#216340000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#216350000000
0!
0'
0/
#216360000000
1!
1'
1/
#216370000000
0!
0'
0/
#216380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#216390000000
0!
0'
0/
#216400000000
1!
1'
1/
#216410000000
0!
1"
0'
1(
0/
10
#216420000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#216430000000
0!
1$
0'
1+
0/
#216440000000
1!
1'
1/
#216450000000
0!
0'
0/
#216460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#216470000000
0!
0'
0/
#216480000000
1!
1'
1/
#216490000000
0!
0'
0/
#216500000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#216510000000
0!
0'
0/
#216520000000
1!
1'
1/
#216530000000
0!
0'
0/
#216540000000
1!
1'
1/
#216550000000
0!
0'
0/
#216560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#216570000000
0!
0'
0/
#216580000000
1!
1'
1/
#216590000000
0!
0'
0/
#216600000000
1!
1'
1/
#216610000000
0!
0'
0/
#216620000000
1!
1'
1/
#216630000000
0!
0'
0/
#216640000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#216650000000
0!
0'
0/
#216660000000
1!
1'
1/
#216670000000
0!
0'
0/
#216680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#216690000000
0!
0'
0/
#216700000000
1!
1'
1/
#216710000000
0!
0'
0/
#216720000000
#216730000000
1!
1'
1/
#216740000000
0!
0'
0/
#216750000000
1!
1'
1/
#216760000000
0!
1"
0'
1(
0/
10
#216770000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#216780000000
0!
0'
0/
#216790000000
1!
1'
1/
#216800000000
0!
0'
0/
#216810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#216820000000
0!
0'
0/
#216830000000
1!
1'
1/
#216840000000
0!
1"
0'
1(
0/
10
#216850000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#216860000000
0!
1$
0'
1+
0/
#216870000000
1!
1'
1/
#216880000000
0!
0'
0/
#216890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#216900000000
0!
0'
0/
#216910000000
1!
1'
1/
#216920000000
0!
0'
0/
#216930000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#216940000000
0!
0'
0/
#216950000000
1!
1'
1/
#216960000000
0!
0'
0/
#216970000000
1!
1'
1/
#216980000000
0!
0'
0/
#216990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#217000000000
0!
0'
0/
#217010000000
1!
1'
1/
#217020000000
0!
0'
0/
#217030000000
1!
1'
1/
#217040000000
0!
0'
0/
#217050000000
1!
1'
1/
#217060000000
0!
0'
0/
#217070000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#217080000000
0!
0'
0/
#217090000000
1!
1'
1/
#217100000000
0!
0'
0/
#217110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#217120000000
0!
0'
0/
#217130000000
1!
1'
1/
#217140000000
0!
0'
0/
#217150000000
#217160000000
1!
1'
1/
#217170000000
0!
0'
0/
#217180000000
1!
1'
1/
#217190000000
0!
1"
0'
1(
0/
10
#217200000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#217210000000
0!
0'
0/
#217220000000
1!
1'
1/
#217230000000
0!
0'
0/
#217240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#217250000000
0!
0'
0/
#217260000000
1!
1'
1/
#217270000000
0!
1"
0'
1(
0/
10
#217280000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#217290000000
0!
1$
0'
1+
0/
#217300000000
1!
1'
1/
#217310000000
0!
0'
0/
#217320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#217330000000
0!
0'
0/
#217340000000
1!
1'
1/
#217350000000
0!
0'
0/
#217360000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#217370000000
0!
0'
0/
#217380000000
1!
1'
1/
#217390000000
0!
0'
0/
#217400000000
1!
1'
1/
#217410000000
0!
0'
0/
#217420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#217430000000
0!
0'
0/
#217440000000
1!
1'
1/
#217450000000
0!
0'
0/
#217460000000
1!
1'
1/
#217470000000
0!
0'
0/
#217480000000
1!
1'
1/
#217490000000
0!
0'
0/
#217500000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#217510000000
0!
0'
0/
#217520000000
1!
1'
1/
#217530000000
0!
0'
0/
#217540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#217550000000
0!
0'
0/
#217560000000
1!
1'
1/
#217570000000
0!
0'
0/
#217580000000
#217590000000
1!
1'
1/
#217600000000
0!
0'
0/
#217610000000
1!
1'
1/
#217620000000
0!
1"
0'
1(
0/
10
#217630000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#217640000000
0!
0'
0/
#217650000000
1!
1'
1/
#217660000000
0!
0'
0/
#217670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#217680000000
0!
0'
0/
#217690000000
1!
1'
1/
#217700000000
0!
1"
0'
1(
0/
10
#217710000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#217720000000
0!
1$
0'
1+
0/
#217730000000
1!
1'
1/
#217740000000
0!
0'
0/
#217750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#217760000000
0!
0'
0/
#217770000000
1!
1'
1/
#217780000000
0!
0'
0/
#217790000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#217800000000
0!
0'
0/
#217810000000
1!
1'
1/
#217820000000
0!
0'
0/
#217830000000
1!
1'
1/
#217840000000
0!
0'
0/
#217850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#217860000000
0!
0'
0/
#217870000000
1!
1'
1/
#217880000000
0!
0'
0/
#217890000000
1!
1'
1/
#217900000000
0!
0'
0/
#217910000000
1!
1'
1/
#217920000000
0!
0'
0/
#217930000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#217940000000
0!
0'
0/
#217950000000
1!
1'
1/
#217960000000
0!
0'
0/
#217970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#217980000000
0!
0'
0/
#217990000000
1!
1'
1/
#218000000000
0!
0'
0/
#218010000000
#218020000000
1!
1'
1/
#218030000000
0!
0'
0/
#218040000000
1!
1'
1/
#218050000000
0!
1"
0'
1(
0/
10
#218060000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#218070000000
0!
0'
0/
#218080000000
1!
1'
1/
#218090000000
0!
0'
0/
#218100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#218110000000
0!
0'
0/
#218120000000
1!
1'
1/
#218130000000
0!
1"
0'
1(
0/
10
#218140000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#218150000000
0!
1$
0'
1+
0/
#218160000000
1!
1'
1/
#218170000000
0!
0'
0/
#218180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#218190000000
0!
0'
0/
#218200000000
1!
1'
1/
#218210000000
0!
0'
0/
#218220000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#218230000000
0!
0'
0/
#218240000000
1!
1'
1/
#218250000000
0!
0'
0/
#218260000000
1!
1'
1/
#218270000000
0!
0'
0/
#218280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#218290000000
0!
0'
0/
#218300000000
1!
1'
1/
#218310000000
0!
0'
0/
#218320000000
1!
1'
1/
#218330000000
0!
0'
0/
#218340000000
1!
1'
1/
#218350000000
0!
0'
0/
#218360000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#218370000000
0!
0'
0/
#218380000000
1!
1'
1/
#218390000000
0!
0'
0/
#218400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#218410000000
0!
0'
0/
#218420000000
1!
1'
1/
#218430000000
0!
0'
0/
#218440000000
#218450000000
1!
1'
1/
#218460000000
0!
0'
0/
#218470000000
1!
1'
1/
#218480000000
0!
1"
0'
1(
0/
10
#218490000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#218500000000
0!
0'
0/
#218510000000
1!
1'
1/
#218520000000
0!
0'
0/
#218530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#218540000000
0!
0'
0/
#218550000000
1!
1'
1/
#218560000000
0!
1"
0'
1(
0/
10
#218570000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#218580000000
0!
1$
0'
1+
0/
#218590000000
1!
1'
1/
#218600000000
0!
0'
0/
#218610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#218620000000
0!
0'
0/
#218630000000
1!
1'
1/
#218640000000
0!
0'
0/
#218650000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#218660000000
0!
0'
0/
#218670000000
1!
1'
1/
#218680000000
0!
0'
0/
#218690000000
1!
1'
1/
#218700000000
0!
0'
0/
#218710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#218720000000
0!
0'
0/
#218730000000
1!
1'
1/
#218740000000
0!
0'
0/
#218750000000
1!
1'
1/
#218760000000
0!
0'
0/
#218770000000
1!
1'
1/
#218780000000
0!
0'
0/
#218790000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#218800000000
0!
0'
0/
#218810000000
1!
1'
1/
#218820000000
0!
0'
0/
#218830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#218840000000
0!
0'
0/
#218850000000
1!
1'
1/
#218860000000
0!
0'
0/
#218870000000
#218880000000
1!
1'
1/
#218890000000
0!
0'
0/
#218900000000
1!
1'
1/
#218910000000
0!
1"
0'
1(
0/
10
#218920000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#218930000000
0!
0'
0/
#218940000000
1!
1'
1/
#218950000000
0!
0'
0/
#218960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#218970000000
0!
0'
0/
#218980000000
1!
1'
1/
#218990000000
0!
1"
0'
1(
0/
10
#219000000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#219010000000
0!
1$
0'
1+
0/
#219020000000
1!
1'
1/
#219030000000
0!
0'
0/
#219040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#219050000000
0!
0'
0/
#219060000000
1!
1'
1/
#219070000000
0!
0'
0/
#219080000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#219090000000
0!
0'
0/
#219100000000
1!
1'
1/
#219110000000
0!
0'
0/
#219120000000
1!
1'
1/
#219130000000
0!
0'
0/
#219140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#219150000000
0!
0'
0/
#219160000000
1!
1'
1/
#219170000000
0!
0'
0/
#219180000000
1!
1'
1/
#219190000000
0!
0'
0/
#219200000000
1!
1'
1/
#219210000000
0!
0'
0/
#219220000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#219230000000
0!
0'
0/
#219240000000
1!
1'
1/
#219250000000
0!
0'
0/
#219260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#219270000000
0!
0'
0/
#219280000000
1!
1'
1/
#219290000000
0!
0'
0/
#219300000000
#219310000000
1!
1'
1/
#219320000000
0!
0'
0/
#219330000000
1!
1'
1/
#219340000000
0!
1"
0'
1(
0/
10
#219350000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#219360000000
0!
0'
0/
#219370000000
1!
1'
1/
#219380000000
0!
0'
0/
#219390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#219400000000
0!
0'
0/
#219410000000
1!
1'
1/
#219420000000
0!
1"
0'
1(
0/
10
#219430000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#219440000000
0!
1$
0'
1+
0/
#219450000000
1!
1'
1/
#219460000000
0!
0'
0/
#219470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#219480000000
0!
0'
0/
#219490000000
1!
1'
1/
#219500000000
0!
0'
0/
#219510000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#219520000000
0!
0'
0/
#219530000000
1!
1'
1/
#219540000000
0!
0'
0/
#219550000000
1!
1'
1/
#219560000000
0!
0'
0/
#219570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#219580000000
0!
0'
0/
#219590000000
1!
1'
1/
#219600000000
0!
0'
0/
#219610000000
1!
1'
1/
#219620000000
0!
0'
0/
#219630000000
1!
1'
1/
#219640000000
0!
0'
0/
#219650000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#219660000000
0!
0'
0/
#219670000000
1!
1'
1/
#219680000000
0!
0'
0/
#219690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#219700000000
0!
0'
0/
#219710000000
1!
1'
1/
#219720000000
0!
0'
0/
#219730000000
#219740000000
1!
1'
1/
#219750000000
0!
0'
0/
#219760000000
1!
1'
1/
#219770000000
0!
1"
0'
1(
0/
10
#219780000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#219790000000
0!
0'
0/
#219800000000
1!
1'
1/
#219810000000
0!
0'
0/
#219820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#219830000000
0!
0'
0/
#219840000000
1!
1'
1/
#219850000000
0!
1"
0'
1(
0/
10
#219860000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#219870000000
0!
1$
0'
1+
0/
#219880000000
1!
1'
1/
#219890000000
0!
0'
0/
#219900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#219910000000
0!
0'
0/
#219920000000
1!
1'
1/
#219930000000
0!
0'
0/
#219940000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#219950000000
0!
0'
0/
#219960000000
1!
1'
1/
#219970000000
0!
0'
0/
#219980000000
1!
1'
1/
#219990000000
0!
0'
0/
#220000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#220010000000
0!
0'
0/
#220020000000
1!
1'
1/
#220030000000
0!
0'
0/
#220040000000
1!
1'
1/
#220050000000
0!
0'
0/
#220060000000
1!
1'
1/
#220070000000
0!
0'
0/
#220080000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#220090000000
0!
0'
0/
#220100000000
1!
1'
1/
#220110000000
0!
0'
0/
#220120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#220130000000
0!
0'
0/
#220140000000
1!
1'
1/
#220150000000
0!
0'
0/
#220160000000
#220170000000
1!
1'
1/
#220180000000
0!
0'
0/
#220190000000
1!
1'
1/
#220200000000
0!
1"
0'
1(
0/
10
#220210000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#220220000000
0!
0'
0/
#220230000000
1!
1'
1/
#220240000000
0!
0'
0/
#220250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#220260000000
0!
0'
0/
#220270000000
1!
1'
1/
#220280000000
0!
1"
0'
1(
0/
10
#220290000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#220300000000
0!
1$
0'
1+
0/
#220310000000
1!
1'
1/
#220320000000
0!
0'
0/
#220330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#220340000000
0!
0'
0/
#220350000000
1!
1'
1/
#220360000000
0!
0'
0/
#220370000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#220380000000
0!
0'
0/
#220390000000
1!
1'
1/
#220400000000
0!
0'
0/
#220410000000
1!
1'
1/
#220420000000
0!
0'
0/
#220430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#220440000000
0!
0'
0/
#220450000000
1!
1'
1/
#220460000000
0!
0'
0/
#220470000000
1!
1'
1/
#220480000000
0!
0'
0/
#220490000000
1!
1'
1/
#220500000000
0!
0'
0/
#220510000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#220520000000
0!
0'
0/
#220530000000
1!
1'
1/
#220540000000
0!
0'
0/
#220550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#220560000000
0!
0'
0/
#220570000000
1!
1'
1/
#220580000000
0!
0'
0/
#220590000000
#220600000000
1!
1'
1/
#220610000000
0!
0'
0/
#220620000000
1!
1'
1/
#220630000000
0!
1"
0'
1(
0/
10
#220640000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#220650000000
0!
0'
0/
#220660000000
1!
1'
1/
#220670000000
0!
0'
0/
#220680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#220690000000
0!
0'
0/
#220700000000
1!
1'
1/
#220710000000
0!
1"
0'
1(
0/
10
#220720000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#220730000000
0!
1$
0'
1+
0/
#220740000000
1!
1'
1/
#220750000000
0!
0'
0/
#220760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#220770000000
0!
0'
0/
#220780000000
1!
1'
1/
#220790000000
0!
0'
0/
#220800000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#220810000000
0!
0'
0/
#220820000000
1!
1'
1/
#220830000000
0!
0'
0/
#220840000000
1!
1'
1/
#220850000000
0!
0'
0/
#220860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#220870000000
0!
0'
0/
#220880000000
1!
1'
1/
#220890000000
0!
0'
0/
#220900000000
1!
1'
1/
#220910000000
0!
0'
0/
#220920000000
1!
1'
1/
#220930000000
0!
0'
0/
#220940000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#220950000000
0!
0'
0/
#220960000000
1!
1'
1/
#220970000000
0!
0'
0/
#220980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#220990000000
0!
0'
0/
#221000000000
1!
1'
1/
#221010000000
0!
0'
0/
#221020000000
#221030000000
1!
1'
1/
#221040000000
0!
0'
0/
#221050000000
1!
1'
1/
#221060000000
0!
1"
0'
1(
0/
10
#221070000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#221080000000
0!
0'
0/
#221090000000
1!
1'
1/
#221100000000
0!
0'
0/
#221110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#221120000000
0!
0'
0/
#221130000000
1!
1'
1/
#221140000000
0!
1"
0'
1(
0/
10
#221150000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#221160000000
0!
1$
0'
1+
0/
#221170000000
1!
1'
1/
#221180000000
0!
0'
0/
#221190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#221200000000
0!
0'
0/
#221210000000
1!
1'
1/
#221220000000
0!
0'
0/
#221230000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#221240000000
0!
0'
0/
#221250000000
1!
1'
1/
#221260000000
0!
0'
0/
#221270000000
1!
1'
1/
#221280000000
0!
0'
0/
#221290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#221300000000
0!
0'
0/
#221310000000
1!
1'
1/
#221320000000
0!
0'
0/
#221330000000
1!
1'
1/
#221340000000
0!
0'
0/
#221350000000
1!
1'
1/
#221360000000
0!
0'
0/
#221370000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#221380000000
0!
0'
0/
#221390000000
1!
1'
1/
#221400000000
0!
0'
0/
#221410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#221420000000
0!
0'
0/
#221430000000
1!
1'
1/
#221440000000
0!
0'
0/
#221450000000
#221460000000
1!
1'
1/
#221470000000
0!
0'
0/
#221480000000
1!
1'
1/
#221490000000
0!
1"
0'
1(
0/
10
#221500000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#221510000000
0!
0'
0/
#221520000000
1!
1'
1/
#221530000000
0!
0'
0/
#221540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#221550000000
0!
0'
0/
#221560000000
1!
1'
1/
#221570000000
0!
1"
0'
1(
0/
10
#221580000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#221590000000
0!
1$
0'
1+
0/
#221600000000
1!
1'
1/
#221610000000
0!
0'
0/
#221620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#221630000000
0!
0'
0/
#221640000000
1!
1'
1/
#221650000000
0!
0'
0/
#221660000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#221670000000
0!
0'
0/
#221680000000
1!
1'
1/
#221690000000
0!
0'
0/
#221700000000
1!
1'
1/
#221710000000
0!
0'
0/
#221720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#221730000000
0!
0'
0/
#221740000000
1!
1'
1/
#221750000000
0!
0'
0/
#221760000000
1!
1'
1/
#221770000000
0!
0'
0/
#221780000000
1!
1'
1/
#221790000000
0!
0'
0/
#221800000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#221810000000
0!
0'
0/
#221820000000
1!
1'
1/
#221830000000
0!
0'
0/
#221840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#221850000000
0!
0'
0/
#221860000000
1!
1'
1/
#221870000000
0!
0'
0/
#221880000000
#221890000000
1!
1'
1/
#221900000000
0!
0'
0/
#221910000000
1!
1'
1/
#221920000000
0!
1"
0'
1(
0/
10
#221930000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#221940000000
0!
0'
0/
#221950000000
1!
1'
1/
#221960000000
0!
0'
0/
#221970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#221980000000
0!
0'
0/
#221990000000
1!
1'
1/
#222000000000
0!
1"
0'
1(
0/
10
#222010000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#222020000000
0!
1$
0'
1+
0/
#222030000000
1!
1'
1/
#222040000000
0!
0'
0/
#222050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#222060000000
0!
0'
0/
#222070000000
1!
1'
1/
#222080000000
0!
0'
0/
#222090000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#222100000000
0!
0'
0/
#222110000000
1!
1'
1/
#222120000000
0!
0'
0/
#222130000000
1!
1'
1/
#222140000000
0!
0'
0/
#222150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#222160000000
0!
0'
0/
#222170000000
1!
1'
1/
#222180000000
0!
0'
0/
#222190000000
1!
1'
1/
#222200000000
0!
0'
0/
#222210000000
1!
1'
1/
#222220000000
0!
0'
0/
#222230000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#222240000000
0!
0'
0/
#222250000000
1!
1'
1/
#222260000000
0!
0'
0/
#222270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#222280000000
0!
0'
0/
#222290000000
1!
1'
1/
#222300000000
0!
0'
0/
#222310000000
#222320000000
1!
1'
1/
#222330000000
0!
0'
0/
#222340000000
1!
1'
1/
#222350000000
0!
1"
0'
1(
0/
10
#222360000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#222370000000
0!
0'
0/
#222380000000
1!
1'
1/
#222390000000
0!
0'
0/
#222400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#222410000000
0!
0'
0/
#222420000000
1!
1'
1/
#222430000000
0!
1"
0'
1(
0/
10
#222440000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#222450000000
0!
1$
0'
1+
0/
#222460000000
1!
1'
1/
#222470000000
0!
0'
0/
#222480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#222490000000
0!
0'
0/
#222500000000
1!
1'
1/
#222510000000
0!
0'
0/
#222520000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#222530000000
0!
0'
0/
#222540000000
1!
1'
1/
#222550000000
0!
0'
0/
#222560000000
1!
1'
1/
#222570000000
0!
0'
0/
#222580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#222590000000
0!
0'
0/
#222600000000
1!
1'
1/
#222610000000
0!
0'
0/
#222620000000
1!
1'
1/
#222630000000
0!
0'
0/
#222640000000
1!
1'
1/
#222650000000
0!
0'
0/
#222660000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#222670000000
0!
0'
0/
#222680000000
1!
1'
1/
#222690000000
0!
0'
0/
#222700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#222710000000
0!
0'
0/
#222720000000
1!
1'
1/
#222730000000
0!
0'
0/
#222740000000
#222750000000
1!
1'
1/
#222760000000
0!
0'
0/
#222770000000
1!
1'
1/
#222780000000
0!
1"
0'
1(
0/
10
#222790000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#222800000000
0!
0'
0/
#222810000000
1!
1'
1/
#222820000000
0!
0'
0/
#222830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#222840000000
0!
0'
0/
#222850000000
1!
1'
1/
#222860000000
0!
1"
0'
1(
0/
10
#222870000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#222880000000
0!
1$
0'
1+
0/
#222890000000
1!
1'
1/
#222900000000
0!
0'
0/
#222910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#222920000000
0!
0'
0/
#222930000000
1!
1'
1/
#222940000000
0!
0'
0/
#222950000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#222960000000
0!
0'
0/
#222970000000
1!
1'
1/
#222980000000
0!
0'
0/
#222990000000
1!
1'
1/
#223000000000
0!
0'
0/
#223010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#223020000000
0!
0'
0/
#223030000000
1!
1'
1/
#223040000000
0!
0'
0/
#223050000000
1!
1'
1/
#223060000000
0!
0'
0/
#223070000000
1!
1'
1/
#223080000000
0!
0'
0/
#223090000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#223100000000
0!
0'
0/
#223110000000
1!
1'
1/
#223120000000
0!
0'
0/
#223130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#223140000000
0!
0'
0/
#223150000000
1!
1'
1/
#223160000000
0!
0'
0/
#223170000000
#223180000000
1!
1'
1/
#223190000000
0!
0'
0/
#223200000000
1!
1'
1/
#223210000000
0!
1"
0'
1(
0/
10
#223220000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#223230000000
0!
0'
0/
#223240000000
1!
1'
1/
#223250000000
0!
0'
0/
#223260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#223270000000
0!
0'
0/
#223280000000
1!
1'
1/
#223290000000
0!
1"
0'
1(
0/
10
#223300000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#223310000000
0!
1$
0'
1+
0/
#223320000000
1!
1'
1/
#223330000000
0!
0'
0/
#223340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#223350000000
0!
0'
0/
#223360000000
1!
1'
1/
#223370000000
0!
0'
0/
#223380000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#223390000000
0!
0'
0/
#223400000000
1!
1'
1/
#223410000000
0!
0'
0/
#223420000000
1!
1'
1/
#223430000000
0!
0'
0/
#223440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#223450000000
0!
0'
0/
#223460000000
1!
1'
1/
#223470000000
0!
0'
0/
#223480000000
1!
1'
1/
#223490000000
0!
0'
0/
#223500000000
1!
1'
1/
#223510000000
0!
0'
0/
#223520000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#223530000000
0!
0'
0/
#223540000000
1!
1'
1/
#223550000000
0!
0'
0/
#223560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#223570000000
0!
0'
0/
#223580000000
1!
1'
1/
#223590000000
0!
0'
0/
#223600000000
#223610000000
1!
1'
1/
#223620000000
0!
0'
0/
#223630000000
1!
1'
1/
#223640000000
0!
1"
0'
1(
0/
10
#223650000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#223660000000
0!
0'
0/
#223670000000
1!
1'
1/
#223680000000
0!
0'
0/
#223690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#223700000000
0!
0'
0/
#223710000000
1!
1'
1/
#223720000000
0!
1"
0'
1(
0/
10
#223730000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#223740000000
0!
1$
0'
1+
0/
#223750000000
1!
1'
1/
#223760000000
0!
0'
0/
#223770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#223780000000
0!
0'
0/
#223790000000
1!
1'
1/
#223800000000
0!
0'
0/
#223810000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#223820000000
0!
0'
0/
#223830000000
1!
1'
1/
#223840000000
0!
0'
0/
#223850000000
1!
1'
1/
#223860000000
0!
0'
0/
#223870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#223880000000
0!
0'
0/
#223890000000
1!
1'
1/
#223900000000
0!
0'
0/
#223910000000
1!
1'
1/
#223920000000
0!
0'
0/
#223930000000
1!
1'
1/
#223940000000
0!
0'
0/
#223950000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#223960000000
0!
0'
0/
#223970000000
1!
1'
1/
#223980000000
0!
0'
0/
#223990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#224000000000
0!
0'
0/
#224010000000
1!
1'
1/
#224020000000
0!
0'
0/
#224030000000
#224040000000
1!
1'
1/
#224050000000
0!
0'
0/
#224060000000
1!
1'
1/
#224070000000
0!
1"
0'
1(
0/
10
#224080000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#224090000000
0!
0'
0/
#224100000000
1!
1'
1/
#224110000000
0!
0'
0/
#224120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#224130000000
0!
0'
0/
#224140000000
1!
1'
1/
#224150000000
0!
1"
0'
1(
0/
10
#224160000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#224170000000
0!
1$
0'
1+
0/
#224180000000
1!
1'
1/
#224190000000
0!
0'
0/
#224200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#224210000000
0!
0'
0/
#224220000000
1!
1'
1/
#224230000000
0!
0'
0/
#224240000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#224250000000
0!
0'
0/
#224260000000
1!
1'
1/
#224270000000
0!
0'
0/
#224280000000
1!
1'
1/
#224290000000
0!
0'
0/
#224300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#224310000000
0!
0'
0/
#224320000000
1!
1'
1/
#224330000000
0!
0'
0/
#224340000000
1!
1'
1/
#224350000000
0!
0'
0/
#224360000000
1!
1'
1/
#224370000000
0!
0'
0/
#224380000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#224390000000
0!
0'
0/
#224400000000
1!
1'
1/
#224410000000
0!
0'
0/
#224420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#224430000000
0!
0'
0/
#224440000000
1!
1'
1/
#224450000000
0!
0'
0/
#224460000000
#224470000000
1!
1'
1/
#224480000000
0!
0'
0/
#224490000000
1!
1'
1/
#224500000000
0!
1"
0'
1(
0/
10
#224510000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#224520000000
0!
0'
0/
#224530000000
1!
1'
1/
#224540000000
0!
0'
0/
#224550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#224560000000
0!
0'
0/
#224570000000
1!
1'
1/
#224580000000
0!
1"
0'
1(
0/
10
#224590000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#224600000000
0!
1$
0'
1+
0/
#224610000000
1!
1'
1/
#224620000000
0!
0'
0/
#224630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#224640000000
0!
0'
0/
#224650000000
1!
1'
1/
#224660000000
0!
0'
0/
#224670000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#224680000000
0!
0'
0/
#224690000000
1!
1'
1/
#224700000000
0!
0'
0/
#224710000000
1!
1'
1/
#224720000000
0!
0'
0/
#224730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#224740000000
0!
0'
0/
#224750000000
1!
1'
1/
#224760000000
0!
0'
0/
#224770000000
1!
1'
1/
#224780000000
0!
0'
0/
#224790000000
1!
1'
1/
#224800000000
0!
0'
0/
#224810000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#224820000000
0!
0'
0/
#224830000000
1!
1'
1/
#224840000000
0!
0'
0/
#224850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#224860000000
0!
0'
0/
#224870000000
1!
1'
1/
#224880000000
0!
0'
0/
#224890000000
#224900000000
1!
1'
1/
#224910000000
0!
0'
0/
#224920000000
1!
1'
1/
#224930000000
0!
1"
0'
1(
0/
10
#224940000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#224950000000
0!
0'
0/
#224960000000
1!
1'
1/
#224970000000
0!
0'
0/
#224980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#224990000000
0!
0'
0/
#225000000000
1!
1'
1/
#225010000000
0!
1"
0'
1(
0/
10
#225020000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#225030000000
0!
1$
0'
1+
0/
#225040000000
1!
1'
1/
#225050000000
0!
0'
0/
#225060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#225070000000
0!
0'
0/
#225080000000
1!
1'
1/
#225090000000
0!
0'
0/
#225100000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#225110000000
0!
0'
0/
#225120000000
1!
1'
1/
#225130000000
0!
0'
0/
#225140000000
1!
1'
1/
#225150000000
0!
0'
0/
#225160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#225170000000
0!
0'
0/
#225180000000
1!
1'
1/
#225190000000
0!
0'
0/
#225200000000
1!
1'
1/
#225210000000
0!
0'
0/
#225220000000
1!
1'
1/
#225230000000
0!
0'
0/
#225240000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#225250000000
0!
0'
0/
#225260000000
1!
1'
1/
#225270000000
0!
0'
0/
#225280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#225290000000
0!
0'
0/
#225300000000
1!
1'
1/
#225310000000
0!
0'
0/
#225320000000
#225330000000
1!
1'
1/
#225340000000
0!
0'
0/
#225350000000
1!
1'
1/
#225360000000
0!
1"
0'
1(
0/
10
#225370000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#225380000000
0!
0'
0/
#225390000000
1!
1'
1/
#225400000000
0!
0'
0/
#225410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#225420000000
0!
0'
0/
#225430000000
1!
1'
1/
#225440000000
0!
1"
0'
1(
0/
10
#225450000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#225460000000
0!
1$
0'
1+
0/
#225470000000
1!
1'
1/
#225480000000
0!
0'
0/
#225490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#225500000000
0!
0'
0/
#225510000000
1!
1'
1/
#225520000000
0!
0'
0/
#225530000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#225540000000
0!
0'
0/
#225550000000
1!
1'
1/
#225560000000
0!
0'
0/
#225570000000
1!
1'
1/
#225580000000
0!
0'
0/
#225590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#225600000000
0!
0'
0/
#225610000000
1!
1'
1/
#225620000000
0!
0'
0/
#225630000000
1!
1'
1/
#225640000000
0!
0'
0/
#225650000000
1!
1'
1/
#225660000000
0!
0'
0/
#225670000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#225680000000
0!
0'
0/
#225690000000
1!
1'
1/
#225700000000
0!
0'
0/
#225710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#225720000000
0!
0'
0/
#225730000000
1!
1'
1/
#225740000000
0!
0'
0/
#225750000000
#225760000000
1!
1'
1/
#225770000000
0!
0'
0/
#225780000000
1!
1'
1/
#225790000000
0!
1"
0'
1(
0/
10
#225800000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#225810000000
0!
0'
0/
#225820000000
1!
1'
1/
#225830000000
0!
0'
0/
#225840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#225850000000
0!
0'
0/
#225860000000
1!
1'
1/
#225870000000
0!
1"
0'
1(
0/
10
#225880000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#225890000000
0!
1$
0'
1+
0/
#225900000000
1!
1'
1/
#225910000000
0!
0'
0/
#225920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#225930000000
0!
0'
0/
#225940000000
1!
1'
1/
#225950000000
0!
0'
0/
#225960000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#225970000000
0!
0'
0/
#225980000000
1!
1'
1/
#225990000000
0!
0'
0/
#226000000000
1!
1'
1/
#226010000000
0!
0'
0/
#226020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#226030000000
0!
0'
0/
#226040000000
1!
1'
1/
#226050000000
0!
0'
0/
#226060000000
1!
1'
1/
#226070000000
0!
0'
0/
#226080000000
1!
1'
1/
#226090000000
0!
0'
0/
#226100000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#226110000000
0!
0'
0/
#226120000000
1!
1'
1/
#226130000000
0!
0'
0/
#226140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#226150000000
0!
0'
0/
#226160000000
1!
1'
1/
#226170000000
0!
0'
0/
#226180000000
#226190000000
1!
1'
1/
#226200000000
0!
0'
0/
#226210000000
1!
1'
1/
#226220000000
0!
1"
0'
1(
0/
10
#226230000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#226240000000
0!
0'
0/
#226250000000
1!
1'
1/
#226260000000
0!
0'
0/
#226270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#226280000000
0!
0'
0/
#226290000000
1!
1'
1/
#226300000000
0!
1"
0'
1(
0/
10
#226310000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#226320000000
0!
1$
0'
1+
0/
#226330000000
1!
1'
1/
#226340000000
0!
0'
0/
#226350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#226360000000
0!
0'
0/
#226370000000
1!
1'
1/
#226380000000
0!
0'
0/
#226390000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#226400000000
0!
0'
0/
#226410000000
1!
1'
1/
#226420000000
0!
0'
0/
#226430000000
1!
1'
1/
#226440000000
0!
0'
0/
#226450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#226460000000
0!
0'
0/
#226470000000
1!
1'
1/
#226480000000
0!
0'
0/
#226490000000
1!
1'
1/
#226500000000
0!
0'
0/
#226510000000
1!
1'
1/
#226520000000
0!
0'
0/
#226530000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#226540000000
0!
0'
0/
#226550000000
1!
1'
1/
#226560000000
0!
0'
0/
#226570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#226580000000
0!
0'
0/
#226590000000
1!
1'
1/
#226600000000
0!
0'
0/
#226610000000
#226620000000
1!
1'
1/
#226630000000
0!
0'
0/
#226640000000
1!
1'
1/
#226650000000
0!
1"
0'
1(
0/
10
#226660000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#226670000000
0!
0'
0/
#226680000000
1!
1'
1/
#226690000000
0!
0'
0/
#226700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#226710000000
0!
0'
0/
#226720000000
1!
1'
1/
#226730000000
0!
1"
0'
1(
0/
10
#226740000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#226750000000
0!
1$
0'
1+
0/
#226760000000
1!
1'
1/
#226770000000
0!
0'
0/
#226780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#226790000000
0!
0'
0/
#226800000000
1!
1'
1/
#226810000000
0!
0'
0/
#226820000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#226830000000
0!
0'
0/
#226840000000
1!
1'
1/
#226850000000
0!
0'
0/
#226860000000
1!
1'
1/
#226870000000
0!
0'
0/
#226880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#226890000000
0!
0'
0/
#226900000000
1!
1'
1/
#226910000000
0!
0'
0/
#226920000000
1!
1'
1/
#226930000000
0!
0'
0/
#226940000000
1!
1'
1/
#226950000000
0!
0'
0/
#226960000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#226970000000
0!
0'
0/
#226980000000
1!
1'
1/
#226990000000
0!
0'
0/
#227000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#227010000000
0!
0'
0/
#227020000000
1!
1'
1/
#227030000000
0!
0'
0/
#227040000000
#227050000000
1!
1'
1/
#227060000000
0!
0'
0/
#227070000000
1!
1'
1/
#227080000000
0!
1"
0'
1(
0/
10
#227090000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#227100000000
0!
0'
0/
#227110000000
1!
1'
1/
#227120000000
0!
0'
0/
#227130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#227140000000
0!
0'
0/
#227150000000
1!
1'
1/
#227160000000
0!
1"
0'
1(
0/
10
#227170000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#227180000000
0!
1$
0'
1+
0/
#227190000000
1!
1'
1/
#227200000000
0!
0'
0/
#227210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#227220000000
0!
0'
0/
#227230000000
1!
1'
1/
#227240000000
0!
0'
0/
#227250000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#227260000000
0!
0'
0/
#227270000000
1!
1'
1/
#227280000000
0!
0'
0/
#227290000000
1!
1'
1/
#227300000000
0!
0'
0/
#227310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#227320000000
0!
0'
0/
#227330000000
1!
1'
1/
#227340000000
0!
0'
0/
#227350000000
1!
1'
1/
#227360000000
0!
0'
0/
#227370000000
1!
1'
1/
#227380000000
0!
0'
0/
#227390000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#227400000000
0!
0'
0/
#227410000000
1!
1'
1/
#227420000000
0!
0'
0/
#227430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#227440000000
0!
0'
0/
#227450000000
1!
1'
1/
#227460000000
0!
0'
0/
#227470000000
#227480000000
1!
1'
1/
#227490000000
0!
0'
0/
#227500000000
1!
1'
1/
#227510000000
0!
1"
0'
1(
0/
10
#227520000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#227530000000
0!
0'
0/
#227540000000
1!
1'
1/
#227550000000
0!
0'
0/
#227560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#227570000000
0!
0'
0/
#227580000000
1!
1'
1/
#227590000000
0!
1"
0'
1(
0/
10
#227600000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#227610000000
0!
1$
0'
1+
0/
#227620000000
1!
1'
1/
#227630000000
0!
0'
0/
#227640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#227650000000
0!
0'
0/
#227660000000
1!
1'
1/
#227670000000
0!
0'
0/
#227680000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#227690000000
0!
0'
0/
#227700000000
1!
1'
1/
#227710000000
0!
0'
0/
#227720000000
1!
1'
1/
#227730000000
0!
0'
0/
#227740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#227750000000
0!
0'
0/
#227760000000
1!
1'
1/
#227770000000
0!
0'
0/
#227780000000
1!
1'
1/
#227790000000
0!
0'
0/
#227800000000
1!
1'
1/
#227810000000
0!
0'
0/
#227820000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#227830000000
0!
0'
0/
#227840000000
1!
1'
1/
#227850000000
0!
0'
0/
#227860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#227870000000
0!
0'
0/
#227880000000
1!
1'
1/
#227890000000
0!
0'
0/
#227900000000
#227910000000
1!
1'
1/
#227920000000
0!
0'
0/
#227930000000
1!
1'
1/
#227940000000
0!
1"
0'
1(
0/
10
#227950000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#227960000000
0!
0'
0/
#227970000000
1!
1'
1/
#227980000000
0!
0'
0/
#227990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#228000000000
0!
0'
0/
#228010000000
1!
1'
1/
#228020000000
0!
1"
0'
1(
0/
10
#228030000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#228040000000
0!
1$
0'
1+
0/
#228050000000
1!
1'
1/
#228060000000
0!
0'
0/
#228070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#228080000000
0!
0'
0/
#228090000000
1!
1'
1/
#228100000000
0!
0'
0/
#228110000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#228120000000
0!
0'
0/
#228130000000
1!
1'
1/
#228140000000
0!
0'
0/
#228150000000
1!
1'
1/
#228160000000
0!
0'
0/
#228170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#228180000000
0!
0'
0/
#228190000000
1!
1'
1/
#228200000000
0!
0'
0/
#228210000000
1!
1'
1/
#228220000000
0!
0'
0/
#228230000000
1!
1'
1/
#228240000000
0!
0'
0/
#228250000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#228260000000
0!
0'
0/
#228270000000
1!
1'
1/
#228280000000
0!
0'
0/
#228290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#228300000000
0!
0'
0/
#228310000000
1!
1'
1/
#228320000000
0!
0'
0/
#228330000000
#228340000000
1!
1'
1/
#228350000000
0!
0'
0/
#228360000000
1!
1'
1/
#228370000000
0!
1"
0'
1(
0/
10
#228380000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#228390000000
0!
0'
0/
#228400000000
1!
1'
1/
#228410000000
0!
0'
0/
#228420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#228430000000
0!
0'
0/
#228440000000
1!
1'
1/
#228450000000
0!
1"
0'
1(
0/
10
#228460000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#228470000000
0!
1$
0'
1+
0/
#228480000000
1!
1'
1/
#228490000000
0!
0'
0/
#228500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#228510000000
0!
0'
0/
#228520000000
1!
1'
1/
#228530000000
0!
0'
0/
#228540000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#228550000000
0!
0'
0/
#228560000000
1!
1'
1/
#228570000000
0!
0'
0/
#228580000000
1!
1'
1/
#228590000000
0!
0'
0/
#228600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#228610000000
0!
0'
0/
#228620000000
1!
1'
1/
#228630000000
0!
0'
0/
#228640000000
1!
1'
1/
#228650000000
0!
0'
0/
#228660000000
1!
1'
1/
#228670000000
0!
0'
0/
#228680000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#228690000000
0!
0'
0/
#228700000000
1!
1'
1/
#228710000000
0!
0'
0/
#228720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#228730000000
0!
0'
0/
#228740000000
1!
1'
1/
#228750000000
0!
0'
0/
#228760000000
#228770000000
1!
1'
1/
#228780000000
0!
0'
0/
#228790000000
1!
1'
1/
#228800000000
0!
1"
0'
1(
0/
10
#228810000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#228820000000
0!
0'
0/
#228830000000
1!
1'
1/
#228840000000
0!
0'
0/
#228850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#228860000000
0!
0'
0/
#228870000000
1!
1'
1/
#228880000000
0!
1"
0'
1(
0/
10
#228890000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#228900000000
0!
1$
0'
1+
0/
#228910000000
1!
1'
1/
#228920000000
0!
0'
0/
#228930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#228940000000
0!
0'
0/
#228950000000
1!
1'
1/
#228960000000
0!
0'
0/
#228970000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#228980000000
0!
0'
0/
#228990000000
1!
1'
1/
#229000000000
0!
0'
0/
#229010000000
1!
1'
1/
#229020000000
0!
0'
0/
#229030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#229040000000
0!
0'
0/
#229050000000
1!
1'
1/
#229060000000
0!
0'
0/
#229070000000
1!
1'
1/
#229080000000
0!
0'
0/
#229090000000
1!
1'
1/
#229100000000
0!
0'
0/
#229110000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#229120000000
0!
0'
0/
#229130000000
1!
1'
1/
#229140000000
0!
0'
0/
#229150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#229160000000
0!
0'
0/
#229170000000
1!
1'
1/
#229180000000
0!
0'
0/
#229190000000
#229200000000
1!
1'
1/
#229210000000
0!
0'
0/
#229220000000
1!
1'
1/
#229230000000
0!
1"
0'
1(
0/
10
#229240000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#229250000000
0!
0'
0/
#229260000000
1!
1'
1/
#229270000000
0!
0'
0/
#229280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#229290000000
0!
0'
0/
#229300000000
1!
1'
1/
#229310000000
0!
1"
0'
1(
0/
10
#229320000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#229330000000
0!
1$
0'
1+
0/
#229340000000
1!
1'
1/
#229350000000
0!
0'
0/
#229360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#229370000000
0!
0'
0/
#229380000000
1!
1'
1/
#229390000000
0!
0'
0/
#229400000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#229410000000
0!
0'
0/
#229420000000
1!
1'
1/
#229430000000
0!
0'
0/
#229440000000
1!
1'
1/
#229450000000
0!
0'
0/
#229460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#229470000000
0!
0'
0/
#229480000000
1!
1'
1/
#229490000000
0!
0'
0/
#229500000000
1!
1'
1/
#229510000000
0!
0'
0/
#229520000000
1!
1'
1/
#229530000000
0!
0'
0/
#229540000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#229550000000
0!
0'
0/
#229560000000
1!
1'
1/
#229570000000
0!
0'
0/
#229580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#229590000000
0!
0'
0/
#229600000000
1!
1'
1/
#229610000000
0!
0'
0/
#229620000000
#229630000000
1!
1'
1/
#229640000000
0!
0'
0/
#229650000000
1!
1'
1/
#229660000000
0!
1"
0'
1(
0/
10
#229670000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#229680000000
0!
0'
0/
#229690000000
1!
1'
1/
#229700000000
0!
0'
0/
#229710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#229720000000
0!
0'
0/
#229730000000
1!
1'
1/
#229740000000
0!
1"
0'
1(
0/
10
#229750000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#229760000000
0!
1$
0'
1+
0/
#229770000000
1!
1'
1/
#229780000000
0!
0'
0/
#229790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#229800000000
0!
0'
0/
#229810000000
1!
1'
1/
#229820000000
0!
0'
0/
#229830000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#229840000000
0!
0'
0/
#229850000000
1!
1'
1/
#229860000000
0!
0'
0/
#229870000000
1!
1'
1/
#229880000000
0!
0'
0/
#229890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#229900000000
0!
0'
0/
#229910000000
1!
1'
1/
#229920000000
0!
0'
0/
#229930000000
1!
1'
1/
#229940000000
0!
0'
0/
#229950000000
1!
1'
1/
#229960000000
0!
0'
0/
#229970000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#229980000000
0!
0'
0/
#229990000000
1!
1'
1/
#230000000000
0!
0'
0/
#230010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#230020000000
0!
0'
0/
#230030000000
1!
1'
1/
#230040000000
0!
0'
0/
#230050000000
#230060000000
1!
1'
1/
#230070000000
0!
0'
0/
#230080000000
1!
1'
1/
#230090000000
0!
1"
0'
1(
0/
10
#230100000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#230110000000
0!
0'
0/
#230120000000
1!
1'
1/
#230130000000
0!
0'
0/
#230140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#230150000000
0!
0'
0/
#230160000000
1!
1'
1/
#230170000000
0!
1"
0'
1(
0/
10
#230180000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#230190000000
0!
1$
0'
1+
0/
#230200000000
1!
1'
1/
#230210000000
0!
0'
0/
#230220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#230230000000
0!
0'
0/
#230240000000
1!
1'
1/
#230250000000
0!
0'
0/
#230260000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#230270000000
0!
0'
0/
#230280000000
1!
1'
1/
#230290000000
0!
0'
0/
#230300000000
1!
1'
1/
#230310000000
0!
0'
0/
#230320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#230330000000
0!
0'
0/
#230340000000
1!
1'
1/
#230350000000
0!
0'
0/
#230360000000
1!
1'
1/
#230370000000
0!
0'
0/
#230380000000
1!
1'
1/
#230390000000
0!
0'
0/
#230400000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#230410000000
0!
0'
0/
#230420000000
1!
1'
1/
#230430000000
0!
0'
0/
#230440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#230450000000
0!
0'
0/
#230460000000
1!
1'
1/
#230470000000
0!
0'
0/
#230480000000
#230490000000
1!
1'
1/
#230500000000
0!
0'
0/
#230510000000
1!
1'
1/
#230520000000
0!
1"
0'
1(
0/
10
#230530000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#230540000000
0!
0'
0/
#230550000000
1!
1'
1/
#230560000000
0!
0'
0/
#230570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#230580000000
0!
0'
0/
#230590000000
1!
1'
1/
#230600000000
0!
1"
0'
1(
0/
10
#230610000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#230620000000
0!
1$
0'
1+
0/
#230630000000
1!
1'
1/
#230640000000
0!
0'
0/
#230650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#230660000000
0!
0'
0/
#230670000000
1!
1'
1/
#230680000000
0!
0'
0/
#230690000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#230700000000
0!
0'
0/
#230710000000
1!
1'
1/
#230720000000
0!
0'
0/
#230730000000
1!
1'
1/
#230740000000
0!
0'
0/
#230750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#230760000000
0!
0'
0/
#230770000000
1!
1'
1/
#230780000000
0!
0'
0/
#230790000000
1!
1'
1/
#230800000000
0!
0'
0/
#230810000000
1!
1'
1/
#230820000000
0!
0'
0/
#230830000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#230840000000
0!
0'
0/
#230850000000
1!
1'
1/
#230860000000
0!
0'
0/
#230870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#230880000000
0!
0'
0/
#230890000000
1!
1'
1/
#230900000000
0!
0'
0/
#230910000000
#230920000000
1!
1'
1/
#230930000000
0!
0'
0/
#230940000000
1!
1'
1/
#230950000000
0!
1"
0'
1(
0/
10
#230960000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#230970000000
0!
0'
0/
#230980000000
1!
1'
1/
#230990000000
0!
0'
0/
#231000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#231010000000
0!
0'
0/
#231020000000
1!
1'
1/
#231030000000
0!
1"
0'
1(
0/
10
#231040000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#231050000000
0!
1$
0'
1+
0/
#231060000000
1!
1'
1/
#231070000000
0!
0'
0/
#231080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#231090000000
0!
0'
0/
#231100000000
1!
1'
1/
#231110000000
0!
0'
0/
#231120000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#231130000000
0!
0'
0/
#231140000000
1!
1'
1/
#231150000000
0!
0'
0/
#231160000000
1!
1'
1/
#231170000000
0!
0'
0/
#231180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#231190000000
0!
0'
0/
#231200000000
1!
1'
1/
#231210000000
0!
0'
0/
#231220000000
1!
1'
1/
#231230000000
0!
0'
0/
#231240000000
1!
1'
1/
#231250000000
0!
0'
0/
#231260000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#231270000000
0!
0'
0/
#231280000000
1!
1'
1/
#231290000000
0!
0'
0/
#231300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#231310000000
0!
0'
0/
#231320000000
1!
1'
1/
#231330000000
0!
0'
0/
#231340000000
#231350000000
1!
1'
1/
#231360000000
0!
0'
0/
#231370000000
1!
1'
1/
#231380000000
0!
1"
0'
1(
0/
10
#231390000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#231400000000
0!
0'
0/
#231410000000
1!
1'
1/
#231420000000
0!
0'
0/
#231430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#231440000000
0!
0'
0/
#231450000000
1!
1'
1/
#231460000000
0!
1"
0'
1(
0/
10
#231470000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#231480000000
0!
1$
0'
1+
0/
#231490000000
1!
1'
1/
#231500000000
0!
0'
0/
#231510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#231520000000
0!
0'
0/
#231530000000
1!
1'
1/
#231540000000
0!
0'
0/
#231550000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#231560000000
0!
0'
0/
#231570000000
1!
1'
1/
#231580000000
0!
0'
0/
#231590000000
1!
1'
1/
#231600000000
0!
0'
0/
#231610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#231620000000
0!
0'
0/
#231630000000
1!
1'
1/
#231640000000
0!
0'
0/
#231650000000
1!
1'
1/
#231660000000
0!
0'
0/
#231670000000
1!
1'
1/
#231680000000
0!
0'
0/
#231690000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#231700000000
0!
0'
0/
#231710000000
1!
1'
1/
#231720000000
0!
0'
0/
#231730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#231740000000
0!
0'
0/
#231750000000
1!
1'
1/
#231760000000
0!
0'
0/
#231770000000
#231780000000
1!
1'
1/
#231790000000
0!
0'
0/
#231800000000
1!
1'
1/
#231810000000
0!
1"
0'
1(
0/
10
#231820000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#231830000000
0!
0'
0/
#231840000000
1!
1'
1/
#231850000000
0!
0'
0/
#231860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#231870000000
0!
0'
0/
#231880000000
1!
1'
1/
#231890000000
0!
1"
0'
1(
0/
10
#231900000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#231910000000
0!
1$
0'
1+
0/
#231920000000
1!
1'
1/
#231930000000
0!
0'
0/
#231940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#231950000000
0!
0'
0/
#231960000000
1!
1'
1/
#231970000000
0!
0'
0/
#231980000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#231990000000
0!
0'
0/
#232000000000
1!
1'
1/
#232010000000
0!
0'
0/
#232020000000
1!
1'
1/
#232030000000
0!
0'
0/
#232040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#232050000000
0!
0'
0/
#232060000000
1!
1'
1/
#232070000000
0!
0'
0/
#232080000000
1!
1'
1/
#232090000000
0!
0'
0/
#232100000000
1!
1'
1/
#232110000000
0!
0'
0/
#232120000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#232130000000
0!
0'
0/
#232140000000
1!
1'
1/
#232150000000
0!
0'
0/
#232160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#232170000000
0!
0'
0/
#232180000000
1!
1'
1/
#232190000000
0!
0'
0/
#232200000000
#232210000000
1!
1'
1/
#232220000000
0!
0'
0/
#232230000000
1!
1'
1/
#232240000000
0!
1"
0'
1(
0/
10
#232250000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#232260000000
0!
0'
0/
#232270000000
1!
1'
1/
#232280000000
0!
0'
0/
#232290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#232300000000
0!
0'
0/
#232310000000
1!
1'
1/
#232320000000
0!
1"
0'
1(
0/
10
#232330000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#232340000000
0!
1$
0'
1+
0/
#232350000000
1!
1'
1/
#232360000000
0!
0'
0/
#232370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#232380000000
0!
0'
0/
#232390000000
1!
1'
1/
#232400000000
0!
0'
0/
#232410000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#232420000000
0!
0'
0/
#232430000000
1!
1'
1/
#232440000000
0!
0'
0/
#232450000000
1!
1'
1/
#232460000000
0!
0'
0/
#232470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#232480000000
0!
0'
0/
#232490000000
1!
1'
1/
#232500000000
0!
0'
0/
#232510000000
1!
1'
1/
#232520000000
0!
0'
0/
#232530000000
1!
1'
1/
#232540000000
0!
0'
0/
#232550000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#232560000000
0!
0'
0/
#232570000000
1!
1'
1/
#232580000000
0!
0'
0/
#232590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#232600000000
0!
0'
0/
#232610000000
1!
1'
1/
#232620000000
0!
0'
0/
#232630000000
#232640000000
1!
1'
1/
#232650000000
0!
0'
0/
#232660000000
1!
1'
1/
#232670000000
0!
1"
0'
1(
0/
10
#232680000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#232690000000
0!
0'
0/
#232700000000
1!
1'
1/
#232710000000
0!
0'
0/
#232720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#232730000000
0!
0'
0/
#232740000000
1!
1'
1/
#232750000000
0!
1"
0'
1(
0/
10
#232760000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#232770000000
0!
1$
0'
1+
0/
#232780000000
1!
1'
1/
#232790000000
0!
0'
0/
#232800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#232810000000
0!
0'
0/
#232820000000
1!
1'
1/
#232830000000
0!
0'
0/
#232840000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#232850000000
0!
0'
0/
#232860000000
1!
1'
1/
#232870000000
0!
0'
0/
#232880000000
1!
1'
1/
#232890000000
0!
0'
0/
#232900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#232910000000
0!
0'
0/
#232920000000
1!
1'
1/
#232930000000
0!
0'
0/
#232940000000
1!
1'
1/
#232950000000
0!
0'
0/
#232960000000
1!
1'
1/
#232970000000
0!
0'
0/
#232980000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#232990000000
0!
0'
0/
#233000000000
1!
1'
1/
#233010000000
0!
0'
0/
#233020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#233030000000
0!
0'
0/
#233040000000
1!
1'
1/
#233050000000
0!
0'
0/
#233060000000
#233070000000
1!
1'
1/
#233080000000
0!
0'
0/
#233090000000
1!
1'
1/
#233100000000
0!
1"
0'
1(
0/
10
#233110000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#233120000000
0!
0'
0/
#233130000000
1!
1'
1/
#233140000000
0!
0'
0/
#233150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#233160000000
0!
0'
0/
#233170000000
1!
1'
1/
#233180000000
0!
1"
0'
1(
0/
10
#233190000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#233200000000
0!
1$
0'
1+
0/
#233210000000
1!
1'
1/
#233220000000
0!
0'
0/
#233230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#233240000000
0!
0'
0/
#233250000000
1!
1'
1/
#233260000000
0!
0'
0/
#233270000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#233280000000
0!
0'
0/
#233290000000
1!
1'
1/
#233300000000
0!
0'
0/
#233310000000
1!
1'
1/
#233320000000
0!
0'
0/
#233330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#233340000000
0!
0'
0/
#233350000000
1!
1'
1/
#233360000000
0!
0'
0/
#233370000000
1!
1'
1/
#233380000000
0!
0'
0/
#233390000000
1!
1'
1/
#233400000000
0!
0'
0/
#233410000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#233420000000
0!
0'
0/
#233430000000
1!
1'
1/
#233440000000
0!
0'
0/
#233450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#233460000000
0!
0'
0/
#233470000000
1!
1'
1/
#233480000000
0!
0'
0/
#233490000000
#233500000000
1!
1'
1/
#233510000000
0!
0'
0/
#233520000000
1!
1'
1/
#233530000000
0!
1"
0'
1(
0/
10
#233540000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#233550000000
0!
0'
0/
#233560000000
1!
1'
1/
#233570000000
0!
0'
0/
#233580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#233590000000
0!
0'
0/
#233600000000
1!
1'
1/
#233610000000
0!
1"
0'
1(
0/
10
#233620000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#233630000000
0!
1$
0'
1+
0/
#233640000000
1!
1'
1/
#233650000000
0!
0'
0/
#233660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#233670000000
0!
0'
0/
#233680000000
1!
1'
1/
#233690000000
0!
0'
0/
#233700000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#233710000000
0!
0'
0/
#233720000000
1!
1'
1/
#233730000000
0!
0'
0/
#233740000000
1!
1'
1/
#233750000000
0!
0'
0/
#233760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#233770000000
0!
0'
0/
#233780000000
1!
1'
1/
#233790000000
0!
0'
0/
#233800000000
1!
1'
1/
#233810000000
0!
0'
0/
#233820000000
1!
1'
1/
#233830000000
0!
0'
0/
#233840000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#233850000000
0!
0'
0/
#233860000000
1!
1'
1/
#233870000000
0!
0'
0/
#233880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#233890000000
0!
0'
0/
#233900000000
1!
1'
1/
#233910000000
0!
0'
0/
#233920000000
#233930000000
1!
1'
1/
#233940000000
0!
0'
0/
#233950000000
1!
1'
1/
#233960000000
0!
1"
0'
1(
0/
10
#233970000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#233980000000
0!
0'
0/
#233990000000
1!
1'
1/
#234000000000
0!
0'
0/
#234010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#234020000000
0!
0'
0/
#234030000000
1!
1'
1/
#234040000000
0!
1"
0'
1(
0/
10
#234050000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#234060000000
0!
1$
0'
1+
0/
#234070000000
1!
1'
1/
#234080000000
0!
0'
0/
#234090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#234100000000
0!
0'
0/
#234110000000
1!
1'
1/
#234120000000
0!
0'
0/
#234130000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#234140000000
0!
0'
0/
#234150000000
1!
1'
1/
#234160000000
0!
0'
0/
#234170000000
1!
1'
1/
#234180000000
0!
0'
0/
#234190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#234200000000
0!
0'
0/
#234210000000
1!
1'
1/
#234220000000
0!
0'
0/
#234230000000
1!
1'
1/
#234240000000
0!
0'
0/
#234250000000
1!
1'
1/
#234260000000
0!
0'
0/
#234270000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#234280000000
0!
0'
0/
#234290000000
1!
1'
1/
#234300000000
0!
0'
0/
#234310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#234320000000
0!
0'
0/
#234330000000
1!
1'
1/
#234340000000
0!
0'
0/
#234350000000
#234360000000
1!
1'
1/
#234370000000
0!
0'
0/
#234380000000
1!
1'
1/
#234390000000
0!
1"
0'
1(
0/
10
#234400000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#234410000000
0!
0'
0/
#234420000000
1!
1'
1/
#234430000000
0!
0'
0/
#234440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#234450000000
0!
0'
0/
#234460000000
1!
1'
1/
#234470000000
0!
1"
0'
1(
0/
10
#234480000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#234490000000
0!
1$
0'
1+
0/
#234500000000
1!
1'
1/
#234510000000
0!
0'
0/
#234520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#234530000000
0!
0'
0/
#234540000000
1!
1'
1/
#234550000000
0!
0'
0/
#234560000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#234570000000
0!
0'
0/
#234580000000
1!
1'
1/
#234590000000
0!
0'
0/
#234600000000
1!
1'
1/
#234610000000
0!
0'
0/
#234620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#234630000000
0!
0'
0/
#234640000000
1!
1'
1/
#234650000000
0!
0'
0/
#234660000000
1!
1'
1/
#234670000000
0!
0'
0/
#234680000000
1!
1'
1/
#234690000000
0!
0'
0/
#234700000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#234710000000
0!
0'
0/
#234720000000
1!
1'
1/
#234730000000
0!
0'
0/
#234740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#234750000000
0!
0'
0/
#234760000000
1!
1'
1/
#234770000000
0!
0'
0/
#234780000000
#234790000000
1!
1'
1/
#234800000000
0!
0'
0/
#234810000000
1!
1'
1/
#234820000000
0!
1"
0'
1(
0/
10
#234830000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#234840000000
0!
0'
0/
#234850000000
1!
1'
1/
#234860000000
0!
0'
0/
#234870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#234880000000
0!
0'
0/
#234890000000
1!
1'
1/
#234900000000
0!
1"
0'
1(
0/
10
#234910000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#234920000000
0!
1$
0'
1+
0/
#234930000000
1!
1'
1/
#234940000000
0!
0'
0/
#234950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#234960000000
0!
0'
0/
#234970000000
1!
1'
1/
#234980000000
0!
0'
0/
#234990000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#235000000000
0!
0'
0/
#235010000000
1!
1'
1/
#235020000000
0!
0'
0/
#235030000000
1!
1'
1/
#235040000000
0!
0'
0/
#235050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#235060000000
0!
0'
0/
#235070000000
1!
1'
1/
#235080000000
0!
0'
0/
#235090000000
1!
1'
1/
#235100000000
0!
0'
0/
#235110000000
1!
1'
1/
#235120000000
0!
0'
0/
#235130000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#235140000000
0!
0'
0/
#235150000000
1!
1'
1/
#235160000000
0!
0'
0/
#235170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#235180000000
0!
0'
0/
#235190000000
1!
1'
1/
#235200000000
0!
0'
0/
#235210000000
#235220000000
1!
1'
1/
#235230000000
0!
0'
0/
#235240000000
1!
1'
1/
#235250000000
0!
1"
0'
1(
0/
10
#235260000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#235270000000
0!
0'
0/
#235280000000
1!
1'
1/
#235290000000
0!
0'
0/
#235300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#235310000000
0!
0'
0/
#235320000000
1!
1'
1/
#235330000000
0!
1"
0'
1(
0/
10
#235340000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#235350000000
0!
1$
0'
1+
0/
#235360000000
1!
1'
1/
#235370000000
0!
0'
0/
#235380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#235390000000
0!
0'
0/
#235400000000
1!
1'
1/
#235410000000
0!
0'
0/
#235420000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#235430000000
0!
0'
0/
#235440000000
1!
1'
1/
#235450000000
0!
0'
0/
#235460000000
1!
1'
1/
#235470000000
0!
0'
0/
#235480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#235490000000
0!
0'
0/
#235500000000
1!
1'
1/
#235510000000
0!
0'
0/
#235520000000
1!
1'
1/
#235530000000
0!
0'
0/
#235540000000
1!
1'
1/
#235550000000
0!
0'
0/
#235560000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#235570000000
0!
0'
0/
#235580000000
1!
1'
1/
#235590000000
0!
0'
0/
#235600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#235610000000
0!
0'
0/
#235620000000
1!
1'
1/
#235630000000
0!
0'
0/
#235640000000
#235650000000
1!
1'
1/
#235660000000
0!
0'
0/
#235670000000
1!
1'
1/
#235680000000
0!
1"
0'
1(
0/
10
#235690000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#235700000000
0!
0'
0/
#235710000000
1!
1'
1/
#235720000000
0!
0'
0/
#235730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#235740000000
0!
0'
0/
#235750000000
1!
1'
1/
#235760000000
0!
1"
0'
1(
0/
10
#235770000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#235780000000
0!
1$
0'
1+
0/
#235790000000
1!
1'
1/
#235800000000
0!
0'
0/
#235810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#235820000000
0!
0'
0/
#235830000000
1!
1'
1/
#235840000000
0!
0'
0/
#235850000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#235860000000
0!
0'
0/
#235870000000
1!
1'
1/
#235880000000
0!
0'
0/
#235890000000
1!
1'
1/
#235900000000
0!
0'
0/
#235910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#235920000000
0!
0'
0/
#235930000000
1!
1'
1/
#235940000000
0!
0'
0/
#235950000000
1!
1'
1/
#235960000000
0!
0'
0/
#235970000000
1!
1'
1/
#235980000000
0!
0'
0/
#235990000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#236000000000
0!
0'
0/
#236010000000
1!
1'
1/
#236020000000
0!
0'
0/
#236030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#236040000000
0!
0'
0/
#236050000000
1!
1'
1/
#236060000000
0!
0'
0/
#236070000000
#236080000000
1!
1'
1/
#236090000000
0!
0'
0/
#236100000000
1!
1'
1/
#236110000000
0!
1"
0'
1(
0/
10
#236120000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#236130000000
0!
0'
0/
#236140000000
1!
1'
1/
#236150000000
0!
0'
0/
#236160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#236170000000
0!
0'
0/
#236180000000
1!
1'
1/
#236190000000
0!
1"
0'
1(
0/
10
#236200000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#236210000000
0!
1$
0'
1+
0/
#236220000000
1!
1'
1/
#236230000000
0!
0'
0/
#236240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#236250000000
0!
0'
0/
#236260000000
1!
1'
1/
#236270000000
0!
0'
0/
#236280000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#236290000000
0!
0'
0/
#236300000000
1!
1'
1/
#236310000000
0!
0'
0/
#236320000000
1!
1'
1/
#236330000000
0!
0'
0/
#236340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#236350000000
0!
0'
0/
#236360000000
1!
1'
1/
#236370000000
0!
0'
0/
#236380000000
1!
1'
1/
#236390000000
0!
0'
0/
#236400000000
1!
1'
1/
#236410000000
0!
0'
0/
#236420000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#236430000000
0!
0'
0/
#236440000000
1!
1'
1/
#236450000000
0!
0'
0/
#236460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#236470000000
0!
0'
0/
#236480000000
1!
1'
1/
#236490000000
0!
0'
0/
#236500000000
#236510000000
1!
1'
1/
#236520000000
0!
0'
0/
#236530000000
1!
1'
1/
#236540000000
0!
1"
0'
1(
0/
10
#236550000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#236560000000
0!
0'
0/
#236570000000
1!
1'
1/
#236580000000
0!
0'
0/
#236590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#236600000000
0!
0'
0/
#236610000000
1!
1'
1/
#236620000000
0!
1"
0'
1(
0/
10
#236630000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#236640000000
0!
1$
0'
1+
0/
#236650000000
1!
1'
1/
#236660000000
0!
0'
0/
#236670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#236680000000
0!
0'
0/
#236690000000
1!
1'
1/
#236700000000
0!
0'
0/
#236710000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#236720000000
0!
0'
0/
#236730000000
1!
1'
1/
#236740000000
0!
0'
0/
#236750000000
1!
1'
1/
#236760000000
0!
0'
0/
#236770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#236780000000
0!
0'
0/
#236790000000
1!
1'
1/
#236800000000
0!
0'
0/
#236810000000
1!
1'
1/
#236820000000
0!
0'
0/
#236830000000
1!
1'
1/
#236840000000
0!
0'
0/
#236850000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#236860000000
0!
0'
0/
#236870000000
1!
1'
1/
#236880000000
0!
0'
0/
#236890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#236900000000
0!
0'
0/
#236910000000
1!
1'
1/
#236920000000
0!
0'
0/
#236930000000
#236940000000
1!
1'
1/
#236950000000
0!
0'
0/
#236960000000
1!
1'
1/
#236970000000
0!
1"
0'
1(
0/
10
#236980000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#236990000000
0!
0'
0/
#237000000000
1!
1'
1/
#237010000000
0!
0'
0/
#237020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#237030000000
0!
0'
0/
#237040000000
1!
1'
1/
#237050000000
0!
1"
0'
1(
0/
10
#237060000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#237070000000
0!
1$
0'
1+
0/
#237080000000
1!
1'
1/
#237090000000
0!
0'
0/
#237100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#237110000000
0!
0'
0/
#237120000000
1!
1'
1/
#237130000000
0!
0'
0/
#237140000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#237150000000
0!
0'
0/
#237160000000
1!
1'
1/
#237170000000
0!
0'
0/
#237180000000
1!
1'
1/
#237190000000
0!
0'
0/
#237200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#237210000000
0!
0'
0/
#237220000000
1!
1'
1/
#237230000000
0!
0'
0/
#237240000000
1!
1'
1/
#237250000000
0!
0'
0/
#237260000000
1!
1'
1/
#237270000000
0!
0'
0/
#237280000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#237290000000
0!
0'
0/
#237300000000
1!
1'
1/
#237310000000
0!
0'
0/
#237320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#237330000000
0!
0'
0/
#237340000000
1!
1'
1/
#237350000000
0!
0'
0/
#237360000000
#237370000000
1!
1'
1/
#237380000000
0!
0'
0/
#237390000000
1!
1'
1/
#237400000000
0!
1"
0'
1(
0/
10
#237410000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#237420000000
0!
0'
0/
#237430000000
1!
1'
1/
#237440000000
0!
0'
0/
#237450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#237460000000
0!
0'
0/
#237470000000
1!
1'
1/
#237480000000
0!
1"
0'
1(
0/
10
#237490000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#237500000000
0!
1$
0'
1+
0/
#237510000000
1!
1'
1/
#237520000000
0!
0'
0/
#237530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#237540000000
0!
0'
0/
#237550000000
1!
1'
1/
#237560000000
0!
0'
0/
#237570000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#237580000000
0!
0'
0/
#237590000000
1!
1'
1/
#237600000000
0!
0'
0/
#237610000000
1!
1'
1/
#237620000000
0!
0'
0/
#237630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#237640000000
0!
0'
0/
#237650000000
1!
1'
1/
#237660000000
0!
0'
0/
#237670000000
1!
1'
1/
#237680000000
0!
0'
0/
#237690000000
1!
1'
1/
#237700000000
0!
0'
0/
#237710000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#237720000000
0!
0'
0/
#237730000000
1!
1'
1/
#237740000000
0!
0'
0/
#237750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#237760000000
0!
0'
0/
#237770000000
1!
1'
1/
#237780000000
0!
0'
0/
#237790000000
#237800000000
1!
1'
1/
#237810000000
0!
0'
0/
#237820000000
1!
1'
1/
#237830000000
0!
1"
0'
1(
0/
10
#237840000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#237850000000
0!
0'
0/
#237860000000
1!
1'
1/
#237870000000
0!
0'
0/
#237880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#237890000000
0!
0'
0/
#237900000000
1!
1'
1/
#237910000000
0!
1"
0'
1(
0/
10
#237920000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#237930000000
0!
1$
0'
1+
0/
#237940000000
1!
1'
1/
#237950000000
0!
0'
0/
#237960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#237970000000
0!
0'
0/
#237980000000
1!
1'
1/
#237990000000
0!
0'
0/
#238000000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#238010000000
0!
0'
0/
#238020000000
1!
1'
1/
#238030000000
0!
0'
0/
#238040000000
1!
1'
1/
#238050000000
0!
0'
0/
#238060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#238070000000
0!
0'
0/
#238080000000
1!
1'
1/
#238090000000
0!
0'
0/
#238100000000
1!
1'
1/
#238110000000
0!
0'
0/
#238120000000
1!
1'
1/
#238130000000
0!
0'
0/
#238140000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#238150000000
0!
0'
0/
#238160000000
1!
1'
1/
#238170000000
0!
0'
0/
#238180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#238190000000
0!
0'
0/
#238200000000
1!
1'
1/
#238210000000
0!
0'
0/
#238220000000
#238230000000
1!
1'
1/
#238240000000
0!
0'
0/
#238250000000
1!
1'
1/
#238260000000
0!
1"
0'
1(
0/
10
#238270000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#238280000000
0!
0'
0/
#238290000000
1!
1'
1/
#238300000000
0!
0'
0/
#238310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#238320000000
0!
0'
0/
#238330000000
1!
1'
1/
#238340000000
0!
1"
0'
1(
0/
10
#238350000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#238360000000
0!
1$
0'
1+
0/
#238370000000
1!
1'
1/
#238380000000
0!
0'
0/
#238390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#238400000000
0!
0'
0/
#238410000000
1!
1'
1/
#238420000000
0!
0'
0/
#238430000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#238440000000
0!
0'
0/
#238450000000
1!
1'
1/
#238460000000
0!
0'
0/
#238470000000
1!
1'
1/
#238480000000
0!
0'
0/
#238490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#238500000000
0!
0'
0/
#238510000000
1!
1'
1/
#238520000000
0!
0'
0/
#238530000000
1!
1'
1/
#238540000000
0!
0'
0/
#238550000000
1!
1'
1/
#238560000000
0!
0'
0/
#238570000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#238580000000
0!
0'
0/
#238590000000
1!
1'
1/
#238600000000
0!
0'
0/
#238610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#238620000000
0!
0'
0/
#238630000000
1!
1'
1/
#238640000000
0!
0'
0/
#238650000000
#238660000000
1!
1'
1/
#238670000000
0!
0'
0/
#238680000000
1!
1'
1/
#238690000000
0!
1"
0'
1(
0/
10
#238700000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#238710000000
0!
0'
0/
#238720000000
1!
1'
1/
#238730000000
0!
0'
0/
#238740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#238750000000
0!
0'
0/
#238760000000
1!
1'
1/
#238770000000
0!
1"
0'
1(
0/
10
#238780000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#238790000000
0!
1$
0'
1+
0/
#238800000000
1!
1'
1/
#238810000000
0!
0'
0/
#238820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#238830000000
0!
0'
0/
#238840000000
1!
1'
1/
#238850000000
0!
0'
0/
#238860000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#238870000000
0!
0'
0/
#238880000000
1!
1'
1/
#238890000000
0!
0'
0/
#238900000000
1!
1'
1/
#238910000000
0!
0'
0/
#238920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#238930000000
0!
0'
0/
#238940000000
1!
1'
1/
#238950000000
0!
0'
0/
#238960000000
1!
1'
1/
#238970000000
0!
0'
0/
#238980000000
1!
1'
1/
#238990000000
0!
0'
0/
#239000000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#239010000000
0!
0'
0/
#239020000000
1!
1'
1/
#239030000000
0!
0'
0/
#239040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#239050000000
0!
0'
0/
#239060000000
1!
1'
1/
#239070000000
0!
0'
0/
#239080000000
#239090000000
1!
1'
1/
#239100000000
0!
0'
0/
#239110000000
1!
1'
1/
#239120000000
0!
1"
0'
1(
0/
10
#239130000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#239140000000
0!
0'
0/
#239150000000
1!
1'
1/
#239160000000
0!
0'
0/
#239170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#239180000000
0!
0'
0/
#239190000000
1!
1'
1/
#239200000000
0!
1"
0'
1(
0/
10
#239210000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#239220000000
0!
1$
0'
1+
0/
#239230000000
1!
1'
1/
#239240000000
0!
0'
0/
#239250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#239260000000
0!
0'
0/
#239270000000
1!
1'
1/
#239280000000
0!
0'
0/
#239290000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#239300000000
0!
0'
0/
#239310000000
1!
1'
1/
#239320000000
0!
0'
0/
#239330000000
1!
1'
1/
#239340000000
0!
0'
0/
#239350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#239360000000
0!
0'
0/
#239370000000
1!
1'
1/
#239380000000
0!
0'
0/
#239390000000
1!
1'
1/
#239400000000
0!
0'
0/
#239410000000
1!
1'
1/
#239420000000
0!
0'
0/
#239430000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#239440000000
0!
0'
0/
#239450000000
1!
1'
1/
#239460000000
0!
0'
0/
#239470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#239480000000
0!
0'
0/
#239490000000
1!
1'
1/
#239500000000
0!
0'
0/
#239510000000
#239520000000
1!
1'
1/
#239530000000
0!
0'
0/
#239540000000
1!
1'
1/
#239550000000
0!
1"
0'
1(
0/
10
#239560000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#239570000000
0!
0'
0/
#239580000000
1!
1'
1/
#239590000000
0!
0'
0/
#239600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#239610000000
0!
0'
0/
#239620000000
1!
1'
1/
#239630000000
0!
1"
0'
1(
0/
10
#239640000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#239650000000
0!
1$
0'
1+
0/
#239660000000
1!
1'
1/
#239670000000
0!
0'
0/
#239680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#239690000000
0!
0'
0/
#239700000000
1!
1'
1/
#239710000000
0!
0'
0/
#239720000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#239730000000
0!
0'
0/
#239740000000
1!
1'
1/
#239750000000
0!
0'
0/
#239760000000
1!
1'
1/
#239770000000
0!
0'
0/
#239780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#239790000000
0!
0'
0/
#239800000000
1!
1'
1/
#239810000000
0!
0'
0/
#239820000000
1!
1'
1/
#239830000000
0!
0'
0/
#239840000000
1!
1'
1/
#239850000000
0!
0'
0/
#239860000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#239870000000
0!
0'
0/
#239880000000
1!
1'
1/
#239890000000
0!
0'
0/
#239900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#239910000000
0!
0'
0/
#239920000000
1!
1'
1/
#239930000000
0!
0'
0/
#239940000000
#239950000000
1!
1'
1/
#239960000000
0!
0'
0/
#239970000000
1!
1'
1/
#239980000000
0!
1"
0'
1(
0/
10
#239990000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#240000000000
0!
0'
0/
#240010000000
1!
1'
1/
#240020000000
0!
0'
0/
#240030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#240040000000
0!
0'
0/
#240050000000
1!
1'
1/
#240060000000
0!
1"
0'
1(
0/
10
#240070000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#240080000000
0!
1$
0'
1+
0/
#240090000000
1!
1'
1/
#240100000000
0!
0'
0/
#240110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#240120000000
0!
0'
0/
#240130000000
1!
1'
1/
#240140000000
0!
0'
0/
#240150000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#240160000000
0!
0'
0/
#240170000000
1!
1'
1/
#240180000000
0!
0'
0/
#240190000000
1!
1'
1/
#240200000000
0!
0'
0/
#240210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#240220000000
0!
0'
0/
#240230000000
1!
1'
1/
#240240000000
0!
0'
0/
#240250000000
1!
1'
1/
#240260000000
0!
0'
0/
#240270000000
1!
1'
1/
#240280000000
0!
0'
0/
#240290000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#240300000000
0!
0'
0/
#240310000000
1!
1'
1/
#240320000000
0!
0'
0/
#240330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#240340000000
0!
0'
0/
#240350000000
1!
1'
1/
#240360000000
0!
0'
0/
#240370000000
#240380000000
1!
1'
1/
#240390000000
0!
0'
0/
#240400000000
1!
1'
1/
#240410000000
0!
1"
0'
1(
0/
10
#240420000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#240430000000
0!
0'
0/
#240440000000
1!
1'
1/
#240450000000
0!
0'
0/
#240460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#240470000000
0!
0'
0/
#240480000000
1!
1'
1/
#240490000000
0!
1"
0'
1(
0/
10
#240500000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#240510000000
0!
1$
0'
1+
0/
#240520000000
1!
1'
1/
#240530000000
0!
0'
0/
#240540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#240550000000
0!
0'
0/
#240560000000
1!
1'
1/
#240570000000
0!
0'
0/
#240580000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#240590000000
0!
0'
0/
#240600000000
1!
1'
1/
#240610000000
0!
0'
0/
#240620000000
1!
1'
1/
#240630000000
0!
0'
0/
#240640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#240650000000
0!
0'
0/
#240660000000
1!
1'
1/
#240670000000
0!
0'
0/
#240680000000
1!
1'
1/
#240690000000
0!
0'
0/
#240700000000
1!
1'
1/
#240710000000
0!
0'
0/
#240720000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#240730000000
0!
0'
0/
#240740000000
1!
1'
1/
#240750000000
0!
0'
0/
#240760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#240770000000
0!
0'
0/
#240780000000
1!
1'
1/
#240790000000
0!
0'
0/
#240800000000
#240810000000
1!
1'
1/
#240820000000
0!
0'
0/
#240830000000
1!
1'
1/
#240840000000
0!
1"
0'
1(
0/
10
#240850000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#240860000000
0!
0'
0/
#240870000000
1!
1'
1/
#240880000000
0!
0'
0/
#240890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#240900000000
0!
0'
0/
#240910000000
1!
1'
1/
#240920000000
0!
1"
0'
1(
0/
10
#240930000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#240940000000
0!
1$
0'
1+
0/
#240950000000
1!
1'
1/
#240960000000
0!
0'
0/
#240970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#240980000000
0!
0'
0/
#240990000000
1!
1'
1/
#241000000000
0!
0'
0/
#241010000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#241020000000
0!
0'
0/
#241030000000
1!
1'
1/
#241040000000
0!
0'
0/
#241050000000
1!
1'
1/
#241060000000
0!
0'
0/
#241070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#241080000000
0!
0'
0/
#241090000000
1!
1'
1/
#241100000000
0!
0'
0/
#241110000000
1!
1'
1/
#241120000000
0!
0'
0/
#241130000000
1!
1'
1/
#241140000000
0!
0'
0/
#241150000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#241160000000
0!
0'
0/
#241170000000
1!
1'
1/
#241180000000
0!
0'
0/
#241190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#241200000000
0!
0'
0/
#241210000000
1!
1'
1/
#241220000000
0!
0'
0/
#241230000000
#241240000000
1!
1'
1/
#241250000000
0!
0'
0/
#241260000000
1!
1'
1/
#241270000000
0!
1"
0'
1(
0/
10
#241280000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#241290000000
0!
0'
0/
#241300000000
1!
1'
1/
#241310000000
0!
0'
0/
#241320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#241330000000
0!
0'
0/
#241340000000
1!
1'
1/
#241350000000
0!
1"
0'
1(
0/
10
#241360000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#241370000000
0!
1$
0'
1+
0/
#241380000000
1!
1'
1/
#241390000000
0!
0'
0/
#241400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#241410000000
0!
0'
0/
#241420000000
1!
1'
1/
#241430000000
0!
0'
0/
#241440000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#241450000000
0!
0'
0/
#241460000000
1!
1'
1/
#241470000000
0!
0'
0/
#241480000000
1!
1'
1/
#241490000000
0!
0'
0/
#241500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#241510000000
0!
0'
0/
#241520000000
1!
1'
1/
#241530000000
0!
0'
0/
#241540000000
1!
1'
1/
#241550000000
0!
0'
0/
#241560000000
1!
1'
1/
#241570000000
0!
0'
0/
#241580000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#241590000000
0!
0'
0/
#241600000000
1!
1'
1/
#241610000000
0!
0'
0/
#241620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#241630000000
0!
0'
0/
#241640000000
1!
1'
1/
#241650000000
0!
0'
0/
#241660000000
#241670000000
1!
1'
1/
#241680000000
0!
0'
0/
#241690000000
1!
1'
1/
#241700000000
0!
1"
0'
1(
0/
10
#241710000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#241720000000
0!
0'
0/
#241730000000
1!
1'
1/
#241740000000
0!
0'
0/
#241750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#241760000000
0!
0'
0/
#241770000000
1!
1'
1/
#241780000000
0!
1"
0'
1(
0/
10
#241790000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#241800000000
0!
1$
0'
1+
0/
#241810000000
1!
1'
1/
#241820000000
0!
0'
0/
#241830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#241840000000
0!
0'
0/
#241850000000
1!
1'
1/
#241860000000
0!
0'
0/
#241870000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#241880000000
0!
0'
0/
#241890000000
1!
1'
1/
#241900000000
0!
0'
0/
#241910000000
1!
1'
1/
#241920000000
0!
0'
0/
#241930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#241940000000
0!
0'
0/
#241950000000
1!
1'
1/
#241960000000
0!
0'
0/
#241970000000
1!
1'
1/
#241980000000
0!
0'
0/
#241990000000
1!
1'
1/
#242000000000
0!
0'
0/
#242010000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#242020000000
0!
0'
0/
#242030000000
1!
1'
1/
#242040000000
0!
0'
0/
#242050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#242060000000
0!
0'
0/
#242070000000
1!
1'
1/
#242080000000
0!
0'
0/
#242090000000
#242100000000
1!
1'
1/
#242110000000
0!
0'
0/
#242120000000
1!
1'
1/
#242130000000
0!
1"
0'
1(
0/
10
#242140000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#242150000000
0!
0'
0/
#242160000000
1!
1'
1/
#242170000000
0!
0'
0/
#242180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#242190000000
0!
0'
0/
#242200000000
1!
1'
1/
#242210000000
0!
1"
0'
1(
0/
10
#242220000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#242230000000
0!
1$
0'
1+
0/
#242240000000
1!
1'
1/
#242250000000
0!
0'
0/
#242260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#242270000000
0!
0'
0/
#242280000000
1!
1'
1/
#242290000000
0!
0'
0/
#242300000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#242310000000
0!
0'
0/
#242320000000
1!
1'
1/
#242330000000
0!
0'
0/
#242340000000
1!
1'
1/
#242350000000
0!
0'
0/
#242360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#242370000000
0!
0'
0/
#242380000000
1!
1'
1/
#242390000000
0!
0'
0/
#242400000000
1!
1'
1/
#242410000000
0!
0'
0/
#242420000000
1!
1'
1/
#242430000000
0!
0'
0/
#242440000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#242450000000
0!
0'
0/
#242460000000
1!
1'
1/
#242470000000
0!
0'
0/
#242480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#242490000000
0!
0'
0/
#242500000000
1!
1'
1/
#242510000000
0!
0'
0/
#242520000000
#242530000000
1!
1'
1/
#242540000000
0!
0'
0/
#242550000000
1!
1'
1/
#242560000000
0!
1"
0'
1(
0/
10
#242570000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#242580000000
0!
0'
0/
#242590000000
1!
1'
1/
#242600000000
0!
0'
0/
#242610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#242620000000
0!
0'
0/
#242630000000
1!
1'
1/
#242640000000
0!
1"
0'
1(
0/
10
#242650000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#242660000000
0!
1$
0'
1+
0/
#242670000000
1!
1'
1/
#242680000000
0!
0'
0/
#242690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#242700000000
0!
0'
0/
#242710000000
1!
1'
1/
#242720000000
0!
0'
0/
#242730000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#242740000000
0!
0'
0/
#242750000000
1!
1'
1/
#242760000000
0!
0'
0/
#242770000000
1!
1'
1/
#242780000000
0!
0'
0/
#242790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#242800000000
0!
0'
0/
#242810000000
1!
1'
1/
#242820000000
0!
0'
0/
#242830000000
1!
1'
1/
#242840000000
0!
0'
0/
#242850000000
1!
1'
1/
#242860000000
0!
0'
0/
#242870000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#242880000000
0!
0'
0/
#242890000000
1!
1'
1/
#242900000000
0!
0'
0/
#242910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#242920000000
0!
0'
0/
#242930000000
1!
1'
1/
#242940000000
0!
0'
0/
#242950000000
#242960000000
1!
1'
1/
#242970000000
0!
0'
0/
#242980000000
1!
1'
1/
#242990000000
0!
1"
0'
1(
0/
10
#243000000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#243010000000
0!
0'
0/
#243020000000
1!
1'
1/
#243030000000
0!
0'
0/
#243040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#243050000000
0!
0'
0/
#243060000000
1!
1'
1/
#243070000000
0!
1"
0'
1(
0/
10
#243080000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#243090000000
0!
1$
0'
1+
0/
#243100000000
1!
1'
1/
#243110000000
0!
0'
0/
#243120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#243130000000
0!
0'
0/
#243140000000
1!
1'
1/
#243150000000
0!
0'
0/
#243160000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#243170000000
0!
0'
0/
#243180000000
1!
1'
1/
#243190000000
0!
0'
0/
#243200000000
1!
1'
1/
#243210000000
0!
0'
0/
#243220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#243230000000
0!
0'
0/
#243240000000
1!
1'
1/
#243250000000
0!
0'
0/
#243260000000
1!
1'
1/
#243270000000
0!
0'
0/
#243280000000
1!
1'
1/
#243290000000
0!
0'
0/
#243300000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#243310000000
0!
0'
0/
#243320000000
1!
1'
1/
#243330000000
0!
0'
0/
#243340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#243350000000
0!
0'
0/
#243360000000
1!
1'
1/
#243370000000
0!
0'
0/
#243380000000
#243390000000
1!
1'
1/
#243400000000
0!
0'
0/
#243410000000
1!
1'
1/
#243420000000
0!
1"
0'
1(
0/
10
#243430000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#243440000000
0!
0'
0/
#243450000000
1!
1'
1/
#243460000000
0!
0'
0/
#243470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#243480000000
0!
0'
0/
#243490000000
1!
1'
1/
#243500000000
0!
1"
0'
1(
0/
10
#243510000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#243520000000
0!
1$
0'
1+
0/
#243530000000
1!
1'
1/
#243540000000
0!
0'
0/
#243550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#243560000000
0!
0'
0/
#243570000000
1!
1'
1/
#243580000000
0!
0'
0/
#243590000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#243600000000
0!
0'
0/
#243610000000
1!
1'
1/
#243620000000
0!
0'
0/
#243630000000
1!
1'
1/
#243640000000
0!
0'
0/
#243650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#243660000000
0!
0'
0/
#243670000000
1!
1'
1/
#243680000000
0!
0'
0/
#243690000000
1!
1'
1/
#243700000000
0!
0'
0/
#243710000000
1!
1'
1/
#243720000000
0!
0'
0/
#243730000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#243740000000
0!
0'
0/
#243750000000
1!
1'
1/
#243760000000
0!
0'
0/
#243770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#243780000000
0!
0'
0/
#243790000000
1!
1'
1/
#243800000000
0!
0'
0/
#243810000000
#243820000000
1!
1'
1/
#243830000000
0!
0'
0/
#243840000000
1!
1'
1/
#243850000000
0!
1"
0'
1(
0/
10
#243860000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#243870000000
0!
0'
0/
#243880000000
1!
1'
1/
#243890000000
0!
0'
0/
#243900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#243910000000
0!
0'
0/
#243920000000
1!
1'
1/
#243930000000
0!
1"
0'
1(
0/
10
#243940000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#243950000000
0!
1$
0'
1+
0/
#243960000000
1!
1'
1/
#243970000000
0!
0'
0/
#243980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#243990000000
0!
0'
0/
#244000000000
1!
1'
1/
#244010000000
0!
0'
0/
#244020000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#244030000000
0!
0'
0/
#244040000000
1!
1'
1/
#244050000000
0!
0'
0/
#244060000000
1!
1'
1/
#244070000000
0!
0'
0/
#244080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#244090000000
0!
0'
0/
#244100000000
1!
1'
1/
#244110000000
0!
0'
0/
#244120000000
1!
1'
1/
#244130000000
0!
0'
0/
#244140000000
1!
1'
1/
#244150000000
0!
0'
0/
#244160000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#244170000000
0!
0'
0/
#244180000000
1!
1'
1/
#244190000000
0!
0'
0/
#244200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#244210000000
0!
0'
0/
#244220000000
1!
1'
1/
#244230000000
0!
0'
0/
#244240000000
#244250000000
1!
1'
1/
#244260000000
0!
0'
0/
#244270000000
1!
1'
1/
#244280000000
0!
1"
0'
1(
0/
10
#244290000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#244300000000
0!
0'
0/
#244310000000
1!
1'
1/
#244320000000
0!
0'
0/
#244330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#244340000000
0!
0'
0/
#244350000000
1!
1'
1/
#244360000000
0!
1"
0'
1(
0/
10
#244370000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#244380000000
0!
1$
0'
1+
0/
#244390000000
1!
1'
1/
#244400000000
0!
0'
0/
#244410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#244420000000
0!
0'
0/
#244430000000
1!
1'
1/
#244440000000
0!
0'
0/
#244450000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#244460000000
0!
0'
0/
#244470000000
1!
1'
1/
#244480000000
0!
0'
0/
#244490000000
1!
1'
1/
#244500000000
0!
0'
0/
#244510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#244520000000
0!
0'
0/
#244530000000
1!
1'
1/
#244540000000
0!
0'
0/
#244550000000
1!
1'
1/
#244560000000
0!
0'
0/
#244570000000
1!
1'
1/
#244580000000
0!
0'
0/
#244590000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#244600000000
0!
0'
0/
#244610000000
1!
1'
1/
#244620000000
0!
0'
0/
#244630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#244640000000
0!
0'
0/
#244650000000
1!
1'
1/
#244660000000
0!
0'
0/
#244670000000
#244680000000
1!
1'
1/
#244690000000
0!
0'
0/
#244700000000
1!
1'
1/
#244710000000
0!
1"
0'
1(
0/
10
#244720000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#244730000000
0!
0'
0/
#244740000000
1!
1'
1/
#244750000000
0!
0'
0/
#244760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#244770000000
0!
0'
0/
#244780000000
1!
1'
1/
#244790000000
0!
1"
0'
1(
0/
10
#244800000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#244810000000
0!
1$
0'
1+
0/
#244820000000
1!
1'
1/
#244830000000
0!
0'
0/
#244840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#244850000000
0!
0'
0/
#244860000000
1!
1'
1/
#244870000000
0!
0'
0/
#244880000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#244890000000
0!
0'
0/
#244900000000
1!
1'
1/
#244910000000
0!
0'
0/
#244920000000
1!
1'
1/
#244930000000
0!
0'
0/
#244940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#244950000000
0!
0'
0/
#244960000000
1!
1'
1/
#244970000000
0!
0'
0/
#244980000000
1!
1'
1/
#244990000000
0!
0'
0/
#245000000000
1!
1'
1/
#245010000000
0!
0'
0/
#245020000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#245030000000
0!
0'
0/
#245040000000
1!
1'
1/
#245050000000
0!
0'
0/
#245060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#245070000000
0!
0'
0/
#245080000000
1!
1'
1/
#245090000000
0!
0'
0/
#245100000000
#245110000000
1!
1'
1/
#245120000000
0!
0'
0/
#245130000000
1!
1'
1/
#245140000000
0!
1"
0'
1(
0/
10
#245150000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#245160000000
0!
0'
0/
#245170000000
1!
1'
1/
#245180000000
0!
0'
0/
#245190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#245200000000
0!
0'
0/
#245210000000
1!
1'
1/
#245220000000
0!
1"
0'
1(
0/
10
#245230000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#245240000000
0!
1$
0'
1+
0/
#245250000000
1!
1'
1/
#245260000000
0!
0'
0/
#245270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#245280000000
0!
0'
0/
#245290000000
1!
1'
1/
#245300000000
0!
0'
0/
#245310000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#245320000000
0!
0'
0/
#245330000000
1!
1'
1/
#245340000000
0!
0'
0/
#245350000000
1!
1'
1/
#245360000000
0!
0'
0/
#245370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#245380000000
0!
0'
0/
#245390000000
1!
1'
1/
#245400000000
0!
0'
0/
#245410000000
1!
1'
1/
#245420000000
0!
0'
0/
#245430000000
1!
1'
1/
#245440000000
0!
0'
0/
#245450000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#245460000000
0!
0'
0/
#245470000000
1!
1'
1/
#245480000000
0!
0'
0/
#245490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#245500000000
0!
0'
0/
#245510000000
1!
1'
1/
#245520000000
0!
0'
0/
#245530000000
#245540000000
1!
1'
1/
#245550000000
0!
0'
0/
#245560000000
1!
1'
1/
#245570000000
0!
1"
0'
1(
0/
10
#245580000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#245590000000
0!
0'
0/
#245600000000
1!
1'
1/
#245610000000
0!
0'
0/
#245620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#245630000000
0!
0'
0/
#245640000000
1!
1'
1/
#245650000000
0!
1"
0'
1(
0/
10
#245660000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#245670000000
0!
1$
0'
1+
0/
#245680000000
1!
1'
1/
#245690000000
0!
0'
0/
#245700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#245710000000
0!
0'
0/
#245720000000
1!
1'
1/
#245730000000
0!
0'
0/
#245740000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#245750000000
0!
0'
0/
#245760000000
1!
1'
1/
#245770000000
0!
0'
0/
#245780000000
1!
1'
1/
#245790000000
0!
0'
0/
#245800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#245810000000
0!
0'
0/
#245820000000
1!
1'
1/
#245830000000
0!
0'
0/
#245840000000
1!
1'
1/
#245850000000
0!
0'
0/
#245860000000
1!
1'
1/
#245870000000
0!
0'
0/
#245880000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#245890000000
0!
0'
0/
#245900000000
1!
1'
1/
#245910000000
0!
0'
0/
#245920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#245930000000
0!
0'
0/
#245940000000
1!
1'
1/
#245950000000
0!
0'
0/
#245960000000
#245970000000
1!
1'
1/
#245980000000
0!
0'
0/
#245990000000
1!
1'
1/
#246000000000
0!
1"
0'
1(
0/
10
#246010000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#246020000000
0!
0'
0/
#246030000000
1!
1'
1/
#246040000000
0!
0'
0/
#246050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#246060000000
0!
0'
0/
#246070000000
1!
1'
1/
#246080000000
0!
1"
0'
1(
0/
10
#246090000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#246100000000
0!
1$
0'
1+
0/
#246110000000
1!
1'
1/
#246120000000
0!
0'
0/
#246130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#246140000000
0!
0'
0/
#246150000000
1!
1'
1/
#246160000000
0!
0'
0/
#246170000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#246180000000
0!
0'
0/
#246190000000
1!
1'
1/
#246200000000
0!
0'
0/
#246210000000
1!
1'
1/
#246220000000
0!
0'
0/
#246230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#246240000000
0!
0'
0/
#246250000000
1!
1'
1/
#246260000000
0!
0'
0/
#246270000000
1!
1'
1/
#246280000000
0!
0'
0/
#246290000000
1!
1'
1/
#246300000000
0!
0'
0/
#246310000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#246320000000
0!
0'
0/
#246330000000
1!
1'
1/
#246340000000
0!
0'
0/
#246350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#246360000000
0!
0'
0/
#246370000000
1!
1'
1/
#246380000000
0!
0'
0/
#246390000000
#246400000000
1!
1'
1/
#246410000000
0!
0'
0/
#246420000000
1!
1'
1/
#246430000000
0!
1"
0'
1(
0/
10
#246440000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#246450000000
0!
0'
0/
#246460000000
1!
1'
1/
#246470000000
0!
0'
0/
#246480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#246490000000
0!
0'
0/
#246500000000
1!
1'
1/
#246510000000
0!
1"
0'
1(
0/
10
#246520000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#246530000000
0!
1$
0'
1+
0/
#246540000000
1!
1'
1/
#246550000000
0!
0'
0/
#246560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#246570000000
0!
0'
0/
#246580000000
1!
1'
1/
#246590000000
0!
0'
0/
#246600000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#246610000000
0!
0'
0/
#246620000000
1!
1'
1/
#246630000000
0!
0'
0/
#246640000000
1!
1'
1/
#246650000000
0!
0'
0/
#246660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#246670000000
0!
0'
0/
#246680000000
1!
1'
1/
#246690000000
0!
0'
0/
#246700000000
1!
1'
1/
#246710000000
0!
0'
0/
#246720000000
1!
1'
1/
#246730000000
0!
0'
0/
#246740000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#246750000000
0!
0'
0/
#246760000000
1!
1'
1/
#246770000000
0!
0'
0/
#246780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#246790000000
0!
0'
0/
#246800000000
1!
1'
1/
#246810000000
0!
0'
0/
#246820000000
#246830000000
1!
1'
1/
#246840000000
0!
0'
0/
#246850000000
1!
1'
1/
#246860000000
0!
1"
0'
1(
0/
10
#246870000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#246880000000
0!
0'
0/
#246890000000
1!
1'
1/
#246900000000
0!
0'
0/
#246910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#246920000000
0!
0'
0/
#246930000000
1!
1'
1/
#246940000000
0!
1"
0'
1(
0/
10
#246950000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#246960000000
0!
1$
0'
1+
0/
#246970000000
1!
1'
1/
#246980000000
0!
0'
0/
#246990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#247000000000
0!
0'
0/
#247010000000
1!
1'
1/
#247020000000
0!
0'
0/
#247030000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#247040000000
0!
0'
0/
#247050000000
1!
1'
1/
#247060000000
0!
0'
0/
#247070000000
1!
1'
1/
#247080000000
0!
0'
0/
#247090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#247100000000
0!
0'
0/
#247110000000
1!
1'
1/
#247120000000
0!
0'
0/
#247130000000
1!
1'
1/
#247140000000
0!
0'
0/
#247150000000
1!
1'
1/
#247160000000
0!
0'
0/
#247170000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#247180000000
0!
0'
0/
#247190000000
1!
1'
1/
#247200000000
0!
0'
0/
#247210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#247220000000
0!
0'
0/
#247230000000
1!
1'
1/
#247240000000
0!
0'
0/
#247250000000
#247260000000
1!
1'
1/
#247270000000
0!
0'
0/
#247280000000
1!
1'
1/
#247290000000
0!
1"
0'
1(
0/
10
#247300000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#247310000000
0!
0'
0/
#247320000000
1!
1'
1/
#247330000000
0!
0'
0/
#247340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#247350000000
0!
0'
0/
#247360000000
1!
1'
1/
#247370000000
0!
1"
0'
1(
0/
10
#247380000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#247390000000
0!
1$
0'
1+
0/
#247400000000
1!
1'
1/
#247410000000
0!
0'
0/
#247420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#247430000000
0!
0'
0/
#247440000000
1!
1'
1/
#247450000000
0!
0'
0/
#247460000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#247470000000
0!
0'
0/
#247480000000
1!
1'
1/
#247490000000
0!
0'
0/
#247500000000
1!
1'
1/
#247510000000
0!
0'
0/
#247520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#247530000000
0!
0'
0/
#247540000000
1!
1'
1/
#247550000000
0!
0'
0/
#247560000000
1!
1'
1/
#247570000000
0!
0'
0/
#247580000000
1!
1'
1/
#247590000000
0!
0'
0/
#247600000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#247610000000
0!
0'
0/
#247620000000
1!
1'
1/
#247630000000
0!
0'
0/
#247640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#247650000000
0!
0'
0/
#247660000000
1!
1'
1/
#247670000000
0!
0'
0/
#247680000000
#247690000000
1!
1'
1/
#247700000000
0!
0'
0/
#247710000000
1!
1'
1/
#247720000000
0!
1"
0'
1(
0/
10
#247730000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#247740000000
0!
0'
0/
#247750000000
1!
1'
1/
#247760000000
0!
0'
0/
#247770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#247780000000
0!
0'
0/
#247790000000
1!
1'
1/
#247800000000
0!
1"
0'
1(
0/
10
#247810000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#247820000000
0!
1$
0'
1+
0/
#247830000000
1!
1'
1/
#247840000000
0!
0'
0/
#247850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#247860000000
0!
0'
0/
#247870000000
1!
1'
1/
#247880000000
0!
0'
0/
#247890000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#247900000000
0!
0'
0/
#247910000000
1!
1'
1/
#247920000000
0!
0'
0/
#247930000000
1!
1'
1/
#247940000000
0!
0'
0/
#247950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#247960000000
0!
0'
0/
#247970000000
1!
1'
1/
#247980000000
0!
0'
0/
#247990000000
1!
1'
1/
#248000000000
0!
0'
0/
#248010000000
1!
1'
1/
#248020000000
0!
0'
0/
#248030000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#248040000000
0!
0'
0/
#248050000000
1!
1'
1/
#248060000000
0!
0'
0/
#248070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#248080000000
0!
0'
0/
#248090000000
1!
1'
1/
#248100000000
0!
0'
0/
#248110000000
#248120000000
1!
1'
1/
#248130000000
0!
0'
0/
#248140000000
1!
1'
1/
#248150000000
0!
1"
0'
1(
0/
10
#248160000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#248170000000
0!
0'
0/
#248180000000
1!
1'
1/
#248190000000
0!
0'
0/
#248200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#248210000000
0!
0'
0/
#248220000000
1!
1'
1/
#248230000000
0!
1"
0'
1(
0/
10
#248240000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#248250000000
0!
1$
0'
1+
0/
#248260000000
1!
1'
1/
#248270000000
0!
0'
0/
#248280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#248290000000
0!
0'
0/
#248300000000
1!
1'
1/
#248310000000
0!
0'
0/
#248320000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#248330000000
0!
0'
0/
#248340000000
1!
1'
1/
#248350000000
0!
0'
0/
#248360000000
1!
1'
1/
#248370000000
0!
0'
0/
#248380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#248390000000
0!
0'
0/
#248400000000
1!
1'
1/
#248410000000
0!
0'
0/
#248420000000
1!
1'
1/
#248430000000
0!
0'
0/
#248440000000
1!
1'
1/
#248450000000
0!
0'
0/
#248460000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#248470000000
0!
0'
0/
#248480000000
1!
1'
1/
#248490000000
0!
0'
0/
#248500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#248510000000
0!
0'
0/
#248520000000
1!
1'
1/
#248530000000
0!
0'
0/
#248540000000
#248550000000
1!
1'
1/
#248560000000
0!
0'
0/
#248570000000
1!
1'
1/
#248580000000
0!
1"
0'
1(
0/
10
#248590000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#248600000000
0!
0'
0/
#248610000000
1!
1'
1/
#248620000000
0!
0'
0/
#248630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#248640000000
0!
0'
0/
#248650000000
1!
1'
1/
#248660000000
0!
1"
0'
1(
0/
10
#248670000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#248680000000
0!
1$
0'
1+
0/
#248690000000
1!
1'
1/
#248700000000
0!
0'
0/
#248710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#248720000000
0!
0'
0/
#248730000000
1!
1'
1/
#248740000000
0!
0'
0/
#248750000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#248760000000
0!
0'
0/
#248770000000
1!
1'
1/
#248780000000
0!
0'
0/
#248790000000
1!
1'
1/
#248800000000
0!
0'
0/
#248810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#248820000000
0!
0'
0/
#248830000000
1!
1'
1/
#248840000000
0!
0'
0/
#248850000000
1!
1'
1/
#248860000000
0!
0'
0/
#248870000000
1!
1'
1/
#248880000000
0!
0'
0/
#248890000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#248900000000
0!
0'
0/
#248910000000
1!
1'
1/
#248920000000
0!
0'
0/
#248930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#248940000000
0!
0'
0/
#248950000000
1!
1'
1/
#248960000000
0!
0'
0/
#248970000000
#248980000000
1!
1'
1/
#248990000000
0!
0'
0/
#249000000000
1!
1'
1/
#249010000000
0!
1"
0'
1(
0/
10
#249020000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#249030000000
0!
0'
0/
#249040000000
1!
1'
1/
#249050000000
0!
0'
0/
#249060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#249070000000
0!
0'
0/
#249080000000
1!
1'
1/
#249090000000
0!
1"
0'
1(
0/
10
#249100000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#249110000000
0!
1$
0'
1+
0/
#249120000000
1!
1'
1/
#249130000000
0!
0'
0/
#249140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#249150000000
0!
0'
0/
#249160000000
1!
1'
1/
#249170000000
0!
0'
0/
#249180000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#249190000000
0!
0'
0/
#249200000000
1!
1'
1/
#249210000000
0!
0'
0/
#249220000000
1!
1'
1/
#249230000000
0!
0'
0/
#249240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#249250000000
0!
0'
0/
#249260000000
1!
1'
1/
#249270000000
0!
0'
0/
#249280000000
1!
1'
1/
#249290000000
0!
0'
0/
#249300000000
1!
1'
1/
#249310000000
0!
0'
0/
#249320000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#249330000000
0!
0'
0/
#249340000000
1!
1'
1/
#249350000000
0!
0'
0/
#249360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#249370000000
0!
0'
0/
#249380000000
1!
1'
1/
#249390000000
0!
0'
0/
#249400000000
#249410000000
1!
1'
1/
#249420000000
0!
0'
0/
#249430000000
1!
1'
1/
#249440000000
0!
1"
0'
1(
0/
10
#249450000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#249460000000
0!
0'
0/
#249470000000
1!
1'
1/
#249480000000
0!
0'
0/
#249490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#249500000000
0!
0'
0/
#249510000000
1!
1'
1/
#249520000000
0!
1"
0'
1(
0/
10
#249530000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#249540000000
0!
1$
0'
1+
0/
#249550000000
1!
1'
1/
#249560000000
0!
0'
0/
#249570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#249580000000
0!
0'
0/
#249590000000
1!
1'
1/
#249600000000
0!
0'
0/
#249610000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#249620000000
0!
0'
0/
#249630000000
1!
1'
1/
#249640000000
0!
0'
0/
#249650000000
1!
1'
1/
#249660000000
0!
0'
0/
#249670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#249680000000
0!
0'
0/
#249690000000
1!
1'
1/
#249700000000
0!
0'
0/
#249710000000
1!
1'
1/
#249720000000
0!
0'
0/
#249730000000
1!
1'
1/
#249740000000
0!
0'
0/
#249750000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#249760000000
0!
0'
0/
#249770000000
1!
1'
1/
#249780000000
0!
0'
0/
#249790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#249800000000
0!
0'
0/
#249810000000
1!
1'
1/
#249820000000
0!
0'
0/
#249830000000
#249840000000
1!
1'
1/
#249850000000
0!
0'
0/
#249860000000
1!
1'
1/
#249870000000
0!
1"
0'
1(
0/
10
#249880000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#249890000000
0!
0'
0/
#249900000000
1!
1'
1/
#249910000000
0!
0'
0/
#249920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#249930000000
0!
0'
0/
#249940000000
1!
1'
1/
#249950000000
0!
1"
0'
1(
0/
10
#249960000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#249970000000
0!
1$
0'
1+
0/
#249980000000
1!
1'
1/
#249990000000
0!
0'
0/
#250000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#250010000000
0!
0'
0/
#250020000000
1!
1'
1/
#250030000000
0!
0'
0/
#250040000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#250050000000
0!
0'
0/
#250060000000
1!
1'
1/
#250070000000
0!
0'
0/
#250080000000
1!
1'
1/
#250090000000
0!
0'
0/
#250100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#250110000000
0!
0'
0/
#250120000000
1!
1'
1/
#250130000000
0!
0'
0/
#250140000000
1!
1'
1/
#250150000000
0!
0'
0/
#250160000000
1!
1'
1/
#250170000000
0!
0'
0/
#250180000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#250190000000
0!
0'
0/
#250200000000
1!
1'
1/
#250210000000
0!
0'
0/
#250220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#250230000000
0!
0'
0/
#250240000000
1!
1'
1/
#250250000000
0!
0'
0/
#250260000000
#250270000000
1!
1'
1/
#250280000000
0!
0'
0/
#250290000000
1!
1'
1/
#250300000000
0!
1"
0'
1(
0/
10
#250310000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#250320000000
0!
0'
0/
#250330000000
1!
1'
1/
#250340000000
0!
0'
0/
#250350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#250360000000
0!
0'
0/
#250370000000
1!
1'
1/
#250380000000
0!
1"
0'
1(
0/
10
#250390000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#250400000000
0!
1$
0'
1+
0/
#250410000000
1!
1'
1/
#250420000000
0!
0'
0/
#250430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#250440000000
0!
0'
0/
#250450000000
1!
1'
1/
#250460000000
0!
0'
0/
#250470000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#250480000000
0!
0'
0/
#250490000000
1!
1'
1/
#250500000000
0!
0'
0/
#250510000000
1!
1'
1/
#250520000000
0!
0'
0/
#250530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#250540000000
0!
0'
0/
#250550000000
1!
1'
1/
#250560000000
0!
0'
0/
#250570000000
1!
1'
1/
#250580000000
0!
0'
0/
#250590000000
1!
1'
1/
#250600000000
0!
0'
0/
#250610000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#250620000000
0!
0'
0/
#250630000000
1!
1'
1/
#250640000000
0!
0'
0/
#250650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#250660000000
0!
0'
0/
#250670000000
1!
1'
1/
#250680000000
0!
0'
0/
#250690000000
#250700000000
1!
1'
1/
#250710000000
0!
0'
0/
#250720000000
1!
1'
1/
#250730000000
0!
1"
0'
1(
0/
10
#250740000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#250750000000
0!
0'
0/
#250760000000
1!
1'
1/
#250770000000
0!
0'
0/
#250780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#250790000000
0!
0'
0/
#250800000000
1!
1'
1/
#250810000000
0!
1"
0'
1(
0/
10
#250820000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#250830000000
0!
1$
0'
1+
0/
#250840000000
1!
1'
1/
#250850000000
0!
0'
0/
#250860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#250870000000
0!
0'
0/
#250880000000
1!
1'
1/
#250890000000
0!
0'
0/
#250900000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#250910000000
0!
0'
0/
#250920000000
1!
1'
1/
#250930000000
0!
0'
0/
#250940000000
1!
1'
1/
#250950000000
0!
0'
0/
#250960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#250970000000
0!
0'
0/
#250980000000
1!
1'
1/
#250990000000
0!
0'
0/
#251000000000
1!
1'
1/
#251010000000
0!
0'
0/
#251020000000
1!
1'
1/
#251030000000
0!
0'
0/
#251040000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#251050000000
0!
0'
0/
#251060000000
1!
1'
1/
#251070000000
0!
0'
0/
#251080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#251090000000
0!
0'
0/
#251100000000
1!
1'
1/
#251110000000
0!
0'
0/
#251120000000
#251130000000
1!
1'
1/
#251140000000
0!
0'
0/
#251150000000
1!
1'
1/
#251160000000
0!
1"
0'
1(
0/
10
#251170000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#251180000000
0!
0'
0/
#251190000000
1!
1'
1/
#251200000000
0!
0'
0/
#251210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#251220000000
0!
0'
0/
#251230000000
1!
1'
1/
#251240000000
0!
1"
0'
1(
0/
10
#251250000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#251260000000
0!
1$
0'
1+
0/
#251270000000
1!
1'
1/
#251280000000
0!
0'
0/
#251290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#251300000000
0!
0'
0/
#251310000000
1!
1'
1/
#251320000000
0!
0'
0/
#251330000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#251340000000
0!
0'
0/
#251350000000
1!
1'
1/
#251360000000
0!
0'
0/
#251370000000
1!
1'
1/
#251380000000
0!
0'
0/
#251390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#251400000000
0!
0'
0/
#251410000000
1!
1'
1/
#251420000000
0!
0'
0/
#251430000000
1!
1'
1/
#251440000000
0!
0'
0/
#251450000000
1!
1'
1/
#251460000000
0!
0'
0/
#251470000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#251480000000
0!
0'
0/
#251490000000
1!
1'
1/
#251500000000
0!
0'
0/
#251510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#251520000000
0!
0'
0/
#251530000000
1!
1'
1/
#251540000000
0!
0'
0/
#251550000000
#251560000000
1!
1'
1/
#251570000000
0!
0'
0/
#251580000000
1!
1'
1/
#251590000000
0!
1"
0'
1(
0/
10
#251600000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#251610000000
0!
0'
0/
#251620000000
1!
1'
1/
#251630000000
0!
0'
0/
#251640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#251650000000
0!
0'
0/
#251660000000
1!
1'
1/
#251670000000
0!
1"
0'
1(
0/
10
#251680000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#251690000000
0!
1$
0'
1+
0/
#251700000000
1!
1'
1/
#251710000000
0!
0'
0/
#251720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#251730000000
0!
0'
0/
#251740000000
1!
1'
1/
#251750000000
0!
0'
0/
#251760000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#251770000000
0!
0'
0/
#251780000000
1!
1'
1/
#251790000000
0!
0'
0/
#251800000000
1!
1'
1/
#251810000000
0!
0'
0/
#251820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#251830000000
0!
0'
0/
#251840000000
1!
1'
1/
#251850000000
0!
0'
0/
#251860000000
1!
1'
1/
#251870000000
0!
0'
0/
#251880000000
1!
1'
1/
#251890000000
0!
0'
0/
#251900000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#251910000000
0!
0'
0/
#251920000000
1!
1'
1/
#251930000000
0!
0'
0/
#251940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#251950000000
0!
0'
0/
#251960000000
1!
1'
1/
#251970000000
0!
0'
0/
#251980000000
#251990000000
1!
1'
1/
#252000000000
0!
0'
0/
#252010000000
1!
1'
1/
#252020000000
0!
1"
0'
1(
0/
10
#252030000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#252040000000
0!
0'
0/
#252050000000
1!
1'
1/
#252060000000
0!
0'
0/
#252070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#252080000000
0!
0'
0/
#252090000000
1!
1'
1/
#252100000000
0!
1"
0'
1(
0/
10
#252110000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#252120000000
0!
1$
0'
1+
0/
#252130000000
1!
1'
1/
#252140000000
0!
0'
0/
#252150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#252160000000
0!
0'
0/
#252170000000
1!
1'
1/
#252180000000
0!
0'
0/
#252190000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#252200000000
0!
0'
0/
#252210000000
1!
1'
1/
#252220000000
0!
0'
0/
#252230000000
1!
1'
1/
#252240000000
0!
0'
0/
#252250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#252260000000
0!
0'
0/
#252270000000
1!
1'
1/
#252280000000
0!
0'
0/
#252290000000
1!
1'
1/
#252300000000
0!
0'
0/
#252310000000
1!
1'
1/
#252320000000
0!
0'
0/
#252330000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#252340000000
0!
0'
0/
#252350000000
1!
1'
1/
#252360000000
0!
0'
0/
#252370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#252380000000
0!
0'
0/
#252390000000
1!
1'
1/
#252400000000
0!
0'
0/
#252410000000
#252420000000
1!
1'
1/
#252430000000
0!
0'
0/
#252440000000
1!
1'
1/
#252450000000
0!
1"
0'
1(
0/
10
#252460000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#252470000000
0!
0'
0/
#252480000000
1!
1'
1/
#252490000000
0!
0'
0/
#252500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#252510000000
0!
0'
0/
#252520000000
1!
1'
1/
#252530000000
0!
1"
0'
1(
0/
10
#252540000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#252550000000
0!
1$
0'
1+
0/
#252560000000
1!
1'
1/
#252570000000
0!
0'
0/
#252580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#252590000000
0!
0'
0/
#252600000000
1!
1'
1/
#252610000000
0!
0'
0/
#252620000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#252630000000
0!
0'
0/
#252640000000
1!
1'
1/
#252650000000
0!
0'
0/
#252660000000
1!
1'
1/
#252670000000
0!
0'
0/
#252680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#252690000000
0!
0'
0/
#252700000000
1!
1'
1/
#252710000000
0!
0'
0/
#252720000000
1!
1'
1/
#252730000000
0!
0'
0/
#252740000000
1!
1'
1/
#252750000000
0!
0'
0/
#252760000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#252770000000
0!
0'
0/
#252780000000
1!
1'
1/
#252790000000
0!
0'
0/
#252800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#252810000000
0!
0'
0/
#252820000000
1!
1'
1/
#252830000000
0!
0'
0/
#252840000000
#252850000000
1!
1'
1/
#252860000000
0!
0'
0/
#252870000000
1!
1'
1/
#252880000000
0!
1"
0'
1(
0/
10
#252890000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#252900000000
0!
0'
0/
#252910000000
1!
1'
1/
#252920000000
0!
0'
0/
#252930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#252940000000
0!
0'
0/
#252950000000
1!
1'
1/
#252960000000
0!
1"
0'
1(
0/
10
#252970000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#252980000000
0!
1$
0'
1+
0/
#252990000000
1!
1'
1/
#253000000000
0!
0'
0/
#253010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#253020000000
0!
0'
0/
#253030000000
1!
1'
1/
#253040000000
0!
0'
0/
#253050000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#253060000000
0!
0'
0/
#253070000000
1!
1'
1/
#253080000000
0!
0'
0/
#253090000000
1!
1'
1/
#253100000000
0!
0'
0/
#253110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#253120000000
0!
0'
0/
#253130000000
1!
1'
1/
#253140000000
0!
0'
0/
#253150000000
1!
1'
1/
#253160000000
0!
0'
0/
#253170000000
1!
1'
1/
#253180000000
0!
0'
0/
#253190000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#253200000000
0!
0'
0/
#253210000000
1!
1'
1/
#253220000000
0!
0'
0/
#253230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#253240000000
0!
0'
0/
#253250000000
1!
1'
1/
#253260000000
0!
0'
0/
#253270000000
#253280000000
1!
1'
1/
#253290000000
0!
0'
0/
#253300000000
1!
1'
1/
#253310000000
0!
1"
0'
1(
0/
10
#253320000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#253330000000
0!
0'
0/
#253340000000
1!
1'
1/
#253350000000
0!
0'
0/
#253360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#253370000000
0!
0'
0/
#253380000000
1!
1'
1/
#253390000000
0!
1"
0'
1(
0/
10
#253400000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#253410000000
0!
1$
0'
1+
0/
#253420000000
1!
1'
1/
#253430000000
0!
0'
0/
#253440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#253450000000
0!
0'
0/
#253460000000
1!
1'
1/
#253470000000
0!
0'
0/
#253480000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#253490000000
0!
0'
0/
#253500000000
1!
1'
1/
#253510000000
0!
0'
0/
#253520000000
1!
1'
1/
#253530000000
0!
0'
0/
#253540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#253550000000
0!
0'
0/
#253560000000
1!
1'
1/
#253570000000
0!
0'
0/
#253580000000
1!
1'
1/
#253590000000
0!
0'
0/
#253600000000
1!
1'
1/
#253610000000
0!
0'
0/
#253620000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#253630000000
0!
0'
0/
#253640000000
1!
1'
1/
#253650000000
0!
0'
0/
#253660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#253670000000
0!
0'
0/
#253680000000
1!
1'
1/
#253690000000
0!
0'
0/
#253700000000
#253710000000
1!
1'
1/
#253720000000
0!
0'
0/
#253730000000
1!
1'
1/
#253740000000
0!
1"
0'
1(
0/
10
#253750000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#253760000000
0!
0'
0/
#253770000000
1!
1'
1/
#253780000000
0!
0'
0/
#253790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#253800000000
0!
0'
0/
#253810000000
1!
1'
1/
#253820000000
0!
1"
0'
1(
0/
10
#253830000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#253840000000
0!
1$
0'
1+
0/
#253850000000
1!
1'
1/
#253860000000
0!
0'
0/
#253870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#253880000000
0!
0'
0/
#253890000000
1!
1'
1/
#253900000000
0!
0'
0/
#253910000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#253920000000
0!
0'
0/
#253930000000
1!
1'
1/
#253940000000
0!
0'
0/
#253950000000
1!
1'
1/
#253960000000
0!
0'
0/
#253970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#253980000000
0!
0'
0/
#253990000000
1!
1'
1/
#254000000000
0!
0'
0/
#254010000000
1!
1'
1/
#254020000000
0!
0'
0/
#254030000000
1!
1'
1/
#254040000000
0!
0'
0/
#254050000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#254060000000
0!
0'
0/
#254070000000
1!
1'
1/
#254080000000
0!
0'
0/
#254090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#254100000000
0!
0'
0/
#254110000000
1!
1'
1/
#254120000000
0!
0'
0/
#254130000000
#254140000000
1!
1'
1/
#254150000000
0!
0'
0/
#254160000000
1!
1'
1/
#254170000000
0!
1"
0'
1(
0/
10
#254180000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#254190000000
0!
0'
0/
#254200000000
1!
1'
1/
#254210000000
0!
0'
0/
#254220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#254230000000
0!
0'
0/
#254240000000
1!
1'
1/
#254250000000
0!
1"
0'
1(
0/
10
#254260000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#254270000000
0!
1$
0'
1+
0/
#254280000000
1!
1'
1/
#254290000000
0!
0'
0/
#254300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#254310000000
0!
0'
0/
#254320000000
1!
1'
1/
#254330000000
0!
0'
0/
#254340000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#254350000000
0!
0'
0/
#254360000000
1!
1'
1/
#254370000000
0!
0'
0/
#254380000000
1!
1'
1/
#254390000000
0!
0'
0/
#254400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#254410000000
0!
0'
0/
#254420000000
1!
1'
1/
#254430000000
0!
0'
0/
#254440000000
1!
1'
1/
#254450000000
0!
0'
0/
#254460000000
1!
1'
1/
#254470000000
0!
0'
0/
#254480000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#254490000000
0!
0'
0/
#254500000000
1!
1'
1/
#254510000000
0!
0'
0/
#254520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#254530000000
0!
0'
0/
#254540000000
1!
1'
1/
#254550000000
0!
0'
0/
#254560000000
#254570000000
1!
1'
1/
#254580000000
0!
0'
0/
#254590000000
1!
1'
1/
#254600000000
0!
1"
0'
1(
0/
10
#254610000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#254620000000
0!
0'
0/
#254630000000
1!
1'
1/
#254640000000
0!
0'
0/
#254650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#254660000000
0!
0'
0/
#254670000000
1!
1'
1/
#254680000000
0!
1"
0'
1(
0/
10
#254690000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#254700000000
0!
1$
0'
1+
0/
#254710000000
1!
1'
1/
#254720000000
0!
0'
0/
#254730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#254740000000
0!
0'
0/
#254750000000
1!
1'
1/
#254760000000
0!
0'
0/
#254770000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#254780000000
0!
0'
0/
#254790000000
1!
1'
1/
#254800000000
0!
0'
0/
#254810000000
1!
1'
1/
#254820000000
0!
0'
0/
#254830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#254840000000
0!
0'
0/
#254850000000
1!
1'
1/
#254860000000
0!
0'
0/
#254870000000
1!
1'
1/
#254880000000
0!
0'
0/
#254890000000
1!
1'
1/
#254900000000
0!
0'
0/
#254910000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#254920000000
0!
0'
0/
#254930000000
1!
1'
1/
#254940000000
0!
0'
0/
#254950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#254960000000
0!
0'
0/
#254970000000
1!
1'
1/
#254980000000
0!
0'
0/
#254990000000
#255000000000
1!
1'
1/
#255010000000
0!
0'
0/
#255020000000
1!
1'
1/
#255030000000
0!
1"
0'
1(
0/
10
#255040000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#255050000000
0!
0'
0/
#255060000000
1!
1'
1/
#255070000000
0!
0'
0/
#255080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#255090000000
0!
0'
0/
#255100000000
1!
1'
1/
#255110000000
0!
1"
0'
1(
0/
10
#255120000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#255130000000
0!
1$
0'
1+
0/
#255140000000
1!
1'
1/
#255150000000
0!
0'
0/
#255160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#255170000000
0!
0'
0/
#255180000000
1!
1'
1/
#255190000000
0!
0'
0/
#255200000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#255210000000
0!
0'
0/
#255220000000
1!
1'
1/
#255230000000
0!
0'
0/
#255240000000
1!
1'
1/
#255250000000
0!
0'
0/
#255260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#255270000000
0!
0'
0/
#255280000000
1!
1'
1/
#255290000000
0!
0'
0/
#255300000000
1!
1'
1/
#255310000000
0!
0'
0/
#255320000000
1!
1'
1/
#255330000000
0!
0'
0/
#255340000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#255350000000
0!
0'
0/
#255360000000
1!
1'
1/
#255370000000
0!
0'
0/
#255380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#255390000000
0!
0'
0/
#255400000000
1!
1'
1/
#255410000000
0!
0'
0/
#255420000000
#255430000000
1!
1'
1/
#255440000000
0!
0'
0/
#255450000000
1!
1'
1/
#255460000000
0!
1"
0'
1(
0/
10
#255470000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#255480000000
0!
0'
0/
#255490000000
1!
1'
1/
#255500000000
0!
0'
0/
#255510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#255520000000
0!
0'
0/
#255530000000
1!
1'
1/
#255540000000
0!
1"
0'
1(
0/
10
#255550000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#255560000000
0!
1$
0'
1+
0/
#255570000000
1!
1'
1/
#255580000000
0!
0'
0/
#255590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#255600000000
0!
0'
0/
#255610000000
1!
1'
1/
#255620000000
0!
0'
0/
#255630000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#255640000000
0!
0'
0/
#255650000000
1!
1'
1/
#255660000000
0!
0'
0/
#255670000000
1!
1'
1/
#255680000000
0!
0'
0/
#255690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#255700000000
0!
0'
0/
#255710000000
1!
1'
1/
#255720000000
0!
0'
0/
#255730000000
1!
1'
1/
#255740000000
0!
0'
0/
#255750000000
1!
1'
1/
#255760000000
0!
0'
0/
#255770000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#255780000000
0!
0'
0/
#255790000000
1!
1'
1/
#255800000000
0!
0'
0/
#255810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#255820000000
0!
0'
0/
#255830000000
1!
1'
1/
#255840000000
0!
0'
0/
#255850000000
#255860000000
1!
1'
1/
#255870000000
0!
0'
0/
#255880000000
1!
1'
1/
#255890000000
0!
1"
0'
1(
0/
10
#255900000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#255910000000
0!
0'
0/
#255920000000
1!
1'
1/
#255930000000
0!
0'
0/
#255940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#255950000000
0!
0'
0/
#255960000000
1!
1'
1/
#255970000000
0!
1"
0'
1(
0/
10
#255980000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#255990000000
0!
1$
0'
1+
0/
#256000000000
1!
1'
1/
#256010000000
0!
0'
0/
#256020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#256030000000
0!
0'
0/
#256040000000
1!
1'
1/
#256050000000
0!
0'
0/
#256060000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#256070000000
0!
0'
0/
#256080000000
1!
1'
1/
#256090000000
0!
0'
0/
#256100000000
1!
1'
1/
#256110000000
0!
0'
0/
#256120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#256130000000
0!
0'
0/
#256140000000
1!
1'
1/
#256150000000
0!
0'
0/
#256160000000
1!
1'
1/
#256170000000
0!
0'
0/
#256180000000
1!
1'
1/
#256190000000
0!
0'
0/
#256200000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#256210000000
0!
0'
0/
#256220000000
1!
1'
1/
#256230000000
0!
0'
0/
#256240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#256250000000
0!
0'
0/
#256260000000
1!
1'
1/
#256270000000
0!
0'
0/
#256280000000
#256290000000
1!
1'
1/
#256300000000
0!
0'
0/
#256310000000
1!
1'
1/
#256320000000
0!
1"
0'
1(
0/
10
#256330000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#256340000000
0!
0'
0/
#256350000000
1!
1'
1/
#256360000000
0!
0'
0/
#256370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#256380000000
0!
0'
0/
#256390000000
1!
1'
1/
#256400000000
0!
1"
0'
1(
0/
10
#256410000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#256420000000
0!
1$
0'
1+
0/
#256430000000
1!
1'
1/
#256440000000
0!
0'
0/
#256450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#256460000000
0!
0'
0/
#256470000000
1!
1'
1/
#256480000000
0!
0'
0/
#256490000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#256500000000
0!
0'
0/
#256510000000
1!
1'
1/
#256520000000
0!
0'
0/
#256530000000
1!
1'
1/
#256540000000
0!
0'
0/
#256550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#256560000000
0!
0'
0/
#256570000000
1!
1'
1/
#256580000000
0!
0'
0/
#256590000000
1!
1'
1/
#256600000000
0!
0'
0/
#256610000000
1!
1'
1/
#256620000000
0!
0'
0/
#256630000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#256640000000
0!
0'
0/
#256650000000
1!
1'
1/
#256660000000
0!
0'
0/
#256670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#256680000000
0!
0'
0/
#256690000000
1!
1'
1/
#256700000000
0!
0'
0/
#256710000000
#256720000000
1!
1'
1/
#256730000000
0!
0'
0/
#256740000000
1!
1'
1/
#256750000000
0!
1"
0'
1(
0/
10
#256760000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#256770000000
0!
0'
0/
#256780000000
1!
1'
1/
#256790000000
0!
0'
0/
#256800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#256810000000
0!
0'
0/
#256820000000
1!
1'
1/
#256830000000
0!
1"
0'
1(
0/
10
#256840000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#256850000000
0!
1$
0'
1+
0/
#256860000000
1!
1'
1/
#256870000000
0!
0'
0/
#256880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#256890000000
0!
0'
0/
#256900000000
1!
1'
1/
#256910000000
0!
0'
0/
#256920000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#256930000000
0!
0'
0/
#256940000000
1!
1'
1/
#256950000000
0!
0'
0/
#256960000000
1!
1'
1/
#256970000000
0!
0'
0/
#256980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#256990000000
0!
0'
0/
#257000000000
1!
1'
1/
#257010000000
0!
0'
0/
#257020000000
1!
1'
1/
#257030000000
0!
0'
0/
#257040000000
1!
1'
1/
#257050000000
0!
0'
0/
#257060000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#257070000000
0!
0'
0/
#257080000000
1!
1'
1/
#257090000000
0!
0'
0/
#257100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#257110000000
0!
0'
0/
#257120000000
1!
1'
1/
#257130000000
0!
0'
0/
#257140000000
#257150000000
1!
1'
1/
#257160000000
0!
0'
0/
#257170000000
1!
1'
1/
#257180000000
0!
1"
0'
1(
0/
10
#257190000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#257200000000
0!
0'
0/
#257210000000
1!
1'
1/
#257220000000
0!
0'
0/
#257230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#257240000000
0!
0'
0/
#257250000000
1!
1'
1/
#257260000000
0!
1"
0'
1(
0/
10
#257270000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#257280000000
0!
1$
0'
1+
0/
#257290000000
1!
1'
1/
#257300000000
0!
0'
0/
#257310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#257320000000
0!
0'
0/
#257330000000
1!
1'
1/
#257340000000
0!
0'
0/
#257350000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#257360000000
0!
0'
0/
#257370000000
1!
1'
1/
#257380000000
0!
0'
0/
#257390000000
1!
1'
1/
#257400000000
0!
0'
0/
#257410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#257420000000
0!
0'
0/
#257430000000
1!
1'
1/
#257440000000
0!
0'
0/
#257450000000
1!
1'
1/
#257460000000
0!
0'
0/
#257470000000
1!
1'
1/
#257480000000
0!
0'
0/
#257490000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#257500000000
0!
0'
0/
#257510000000
1!
1'
1/
#257520000000
0!
0'
0/
#257530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#257540000000
0!
0'
0/
#257550000000
1!
1'
1/
#257560000000
0!
0'
0/
#257570000000
#257580000000
1!
1'
1/
#257590000000
0!
0'
0/
#257600000000
1!
1'
1/
#257610000000
0!
1"
0'
1(
0/
10
#257620000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#257630000000
0!
0'
0/
#257640000000
1!
1'
1/
#257650000000
0!
0'
0/
#257660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#257670000000
0!
0'
0/
#257680000000
1!
1'
1/
#257690000000
0!
1"
0'
1(
0/
10
#257700000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#257710000000
0!
1$
0'
1+
0/
#257720000000
1!
1'
1/
#257730000000
0!
0'
0/
#257740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#257750000000
0!
0'
0/
#257760000000
1!
1'
1/
#257770000000
0!
0'
0/
#257780000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#257790000000
0!
0'
0/
#257800000000
1!
1'
1/
#257810000000
0!
0'
0/
#257820000000
1!
1'
1/
#257830000000
0!
0'
0/
#257840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#257850000000
0!
0'
0/
#257860000000
1!
1'
1/
#257870000000
0!
0'
0/
#257880000000
1!
1'
1/
#257890000000
0!
0'
0/
#257900000000
1!
1'
1/
#257910000000
0!
0'
0/
#257920000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#257930000000
0!
0'
0/
#257940000000
1!
1'
1/
#257950000000
0!
0'
0/
#257960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#257970000000
0!
0'
0/
#257980000000
1!
1'
1/
#257990000000
0!
0'
0/
#258000000000
#258010000000
1!
1'
1/
#258020000000
0!
0'
0/
#258030000000
1!
1'
1/
#258040000000
0!
1"
0'
1(
0/
10
#258050000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#258060000000
0!
0'
0/
#258070000000
1!
1'
1/
#258080000000
0!
0'
0/
#258090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#258100000000
0!
0'
0/
#258110000000
1!
1'
1/
#258120000000
0!
1"
0'
1(
0/
10
#258130000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#258140000000
0!
1$
0'
1+
0/
#258150000000
1!
1'
1/
#258160000000
0!
0'
0/
#258170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#258180000000
0!
0'
0/
#258190000000
1!
1'
1/
#258200000000
0!
0'
0/
#258210000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#258220000000
0!
0'
0/
#258230000000
1!
1'
1/
#258240000000
0!
0'
0/
#258250000000
1!
1'
1/
#258260000000
0!
0'
0/
#258270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#258280000000
0!
0'
0/
#258290000000
1!
1'
1/
#258300000000
0!
0'
0/
#258310000000
1!
1'
1/
#258320000000
0!
0'
0/
#258330000000
1!
1'
1/
#258340000000
0!
0'
0/
#258350000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#258360000000
0!
0'
0/
#258370000000
1!
1'
1/
#258380000000
0!
0'
0/
#258390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#258400000000
0!
0'
0/
#258410000000
1!
1'
1/
#258420000000
0!
0'
0/
#258430000000
#258440000000
1!
1'
1/
#258450000000
0!
0'
0/
#258460000000
1!
1'
1/
#258470000000
0!
1"
0'
1(
0/
10
#258480000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#258490000000
0!
0'
0/
#258500000000
1!
1'
1/
#258510000000
0!
0'
0/
#258520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#258530000000
0!
0'
0/
#258540000000
1!
1'
1/
#258550000000
0!
1"
0'
1(
0/
10
#258560000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#258570000000
0!
1$
0'
1+
0/
#258580000000
1!
1'
1/
#258590000000
0!
0'
0/
#258600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#258610000000
0!
0'
0/
#258620000000
1!
1'
1/
#258630000000
0!
0'
0/
#258640000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#258650000000
0!
0'
0/
#258660000000
1!
1'
1/
#258670000000
0!
0'
0/
#258680000000
1!
1'
1/
#258690000000
0!
0'
0/
#258700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#258710000000
0!
0'
0/
#258720000000
1!
1'
1/
#258730000000
0!
0'
0/
#258740000000
1!
1'
1/
#258750000000
0!
0'
0/
#258760000000
1!
1'
1/
#258770000000
0!
0'
0/
#258780000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#258790000000
0!
0'
0/
#258800000000
1!
1'
1/
#258810000000
0!
0'
0/
#258820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#258830000000
0!
0'
0/
#258840000000
1!
1'
1/
#258850000000
0!
0'
0/
#258860000000
#258870000000
1!
1'
1/
#258880000000
0!
0'
0/
#258890000000
1!
1'
1/
#258900000000
0!
1"
0'
1(
0/
10
#258910000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#258920000000
0!
0'
0/
#258930000000
1!
1'
1/
#258940000000
0!
0'
0/
#258950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#258960000000
0!
0'
0/
#258970000000
1!
1'
1/
#258980000000
0!
1"
0'
1(
0/
10
#258990000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#259000000000
0!
1$
0'
1+
0/
#259010000000
1!
1'
1/
#259020000000
0!
0'
0/
#259030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#259040000000
0!
0'
0/
#259050000000
1!
1'
1/
#259060000000
0!
0'
0/
#259070000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#259080000000
0!
0'
0/
#259090000000
1!
1'
1/
#259100000000
0!
0'
0/
#259110000000
1!
1'
1/
#259120000000
0!
0'
0/
#259130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#259140000000
0!
0'
0/
#259150000000
1!
1'
1/
#259160000000
0!
0'
0/
#259170000000
1!
1'
1/
#259180000000
0!
0'
0/
#259190000000
1!
1'
1/
#259200000000
0!
0'
0/
#259210000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#259220000000
0!
0'
0/
#259230000000
1!
1'
1/
#259240000000
0!
0'
0/
#259250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#259260000000
0!
0'
0/
#259270000000
1!
1'
1/
#259280000000
0!
0'
0/
#259290000000
#259300000000
1!
1'
1/
#259310000000
0!
0'
0/
#259320000000
1!
1'
1/
#259330000000
0!
1"
0'
1(
0/
10
#259340000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#259350000000
0!
0'
0/
#259360000000
1!
1'
1/
#259370000000
0!
0'
0/
#259380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#259390000000
0!
0'
0/
#259400000000
1!
1'
1/
#259410000000
0!
1"
0'
1(
0/
10
#259420000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#259430000000
0!
1$
0'
1+
0/
#259440000000
1!
1'
1/
#259450000000
0!
0'
0/
#259460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#259470000000
0!
0'
0/
#259480000000
1!
1'
1/
#259490000000
0!
0'
0/
#259500000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#259510000000
0!
0'
0/
#259520000000
1!
1'
1/
#259530000000
0!
0'
0/
#259540000000
1!
1'
1/
#259550000000
0!
0'
0/
#259560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#259570000000
0!
0'
0/
#259580000000
1!
1'
1/
#259590000000
0!
0'
0/
#259600000000
1!
1'
1/
#259610000000
0!
0'
0/
#259620000000
1!
1'
1/
#259630000000
0!
0'
0/
#259640000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#259650000000
0!
0'
0/
#259660000000
1!
1'
1/
#259670000000
0!
0'
0/
#259680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#259690000000
0!
0'
0/
#259700000000
1!
1'
1/
#259710000000
0!
0'
0/
#259720000000
#259730000000
1!
1'
1/
#259740000000
0!
0'
0/
#259750000000
1!
1'
1/
#259760000000
0!
1"
0'
1(
0/
10
#259770000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#259780000000
0!
0'
0/
#259790000000
1!
1'
1/
#259800000000
0!
0'
0/
#259810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#259820000000
0!
0'
0/
#259830000000
1!
1'
1/
#259840000000
0!
1"
0'
1(
0/
10
#259850000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#259860000000
0!
1$
0'
1+
0/
#259870000000
1!
1'
1/
#259880000000
0!
0'
0/
#259890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#259900000000
0!
0'
0/
#259910000000
1!
1'
1/
#259920000000
0!
0'
0/
#259930000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#259940000000
0!
0'
0/
#259950000000
1!
1'
1/
#259960000000
0!
0'
0/
#259970000000
1!
1'
1/
#259980000000
0!
0'
0/
#259990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#260000000000
0!
0'
0/
#260010000000
1!
1'
1/
#260020000000
0!
0'
0/
#260030000000
1!
1'
1/
#260040000000
0!
0'
0/
#260050000000
1!
1'
1/
#260060000000
0!
0'
0/
#260070000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#260080000000
0!
0'
0/
#260090000000
1!
1'
1/
#260100000000
0!
0'
0/
#260110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#260120000000
0!
0'
0/
#260130000000
1!
1'
1/
#260140000000
0!
0'
0/
#260150000000
#260160000000
1!
1'
1/
#260170000000
0!
0'
0/
#260180000000
1!
1'
1/
#260190000000
0!
1"
0'
1(
0/
10
#260200000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#260210000000
0!
0'
0/
#260220000000
1!
1'
1/
#260230000000
0!
0'
0/
#260240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#260250000000
0!
0'
0/
#260260000000
1!
1'
1/
#260270000000
0!
1"
0'
1(
0/
10
#260280000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#260290000000
0!
1$
0'
1+
0/
#260300000000
1!
1'
1/
#260310000000
0!
0'
0/
#260320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#260330000000
0!
0'
0/
#260340000000
1!
1'
1/
#260350000000
0!
0'
0/
#260360000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#260370000000
0!
0'
0/
#260380000000
1!
1'
1/
#260390000000
0!
0'
0/
#260400000000
1!
1'
1/
#260410000000
0!
0'
0/
#260420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#260430000000
0!
0'
0/
#260440000000
1!
1'
1/
#260450000000
0!
0'
0/
#260460000000
1!
1'
1/
#260470000000
0!
0'
0/
#260480000000
1!
1'
1/
#260490000000
0!
0'
0/
#260500000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#260510000000
0!
0'
0/
#260520000000
1!
1'
1/
#260530000000
0!
0'
0/
#260540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#260550000000
0!
0'
0/
#260560000000
1!
1'
1/
#260570000000
0!
0'
0/
#260580000000
#260590000000
1!
1'
1/
#260600000000
0!
0'
0/
#260610000000
1!
1'
1/
#260620000000
0!
1"
0'
1(
0/
10
#260630000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#260640000000
0!
0'
0/
#260650000000
1!
1'
1/
#260660000000
0!
0'
0/
#260670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#260680000000
0!
0'
0/
#260690000000
1!
1'
1/
#260700000000
0!
1"
0'
1(
0/
10
#260710000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#260720000000
0!
1$
0'
1+
0/
#260730000000
1!
1'
1/
#260740000000
0!
0'
0/
#260750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#260760000000
0!
0'
0/
#260770000000
1!
1'
1/
#260780000000
0!
0'
0/
#260790000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#260800000000
0!
0'
0/
#260810000000
1!
1'
1/
#260820000000
0!
0'
0/
#260830000000
1!
1'
1/
#260840000000
0!
0'
0/
#260850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#260860000000
0!
0'
0/
#260870000000
1!
1'
1/
#260880000000
0!
0'
0/
#260890000000
1!
1'
1/
#260900000000
0!
0'
0/
#260910000000
1!
1'
1/
#260920000000
0!
0'
0/
#260930000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#260940000000
0!
0'
0/
#260950000000
1!
1'
1/
#260960000000
0!
0'
0/
#260970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#260980000000
0!
0'
0/
#260990000000
1!
1'
1/
#261000000000
0!
0'
0/
#261010000000
#261020000000
1!
1'
1/
#261030000000
0!
0'
0/
#261040000000
1!
1'
1/
#261050000000
0!
1"
0'
1(
0/
10
#261060000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#261070000000
0!
0'
0/
#261080000000
1!
1'
1/
#261090000000
0!
0'
0/
#261100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#261110000000
0!
0'
0/
#261120000000
1!
1'
1/
#261130000000
0!
1"
0'
1(
0/
10
#261140000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#261150000000
0!
1$
0'
1+
0/
#261160000000
1!
1'
1/
#261170000000
0!
0'
0/
#261180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#261190000000
0!
0'
0/
#261200000000
1!
1'
1/
#261210000000
0!
0'
0/
#261220000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#261230000000
0!
0'
0/
#261240000000
1!
1'
1/
#261250000000
0!
0'
0/
#261260000000
1!
1'
1/
#261270000000
0!
0'
0/
#261280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#261290000000
0!
0'
0/
#261300000000
1!
1'
1/
#261310000000
0!
0'
0/
#261320000000
1!
1'
1/
#261330000000
0!
0'
0/
#261340000000
1!
1'
1/
#261350000000
0!
0'
0/
#261360000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#261370000000
0!
0'
0/
#261380000000
1!
1'
1/
#261390000000
0!
0'
0/
#261400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#261410000000
0!
0'
0/
#261420000000
1!
1'
1/
#261430000000
0!
0'
0/
#261440000000
#261450000000
1!
1'
1/
#261460000000
0!
0'
0/
#261470000000
1!
1'
1/
#261480000000
0!
1"
0'
1(
0/
10
#261490000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#261500000000
0!
0'
0/
#261510000000
1!
1'
1/
#261520000000
0!
0'
0/
#261530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#261540000000
0!
0'
0/
#261550000000
1!
1'
1/
#261560000000
0!
1"
0'
1(
0/
10
#261570000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#261580000000
0!
1$
0'
1+
0/
#261590000000
1!
1'
1/
#261600000000
0!
0'
0/
#261610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#261620000000
0!
0'
0/
#261630000000
1!
1'
1/
#261640000000
0!
0'
0/
#261650000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#261660000000
0!
0'
0/
#261670000000
1!
1'
1/
#261680000000
0!
0'
0/
#261690000000
1!
1'
1/
#261700000000
0!
0'
0/
#261710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#261720000000
0!
0'
0/
#261730000000
1!
1'
1/
#261740000000
0!
0'
0/
#261750000000
1!
1'
1/
#261760000000
0!
0'
0/
#261770000000
1!
1'
1/
#261780000000
0!
0'
0/
#261790000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#261800000000
0!
0'
0/
#261810000000
1!
1'
1/
#261820000000
0!
0'
0/
#261830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#261840000000
0!
0'
0/
#261850000000
1!
1'
1/
#261860000000
0!
0'
0/
#261870000000
#261880000000
1!
1'
1/
#261890000000
0!
0'
0/
#261900000000
1!
1'
1/
#261910000000
0!
1"
0'
1(
0/
10
#261920000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#261930000000
0!
0'
0/
#261940000000
1!
1'
1/
#261950000000
0!
0'
0/
#261960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#261970000000
0!
0'
0/
#261980000000
1!
1'
1/
#261990000000
0!
1"
0'
1(
0/
10
#262000000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#262010000000
0!
1$
0'
1+
0/
#262020000000
1!
1'
1/
#262030000000
0!
0'
0/
#262040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#262050000000
0!
0'
0/
#262060000000
1!
1'
1/
#262070000000
0!
0'
0/
#262080000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#262090000000
0!
0'
0/
#262100000000
1!
1'
1/
#262110000000
0!
0'
0/
#262120000000
1!
1'
1/
#262130000000
0!
0'
0/
#262140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#262150000000
0!
0'
0/
#262160000000
1!
1'
1/
#262170000000
0!
0'
0/
#262180000000
1!
1'
1/
#262190000000
0!
0'
0/
#262200000000
1!
1'
1/
#262210000000
0!
0'
0/
#262220000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#262230000000
0!
0'
0/
#262240000000
1!
1'
1/
#262250000000
0!
0'
0/
#262260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#262270000000
0!
0'
0/
#262280000000
1!
1'
1/
#262290000000
0!
0'
0/
#262300000000
#262310000000
1!
1'
1/
#262320000000
0!
0'
0/
#262330000000
1!
1'
1/
#262340000000
0!
1"
0'
1(
0/
10
#262350000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#262360000000
0!
0'
0/
#262370000000
1!
1'
1/
#262380000000
0!
0'
0/
#262390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#262400000000
0!
0'
0/
#262410000000
1!
1'
1/
#262420000000
0!
1"
0'
1(
0/
10
#262430000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#262440000000
0!
1$
0'
1+
0/
#262450000000
1!
1'
1/
#262460000000
0!
0'
0/
#262470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#262480000000
0!
0'
0/
#262490000000
1!
1'
1/
#262500000000
0!
0'
0/
#262510000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#262520000000
0!
0'
0/
#262530000000
1!
1'
1/
#262540000000
0!
0'
0/
#262550000000
1!
1'
1/
#262560000000
0!
0'
0/
#262570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#262580000000
0!
0'
0/
#262590000000
1!
1'
1/
#262600000000
0!
0'
0/
#262610000000
1!
1'
1/
#262620000000
0!
0'
0/
#262630000000
1!
1'
1/
#262640000000
0!
0'
0/
#262650000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#262660000000
0!
0'
0/
#262670000000
1!
1'
1/
#262680000000
0!
0'
0/
#262690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#262700000000
0!
0'
0/
#262710000000
1!
1'
1/
#262720000000
0!
0'
0/
#262730000000
#262740000000
1!
1'
1/
#262750000000
0!
0'
0/
#262760000000
1!
1'
1/
#262770000000
0!
1"
0'
1(
0/
10
#262780000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#262790000000
0!
0'
0/
#262800000000
1!
1'
1/
#262810000000
0!
0'
0/
#262820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#262830000000
0!
0'
0/
#262840000000
1!
1'
1/
#262850000000
0!
1"
0'
1(
0/
10
#262860000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#262870000000
0!
1$
0'
1+
0/
#262880000000
1!
1'
1/
#262890000000
0!
0'
0/
#262900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#262910000000
0!
0'
0/
#262920000000
1!
1'
1/
#262930000000
0!
0'
0/
#262940000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#262950000000
0!
0'
0/
#262960000000
1!
1'
1/
#262970000000
0!
0'
0/
#262980000000
1!
1'
1/
#262990000000
0!
0'
0/
#263000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#263010000000
0!
0'
0/
#263020000000
1!
1'
1/
#263030000000
0!
0'
0/
#263040000000
1!
1'
1/
#263050000000
0!
0'
0/
#263060000000
1!
1'
1/
#263070000000
0!
0'
0/
#263080000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#263090000000
0!
0'
0/
#263100000000
1!
1'
1/
#263110000000
0!
0'
0/
#263120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#263130000000
0!
0'
0/
#263140000000
1!
1'
1/
#263150000000
0!
0'
0/
#263160000000
#263170000000
1!
1'
1/
#263180000000
0!
0'
0/
#263190000000
1!
1'
1/
#263200000000
0!
1"
0'
1(
0/
10
#263210000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#263220000000
0!
0'
0/
#263230000000
1!
1'
1/
#263240000000
0!
0'
0/
#263250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#263260000000
0!
0'
0/
#263270000000
1!
1'
1/
#263280000000
0!
1"
0'
1(
0/
10
#263290000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#263300000000
0!
1$
0'
1+
0/
#263310000000
1!
1'
1/
#263320000000
0!
0'
0/
#263330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#263340000000
0!
0'
0/
#263350000000
1!
1'
1/
#263360000000
0!
0'
0/
#263370000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#263380000000
0!
0'
0/
#263390000000
1!
1'
1/
#263400000000
0!
0'
0/
#263410000000
1!
1'
1/
#263420000000
0!
0'
0/
#263430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#263440000000
0!
0'
0/
#263450000000
1!
1'
1/
#263460000000
0!
0'
0/
#263470000000
1!
1'
1/
#263480000000
0!
0'
0/
#263490000000
1!
1'
1/
#263500000000
0!
0'
0/
#263510000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#263520000000
0!
0'
0/
#263530000000
1!
1'
1/
#263540000000
0!
0'
0/
#263550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#263560000000
0!
0'
0/
#263570000000
1!
1'
1/
#263580000000
0!
0'
0/
#263590000000
#263600000000
1!
1'
1/
#263610000000
0!
0'
0/
#263620000000
1!
1'
1/
#263630000000
0!
1"
0'
1(
0/
10
#263640000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#263650000000
0!
0'
0/
#263660000000
1!
1'
1/
#263670000000
0!
0'
0/
#263680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#263690000000
0!
0'
0/
#263700000000
1!
1'
1/
#263710000000
0!
1"
0'
1(
0/
10
#263720000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#263730000000
0!
1$
0'
1+
0/
#263740000000
1!
1'
1/
#263750000000
0!
0'
0/
#263760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#263770000000
0!
0'
0/
#263780000000
1!
1'
1/
#263790000000
0!
0'
0/
#263800000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#263810000000
0!
0'
0/
#263820000000
1!
1'
1/
#263830000000
0!
0'
0/
#263840000000
1!
1'
1/
#263850000000
0!
0'
0/
#263860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#263870000000
0!
0'
0/
#263880000000
1!
1'
1/
#263890000000
0!
0'
0/
#263900000000
1!
1'
1/
#263910000000
0!
0'
0/
#263920000000
1!
1'
1/
#263930000000
0!
0'
0/
#263940000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#263950000000
0!
0'
0/
#263960000000
1!
1'
1/
#263970000000
0!
0'
0/
#263980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#263990000000
0!
0'
0/
#264000000000
1!
1'
1/
#264010000000
0!
0'
0/
#264020000000
#264030000000
1!
1'
1/
#264040000000
0!
0'
0/
#264050000000
1!
1'
1/
#264060000000
0!
1"
0'
1(
0/
10
#264070000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#264080000000
0!
0'
0/
#264090000000
1!
1'
1/
#264100000000
0!
0'
0/
#264110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#264120000000
0!
0'
0/
#264130000000
1!
1'
1/
#264140000000
0!
1"
0'
1(
0/
10
#264150000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#264160000000
0!
1$
0'
1+
0/
#264170000000
1!
1'
1/
#264180000000
0!
0'
0/
#264190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#264200000000
0!
0'
0/
#264210000000
1!
1'
1/
#264220000000
0!
0'
0/
#264230000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#264240000000
0!
0'
0/
#264250000000
1!
1'
1/
#264260000000
0!
0'
0/
#264270000000
1!
1'
1/
#264280000000
0!
0'
0/
#264290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#264300000000
0!
0'
0/
#264310000000
1!
1'
1/
#264320000000
0!
0'
0/
#264330000000
1!
1'
1/
#264340000000
0!
0'
0/
#264350000000
1!
1'
1/
#264360000000
0!
0'
0/
#264370000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#264380000000
0!
0'
0/
#264390000000
1!
1'
1/
#264400000000
0!
0'
0/
#264410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#264420000000
0!
0'
0/
#264430000000
1!
1'
1/
#264440000000
0!
0'
0/
#264450000000
#264460000000
1!
1'
1/
#264470000000
0!
0'
0/
#264480000000
1!
1'
1/
#264490000000
0!
1"
0'
1(
0/
10
#264500000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#264510000000
0!
0'
0/
#264520000000
1!
1'
1/
#264530000000
0!
0'
0/
#264540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#264550000000
0!
0'
0/
#264560000000
1!
1'
1/
#264570000000
0!
1"
0'
1(
0/
10
#264580000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#264590000000
0!
1$
0'
1+
0/
#264600000000
1!
1'
1/
#264610000000
0!
0'
0/
#264620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#264630000000
0!
0'
0/
#264640000000
1!
1'
1/
#264650000000
0!
0'
0/
#264660000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#264670000000
0!
0'
0/
#264680000000
1!
1'
1/
#264690000000
0!
0'
0/
#264700000000
1!
1'
1/
#264710000000
0!
0'
0/
#264720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#264730000000
0!
0'
0/
#264740000000
1!
1'
1/
#264750000000
0!
0'
0/
#264760000000
1!
1'
1/
#264770000000
0!
0'
0/
#264780000000
1!
1'
1/
#264790000000
0!
0'
0/
#264800000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#264810000000
0!
0'
0/
#264820000000
1!
1'
1/
#264830000000
0!
0'
0/
#264840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#264850000000
0!
0'
0/
#264860000000
1!
1'
1/
#264870000000
0!
0'
0/
#264880000000
#264890000000
1!
1'
1/
#264900000000
0!
0'
0/
#264910000000
1!
1'
1/
#264920000000
0!
1"
0'
1(
0/
10
#264930000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#264940000000
0!
0'
0/
#264950000000
1!
1'
1/
#264960000000
0!
0'
0/
#264970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#264980000000
0!
0'
0/
#264990000000
1!
1'
1/
#265000000000
0!
1"
0'
1(
0/
10
#265010000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#265020000000
0!
1$
0'
1+
0/
#265030000000
1!
1'
1/
#265040000000
0!
0'
0/
#265050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#265060000000
0!
0'
0/
#265070000000
1!
1'
1/
#265080000000
0!
0'
0/
#265090000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#265100000000
0!
0'
0/
#265110000000
1!
1'
1/
#265120000000
0!
0'
0/
#265130000000
1!
1'
1/
#265140000000
0!
0'
0/
#265150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#265160000000
0!
0'
0/
#265170000000
1!
1'
1/
#265180000000
0!
0'
0/
#265190000000
1!
1'
1/
#265200000000
0!
0'
0/
#265210000000
1!
1'
1/
#265220000000
0!
0'
0/
#265230000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#265240000000
0!
0'
0/
#265250000000
1!
1'
1/
#265260000000
0!
0'
0/
#265270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#265280000000
0!
0'
0/
#265290000000
1!
1'
1/
#265300000000
0!
0'
0/
#265310000000
#265320000000
1!
1'
1/
#265330000000
0!
0'
0/
#265340000000
1!
1'
1/
#265350000000
0!
1"
0'
1(
0/
10
#265360000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#265370000000
0!
0'
0/
#265380000000
1!
1'
1/
#265390000000
0!
0'
0/
#265400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#265410000000
0!
0'
0/
#265420000000
1!
1'
1/
#265430000000
0!
1"
0'
1(
0/
10
#265440000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#265450000000
0!
1$
0'
1+
0/
#265460000000
1!
1'
1/
#265470000000
0!
0'
0/
#265480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#265490000000
0!
0'
0/
#265500000000
1!
1'
1/
#265510000000
0!
0'
0/
#265520000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#265530000000
0!
0'
0/
#265540000000
1!
1'
1/
#265550000000
0!
0'
0/
#265560000000
1!
1'
1/
#265570000000
0!
0'
0/
#265580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#265590000000
0!
0'
0/
#265600000000
1!
1'
1/
#265610000000
0!
0'
0/
#265620000000
1!
1'
1/
#265630000000
0!
0'
0/
#265640000000
1!
1'
1/
#265650000000
0!
0'
0/
#265660000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#265670000000
0!
0'
0/
#265680000000
1!
1'
1/
#265690000000
0!
0'
0/
#265700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#265710000000
0!
0'
0/
#265720000000
1!
1'
1/
#265730000000
0!
0'
0/
#265740000000
#265750000000
1!
1'
1/
#265760000000
0!
0'
0/
#265770000000
1!
1'
1/
#265780000000
0!
1"
0'
1(
0/
10
#265790000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#265800000000
0!
0'
0/
#265810000000
1!
1'
1/
#265820000000
0!
0'
0/
#265830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#265840000000
0!
0'
0/
#265850000000
1!
1'
1/
#265860000000
0!
1"
0'
1(
0/
10
#265870000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#265880000000
0!
1$
0'
1+
0/
#265890000000
1!
1'
1/
#265900000000
0!
0'
0/
#265910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#265920000000
0!
0'
0/
#265930000000
1!
1'
1/
#265940000000
0!
0'
0/
#265950000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#265960000000
0!
0'
0/
#265970000000
1!
1'
1/
#265980000000
0!
0'
0/
#265990000000
1!
1'
1/
#266000000000
0!
0'
0/
#266010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#266020000000
0!
0'
0/
#266030000000
1!
1'
1/
#266040000000
0!
0'
0/
#266050000000
1!
1'
1/
#266060000000
0!
0'
0/
#266070000000
1!
1'
1/
#266080000000
0!
0'
0/
#266090000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#266100000000
0!
0'
0/
#266110000000
1!
1'
1/
#266120000000
0!
0'
0/
#266130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#266140000000
0!
0'
0/
#266150000000
1!
1'
1/
#266160000000
0!
0'
0/
#266170000000
#266180000000
1!
1'
1/
#266190000000
0!
0'
0/
#266200000000
1!
1'
1/
#266210000000
0!
1"
0'
1(
0/
10
#266220000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#266230000000
0!
0'
0/
#266240000000
1!
1'
1/
#266250000000
0!
0'
0/
#266260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#266270000000
0!
0'
0/
#266280000000
1!
1'
1/
#266290000000
0!
1"
0'
1(
0/
10
#266300000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#266310000000
0!
1$
0'
1+
0/
#266320000000
1!
1'
1/
#266330000000
0!
0'
0/
#266340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#266350000000
0!
0'
0/
#266360000000
1!
1'
1/
#266370000000
0!
0'
0/
#266380000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#266390000000
0!
0'
0/
#266400000000
1!
1'
1/
#266410000000
0!
0'
0/
#266420000000
1!
1'
1/
#266430000000
0!
0'
0/
#266440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#266450000000
0!
0'
0/
#266460000000
1!
1'
1/
#266470000000
0!
0'
0/
#266480000000
1!
1'
1/
#266490000000
0!
0'
0/
#266500000000
1!
1'
1/
#266510000000
0!
0'
0/
#266520000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#266530000000
0!
0'
0/
#266540000000
1!
1'
1/
#266550000000
0!
0'
0/
#266560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#266570000000
0!
0'
0/
#266580000000
1!
1'
1/
#266590000000
0!
0'
0/
#266600000000
#266610000000
1!
1'
1/
#266620000000
0!
0'
0/
#266630000000
1!
1'
1/
#266640000000
0!
1"
0'
1(
0/
10
#266650000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#266660000000
0!
0'
0/
#266670000000
1!
1'
1/
#266680000000
0!
0'
0/
#266690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#266700000000
0!
0'
0/
#266710000000
1!
1'
1/
#266720000000
0!
1"
0'
1(
0/
10
#266730000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#266740000000
0!
1$
0'
1+
0/
#266750000000
1!
1'
1/
#266760000000
0!
0'
0/
#266770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#266780000000
0!
0'
0/
#266790000000
1!
1'
1/
#266800000000
0!
0'
0/
#266810000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#266820000000
0!
0'
0/
#266830000000
1!
1'
1/
#266840000000
0!
0'
0/
#266850000000
1!
1'
1/
#266860000000
0!
0'
0/
#266870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#266880000000
0!
0'
0/
#266890000000
1!
1'
1/
#266900000000
0!
0'
0/
#266910000000
1!
1'
1/
#266920000000
0!
0'
0/
#266930000000
1!
1'
1/
#266940000000
0!
0'
0/
#266950000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#266960000000
0!
0'
0/
#266970000000
1!
1'
1/
#266980000000
0!
0'
0/
#266990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#267000000000
0!
0'
0/
#267010000000
1!
1'
1/
#267020000000
0!
0'
0/
#267030000000
#267040000000
1!
1'
1/
#267050000000
0!
0'
0/
#267060000000
1!
1'
1/
#267070000000
0!
1"
0'
1(
0/
10
#267080000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#267090000000
0!
0'
0/
#267100000000
1!
1'
1/
#267110000000
0!
0'
0/
#267120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#267130000000
0!
0'
0/
#267140000000
1!
1'
1/
#267150000000
0!
1"
0'
1(
0/
10
#267160000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#267170000000
0!
1$
0'
1+
0/
#267180000000
1!
1'
1/
#267190000000
0!
0'
0/
#267200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#267210000000
0!
0'
0/
#267220000000
1!
1'
1/
#267230000000
0!
0'
0/
#267240000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#267250000000
0!
0'
0/
#267260000000
1!
1'
1/
#267270000000
0!
0'
0/
#267280000000
1!
1'
1/
#267290000000
0!
0'
0/
#267300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#267310000000
0!
0'
0/
#267320000000
1!
1'
1/
#267330000000
0!
0'
0/
#267340000000
1!
1'
1/
#267350000000
0!
0'
0/
#267360000000
1!
1'
1/
#267370000000
0!
0'
0/
#267380000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#267390000000
0!
0'
0/
#267400000000
1!
1'
1/
#267410000000
0!
0'
0/
#267420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#267430000000
0!
0'
0/
#267440000000
1!
1'
1/
#267450000000
0!
0'
0/
#267460000000
#267470000000
1!
1'
1/
#267480000000
0!
0'
0/
#267490000000
1!
1'
1/
#267500000000
0!
1"
0'
1(
0/
10
#267510000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#267520000000
0!
0'
0/
#267530000000
1!
1'
1/
#267540000000
0!
0'
0/
#267550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#267560000000
0!
0'
0/
#267570000000
1!
1'
1/
#267580000000
0!
1"
0'
1(
0/
10
#267590000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#267600000000
0!
1$
0'
1+
0/
#267610000000
1!
1'
1/
#267620000000
0!
0'
0/
#267630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#267640000000
0!
0'
0/
#267650000000
1!
1'
1/
#267660000000
0!
0'
0/
#267670000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#267680000000
0!
0'
0/
#267690000000
1!
1'
1/
#267700000000
0!
0'
0/
#267710000000
1!
1'
1/
#267720000000
0!
0'
0/
#267730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#267740000000
0!
0'
0/
#267750000000
1!
1'
1/
#267760000000
0!
0'
0/
#267770000000
1!
1'
1/
#267780000000
0!
0'
0/
#267790000000
1!
1'
1/
#267800000000
0!
0'
0/
#267810000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#267820000000
0!
0'
0/
#267830000000
1!
1'
1/
#267840000000
0!
0'
0/
#267850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#267860000000
0!
0'
0/
#267870000000
1!
1'
1/
#267880000000
0!
0'
0/
#267890000000
#267900000000
1!
1'
1/
#267910000000
0!
0'
0/
#267920000000
1!
1'
1/
#267930000000
0!
1"
0'
1(
0/
10
#267940000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#267950000000
0!
0'
0/
#267960000000
1!
1'
1/
#267970000000
0!
0'
0/
#267980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#267990000000
0!
0'
0/
#268000000000
1!
1'
1/
#268010000000
0!
1"
0'
1(
0/
10
#268020000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#268030000000
0!
1$
0'
1+
0/
#268040000000
1!
1'
1/
#268050000000
0!
0'
0/
#268060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#268070000000
0!
0'
0/
#268080000000
1!
1'
1/
#268090000000
0!
0'
0/
#268100000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#268110000000
0!
0'
0/
#268120000000
1!
1'
1/
#268130000000
0!
0'
0/
#268140000000
1!
1'
1/
#268150000000
0!
0'
0/
#268160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#268170000000
0!
0'
0/
#268180000000
1!
1'
1/
#268190000000
0!
0'
0/
#268200000000
1!
1'
1/
#268210000000
0!
0'
0/
#268220000000
1!
1'
1/
#268230000000
0!
0'
0/
#268240000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#268250000000
0!
0'
0/
#268260000000
1!
1'
1/
#268270000000
0!
0'
0/
#268280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#268290000000
0!
0'
0/
#268300000000
1!
1'
1/
#268310000000
0!
0'
0/
#268320000000
#268330000000
1!
1'
1/
#268340000000
0!
0'
0/
#268350000000
1!
1'
1/
#268360000000
0!
1"
0'
1(
0/
10
#268370000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#268380000000
0!
0'
0/
#268390000000
1!
1'
1/
#268400000000
0!
0'
0/
#268410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#268420000000
0!
0'
0/
#268430000000
1!
1'
1/
#268440000000
0!
1"
0'
1(
0/
10
#268450000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#268460000000
0!
1$
0'
1+
0/
#268470000000
1!
1'
1/
#268480000000
0!
0'
0/
#268490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#268500000000
0!
0'
0/
#268510000000
1!
1'
1/
#268520000000
0!
0'
0/
#268530000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#268540000000
0!
0'
0/
#268550000000
1!
1'
1/
#268560000000
0!
0'
0/
#268570000000
1!
1'
1/
#268580000000
0!
0'
0/
#268590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#268600000000
0!
0'
0/
#268610000000
1!
1'
1/
#268620000000
0!
0'
0/
#268630000000
1!
1'
1/
#268640000000
0!
0'
0/
#268650000000
1!
1'
1/
#268660000000
0!
0'
0/
#268670000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#268680000000
0!
0'
0/
#268690000000
1!
1'
1/
#268700000000
0!
0'
0/
#268710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#268720000000
0!
0'
0/
#268730000000
1!
1'
1/
#268740000000
0!
0'
0/
#268750000000
#268760000000
1!
1'
1/
#268770000000
0!
0'
0/
#268780000000
1!
1'
1/
#268790000000
0!
1"
0'
1(
0/
10
#268800000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#268810000000
0!
0'
0/
#268820000000
1!
1'
1/
#268830000000
0!
0'
0/
#268840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#268850000000
0!
0'
0/
#268860000000
1!
1'
1/
#268870000000
0!
1"
0'
1(
0/
10
#268880000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#268890000000
0!
1$
0'
1+
0/
#268900000000
1!
1'
1/
#268910000000
0!
0'
0/
#268920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#268930000000
0!
0'
0/
#268940000000
1!
1'
1/
#268950000000
0!
0'
0/
#268960000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#268970000000
0!
0'
0/
#268980000000
1!
1'
1/
#268990000000
0!
0'
0/
#269000000000
1!
1'
1/
#269010000000
0!
0'
0/
#269020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#269030000000
0!
0'
0/
#269040000000
1!
1'
1/
#269050000000
0!
0'
0/
#269060000000
1!
1'
1/
#269070000000
0!
0'
0/
#269080000000
1!
1'
1/
#269090000000
0!
0'
0/
#269100000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#269110000000
0!
0'
0/
#269120000000
1!
1'
1/
#269130000000
0!
0'
0/
#269140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#269150000000
0!
0'
0/
#269160000000
1!
1'
1/
#269170000000
0!
0'
0/
#269180000000
#269190000000
1!
1'
1/
#269200000000
0!
0'
0/
#269210000000
1!
1'
1/
#269220000000
0!
1"
0'
1(
0/
10
#269230000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#269240000000
0!
0'
0/
#269250000000
1!
1'
1/
#269260000000
0!
0'
0/
#269270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#269280000000
0!
0'
0/
#269290000000
1!
1'
1/
#269300000000
0!
1"
0'
1(
0/
10
#269310000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#269320000000
0!
1$
0'
1+
0/
#269330000000
1!
1'
1/
#269340000000
0!
0'
0/
#269350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#269360000000
0!
0'
0/
#269370000000
1!
1'
1/
#269380000000
0!
0'
0/
#269390000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#269400000000
0!
0'
0/
#269410000000
1!
1'
1/
#269420000000
0!
0'
0/
#269430000000
1!
1'
1/
#269440000000
0!
0'
0/
#269450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#269460000000
0!
0'
0/
#269470000000
1!
1'
1/
#269480000000
0!
0'
0/
#269490000000
1!
1'
1/
#269500000000
0!
0'
0/
#269510000000
1!
1'
1/
#269520000000
0!
0'
0/
#269530000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#269540000000
0!
0'
0/
#269550000000
1!
1'
1/
#269560000000
0!
0'
0/
#269570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#269580000000
0!
0'
0/
#269590000000
1!
1'
1/
#269600000000
0!
0'
0/
#269610000000
#269620000000
1!
1'
1/
#269630000000
0!
0'
0/
#269640000000
1!
1'
1/
#269650000000
0!
1"
0'
1(
0/
10
#269660000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#269670000000
0!
0'
0/
#269680000000
1!
1'
1/
#269690000000
0!
0'
0/
#269700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#269710000000
0!
0'
0/
#269720000000
1!
1'
1/
#269730000000
0!
1"
0'
1(
0/
10
#269740000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#269750000000
0!
1$
0'
1+
0/
#269760000000
1!
1'
1/
#269770000000
0!
0'
0/
#269780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#269790000000
0!
0'
0/
#269800000000
1!
1'
1/
#269810000000
0!
0'
0/
#269820000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#269830000000
0!
0'
0/
#269840000000
1!
1'
1/
#269850000000
0!
0'
0/
#269860000000
1!
1'
1/
#269870000000
0!
0'
0/
#269880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#269890000000
0!
0'
0/
#269900000000
1!
1'
1/
#269910000000
0!
0'
0/
#269920000000
1!
1'
1/
#269930000000
0!
0'
0/
#269940000000
1!
1'
1/
#269950000000
0!
0'
0/
#269960000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#269970000000
0!
0'
0/
#269980000000
1!
1'
1/
#269990000000
0!
0'
0/
#270000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#270010000000
0!
0'
0/
#270020000000
1!
1'
1/
#270030000000
0!
0'
0/
#270040000000
#270050000000
1!
1'
1/
#270060000000
0!
0'
0/
#270070000000
1!
1'
1/
#270080000000
0!
1"
0'
1(
0/
10
#270090000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#270100000000
0!
0'
0/
#270110000000
1!
1'
1/
#270120000000
0!
0'
0/
#270130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#270140000000
0!
0'
0/
#270150000000
1!
1'
1/
#270160000000
0!
1"
0'
1(
0/
10
#270170000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#270180000000
0!
1$
0'
1+
0/
#270190000000
1!
1'
1/
#270200000000
0!
0'
0/
#270210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#270220000000
0!
0'
0/
#270230000000
1!
1'
1/
#270240000000
0!
0'
0/
#270250000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#270260000000
0!
0'
0/
#270270000000
1!
1'
1/
#270280000000
0!
0'
0/
#270290000000
1!
1'
1/
#270300000000
0!
0'
0/
#270310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#270320000000
0!
0'
0/
#270330000000
1!
1'
1/
#270340000000
0!
0'
0/
#270350000000
1!
1'
1/
#270360000000
0!
0'
0/
#270370000000
1!
1'
1/
#270380000000
0!
0'
0/
#270390000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#270400000000
0!
0'
0/
#270410000000
1!
1'
1/
#270420000000
0!
0'
0/
#270430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#270440000000
0!
0'
0/
#270450000000
1!
1'
1/
#270460000000
0!
0'
0/
#270470000000
#270480000000
1!
1'
1/
#270490000000
0!
0'
0/
#270500000000
1!
1'
1/
#270510000000
0!
1"
0'
1(
0/
10
#270520000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#270530000000
0!
0'
0/
#270540000000
1!
1'
1/
#270550000000
0!
0'
0/
#270560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#270570000000
0!
0'
0/
#270580000000
1!
1'
1/
#270590000000
0!
1"
0'
1(
0/
10
#270600000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#270610000000
0!
1$
0'
1+
0/
#270620000000
1!
1'
1/
#270630000000
0!
0'
0/
#270640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#270650000000
0!
0'
0/
#270660000000
1!
1'
1/
#270670000000
0!
0'
0/
#270680000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#270690000000
0!
0'
0/
#270700000000
1!
1'
1/
#270710000000
0!
0'
0/
#270720000000
1!
1'
1/
#270730000000
0!
0'
0/
#270740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#270750000000
0!
0'
0/
#270760000000
1!
1'
1/
#270770000000
0!
0'
0/
#270780000000
1!
1'
1/
#270790000000
0!
0'
0/
#270800000000
1!
1'
1/
#270810000000
0!
0'
0/
#270820000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#270830000000
0!
0'
0/
#270840000000
1!
1'
1/
#270850000000
0!
0'
0/
#270860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#270870000000
0!
0'
0/
#270880000000
1!
1'
1/
#270890000000
0!
0'
0/
#270900000000
#270910000000
1!
1'
1/
#270920000000
0!
0'
0/
#270930000000
1!
1'
1/
#270940000000
0!
1"
0'
1(
0/
10
#270950000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#270960000000
0!
0'
0/
#270970000000
1!
1'
1/
#270980000000
0!
0'
0/
#270990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#271000000000
0!
0'
0/
#271010000000
1!
1'
1/
#271020000000
0!
1"
0'
1(
0/
10
#271030000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#271040000000
0!
1$
0'
1+
0/
#271050000000
1!
1'
1/
#271060000000
0!
0'
0/
#271070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#271080000000
0!
0'
0/
#271090000000
1!
1'
1/
#271100000000
0!
0'
0/
#271110000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#271120000000
0!
0'
0/
#271130000000
1!
1'
1/
#271140000000
0!
0'
0/
#271150000000
1!
1'
1/
#271160000000
0!
0'
0/
#271170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#271180000000
0!
0'
0/
#271190000000
1!
1'
1/
#271200000000
0!
0'
0/
#271210000000
1!
1'
1/
#271220000000
0!
0'
0/
#271230000000
1!
1'
1/
#271240000000
0!
0'
0/
#271250000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#271260000000
0!
0'
0/
#271270000000
1!
1'
1/
#271280000000
0!
0'
0/
#271290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#271300000000
0!
0'
0/
#271310000000
1!
1'
1/
#271320000000
0!
0'
0/
#271330000000
#271340000000
1!
1'
1/
#271350000000
0!
0'
0/
#271360000000
1!
1'
1/
#271370000000
0!
1"
0'
1(
0/
10
#271380000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#271390000000
0!
0'
0/
#271400000000
1!
1'
1/
#271410000000
0!
0'
0/
#271420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#271430000000
0!
0'
0/
#271440000000
1!
1'
1/
#271450000000
0!
1"
0'
1(
0/
10
#271460000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#271470000000
0!
1$
0'
1+
0/
#271480000000
1!
1'
1/
#271490000000
0!
0'
0/
#271500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#271510000000
0!
0'
0/
#271520000000
1!
1'
1/
#271530000000
0!
0'
0/
#271540000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#271550000000
0!
0'
0/
#271560000000
1!
1'
1/
#271570000000
0!
0'
0/
#271580000000
1!
1'
1/
#271590000000
0!
0'
0/
#271600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#271610000000
0!
0'
0/
#271620000000
1!
1'
1/
#271630000000
0!
0'
0/
#271640000000
1!
1'
1/
#271650000000
0!
0'
0/
#271660000000
1!
1'
1/
#271670000000
0!
0'
0/
#271680000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#271690000000
0!
0'
0/
#271700000000
1!
1'
1/
#271710000000
0!
0'
0/
#271720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#271730000000
0!
0'
0/
#271740000000
1!
1'
1/
#271750000000
0!
0'
0/
#271760000000
#271770000000
1!
1'
1/
#271780000000
0!
0'
0/
#271790000000
1!
1'
1/
#271800000000
0!
1"
0'
1(
0/
10
#271810000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#271820000000
0!
0'
0/
#271830000000
1!
1'
1/
#271840000000
0!
0'
0/
#271850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#271860000000
0!
0'
0/
#271870000000
1!
1'
1/
#271880000000
0!
1"
0'
1(
0/
10
#271890000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#271900000000
0!
1$
0'
1+
0/
#271910000000
1!
1'
1/
#271920000000
0!
0'
0/
#271930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#271940000000
0!
0'
0/
#271950000000
1!
1'
1/
#271960000000
0!
0'
0/
#271970000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#271980000000
0!
0'
0/
#271990000000
1!
1'
1/
#272000000000
0!
0'
0/
#272010000000
1!
1'
1/
#272020000000
0!
0'
0/
#272030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#272040000000
0!
0'
0/
#272050000000
1!
1'
1/
#272060000000
0!
0'
0/
#272070000000
1!
1'
1/
#272080000000
0!
0'
0/
#272090000000
1!
1'
1/
#272100000000
0!
0'
0/
#272110000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#272120000000
0!
0'
0/
#272130000000
1!
1'
1/
#272140000000
0!
0'
0/
#272150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#272160000000
0!
0'
0/
#272170000000
1!
1'
1/
#272180000000
0!
0'
0/
#272190000000
#272200000000
1!
1'
1/
#272210000000
0!
0'
0/
#272220000000
1!
1'
1/
#272230000000
0!
1"
0'
1(
0/
10
#272240000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#272250000000
0!
0'
0/
#272260000000
1!
1'
1/
#272270000000
0!
0'
0/
#272280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#272290000000
0!
0'
0/
#272300000000
1!
1'
1/
#272310000000
0!
1"
0'
1(
0/
10
#272320000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#272330000000
0!
1$
0'
1+
0/
#272340000000
1!
1'
1/
#272350000000
0!
0'
0/
#272360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#272370000000
0!
0'
0/
#272380000000
1!
1'
1/
#272390000000
0!
0'
0/
#272400000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#272410000000
0!
0'
0/
#272420000000
1!
1'
1/
#272430000000
0!
0'
0/
#272440000000
1!
1'
1/
#272450000000
0!
0'
0/
#272460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#272470000000
0!
0'
0/
#272480000000
1!
1'
1/
#272490000000
0!
0'
0/
#272500000000
1!
1'
1/
#272510000000
0!
0'
0/
#272520000000
1!
1'
1/
#272530000000
0!
0'
0/
#272540000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#272550000000
0!
0'
0/
#272560000000
1!
1'
1/
#272570000000
0!
0'
0/
#272580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#272590000000
0!
0'
0/
#272600000000
1!
1'
1/
#272610000000
0!
0'
0/
#272620000000
#272630000000
1!
1'
1/
#272640000000
0!
0'
0/
#272650000000
1!
1'
1/
#272660000000
0!
1"
0'
1(
0/
10
#272670000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#272680000000
0!
0'
0/
#272690000000
1!
1'
1/
#272700000000
0!
0'
0/
#272710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#272720000000
0!
0'
0/
#272730000000
1!
1'
1/
#272740000000
0!
1"
0'
1(
0/
10
#272750000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#272760000000
0!
1$
0'
1+
0/
#272770000000
1!
1'
1/
#272780000000
0!
0'
0/
#272790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#272800000000
0!
0'
0/
#272810000000
1!
1'
1/
#272820000000
0!
0'
0/
#272830000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#272840000000
0!
0'
0/
#272850000000
1!
1'
1/
#272860000000
0!
0'
0/
#272870000000
1!
1'
1/
#272880000000
0!
0'
0/
#272890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#272900000000
0!
0'
0/
#272910000000
1!
1'
1/
#272920000000
0!
0'
0/
#272930000000
1!
1'
1/
#272940000000
0!
0'
0/
#272950000000
1!
1'
1/
#272960000000
0!
0'
0/
#272970000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#272980000000
0!
0'
0/
#272990000000
1!
1'
1/
#273000000000
0!
0'
0/
#273010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#273020000000
0!
0'
0/
#273030000000
1!
1'
1/
#273040000000
0!
0'
0/
#273050000000
#273060000000
1!
1'
1/
#273070000000
0!
0'
0/
#273080000000
1!
1'
1/
#273090000000
0!
1"
0'
1(
0/
10
#273100000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#273110000000
0!
0'
0/
#273120000000
1!
1'
1/
#273130000000
0!
0'
0/
#273140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#273150000000
0!
0'
0/
#273160000000
1!
1'
1/
#273170000000
0!
1"
0'
1(
0/
10
#273180000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#273190000000
0!
1$
0'
1+
0/
#273200000000
1!
1'
1/
#273210000000
0!
0'
0/
#273220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#273230000000
0!
0'
0/
#273240000000
1!
1'
1/
#273250000000
0!
0'
0/
#273260000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#273270000000
0!
0'
0/
#273280000000
1!
1'
1/
#273290000000
0!
0'
0/
#273300000000
1!
1'
1/
#273310000000
0!
0'
0/
#273320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#273330000000
0!
0'
0/
#273340000000
1!
1'
1/
#273350000000
0!
0'
0/
#273360000000
1!
1'
1/
#273370000000
0!
0'
0/
#273380000000
1!
1'
1/
#273390000000
0!
0'
0/
#273400000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#273410000000
0!
0'
0/
#273420000000
1!
1'
1/
#273430000000
0!
0'
0/
#273440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#273450000000
0!
0'
0/
#273460000000
1!
1'
1/
#273470000000
0!
0'
0/
#273480000000
#273490000000
1!
1'
1/
#273500000000
0!
0'
0/
#273510000000
1!
1'
1/
#273520000000
0!
1"
0'
1(
0/
10
#273530000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#273540000000
0!
0'
0/
#273550000000
1!
1'
1/
#273560000000
0!
0'
0/
#273570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#273580000000
0!
0'
0/
#273590000000
1!
1'
1/
#273600000000
0!
1"
0'
1(
0/
10
#273610000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#273620000000
0!
1$
0'
1+
0/
#273630000000
1!
1'
1/
#273640000000
0!
0'
0/
#273650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#273660000000
0!
0'
0/
#273670000000
1!
1'
1/
#273680000000
0!
0'
0/
#273690000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#273700000000
0!
0'
0/
#273710000000
1!
1'
1/
#273720000000
0!
0'
0/
#273730000000
1!
1'
1/
#273740000000
0!
0'
0/
#273750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#273760000000
0!
0'
0/
#273770000000
1!
1'
1/
#273780000000
0!
0'
0/
#273790000000
1!
1'
1/
#273800000000
0!
0'
0/
#273810000000
1!
1'
1/
#273820000000
0!
0'
0/
#273830000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#273840000000
0!
0'
0/
#273850000000
1!
1'
1/
#273860000000
0!
0'
0/
#273870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#273880000000
0!
0'
0/
#273890000000
1!
1'
1/
#273900000000
0!
0'
0/
#273910000000
#273920000000
1!
1'
1/
#273930000000
0!
0'
0/
#273940000000
1!
1'
1/
#273950000000
0!
1"
0'
1(
0/
10
#273960000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#273970000000
0!
0'
0/
#273980000000
1!
1'
1/
#273990000000
0!
0'
0/
#274000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#274010000000
0!
0'
0/
#274020000000
1!
1'
1/
#274030000000
0!
1"
0'
1(
0/
10
#274040000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#274050000000
0!
1$
0'
1+
0/
#274060000000
1!
1'
1/
#274070000000
0!
0'
0/
#274080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#274090000000
0!
0'
0/
#274100000000
1!
1'
1/
#274110000000
0!
0'
0/
#274120000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#274130000000
0!
0'
0/
#274140000000
1!
1'
1/
#274150000000
0!
0'
0/
#274160000000
1!
1'
1/
#274170000000
0!
0'
0/
#274180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#274190000000
0!
0'
0/
#274200000000
1!
1'
1/
#274210000000
0!
0'
0/
#274220000000
1!
1'
1/
#274230000000
0!
0'
0/
#274240000000
1!
1'
1/
#274250000000
0!
0'
0/
#274260000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#274270000000
0!
0'
0/
#274280000000
1!
1'
1/
#274290000000
0!
0'
0/
#274300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#274310000000
0!
0'
0/
#274320000000
1!
1'
1/
#274330000000
0!
0'
0/
#274340000000
#274350000000
1!
1'
1/
#274360000000
0!
0'
0/
#274370000000
1!
1'
1/
#274380000000
0!
1"
0'
1(
0/
10
#274390000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#274400000000
0!
0'
0/
#274410000000
1!
1'
1/
#274420000000
0!
0'
0/
#274430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#274440000000
0!
0'
0/
#274450000000
1!
1'
1/
#274460000000
0!
1"
0'
1(
0/
10
#274470000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#274480000000
0!
1$
0'
1+
0/
#274490000000
1!
1'
1/
#274500000000
0!
0'
0/
#274510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#274520000000
0!
0'
0/
#274530000000
1!
1'
1/
#274540000000
0!
0'
0/
#274550000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#274560000000
0!
0'
0/
#274570000000
1!
1'
1/
#274580000000
0!
0'
0/
#274590000000
1!
1'
1/
#274600000000
0!
0'
0/
#274610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#274620000000
0!
0'
0/
#274630000000
1!
1'
1/
#274640000000
0!
0'
0/
#274650000000
1!
1'
1/
#274660000000
0!
0'
0/
#274670000000
1!
1'
1/
#274680000000
0!
0'
0/
#274690000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#274700000000
0!
0'
0/
#274710000000
1!
1'
1/
#274720000000
0!
0'
0/
#274730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#274740000000
0!
0'
0/
#274750000000
1!
1'
1/
#274760000000
0!
0'
0/
#274770000000
#274780000000
1!
1'
1/
#274790000000
0!
0'
0/
#274800000000
1!
1'
1/
#274810000000
0!
1"
0'
1(
0/
10
#274820000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#274830000000
0!
0'
0/
#274840000000
1!
1'
1/
#274850000000
0!
0'
0/
#274860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#274870000000
0!
0'
0/
#274880000000
1!
1'
1/
#274890000000
0!
1"
0'
1(
0/
10
#274900000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#274910000000
0!
1$
0'
1+
0/
#274920000000
1!
1'
1/
#274930000000
0!
0'
0/
#274940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#274950000000
0!
0'
0/
#274960000000
1!
1'
1/
#274970000000
0!
0'
0/
#274980000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#274990000000
0!
0'
0/
#275000000000
1!
1'
1/
#275010000000
0!
0'
0/
#275020000000
1!
1'
1/
#275030000000
0!
0'
0/
#275040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#275050000000
0!
0'
0/
#275060000000
1!
1'
1/
#275070000000
0!
0'
0/
#275080000000
1!
1'
1/
#275090000000
0!
0'
0/
#275100000000
1!
1'
1/
#275110000000
0!
0'
0/
#275120000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#275130000000
0!
0'
0/
#275140000000
1!
1'
1/
#275150000000
0!
0'
0/
#275160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#275170000000
0!
0'
0/
#275180000000
1!
1'
1/
#275190000000
0!
0'
0/
#275200000000
#275210000000
1!
1'
1/
#275220000000
0!
0'
0/
#275230000000
1!
1'
1/
#275240000000
0!
1"
0'
1(
0/
10
#275250000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#275260000000
0!
0'
0/
#275270000000
1!
1'
1/
#275280000000
0!
0'
0/
#275290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#275300000000
0!
0'
0/
#275310000000
1!
1'
1/
#275320000000
0!
1"
0'
1(
0/
10
#275330000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#275340000000
0!
1$
0'
1+
0/
#275350000000
1!
1'
1/
#275360000000
0!
0'
0/
#275370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#275380000000
0!
0'
0/
#275390000000
1!
1'
1/
#275400000000
0!
0'
0/
#275410000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#275420000000
0!
0'
0/
#275430000000
1!
1'
1/
#275440000000
0!
0'
0/
#275450000000
1!
1'
1/
#275460000000
0!
0'
0/
#275470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#275480000000
0!
0'
0/
#275490000000
1!
1'
1/
#275500000000
0!
0'
0/
#275510000000
1!
1'
1/
#275520000000
0!
0'
0/
#275530000000
1!
1'
1/
#275540000000
0!
0'
0/
#275550000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#275560000000
0!
0'
0/
#275570000000
1!
1'
1/
#275580000000
0!
0'
0/
#275590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#275600000000
0!
0'
0/
#275610000000
1!
1'
1/
#275620000000
0!
0'
0/
#275630000000
#275640000000
1!
1'
1/
#275650000000
0!
0'
0/
#275660000000
1!
1'
1/
#275670000000
0!
1"
0'
1(
0/
10
#275680000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#275690000000
0!
0'
0/
#275700000000
1!
1'
1/
#275710000000
0!
0'
0/
#275720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#275730000000
0!
0'
0/
#275740000000
1!
1'
1/
#275750000000
0!
1"
0'
1(
0/
10
#275760000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#275770000000
0!
1$
0'
1+
0/
#275780000000
1!
1'
1/
#275790000000
0!
0'
0/
#275800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#275810000000
0!
0'
0/
#275820000000
1!
1'
1/
#275830000000
0!
0'
0/
#275840000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#275850000000
0!
0'
0/
#275860000000
1!
1'
1/
#275870000000
0!
0'
0/
#275880000000
1!
1'
1/
#275890000000
0!
0'
0/
#275900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#275910000000
0!
0'
0/
#275920000000
1!
1'
1/
#275930000000
0!
0'
0/
#275940000000
1!
1'
1/
#275950000000
0!
0'
0/
#275960000000
1!
1'
1/
#275970000000
0!
0'
0/
#275980000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#275990000000
0!
0'
0/
#276000000000
1!
1'
1/
#276010000000
0!
0'
0/
#276020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#276030000000
0!
0'
0/
#276040000000
1!
1'
1/
#276050000000
0!
0'
0/
#276060000000
#276070000000
1!
1'
1/
#276080000000
0!
0'
0/
#276090000000
1!
1'
1/
#276100000000
0!
1"
0'
1(
0/
10
#276110000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#276120000000
0!
0'
0/
#276130000000
1!
1'
1/
#276140000000
0!
0'
0/
#276150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#276160000000
0!
0'
0/
#276170000000
1!
1'
1/
#276180000000
0!
1"
0'
1(
0/
10
#276190000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#276200000000
0!
1$
0'
1+
0/
#276210000000
1!
1'
1/
#276220000000
0!
0'
0/
#276230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#276240000000
0!
0'
0/
#276250000000
1!
1'
1/
#276260000000
0!
0'
0/
#276270000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#276280000000
0!
0'
0/
#276290000000
1!
1'
1/
#276300000000
0!
0'
0/
#276310000000
1!
1'
1/
#276320000000
0!
0'
0/
#276330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#276340000000
0!
0'
0/
#276350000000
1!
1'
1/
#276360000000
0!
0'
0/
#276370000000
1!
1'
1/
#276380000000
0!
0'
0/
#276390000000
1!
1'
1/
#276400000000
0!
0'
0/
#276410000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#276420000000
0!
0'
0/
#276430000000
1!
1'
1/
#276440000000
0!
0'
0/
#276450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#276460000000
0!
0'
0/
#276470000000
1!
1'
1/
#276480000000
0!
0'
0/
#276490000000
#276500000000
1!
1'
1/
#276510000000
0!
0'
0/
#276520000000
1!
1'
1/
#276530000000
0!
1"
0'
1(
0/
10
#276540000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#276550000000
0!
0'
0/
#276560000000
1!
1'
1/
#276570000000
0!
0'
0/
#276580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#276590000000
0!
0'
0/
#276600000000
1!
1'
1/
#276610000000
0!
1"
0'
1(
0/
10
#276620000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#276630000000
0!
1$
0'
1+
0/
#276640000000
1!
1'
1/
#276650000000
0!
0'
0/
#276660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#276670000000
0!
0'
0/
#276680000000
1!
1'
1/
#276690000000
0!
0'
0/
#276700000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#276710000000
0!
0'
0/
#276720000000
1!
1'
1/
#276730000000
0!
0'
0/
#276740000000
1!
1'
1/
#276750000000
0!
0'
0/
#276760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#276770000000
0!
0'
0/
#276780000000
1!
1'
1/
#276790000000
0!
0'
0/
#276800000000
1!
1'
1/
#276810000000
0!
0'
0/
#276820000000
1!
1'
1/
#276830000000
0!
0'
0/
#276840000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#276850000000
0!
0'
0/
#276860000000
1!
1'
1/
#276870000000
0!
0'
0/
#276880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#276890000000
0!
0'
0/
#276900000000
1!
1'
1/
#276910000000
0!
0'
0/
#276920000000
#276930000000
1!
1'
1/
#276940000000
0!
0'
0/
#276950000000
1!
1'
1/
#276960000000
0!
1"
0'
1(
0/
10
#276970000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#276980000000
0!
0'
0/
#276990000000
1!
1'
1/
#277000000000
0!
0'
0/
#277010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#277020000000
0!
0'
0/
#277030000000
1!
1'
1/
#277040000000
0!
1"
0'
1(
0/
10
#277050000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#277060000000
0!
1$
0'
1+
0/
#277070000000
1!
1'
1/
#277080000000
0!
0'
0/
#277090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#277100000000
0!
0'
0/
#277110000000
1!
1'
1/
#277120000000
0!
0'
0/
#277130000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#277140000000
0!
0'
0/
#277150000000
1!
1'
1/
#277160000000
0!
0'
0/
#277170000000
1!
1'
1/
#277180000000
0!
0'
0/
#277190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#277200000000
0!
0'
0/
#277210000000
1!
1'
1/
#277220000000
0!
0'
0/
#277230000000
1!
1'
1/
#277240000000
0!
0'
0/
#277250000000
1!
1'
1/
#277260000000
0!
0'
0/
#277270000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#277280000000
0!
0'
0/
#277290000000
1!
1'
1/
#277300000000
0!
0'
0/
#277310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#277320000000
0!
0'
0/
#277330000000
1!
1'
1/
#277340000000
0!
0'
0/
#277350000000
#277360000000
1!
1'
1/
#277370000000
0!
0'
0/
#277380000000
1!
1'
1/
#277390000000
0!
1"
0'
1(
0/
10
#277400000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#277410000000
0!
0'
0/
#277420000000
1!
1'
1/
#277430000000
0!
0'
0/
#277440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#277450000000
0!
0'
0/
#277460000000
1!
1'
1/
#277470000000
0!
1"
0'
1(
0/
10
#277480000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#277490000000
0!
1$
0'
1+
0/
#277500000000
1!
1'
1/
#277510000000
0!
0'
0/
#277520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#277530000000
0!
0'
0/
#277540000000
1!
1'
1/
#277550000000
0!
0'
0/
#277560000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#277570000000
0!
0'
0/
#277580000000
1!
1'
1/
#277590000000
0!
0'
0/
#277600000000
1!
1'
1/
#277610000000
0!
0'
0/
#277620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#277630000000
0!
0'
0/
#277640000000
1!
1'
1/
#277650000000
0!
0'
0/
#277660000000
1!
1'
1/
#277670000000
0!
0'
0/
#277680000000
1!
1'
1/
#277690000000
0!
0'
0/
#277700000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#277710000000
0!
0'
0/
#277720000000
1!
1'
1/
#277730000000
0!
0'
0/
#277740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#277750000000
0!
0'
0/
#277760000000
1!
1'
1/
#277770000000
0!
0'
0/
#277780000000
#277790000000
1!
1'
1/
#277800000000
0!
0'
0/
#277810000000
1!
1'
1/
#277820000000
0!
1"
0'
1(
0/
10
#277830000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#277840000000
0!
0'
0/
#277850000000
1!
1'
1/
#277860000000
0!
0'
0/
#277870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#277880000000
0!
0'
0/
#277890000000
1!
1'
1/
#277900000000
0!
1"
0'
1(
0/
10
#277910000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#277920000000
0!
1$
0'
1+
0/
#277930000000
1!
1'
1/
#277940000000
0!
0'
0/
#277950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#277960000000
0!
0'
0/
#277970000000
1!
1'
1/
#277980000000
0!
0'
0/
#277990000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#278000000000
0!
0'
0/
#278010000000
1!
1'
1/
#278020000000
0!
0'
0/
#278030000000
1!
1'
1/
#278040000000
0!
0'
0/
#278050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#278060000000
0!
0'
0/
#278070000000
1!
1'
1/
#278080000000
0!
0'
0/
#278090000000
1!
1'
1/
#278100000000
0!
0'
0/
#278110000000
1!
1'
1/
#278120000000
0!
0'
0/
#278130000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#278140000000
0!
0'
0/
#278150000000
1!
1'
1/
#278160000000
0!
0'
0/
#278170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#278180000000
0!
0'
0/
#278190000000
1!
1'
1/
#278200000000
0!
0'
0/
#278210000000
#278220000000
1!
1'
1/
#278230000000
0!
0'
0/
#278240000000
1!
1'
1/
#278250000000
0!
1"
0'
1(
0/
10
#278260000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#278270000000
0!
0'
0/
#278280000000
1!
1'
1/
#278290000000
0!
0'
0/
#278300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#278310000000
0!
0'
0/
#278320000000
1!
1'
1/
#278330000000
0!
1"
0'
1(
0/
10
#278340000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#278350000000
0!
1$
0'
1+
0/
#278360000000
1!
1'
1/
#278370000000
0!
0'
0/
#278380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#278390000000
0!
0'
0/
#278400000000
1!
1'
1/
#278410000000
0!
0'
0/
#278420000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#278430000000
0!
0'
0/
#278440000000
1!
1'
1/
#278450000000
0!
0'
0/
#278460000000
1!
1'
1/
#278470000000
0!
0'
0/
#278480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#278490000000
0!
0'
0/
#278500000000
1!
1'
1/
#278510000000
0!
0'
0/
#278520000000
1!
1'
1/
#278530000000
0!
0'
0/
#278540000000
1!
1'
1/
#278550000000
0!
0'
0/
#278560000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#278570000000
0!
0'
0/
#278580000000
1!
1'
1/
#278590000000
0!
0'
0/
#278600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#278610000000
0!
0'
0/
#278620000000
1!
1'
1/
#278630000000
0!
0'
0/
#278640000000
#278650000000
1!
1'
1/
#278660000000
0!
0'
0/
#278670000000
1!
1'
1/
#278680000000
0!
1"
0'
1(
0/
10
#278690000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#278700000000
0!
0'
0/
#278710000000
1!
1'
1/
#278720000000
0!
0'
0/
#278730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#278740000000
0!
0'
0/
#278750000000
1!
1'
1/
#278760000000
0!
1"
0'
1(
0/
10
#278770000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#278780000000
0!
1$
0'
1+
0/
#278790000000
1!
1'
1/
#278800000000
0!
0'
0/
#278810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#278820000000
0!
0'
0/
#278830000000
1!
1'
1/
#278840000000
0!
0'
0/
#278850000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#278860000000
0!
0'
0/
#278870000000
1!
1'
1/
#278880000000
0!
0'
0/
#278890000000
1!
1'
1/
#278900000000
0!
0'
0/
#278910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#278920000000
0!
0'
0/
#278930000000
1!
1'
1/
#278940000000
0!
0'
0/
#278950000000
1!
1'
1/
#278960000000
0!
0'
0/
#278970000000
1!
1'
1/
#278980000000
0!
0'
0/
#278990000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#279000000000
0!
0'
0/
#279010000000
1!
1'
1/
#279020000000
0!
0'
0/
#279030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#279040000000
0!
0'
0/
#279050000000
1!
1'
1/
#279060000000
0!
0'
0/
#279070000000
#279080000000
1!
1'
1/
#279090000000
0!
0'
0/
#279100000000
1!
1'
1/
#279110000000
0!
1"
0'
1(
0/
10
#279120000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#279130000000
0!
0'
0/
#279140000000
1!
1'
1/
#279150000000
0!
0'
0/
#279160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#279170000000
0!
0'
0/
#279180000000
1!
1'
1/
#279190000000
0!
1"
0'
1(
0/
10
#279200000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#279210000000
0!
1$
0'
1+
0/
#279220000000
1!
1'
1/
#279230000000
0!
0'
0/
#279240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#279250000000
0!
0'
0/
#279260000000
1!
1'
1/
#279270000000
0!
0'
0/
#279280000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#279290000000
0!
0'
0/
#279300000000
1!
1'
1/
#279310000000
0!
0'
0/
#279320000000
1!
1'
1/
#279330000000
0!
0'
0/
#279340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#279350000000
0!
0'
0/
#279360000000
1!
1'
1/
#279370000000
0!
0'
0/
#279380000000
1!
1'
1/
#279390000000
0!
0'
0/
#279400000000
1!
1'
1/
#279410000000
0!
0'
0/
#279420000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#279430000000
0!
0'
0/
#279440000000
1!
1'
1/
#279450000000
0!
0'
0/
#279460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#279470000000
0!
0'
0/
#279480000000
1!
1'
1/
#279490000000
0!
0'
0/
#279500000000
#279510000000
1!
1'
1/
#279520000000
0!
0'
0/
#279530000000
1!
1'
1/
#279540000000
0!
1"
0'
1(
0/
10
#279550000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#279560000000
0!
0'
0/
#279570000000
1!
1'
1/
#279580000000
0!
0'
0/
#279590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#279600000000
0!
0'
0/
#279610000000
1!
1'
1/
#279620000000
0!
1"
0'
1(
0/
10
#279630000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#279640000000
0!
1$
0'
1+
0/
#279650000000
1!
1'
1/
#279660000000
0!
0'
0/
#279670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#279680000000
0!
0'
0/
#279690000000
1!
1'
1/
#279700000000
0!
0'
0/
#279710000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#279720000000
0!
0'
0/
#279730000000
1!
1'
1/
#279740000000
0!
0'
0/
#279750000000
1!
1'
1/
#279760000000
0!
0'
0/
#279770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#279780000000
0!
0'
0/
#279790000000
1!
1'
1/
#279800000000
0!
0'
0/
#279810000000
1!
1'
1/
#279820000000
0!
0'
0/
#279830000000
1!
1'
1/
#279840000000
0!
0'
0/
#279850000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#279860000000
0!
0'
0/
#279870000000
1!
1'
1/
#279880000000
0!
0'
0/
#279890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#279900000000
0!
0'
0/
#279910000000
1!
1'
1/
#279920000000
0!
0'
0/
#279930000000
#279940000000
1!
1'
1/
#279950000000
0!
0'
0/
#279960000000
1!
1'
1/
#279970000000
0!
1"
0'
1(
0/
10
#279980000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#279990000000
0!
0'
0/
#280000000000
1!
1'
1/
#280010000000
0!
0'
0/
#280020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#280030000000
0!
0'
0/
#280040000000
1!
1'
1/
#280050000000
0!
1"
0'
1(
0/
10
#280060000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#280070000000
0!
1$
0'
1+
0/
#280080000000
1!
1'
1/
#280090000000
0!
0'
0/
#280100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#280110000000
0!
0'
0/
#280120000000
1!
1'
1/
#280130000000
0!
0'
0/
#280140000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#280150000000
0!
0'
0/
#280160000000
1!
1'
1/
#280170000000
0!
0'
0/
#280180000000
1!
1'
1/
#280190000000
0!
0'
0/
#280200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#280210000000
0!
0'
0/
#280220000000
1!
1'
1/
#280230000000
0!
0'
0/
#280240000000
1!
1'
1/
#280250000000
0!
0'
0/
#280260000000
1!
1'
1/
#280270000000
0!
0'
0/
#280280000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#280290000000
0!
0'
0/
#280300000000
1!
1'
1/
#280310000000
0!
0'
0/
#280320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#280330000000
0!
0'
0/
#280340000000
1!
1'
1/
#280350000000
0!
0'
0/
#280360000000
#280370000000
1!
1'
1/
#280380000000
0!
0'
0/
#280390000000
1!
1'
1/
#280400000000
0!
1"
0'
1(
0/
10
#280410000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#280420000000
0!
0'
0/
#280430000000
1!
1'
1/
#280440000000
0!
0'
0/
#280450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#280460000000
0!
0'
0/
#280470000000
1!
1'
1/
#280480000000
0!
1"
0'
1(
0/
10
#280490000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#280500000000
0!
1$
0'
1+
0/
#280510000000
1!
1'
1/
#280520000000
0!
0'
0/
#280530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#280540000000
0!
0'
0/
#280550000000
1!
1'
1/
#280560000000
0!
0'
0/
#280570000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#280580000000
0!
0'
0/
#280590000000
1!
1'
1/
#280600000000
0!
0'
0/
#280610000000
1!
1'
1/
#280620000000
0!
0'
0/
#280630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#280640000000
0!
0'
0/
#280650000000
1!
1'
1/
#280660000000
0!
0'
0/
#280670000000
1!
1'
1/
#280680000000
0!
0'
0/
#280690000000
1!
1'
1/
#280700000000
0!
0'
0/
#280710000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#280720000000
0!
0'
0/
#280730000000
1!
1'
1/
#280740000000
0!
0'
0/
#280750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#280760000000
0!
0'
0/
#280770000000
1!
1'
1/
#280780000000
0!
0'
0/
#280790000000
#280800000000
1!
1'
1/
#280810000000
0!
0'
0/
#280820000000
1!
1'
1/
#280830000000
0!
1"
0'
1(
0/
10
#280840000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#280850000000
0!
0'
0/
#280860000000
1!
1'
1/
#280870000000
0!
0'
0/
#280880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#280890000000
0!
0'
0/
#280900000000
1!
1'
1/
#280910000000
0!
1"
0'
1(
0/
10
#280920000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#280930000000
0!
1$
0'
1+
0/
#280940000000
1!
1'
1/
#280950000000
0!
0'
0/
#280960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#280970000000
0!
0'
0/
#280980000000
1!
1'
1/
#280990000000
0!
0'
0/
#281000000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#281010000000
0!
0'
0/
#281020000000
1!
1'
1/
#281030000000
0!
0'
0/
#281040000000
1!
1'
1/
#281050000000
0!
0'
0/
#281060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#281070000000
0!
0'
0/
#281080000000
1!
1'
1/
#281090000000
0!
0'
0/
#281100000000
1!
1'
1/
#281110000000
0!
0'
0/
#281120000000
1!
1'
1/
#281130000000
0!
0'
0/
#281140000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#281150000000
0!
0'
0/
#281160000000
1!
1'
1/
#281170000000
0!
0'
0/
#281180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#281190000000
0!
0'
0/
#281200000000
1!
1'
1/
#281210000000
0!
0'
0/
#281220000000
#281230000000
1!
1'
1/
#281240000000
0!
0'
0/
#281250000000
1!
1'
1/
#281260000000
0!
1"
0'
1(
0/
10
#281270000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#281280000000
0!
0'
0/
#281290000000
1!
1'
1/
#281300000000
0!
0'
0/
#281310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#281320000000
0!
0'
0/
#281330000000
1!
1'
1/
#281340000000
0!
1"
0'
1(
0/
10
#281350000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#281360000000
0!
1$
0'
1+
0/
#281370000000
1!
1'
1/
#281380000000
0!
0'
0/
#281390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#281400000000
0!
0'
0/
#281410000000
1!
1'
1/
#281420000000
0!
0'
0/
#281430000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#281440000000
0!
0'
0/
#281450000000
1!
1'
1/
#281460000000
0!
0'
0/
#281470000000
1!
1'
1/
#281480000000
0!
0'
0/
#281490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#281500000000
0!
0'
0/
#281510000000
1!
1'
1/
#281520000000
0!
0'
0/
#281530000000
1!
1'
1/
#281540000000
0!
0'
0/
#281550000000
1!
1'
1/
#281560000000
0!
0'
0/
#281570000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#281580000000
0!
0'
0/
#281590000000
1!
1'
1/
#281600000000
0!
0'
0/
#281610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#281620000000
0!
0'
0/
#281630000000
1!
1'
1/
#281640000000
0!
0'
0/
#281650000000
#281660000000
1!
1'
1/
#281670000000
0!
0'
0/
#281680000000
1!
1'
1/
#281690000000
0!
1"
0'
1(
0/
10
#281700000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#281710000000
0!
0'
0/
#281720000000
1!
1'
1/
#281730000000
0!
0'
0/
#281740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#281750000000
0!
0'
0/
#281760000000
1!
1'
1/
#281770000000
0!
1"
0'
1(
0/
10
#281780000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#281790000000
0!
1$
0'
1+
0/
#281800000000
1!
1'
1/
#281810000000
0!
0'
0/
#281820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#281830000000
0!
0'
0/
#281840000000
1!
1'
1/
#281850000000
0!
0'
0/
#281860000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#281870000000
0!
0'
0/
#281880000000
1!
1'
1/
#281890000000
0!
0'
0/
#281900000000
1!
1'
1/
#281910000000
0!
0'
0/
#281920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#281930000000
0!
0'
0/
#281940000000
1!
1'
1/
#281950000000
0!
0'
0/
#281960000000
1!
1'
1/
#281970000000
0!
0'
0/
#281980000000
1!
1'
1/
#281990000000
0!
0'
0/
#282000000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#282010000000
0!
0'
0/
#282020000000
1!
1'
1/
#282030000000
0!
0'
0/
#282040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#282050000000
0!
0'
0/
#282060000000
1!
1'
1/
#282070000000
0!
0'
0/
#282080000000
#282090000000
1!
1'
1/
#282100000000
0!
0'
0/
#282110000000
1!
1'
1/
#282120000000
0!
1"
0'
1(
0/
10
#282130000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#282140000000
0!
0'
0/
#282150000000
1!
1'
1/
#282160000000
0!
0'
0/
#282170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#282180000000
0!
0'
0/
#282190000000
1!
1'
1/
#282200000000
0!
1"
0'
1(
0/
10
#282210000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#282220000000
0!
1$
0'
1+
0/
#282230000000
1!
1'
1/
#282240000000
0!
0'
0/
#282250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#282260000000
0!
0'
0/
#282270000000
1!
1'
1/
#282280000000
0!
0'
0/
#282290000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#282300000000
0!
0'
0/
#282310000000
1!
1'
1/
#282320000000
0!
0'
0/
#282330000000
1!
1'
1/
#282340000000
0!
0'
0/
#282350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#282360000000
0!
0'
0/
#282370000000
1!
1'
1/
#282380000000
0!
0'
0/
#282390000000
1!
1'
1/
#282400000000
0!
0'
0/
#282410000000
1!
1'
1/
#282420000000
0!
0'
0/
#282430000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#282440000000
0!
0'
0/
#282450000000
1!
1'
1/
#282460000000
0!
0'
0/
#282470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#282480000000
0!
0'
0/
#282490000000
1!
1'
1/
#282500000000
0!
0'
0/
#282510000000
#282520000000
1!
1'
1/
#282530000000
0!
0'
0/
#282540000000
1!
1'
1/
#282550000000
0!
1"
0'
1(
0/
10
#282560000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#282570000000
0!
0'
0/
#282580000000
1!
1'
1/
#282590000000
0!
0'
0/
#282600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#282610000000
0!
0'
0/
#282620000000
1!
1'
1/
#282630000000
0!
1"
0'
1(
0/
10
#282640000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#282650000000
0!
1$
0'
1+
0/
#282660000000
1!
1'
1/
#282670000000
0!
0'
0/
#282680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#282690000000
0!
0'
0/
#282700000000
1!
1'
1/
#282710000000
0!
0'
0/
#282720000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#282730000000
0!
0'
0/
#282740000000
1!
1'
1/
#282750000000
0!
0'
0/
#282760000000
1!
1'
1/
#282770000000
0!
0'
0/
#282780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#282790000000
0!
0'
0/
#282800000000
1!
1'
1/
#282810000000
0!
0'
0/
#282820000000
1!
1'
1/
#282830000000
0!
0'
0/
#282840000000
1!
1'
1/
#282850000000
0!
0'
0/
#282860000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#282870000000
0!
0'
0/
#282880000000
1!
1'
1/
#282890000000
0!
0'
0/
#282900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#282910000000
0!
0'
0/
#282920000000
1!
1'
1/
#282930000000
0!
0'
0/
#282940000000
#282950000000
1!
1'
1/
#282960000000
0!
0'
0/
#282970000000
1!
1'
1/
#282980000000
0!
1"
0'
1(
0/
10
#282990000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#283000000000
0!
0'
0/
#283010000000
1!
1'
1/
#283020000000
0!
0'
0/
#283030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#283040000000
0!
0'
0/
#283050000000
1!
1'
1/
#283060000000
0!
1"
0'
1(
0/
10
#283070000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#283080000000
0!
1$
0'
1+
0/
#283090000000
1!
1'
1/
#283100000000
0!
0'
0/
#283110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#283120000000
0!
0'
0/
#283130000000
1!
1'
1/
#283140000000
0!
0'
0/
#283150000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#283160000000
0!
0'
0/
#283170000000
1!
1'
1/
#283180000000
0!
0'
0/
#283190000000
1!
1'
1/
#283200000000
0!
0'
0/
#283210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#283220000000
0!
0'
0/
#283230000000
1!
1'
1/
#283240000000
0!
0'
0/
#283250000000
1!
1'
1/
#283260000000
0!
0'
0/
#283270000000
1!
1'
1/
#283280000000
0!
0'
0/
#283290000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#283300000000
0!
0'
0/
#283310000000
1!
1'
1/
#283320000000
0!
0'
0/
#283330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#283340000000
0!
0'
0/
#283350000000
1!
1'
1/
#283360000000
0!
0'
0/
#283370000000
#283380000000
1!
1'
1/
#283390000000
0!
0'
0/
#283400000000
1!
1'
1/
#283410000000
0!
1"
0'
1(
0/
10
#283420000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#283430000000
0!
0'
0/
#283440000000
1!
1'
1/
#283450000000
0!
0'
0/
#283460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#283470000000
0!
0'
0/
#283480000000
1!
1'
1/
#283490000000
0!
1"
0'
1(
0/
10
#283500000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#283510000000
0!
1$
0'
1+
0/
#283520000000
1!
1'
1/
#283530000000
0!
0'
0/
#283540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#283550000000
0!
0'
0/
#283560000000
1!
1'
1/
#283570000000
0!
0'
0/
#283580000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#283590000000
0!
0'
0/
#283600000000
1!
1'
1/
#283610000000
0!
0'
0/
#283620000000
1!
1'
1/
#283630000000
0!
0'
0/
#283640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#283650000000
0!
0'
0/
#283660000000
1!
1'
1/
#283670000000
0!
0'
0/
#283680000000
1!
1'
1/
#283690000000
0!
0'
0/
#283700000000
1!
1'
1/
#283710000000
0!
0'
0/
#283720000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#283730000000
0!
0'
0/
#283740000000
1!
1'
1/
#283750000000
0!
0'
0/
#283760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#283770000000
0!
0'
0/
#283780000000
1!
1'
1/
#283790000000
0!
0'
0/
#283800000000
#283810000000
1!
1'
1/
#283820000000
0!
0'
0/
#283830000000
1!
1'
1/
#283840000000
0!
1"
0'
1(
0/
10
#283850000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#283860000000
0!
0'
0/
#283870000000
1!
1'
1/
#283880000000
0!
0'
0/
#283890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#283900000000
0!
0'
0/
#283910000000
1!
1'
1/
#283920000000
0!
1"
0'
1(
0/
10
#283930000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#283940000000
0!
1$
0'
1+
0/
#283950000000
1!
1'
1/
#283960000000
0!
0'
0/
#283970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#283980000000
0!
0'
0/
#283990000000
1!
1'
1/
#284000000000
0!
0'
0/
#284010000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#284020000000
0!
0'
0/
#284030000000
1!
1'
1/
#284040000000
0!
0'
0/
#284050000000
1!
1'
1/
#284060000000
0!
0'
0/
#284070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#284080000000
0!
0'
0/
#284090000000
1!
1'
1/
#284100000000
0!
0'
0/
#284110000000
1!
1'
1/
#284120000000
0!
0'
0/
#284130000000
1!
1'
1/
#284140000000
0!
0'
0/
#284150000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#284160000000
0!
0'
0/
#284170000000
1!
1'
1/
#284180000000
0!
0'
0/
#284190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#284200000000
0!
0'
0/
#284210000000
1!
1'
1/
#284220000000
0!
0'
0/
#284230000000
#284240000000
1!
1'
1/
#284250000000
0!
0'
0/
#284260000000
1!
1'
1/
#284270000000
0!
1"
0'
1(
0/
10
#284280000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#284290000000
0!
0'
0/
#284300000000
1!
1'
1/
#284310000000
0!
0'
0/
#284320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#284330000000
0!
0'
0/
#284340000000
1!
1'
1/
#284350000000
0!
1"
0'
1(
0/
10
#284360000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#284370000000
0!
1$
0'
1+
0/
#284380000000
1!
1'
1/
#284390000000
0!
0'
0/
#284400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#284410000000
0!
0'
0/
#284420000000
1!
1'
1/
#284430000000
0!
0'
0/
#284440000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#284450000000
0!
0'
0/
#284460000000
1!
1'
1/
#284470000000
0!
0'
0/
#284480000000
1!
1'
1/
#284490000000
0!
0'
0/
#284500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#284510000000
0!
0'
0/
#284520000000
1!
1'
1/
#284530000000
0!
0'
0/
#284540000000
1!
1'
1/
#284550000000
0!
0'
0/
#284560000000
1!
1'
1/
#284570000000
0!
0'
0/
#284580000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#284590000000
0!
0'
0/
#284600000000
1!
1'
1/
#284610000000
0!
0'
0/
#284620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#284630000000
0!
0'
0/
#284640000000
1!
1'
1/
#284650000000
0!
0'
0/
#284660000000
#284670000000
1!
1'
1/
#284680000000
0!
0'
0/
#284690000000
1!
1'
1/
#284700000000
0!
1"
0'
1(
0/
10
#284710000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#284720000000
0!
0'
0/
#284730000000
1!
1'
1/
#284740000000
0!
0'
0/
#284750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#284760000000
0!
0'
0/
#284770000000
1!
1'
1/
#284780000000
0!
1"
0'
1(
0/
10
#284790000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#284800000000
0!
1$
0'
1+
0/
#284810000000
1!
1'
1/
#284820000000
0!
0'
0/
#284830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#284840000000
0!
0'
0/
#284850000000
1!
1'
1/
#284860000000
0!
0'
0/
#284870000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#284880000000
0!
0'
0/
#284890000000
1!
1'
1/
#284900000000
0!
0'
0/
#284910000000
1!
1'
1/
#284920000000
0!
0'
0/
#284930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#284940000000
0!
0'
0/
#284950000000
1!
1'
1/
#284960000000
0!
0'
0/
#284970000000
1!
1'
1/
#284980000000
0!
0'
0/
#284990000000
1!
1'
1/
#285000000000
0!
0'
0/
#285010000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#285020000000
0!
0'
0/
#285030000000
1!
1'
1/
#285040000000
0!
0'
0/
#285050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#285060000000
0!
0'
0/
#285070000000
1!
1'
1/
#285080000000
0!
0'
0/
#285090000000
#285100000000
1!
1'
1/
#285110000000
0!
0'
0/
#285120000000
1!
1'
1/
#285130000000
0!
1"
0'
1(
0/
10
#285140000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#285150000000
0!
0'
0/
#285160000000
1!
1'
1/
#285170000000
0!
0'
0/
#285180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#285190000000
0!
0'
0/
#285200000000
1!
1'
1/
#285210000000
0!
1"
0'
1(
0/
10
#285220000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#285230000000
0!
1$
0'
1+
0/
#285240000000
1!
1'
1/
#285250000000
0!
0'
0/
#285260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#285270000000
0!
0'
0/
#285280000000
1!
1'
1/
#285290000000
0!
0'
0/
#285300000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#285310000000
0!
0'
0/
#285320000000
1!
1'
1/
#285330000000
0!
0'
0/
#285340000000
1!
1'
1/
#285350000000
0!
0'
0/
#285360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#285370000000
0!
0'
0/
#285380000000
1!
1'
1/
#285390000000
0!
0'
0/
#285400000000
1!
1'
1/
#285410000000
0!
0'
0/
#285420000000
1!
1'
1/
#285430000000
0!
0'
0/
#285440000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#285450000000
0!
0'
0/
#285460000000
1!
1'
1/
#285470000000
0!
0'
0/
#285480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#285490000000
0!
0'
0/
#285500000000
1!
1'
1/
#285510000000
0!
0'
0/
#285520000000
#285530000000
1!
1'
1/
#285540000000
0!
0'
0/
#285550000000
1!
1'
1/
#285560000000
0!
1"
0'
1(
0/
10
#285570000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#285580000000
0!
0'
0/
#285590000000
1!
1'
1/
#285600000000
0!
0'
0/
#285610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#285620000000
0!
0'
0/
#285630000000
1!
1'
1/
#285640000000
0!
1"
0'
1(
0/
10
#285650000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#285660000000
0!
1$
0'
1+
0/
#285670000000
1!
1'
1/
#285680000000
0!
0'
0/
#285690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#285700000000
0!
0'
0/
#285710000000
1!
1'
1/
#285720000000
0!
0'
0/
#285730000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#285740000000
0!
0'
0/
#285750000000
1!
1'
1/
#285760000000
0!
0'
0/
#285770000000
1!
1'
1/
#285780000000
0!
0'
0/
#285790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#285800000000
0!
0'
0/
#285810000000
1!
1'
1/
#285820000000
0!
0'
0/
#285830000000
1!
1'
1/
#285840000000
0!
0'
0/
#285850000000
1!
1'
1/
#285860000000
0!
0'
0/
#285870000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#285880000000
0!
0'
0/
#285890000000
1!
1'
1/
#285900000000
0!
0'
0/
#285910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#285920000000
0!
0'
0/
#285930000000
1!
1'
1/
#285940000000
0!
0'
0/
#285950000000
#285960000000
1!
1'
1/
#285970000000
0!
0'
0/
#285980000000
1!
1'
1/
#285990000000
0!
1"
0'
1(
0/
10
#286000000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#286010000000
0!
0'
0/
#286020000000
1!
1'
1/
#286030000000
0!
0'
0/
#286040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#286050000000
0!
0'
0/
#286060000000
1!
1'
1/
#286070000000
0!
1"
0'
1(
0/
10
#286080000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#286090000000
0!
1$
0'
1+
0/
#286100000000
1!
1'
1/
#286110000000
0!
0'
0/
#286120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#286130000000
0!
0'
0/
#286140000000
1!
1'
1/
#286150000000
0!
0'
0/
#286160000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#286170000000
0!
0'
0/
#286180000000
1!
1'
1/
#286190000000
0!
0'
0/
#286200000000
1!
1'
1/
#286210000000
0!
0'
0/
#286220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#286230000000
0!
0'
0/
#286240000000
1!
1'
1/
#286250000000
0!
0'
0/
#286260000000
1!
1'
1/
#286270000000
0!
0'
0/
#286280000000
1!
1'
1/
#286290000000
0!
0'
0/
#286300000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#286310000000
0!
0'
0/
#286320000000
1!
1'
1/
#286330000000
0!
0'
0/
#286340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#286350000000
0!
0'
0/
#286360000000
1!
1'
1/
#286370000000
0!
0'
0/
#286380000000
#286390000000
1!
1'
1/
#286400000000
0!
0'
0/
#286410000000
1!
1'
1/
#286420000000
0!
1"
0'
1(
0/
10
#286430000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#286440000000
0!
0'
0/
#286450000000
1!
1'
1/
#286460000000
0!
0'
0/
#286470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#286480000000
0!
0'
0/
#286490000000
1!
1'
1/
#286500000000
0!
1"
0'
1(
0/
10
#286510000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#286520000000
0!
1$
0'
1+
0/
#286530000000
1!
1'
1/
#286540000000
0!
0'
0/
#286550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#286560000000
0!
0'
0/
#286570000000
1!
1'
1/
#286580000000
0!
0'
0/
#286590000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#286600000000
0!
0'
0/
#286610000000
1!
1'
1/
#286620000000
0!
0'
0/
#286630000000
1!
1'
1/
#286640000000
0!
0'
0/
#286650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#286660000000
0!
0'
0/
#286670000000
1!
1'
1/
#286680000000
0!
0'
0/
#286690000000
1!
1'
1/
#286700000000
0!
0'
0/
#286710000000
1!
1'
1/
#286720000000
0!
0'
0/
#286730000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#286740000000
0!
0'
0/
#286750000000
1!
1'
1/
#286760000000
0!
0'
0/
#286770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#286780000000
0!
0'
0/
#286790000000
1!
1'
1/
#286800000000
0!
0'
0/
#286810000000
#286820000000
1!
1'
1/
#286830000000
0!
0'
0/
#286840000000
1!
1'
1/
#286850000000
0!
1"
0'
1(
0/
10
#286860000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#286870000000
0!
0'
0/
#286880000000
1!
1'
1/
#286890000000
0!
0'
0/
#286900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#286910000000
0!
0'
0/
#286920000000
1!
1'
1/
#286930000000
0!
1"
0'
1(
0/
10
#286940000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#286950000000
0!
1$
0'
1+
0/
#286960000000
1!
1'
1/
#286970000000
0!
0'
0/
#286980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#286990000000
0!
0'
0/
#287000000000
1!
1'
1/
#287010000000
0!
0'
0/
#287020000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#287030000000
0!
0'
0/
#287040000000
1!
1'
1/
#287050000000
0!
0'
0/
#287060000000
1!
1'
1/
#287070000000
0!
0'
0/
#287080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#287090000000
0!
0'
0/
#287100000000
1!
1'
1/
#287110000000
0!
0'
0/
#287120000000
1!
1'
1/
#287130000000
0!
0'
0/
#287140000000
1!
1'
1/
#287150000000
0!
0'
0/
#287160000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#287170000000
0!
0'
0/
#287180000000
1!
1'
1/
#287190000000
0!
0'
0/
#287200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#287210000000
0!
0'
0/
#287220000000
1!
1'
1/
#287230000000
0!
0'
0/
#287240000000
#287250000000
1!
1'
1/
#287260000000
0!
0'
0/
#287270000000
1!
1'
1/
#287280000000
0!
1"
0'
1(
0/
10
#287290000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#287300000000
0!
0'
0/
#287310000000
1!
1'
1/
#287320000000
0!
0'
0/
#287330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#287340000000
0!
0'
0/
#287350000000
1!
1'
1/
#287360000000
0!
1"
0'
1(
0/
10
#287370000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#287380000000
0!
1$
0'
1+
0/
#287390000000
1!
1'
1/
#287400000000
0!
0'
0/
#287410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#287420000000
0!
0'
0/
#287430000000
1!
1'
1/
#287440000000
0!
0'
0/
#287450000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#287460000000
0!
0'
0/
#287470000000
1!
1'
1/
#287480000000
0!
0'
0/
#287490000000
1!
1'
1/
#287500000000
0!
0'
0/
#287510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#287520000000
0!
0'
0/
#287530000000
1!
1'
1/
#287540000000
0!
0'
0/
#287550000000
1!
1'
1/
#287560000000
0!
0'
0/
#287570000000
1!
1'
1/
#287580000000
0!
0'
0/
#287590000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#287600000000
0!
0'
0/
#287610000000
1!
1'
1/
#287620000000
0!
0'
0/
#287630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#287640000000
0!
0'
0/
#287650000000
1!
1'
1/
#287660000000
0!
0'
0/
#287670000000
#287680000000
1!
1'
1/
#287690000000
0!
0'
0/
#287700000000
1!
1'
1/
#287710000000
0!
1"
0'
1(
0/
10
#287720000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#287730000000
0!
0'
0/
#287740000000
1!
1'
1/
#287750000000
0!
0'
0/
#287760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#287770000000
0!
0'
0/
#287780000000
1!
1'
1/
#287790000000
0!
1"
0'
1(
0/
10
#287800000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#287810000000
0!
1$
0'
1+
0/
#287820000000
1!
1'
1/
#287830000000
0!
0'
0/
#287840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#287850000000
0!
0'
0/
#287860000000
1!
1'
1/
#287870000000
0!
0'
0/
#287880000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#287890000000
0!
0'
0/
#287900000000
1!
1'
1/
#287910000000
0!
0'
0/
#287920000000
1!
1'
1/
#287930000000
0!
0'
0/
#287940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#287950000000
0!
0'
0/
#287960000000
1!
1'
1/
#287970000000
0!
0'
0/
#287980000000
1!
1'
1/
#287990000000
0!
0'
0/
#288000000000
1!
1'
1/
#288010000000
0!
0'
0/
#288020000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#288030000000
0!
0'
0/
#288040000000
1!
1'
1/
#288050000000
0!
0'
0/
#288060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#288070000000
0!
0'
0/
#288080000000
1!
1'
1/
#288090000000
0!
0'
0/
#288100000000
#288110000000
1!
1'
1/
#288120000000
0!
0'
0/
#288130000000
1!
1'
1/
#288140000000
0!
1"
0'
1(
0/
10
#288150000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#288160000000
0!
0'
0/
#288170000000
1!
1'
1/
#288180000000
0!
0'
0/
#288190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#288200000000
0!
0'
0/
#288210000000
1!
1'
1/
#288220000000
0!
1"
0'
1(
0/
10
#288230000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#288240000000
0!
1$
0'
1+
0/
#288250000000
1!
1'
1/
#288260000000
0!
0'
0/
#288270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#288280000000
0!
0'
0/
#288290000000
1!
1'
1/
#288300000000
0!
0'
0/
#288310000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#288320000000
0!
0'
0/
#288330000000
1!
1'
1/
#288340000000
0!
0'
0/
#288350000000
1!
1'
1/
#288360000000
0!
0'
0/
#288370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#288380000000
0!
0'
0/
#288390000000
1!
1'
1/
#288400000000
0!
0'
0/
#288410000000
1!
1'
1/
#288420000000
0!
0'
0/
#288430000000
1!
1'
1/
#288440000000
0!
0'
0/
#288450000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#288460000000
0!
0'
0/
#288470000000
1!
1'
1/
#288480000000
0!
0'
0/
#288490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#288500000000
0!
0'
0/
#288510000000
1!
1'
1/
#288520000000
0!
0'
0/
#288530000000
#288540000000
1!
1'
1/
#288550000000
0!
0'
0/
#288560000000
1!
1'
1/
#288570000000
0!
1"
0'
1(
0/
10
#288580000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#288590000000
0!
0'
0/
#288600000000
1!
1'
1/
#288610000000
0!
0'
0/
#288620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#288630000000
0!
0'
0/
#288640000000
1!
1'
1/
#288650000000
0!
1"
0'
1(
0/
10
#288660000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#288670000000
0!
1$
0'
1+
0/
#288680000000
1!
1'
1/
#288690000000
0!
0'
0/
#288700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#288710000000
0!
0'
0/
#288720000000
1!
1'
1/
#288730000000
0!
0'
0/
#288740000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#288750000000
0!
0'
0/
#288760000000
1!
1'
1/
#288770000000
0!
0'
0/
#288780000000
1!
1'
1/
#288790000000
0!
0'
0/
#288800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#288810000000
0!
0'
0/
#288820000000
1!
1'
1/
#288830000000
0!
0'
0/
#288840000000
1!
1'
1/
#288850000000
0!
0'
0/
#288860000000
1!
1'
1/
#288870000000
0!
0'
0/
#288880000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#288890000000
0!
0'
0/
#288900000000
1!
1'
1/
#288910000000
0!
0'
0/
#288920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#288930000000
0!
0'
0/
#288940000000
1!
1'
1/
#288950000000
0!
0'
0/
#288960000000
#288970000000
1!
1'
1/
#288980000000
0!
0'
0/
#288990000000
1!
1'
1/
#289000000000
0!
1"
0'
1(
0/
10
#289010000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#289020000000
0!
0'
0/
#289030000000
1!
1'
1/
#289040000000
0!
0'
0/
#289050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#289060000000
0!
0'
0/
#289070000000
1!
1'
1/
#289080000000
0!
1"
0'
1(
0/
10
#289090000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#289100000000
0!
1$
0'
1+
0/
#289110000000
1!
1'
1/
#289120000000
0!
0'
0/
#289130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#289140000000
0!
0'
0/
#289150000000
1!
1'
1/
#289160000000
0!
0'
0/
#289170000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#289180000000
0!
0'
0/
#289190000000
1!
1'
1/
#289200000000
0!
0'
0/
#289210000000
1!
1'
1/
#289220000000
0!
0'
0/
#289230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#289240000000
0!
0'
0/
#289250000000
1!
1'
1/
#289260000000
0!
0'
0/
#289270000000
1!
1'
1/
#289280000000
0!
0'
0/
#289290000000
1!
1'
1/
#289300000000
0!
0'
0/
#289310000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#289320000000
0!
0'
0/
#289330000000
1!
1'
1/
#289340000000
0!
0'
0/
#289350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#289360000000
0!
0'
0/
#289370000000
1!
1'
1/
#289380000000
0!
0'
0/
#289390000000
#289400000000
1!
1'
1/
#289410000000
0!
0'
0/
#289420000000
1!
1'
1/
#289430000000
0!
1"
0'
1(
0/
10
#289440000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#289450000000
0!
0'
0/
#289460000000
1!
1'
1/
#289470000000
0!
0'
0/
#289480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#289490000000
0!
0'
0/
#289500000000
1!
1'
1/
#289510000000
0!
1"
0'
1(
0/
10
#289520000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#289530000000
0!
1$
0'
1+
0/
#289540000000
1!
1'
1/
#289550000000
0!
0'
0/
#289560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#289570000000
0!
0'
0/
#289580000000
1!
1'
1/
#289590000000
0!
0'
0/
#289600000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#289610000000
0!
0'
0/
#289620000000
1!
1'
1/
#289630000000
0!
0'
0/
#289640000000
1!
1'
1/
#289650000000
0!
0'
0/
#289660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#289670000000
0!
0'
0/
#289680000000
1!
1'
1/
#289690000000
0!
0'
0/
#289700000000
1!
1'
1/
#289710000000
0!
0'
0/
#289720000000
1!
1'
1/
#289730000000
0!
0'
0/
#289740000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#289750000000
0!
0'
0/
#289760000000
1!
1'
1/
#289770000000
0!
0'
0/
#289780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#289790000000
0!
0'
0/
#289800000000
1!
1'
1/
#289810000000
0!
0'
0/
#289820000000
#289830000000
1!
1'
1/
#289840000000
0!
0'
0/
#289850000000
1!
1'
1/
#289860000000
0!
1"
0'
1(
0/
10
#289870000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#289880000000
0!
0'
0/
#289890000000
1!
1'
1/
#289900000000
0!
0'
0/
#289910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#289920000000
0!
0'
0/
#289930000000
1!
1'
1/
#289940000000
0!
1"
0'
1(
0/
10
#289950000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#289960000000
0!
1$
0'
1+
0/
#289970000000
1!
1'
1/
#289980000000
0!
0'
0/
#289990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#290000000000
0!
0'
0/
#290010000000
1!
1'
1/
#290020000000
0!
0'
0/
#290030000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#290040000000
0!
0'
0/
#290050000000
1!
1'
1/
#290060000000
0!
0'
0/
#290070000000
1!
1'
1/
#290080000000
0!
0'
0/
#290090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#290100000000
0!
0'
0/
#290110000000
1!
1'
1/
#290120000000
0!
0'
0/
#290130000000
1!
1'
1/
#290140000000
0!
0'
0/
#290150000000
1!
1'
1/
#290160000000
0!
0'
0/
#290170000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#290180000000
0!
0'
0/
#290190000000
1!
1'
1/
#290200000000
0!
0'
0/
#290210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#290220000000
0!
0'
0/
#290230000000
1!
1'
1/
#290240000000
0!
0'
0/
#290250000000
#290260000000
1!
1'
1/
#290270000000
0!
0'
0/
#290280000000
1!
1'
1/
#290290000000
0!
1"
0'
1(
0/
10
#290300000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#290310000000
0!
0'
0/
#290320000000
1!
1'
1/
#290330000000
0!
0'
0/
#290340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#290350000000
0!
0'
0/
#290360000000
1!
1'
1/
#290370000000
0!
1"
0'
1(
0/
10
#290380000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#290390000000
0!
1$
0'
1+
0/
#290400000000
1!
1'
1/
#290410000000
0!
0'
0/
#290420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#290430000000
0!
0'
0/
#290440000000
1!
1'
1/
#290450000000
0!
0'
0/
#290460000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#290470000000
0!
0'
0/
#290480000000
1!
1'
1/
#290490000000
0!
0'
0/
#290500000000
1!
1'
1/
#290510000000
0!
0'
0/
#290520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#290530000000
0!
0'
0/
#290540000000
1!
1'
1/
#290550000000
0!
0'
0/
#290560000000
1!
1'
1/
#290570000000
0!
0'
0/
#290580000000
1!
1'
1/
#290590000000
0!
0'
0/
#290600000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#290610000000
0!
0'
0/
#290620000000
1!
1'
1/
#290630000000
0!
0'
0/
#290640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#290650000000
0!
0'
0/
#290660000000
1!
1'
1/
#290670000000
0!
0'
0/
#290680000000
#290690000000
1!
1'
1/
#290700000000
0!
0'
0/
#290710000000
1!
1'
1/
#290720000000
0!
1"
0'
1(
0/
10
#290730000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#290740000000
0!
0'
0/
#290750000000
1!
1'
1/
#290760000000
0!
0'
0/
#290770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#290780000000
0!
0'
0/
#290790000000
1!
1'
1/
#290800000000
0!
1"
0'
1(
0/
10
#290810000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#290820000000
0!
1$
0'
1+
0/
#290830000000
1!
1'
1/
#290840000000
0!
0'
0/
#290850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#290860000000
0!
0'
0/
#290870000000
1!
1'
1/
#290880000000
0!
0'
0/
#290890000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#290900000000
0!
0'
0/
#290910000000
1!
1'
1/
#290920000000
0!
0'
0/
#290930000000
1!
1'
1/
#290940000000
0!
0'
0/
#290950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#290960000000
0!
0'
0/
#290970000000
1!
1'
1/
#290980000000
0!
0'
0/
#290990000000
1!
1'
1/
#291000000000
0!
0'
0/
#291010000000
1!
1'
1/
#291020000000
0!
0'
0/
#291030000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#291040000000
0!
0'
0/
#291050000000
1!
1'
1/
#291060000000
0!
0'
0/
#291070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#291080000000
0!
0'
0/
#291090000000
1!
1'
1/
#291100000000
0!
0'
0/
#291110000000
#291120000000
1!
1'
1/
#291130000000
0!
0'
0/
#291140000000
1!
1'
1/
#291150000000
0!
1"
0'
1(
0/
10
#291160000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#291170000000
0!
0'
0/
#291180000000
1!
1'
1/
#291190000000
0!
0'
0/
#291200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#291210000000
0!
0'
0/
#291220000000
1!
1'
1/
#291230000000
0!
1"
0'
1(
0/
10
#291240000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#291250000000
0!
1$
0'
1+
0/
#291260000000
1!
1'
1/
#291270000000
0!
0'
0/
#291280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#291290000000
0!
0'
0/
#291300000000
1!
1'
1/
#291310000000
0!
0'
0/
#291320000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#291330000000
0!
0'
0/
#291340000000
1!
1'
1/
#291350000000
0!
0'
0/
#291360000000
1!
1'
1/
#291370000000
0!
0'
0/
#291380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#291390000000
0!
0'
0/
#291400000000
1!
1'
1/
#291410000000
0!
0'
0/
#291420000000
1!
1'
1/
#291430000000
0!
0'
0/
#291440000000
1!
1'
1/
#291450000000
0!
0'
0/
#291460000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#291470000000
0!
0'
0/
#291480000000
1!
1'
1/
#291490000000
0!
0'
0/
#291500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#291510000000
0!
0'
0/
#291520000000
1!
1'
1/
#291530000000
0!
0'
0/
#291540000000
#291550000000
1!
1'
1/
#291560000000
0!
0'
0/
#291570000000
1!
1'
1/
#291580000000
0!
1"
0'
1(
0/
10
#291590000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#291600000000
0!
0'
0/
#291610000000
1!
1'
1/
#291620000000
0!
0'
0/
#291630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#291640000000
0!
0'
0/
#291650000000
1!
1'
1/
#291660000000
0!
1"
0'
1(
0/
10
#291670000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#291680000000
0!
1$
0'
1+
0/
#291690000000
1!
1'
1/
#291700000000
0!
0'
0/
#291710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#291720000000
0!
0'
0/
#291730000000
1!
1'
1/
#291740000000
0!
0'
0/
#291750000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#291760000000
0!
0'
0/
#291770000000
1!
1'
1/
#291780000000
0!
0'
0/
#291790000000
1!
1'
1/
#291800000000
0!
0'
0/
#291810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#291820000000
0!
0'
0/
#291830000000
1!
1'
1/
#291840000000
0!
0'
0/
#291850000000
1!
1'
1/
#291860000000
0!
0'
0/
#291870000000
1!
1'
1/
#291880000000
0!
0'
0/
#291890000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#291900000000
0!
0'
0/
#291910000000
1!
1'
1/
#291920000000
0!
0'
0/
#291930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#291940000000
0!
0'
0/
#291950000000
1!
1'
1/
#291960000000
0!
0'
0/
#291970000000
#291980000000
1!
1'
1/
#291990000000
0!
0'
0/
#292000000000
1!
1'
1/
#292010000000
0!
1"
0'
1(
0/
10
#292020000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#292030000000
0!
0'
0/
#292040000000
1!
1'
1/
#292050000000
0!
0'
0/
#292060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#292070000000
0!
0'
0/
#292080000000
1!
1'
1/
#292090000000
0!
1"
0'
1(
0/
10
#292100000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#292110000000
0!
1$
0'
1+
0/
#292120000000
1!
1'
1/
#292130000000
0!
0'
0/
#292140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#292150000000
0!
0'
0/
#292160000000
1!
1'
1/
#292170000000
0!
0'
0/
#292180000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#292190000000
0!
0'
0/
#292200000000
1!
1'
1/
#292210000000
0!
0'
0/
#292220000000
1!
1'
1/
#292230000000
0!
0'
0/
#292240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#292250000000
0!
0'
0/
#292260000000
1!
1'
1/
#292270000000
0!
0'
0/
#292280000000
1!
1'
1/
#292290000000
0!
0'
0/
#292300000000
1!
1'
1/
#292310000000
0!
0'
0/
#292320000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#292330000000
0!
0'
0/
#292340000000
1!
1'
1/
#292350000000
0!
0'
0/
#292360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#292370000000
0!
0'
0/
#292380000000
1!
1'
1/
#292390000000
0!
0'
0/
#292400000000
#292410000000
1!
1'
1/
#292420000000
0!
0'
0/
#292430000000
1!
1'
1/
#292440000000
0!
1"
0'
1(
0/
10
#292450000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#292460000000
0!
0'
0/
#292470000000
1!
1'
1/
#292480000000
0!
0'
0/
#292490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#292500000000
0!
0'
0/
#292510000000
1!
1'
1/
#292520000000
0!
1"
0'
1(
0/
10
#292530000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#292540000000
0!
1$
0'
1+
0/
#292550000000
1!
1'
1/
#292560000000
0!
0'
0/
#292570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#292580000000
0!
0'
0/
#292590000000
1!
1'
1/
#292600000000
0!
0'
0/
#292610000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#292620000000
0!
0'
0/
#292630000000
1!
1'
1/
#292640000000
0!
0'
0/
#292650000000
1!
1'
1/
#292660000000
0!
0'
0/
#292670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#292680000000
0!
0'
0/
#292690000000
1!
1'
1/
#292700000000
0!
0'
0/
#292710000000
1!
1'
1/
#292720000000
0!
0'
0/
#292730000000
1!
1'
1/
#292740000000
0!
0'
0/
#292750000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#292760000000
0!
0'
0/
#292770000000
1!
1'
1/
#292780000000
0!
0'
0/
#292790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#292800000000
0!
0'
0/
#292810000000
1!
1'
1/
#292820000000
0!
0'
0/
#292830000000
#292840000000
1!
1'
1/
#292850000000
0!
0'
0/
#292860000000
1!
1'
1/
#292870000000
0!
1"
0'
1(
0/
10
#292880000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#292890000000
0!
0'
0/
#292900000000
1!
1'
1/
#292910000000
0!
0'
0/
#292920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#292930000000
0!
0'
0/
#292940000000
1!
1'
1/
#292950000000
0!
1"
0'
1(
0/
10
#292960000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#292970000000
0!
1$
0'
1+
0/
#292980000000
1!
1'
1/
#292990000000
0!
0'
0/
#293000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#293010000000
0!
0'
0/
#293020000000
1!
1'
1/
#293030000000
0!
0'
0/
#293040000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#293050000000
0!
0'
0/
#293060000000
1!
1'
1/
#293070000000
0!
0'
0/
#293080000000
1!
1'
1/
#293090000000
0!
0'
0/
#293100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#293110000000
0!
0'
0/
#293120000000
1!
1'
1/
#293130000000
0!
0'
0/
#293140000000
1!
1'
1/
#293150000000
0!
0'
0/
#293160000000
1!
1'
1/
#293170000000
0!
0'
0/
#293180000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#293190000000
0!
0'
0/
#293200000000
1!
1'
1/
#293210000000
0!
0'
0/
#293220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#293230000000
0!
0'
0/
#293240000000
1!
1'
1/
#293250000000
0!
0'
0/
#293260000000
#293270000000
1!
1'
1/
#293280000000
0!
0'
0/
#293290000000
1!
1'
1/
#293300000000
0!
1"
0'
1(
0/
10
#293310000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#293320000000
0!
0'
0/
#293330000000
1!
1'
1/
#293340000000
0!
0'
0/
#293350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#293360000000
0!
0'
0/
#293370000000
1!
1'
1/
#293380000000
0!
1"
0'
1(
0/
10
#293390000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#293400000000
0!
1$
0'
1+
0/
#293410000000
1!
1'
1/
#293420000000
0!
0'
0/
#293430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#293440000000
0!
0'
0/
#293450000000
1!
1'
1/
#293460000000
0!
0'
0/
#293470000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#293480000000
0!
0'
0/
#293490000000
1!
1'
1/
#293500000000
0!
0'
0/
#293510000000
1!
1'
1/
#293520000000
0!
0'
0/
#293530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#293540000000
0!
0'
0/
#293550000000
1!
1'
1/
#293560000000
0!
0'
0/
#293570000000
1!
1'
1/
#293580000000
0!
0'
0/
#293590000000
1!
1'
1/
#293600000000
0!
0'
0/
#293610000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#293620000000
0!
0'
0/
#293630000000
1!
1'
1/
#293640000000
0!
0'
0/
#293650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#293660000000
0!
0'
0/
#293670000000
1!
1'
1/
#293680000000
0!
0'
0/
#293690000000
#293700000000
1!
1'
1/
#293710000000
0!
0'
0/
#293720000000
1!
1'
1/
#293730000000
0!
1"
0'
1(
0/
10
#293740000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#293750000000
0!
0'
0/
#293760000000
1!
1'
1/
#293770000000
0!
0'
0/
#293780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#293790000000
0!
0'
0/
#293800000000
1!
1'
1/
#293810000000
0!
1"
0'
1(
0/
10
#293820000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#293830000000
0!
1$
0'
1+
0/
#293840000000
1!
1'
1/
#293850000000
0!
0'
0/
#293860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#293870000000
0!
0'
0/
#293880000000
1!
1'
1/
#293890000000
0!
0'
0/
#293900000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#293910000000
0!
0'
0/
#293920000000
1!
1'
1/
#293930000000
0!
0'
0/
#293940000000
1!
1'
1/
#293950000000
0!
0'
0/
#293960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#293970000000
0!
0'
0/
#293980000000
1!
1'
1/
#293990000000
0!
0'
0/
#294000000000
1!
1'
1/
#294010000000
0!
0'
0/
#294020000000
1!
1'
1/
#294030000000
0!
0'
0/
#294040000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#294050000000
0!
0'
0/
#294060000000
1!
1'
1/
#294070000000
0!
0'
0/
#294080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#294090000000
0!
0'
0/
#294100000000
1!
1'
1/
#294110000000
0!
0'
0/
#294120000000
#294130000000
1!
1'
1/
#294140000000
0!
0'
0/
#294150000000
1!
1'
1/
#294160000000
0!
1"
0'
1(
0/
10
#294170000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#294180000000
0!
0'
0/
#294190000000
1!
1'
1/
#294200000000
0!
0'
0/
#294210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#294220000000
0!
0'
0/
#294230000000
1!
1'
1/
#294240000000
0!
1"
0'
1(
0/
10
#294250000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#294260000000
0!
1$
0'
1+
0/
#294270000000
1!
1'
1/
#294280000000
0!
0'
0/
#294290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#294300000000
0!
0'
0/
#294310000000
1!
1'
1/
#294320000000
0!
0'
0/
#294330000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#294340000000
0!
0'
0/
#294350000000
1!
1'
1/
#294360000000
0!
0'
0/
#294370000000
1!
1'
1/
#294380000000
0!
0'
0/
#294390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#294400000000
0!
0'
0/
#294410000000
1!
1'
1/
#294420000000
0!
0'
0/
#294430000000
1!
1'
1/
#294440000000
0!
0'
0/
#294450000000
1!
1'
1/
#294460000000
0!
0'
0/
#294470000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#294480000000
0!
0'
0/
#294490000000
1!
1'
1/
#294500000000
0!
0'
0/
#294510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#294520000000
0!
0'
0/
#294530000000
1!
1'
1/
#294540000000
0!
0'
0/
#294550000000
#294560000000
1!
1'
1/
#294570000000
0!
0'
0/
#294580000000
1!
1'
1/
#294590000000
0!
1"
0'
1(
0/
10
#294600000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#294610000000
0!
0'
0/
#294620000000
1!
1'
1/
#294630000000
0!
0'
0/
#294640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#294650000000
0!
0'
0/
#294660000000
1!
1'
1/
#294670000000
0!
1"
0'
1(
0/
10
#294680000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#294690000000
0!
1$
0'
1+
0/
#294700000000
1!
1'
1/
#294710000000
0!
0'
0/
#294720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#294730000000
0!
0'
0/
#294740000000
1!
1'
1/
#294750000000
0!
0'
0/
#294760000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#294770000000
0!
0'
0/
#294780000000
1!
1'
1/
#294790000000
0!
0'
0/
#294800000000
1!
1'
1/
#294810000000
0!
0'
0/
#294820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#294830000000
0!
0'
0/
#294840000000
1!
1'
1/
#294850000000
0!
0'
0/
#294860000000
1!
1'
1/
#294870000000
0!
0'
0/
#294880000000
1!
1'
1/
#294890000000
0!
0'
0/
#294900000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#294910000000
0!
0'
0/
#294920000000
1!
1'
1/
#294930000000
0!
0'
0/
#294940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#294950000000
0!
0'
0/
#294960000000
1!
1'
1/
#294970000000
0!
0'
0/
#294980000000
#294990000000
1!
1'
1/
#295000000000
0!
0'
0/
#295010000000
1!
1'
1/
#295020000000
0!
1"
0'
1(
0/
10
#295030000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#295040000000
0!
0'
0/
#295050000000
1!
1'
1/
#295060000000
0!
0'
0/
#295070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#295080000000
0!
0'
0/
#295090000000
1!
1'
1/
#295100000000
0!
1"
0'
1(
0/
10
#295110000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#295120000000
0!
1$
0'
1+
0/
#295130000000
1!
1'
1/
#295140000000
0!
0'
0/
#295150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#295160000000
0!
0'
0/
#295170000000
1!
1'
1/
#295180000000
0!
0'
0/
#295190000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#295200000000
0!
0'
0/
#295210000000
1!
1'
1/
#295220000000
0!
0'
0/
#295230000000
1!
1'
1/
#295240000000
0!
0'
0/
#295250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#295260000000
0!
0'
0/
#295270000000
1!
1'
1/
#295280000000
0!
0'
0/
#295290000000
1!
1'
1/
#295300000000
0!
0'
0/
#295310000000
1!
1'
1/
#295320000000
0!
0'
0/
#295330000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#295340000000
0!
0'
0/
#295350000000
1!
1'
1/
#295360000000
0!
0'
0/
#295370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#295380000000
0!
0'
0/
#295390000000
1!
1'
1/
#295400000000
0!
0'
0/
#295410000000
#295420000000
1!
1'
1/
#295430000000
0!
0'
0/
#295440000000
1!
1'
1/
#295450000000
0!
1"
0'
1(
0/
10
#295460000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#295470000000
0!
0'
0/
#295480000000
1!
1'
1/
#295490000000
0!
0'
0/
#295500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#295510000000
0!
0'
0/
#295520000000
1!
1'
1/
#295530000000
0!
1"
0'
1(
0/
10
#295540000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#295550000000
0!
1$
0'
1+
0/
#295560000000
1!
1'
1/
#295570000000
0!
0'
0/
#295580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#295590000000
0!
0'
0/
#295600000000
1!
1'
1/
#295610000000
0!
0'
0/
#295620000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#295630000000
0!
0'
0/
#295640000000
1!
1'
1/
#295650000000
0!
0'
0/
#295660000000
1!
1'
1/
#295670000000
0!
0'
0/
#295680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#295690000000
0!
0'
0/
#295700000000
1!
1'
1/
#295710000000
0!
0'
0/
#295720000000
1!
1'
1/
#295730000000
0!
0'
0/
#295740000000
1!
1'
1/
#295750000000
0!
0'
0/
#295760000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#295770000000
0!
0'
0/
#295780000000
1!
1'
1/
#295790000000
0!
0'
0/
#295800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#295810000000
0!
0'
0/
#295820000000
1!
1'
1/
#295830000000
0!
0'
0/
#295840000000
#295850000000
1!
1'
1/
#295860000000
0!
0'
0/
#295870000000
1!
1'
1/
#295880000000
0!
1"
0'
1(
0/
10
#295890000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#295900000000
0!
0'
0/
#295910000000
1!
1'
1/
#295920000000
0!
0'
0/
#295930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#295940000000
0!
0'
0/
#295950000000
1!
1'
1/
#295960000000
0!
1"
0'
1(
0/
10
#295970000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#295980000000
0!
1$
0'
1+
0/
#295990000000
1!
1'
1/
#296000000000
0!
0'
0/
#296010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#296020000000
0!
0'
0/
#296030000000
1!
1'
1/
#296040000000
0!
0'
0/
#296050000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#296060000000
0!
0'
0/
#296070000000
1!
1'
1/
#296080000000
0!
0'
0/
#296090000000
1!
1'
1/
#296100000000
0!
0'
0/
#296110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#296120000000
0!
0'
0/
#296130000000
1!
1'
1/
#296140000000
0!
0'
0/
#296150000000
1!
1'
1/
#296160000000
0!
0'
0/
#296170000000
1!
1'
1/
#296180000000
0!
0'
0/
#296190000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#296200000000
0!
0'
0/
#296210000000
1!
1'
1/
#296220000000
0!
0'
0/
#296230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#296240000000
0!
0'
0/
#296250000000
1!
1'
1/
#296260000000
0!
0'
0/
#296270000000
#296280000000
1!
1'
1/
#296290000000
0!
0'
0/
#296300000000
1!
1'
1/
#296310000000
0!
1"
0'
1(
0/
10
#296320000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#296330000000
0!
0'
0/
#296340000000
1!
1'
1/
#296350000000
0!
0'
0/
#296360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#296370000000
0!
0'
0/
#296380000000
1!
1'
1/
#296390000000
0!
1"
0'
1(
0/
10
#296400000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#296410000000
0!
1$
0'
1+
0/
#296420000000
1!
1'
1/
#296430000000
0!
0'
0/
#296440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#296450000000
0!
0'
0/
#296460000000
1!
1'
1/
#296470000000
0!
0'
0/
#296480000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#296490000000
0!
0'
0/
#296500000000
1!
1'
1/
#296510000000
0!
0'
0/
#296520000000
1!
1'
1/
#296530000000
0!
0'
0/
#296540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#296550000000
0!
0'
0/
#296560000000
1!
1'
1/
#296570000000
0!
0'
0/
#296580000000
1!
1'
1/
#296590000000
0!
0'
0/
#296600000000
1!
1'
1/
#296610000000
0!
0'
0/
#296620000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#296630000000
0!
0'
0/
#296640000000
1!
1'
1/
#296650000000
0!
0'
0/
#296660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#296670000000
0!
0'
0/
#296680000000
1!
1'
1/
#296690000000
0!
0'
0/
#296700000000
#296710000000
1!
1'
1/
#296720000000
0!
0'
0/
#296730000000
1!
1'
1/
#296740000000
0!
1"
0'
1(
0/
10
#296750000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#296760000000
0!
0'
0/
#296770000000
1!
1'
1/
#296780000000
0!
0'
0/
#296790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#296800000000
0!
0'
0/
#296810000000
1!
1'
1/
#296820000000
0!
1"
0'
1(
0/
10
#296830000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#296840000000
0!
1$
0'
1+
0/
#296850000000
1!
1'
1/
#296860000000
0!
0'
0/
#296870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#296880000000
0!
0'
0/
#296890000000
1!
1'
1/
#296900000000
0!
0'
0/
#296910000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#296920000000
0!
0'
0/
#296930000000
1!
1'
1/
#296940000000
0!
0'
0/
#296950000000
1!
1'
1/
#296960000000
0!
0'
0/
#296970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#296980000000
0!
0'
0/
#296990000000
1!
1'
1/
#297000000000
0!
0'
0/
#297010000000
1!
1'
1/
#297020000000
0!
0'
0/
#297030000000
1!
1'
1/
#297040000000
0!
0'
0/
#297050000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#297060000000
0!
0'
0/
#297070000000
1!
1'
1/
#297080000000
0!
0'
0/
#297090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#297100000000
0!
0'
0/
#297110000000
1!
1'
1/
#297120000000
0!
0'
0/
#297130000000
#297140000000
1!
1'
1/
#297150000000
0!
0'
0/
#297160000000
1!
1'
1/
#297170000000
0!
1"
0'
1(
0/
10
#297180000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#297190000000
0!
0'
0/
#297200000000
1!
1'
1/
#297210000000
0!
0'
0/
#297220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#297230000000
0!
0'
0/
#297240000000
1!
1'
1/
#297250000000
0!
1"
0'
1(
0/
10
#297260000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#297270000000
0!
1$
0'
1+
0/
#297280000000
1!
1'
1/
#297290000000
0!
0'
0/
#297300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#297310000000
0!
0'
0/
#297320000000
1!
1'
1/
#297330000000
0!
0'
0/
#297340000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#297350000000
0!
0'
0/
#297360000000
1!
1'
1/
#297370000000
0!
0'
0/
#297380000000
1!
1'
1/
#297390000000
0!
0'
0/
#297400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#297410000000
0!
0'
0/
#297420000000
1!
1'
1/
#297430000000
0!
0'
0/
#297440000000
1!
1'
1/
#297450000000
0!
0'
0/
#297460000000
1!
1'
1/
#297470000000
0!
0'
0/
#297480000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#297490000000
0!
0'
0/
#297500000000
1!
1'
1/
#297510000000
0!
0'
0/
#297520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#297530000000
0!
0'
0/
#297540000000
1!
1'
1/
#297550000000
0!
0'
0/
#297560000000
#297570000000
1!
1'
1/
#297580000000
0!
0'
0/
#297590000000
1!
1'
1/
#297600000000
0!
1"
0'
1(
0/
10
#297610000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#297620000000
0!
0'
0/
#297630000000
1!
1'
1/
#297640000000
0!
0'
0/
#297650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#297660000000
0!
0'
0/
#297670000000
1!
1'
1/
#297680000000
0!
1"
0'
1(
0/
10
#297690000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#297700000000
0!
1$
0'
1+
0/
#297710000000
1!
1'
1/
#297720000000
0!
0'
0/
#297730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#297740000000
0!
0'
0/
#297750000000
1!
1'
1/
#297760000000
0!
0'
0/
#297770000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#297780000000
0!
0'
0/
#297790000000
1!
1'
1/
#297800000000
0!
0'
0/
#297810000000
1!
1'
1/
#297820000000
0!
0'
0/
#297830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#297840000000
0!
0'
0/
#297850000000
1!
1'
1/
#297860000000
0!
0'
0/
#297870000000
1!
1'
1/
#297880000000
0!
0'
0/
#297890000000
1!
1'
1/
#297900000000
0!
0'
0/
#297910000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#297920000000
0!
0'
0/
#297930000000
1!
1'
1/
#297940000000
0!
0'
0/
#297950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#297960000000
0!
0'
0/
#297970000000
1!
1'
1/
#297980000000
0!
0'
0/
#297990000000
#298000000000
1!
1'
1/
#298010000000
0!
0'
0/
#298020000000
1!
1'
1/
#298030000000
0!
1"
0'
1(
0/
10
#298040000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#298050000000
0!
0'
0/
#298060000000
1!
1'
1/
#298070000000
0!
0'
0/
#298080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#298090000000
0!
0'
0/
#298100000000
1!
1'
1/
#298110000000
0!
1"
0'
1(
0/
10
#298120000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#298130000000
0!
1$
0'
1+
0/
#298140000000
1!
1'
1/
#298150000000
0!
0'
0/
#298160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#298170000000
0!
0'
0/
#298180000000
1!
1'
1/
#298190000000
0!
0'
0/
#298200000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#298210000000
0!
0'
0/
#298220000000
1!
1'
1/
#298230000000
0!
0'
0/
#298240000000
1!
1'
1/
#298250000000
0!
0'
0/
#298260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#298270000000
0!
0'
0/
#298280000000
1!
1'
1/
#298290000000
0!
0'
0/
#298300000000
1!
1'
1/
#298310000000
0!
0'
0/
#298320000000
1!
1'
1/
#298330000000
0!
0'
0/
#298340000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#298350000000
0!
0'
0/
#298360000000
1!
1'
1/
#298370000000
0!
0'
0/
#298380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#298390000000
0!
0'
0/
#298400000000
1!
1'
1/
#298410000000
0!
0'
0/
#298420000000
#298430000000
1!
1'
1/
#298440000000
0!
0'
0/
#298450000000
1!
1'
1/
#298460000000
0!
1"
0'
1(
0/
10
#298470000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#298480000000
0!
0'
0/
#298490000000
1!
1'
1/
#298500000000
0!
0'
0/
#298510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#298520000000
0!
0'
0/
#298530000000
1!
1'
1/
#298540000000
0!
1"
0'
1(
0/
10
#298550000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#298560000000
0!
1$
0'
1+
0/
#298570000000
1!
1'
1/
#298580000000
0!
0'
0/
#298590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#298600000000
0!
0'
0/
#298610000000
1!
1'
1/
#298620000000
0!
0'
0/
#298630000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#298640000000
0!
0'
0/
#298650000000
1!
1'
1/
#298660000000
0!
0'
0/
#298670000000
1!
1'
1/
#298680000000
0!
0'
0/
#298690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#298700000000
0!
0'
0/
#298710000000
1!
1'
1/
#298720000000
0!
0'
0/
#298730000000
1!
1'
1/
#298740000000
0!
0'
0/
#298750000000
1!
1'
1/
#298760000000
0!
0'
0/
#298770000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#298780000000
0!
0'
0/
#298790000000
1!
1'
1/
#298800000000
0!
0'
0/
#298810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#298820000000
0!
0'
0/
#298830000000
1!
1'
1/
#298840000000
0!
0'
0/
#298850000000
#298860000000
1!
1'
1/
#298870000000
0!
0'
0/
#298880000000
1!
1'
1/
#298890000000
0!
1"
0'
1(
0/
10
#298900000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#298910000000
0!
0'
0/
#298920000000
1!
1'
1/
#298930000000
0!
0'
0/
#298940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#298950000000
0!
0'
0/
#298960000000
1!
1'
1/
#298970000000
0!
1"
0'
1(
0/
10
#298980000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#298990000000
0!
1$
0'
1+
0/
#299000000000
1!
1'
1/
#299010000000
0!
0'
0/
#299020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#299030000000
0!
0'
0/
#299040000000
1!
1'
1/
#299050000000
0!
0'
0/
#299060000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#299070000000
0!
0'
0/
#299080000000
1!
1'
1/
#299090000000
0!
0'
0/
#299100000000
1!
1'
1/
#299110000000
0!
0'
0/
#299120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#299130000000
0!
0'
0/
#299140000000
1!
1'
1/
#299150000000
0!
0'
0/
#299160000000
1!
1'
1/
#299170000000
0!
0'
0/
#299180000000
1!
1'
1/
#299190000000
0!
0'
0/
#299200000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#299210000000
0!
0'
0/
#299220000000
1!
1'
1/
#299230000000
0!
0'
0/
#299240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#299250000000
0!
0'
0/
#299260000000
1!
1'
1/
#299270000000
0!
0'
0/
#299280000000
#299290000000
1!
1'
1/
#299300000000
0!
0'
0/
#299310000000
1!
1'
1/
#299320000000
0!
1"
0'
1(
0/
10
#299330000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#299340000000
0!
0'
0/
#299350000000
1!
1'
1/
#299360000000
0!
0'
0/
#299370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#299380000000
0!
0'
0/
#299390000000
1!
1'
1/
#299400000000
0!
1"
0'
1(
0/
10
#299410000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#299420000000
0!
1$
0'
1+
0/
#299430000000
1!
1'
1/
#299440000000
0!
0'
0/
#299450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#299460000000
0!
0'
0/
#299470000000
1!
1'
1/
#299480000000
0!
0'
0/
#299490000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#299500000000
0!
0'
0/
#299510000000
1!
1'
1/
#299520000000
0!
0'
0/
#299530000000
1!
1'
1/
#299540000000
0!
0'
0/
#299550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#299560000000
0!
0'
0/
#299570000000
1!
1'
1/
#299580000000
0!
0'
0/
#299590000000
1!
1'
1/
#299600000000
0!
0'
0/
#299610000000
1!
1'
1/
#299620000000
0!
0'
0/
#299630000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#299640000000
0!
0'
0/
#299650000000
1!
1'
1/
#299660000000
0!
0'
0/
#299670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#299680000000
0!
0'
0/
#299690000000
1!
1'
1/
#299700000000
0!
0'
0/
#299710000000
#299720000000
1!
1'
1/
#299730000000
0!
0'
0/
#299740000000
1!
1'
1/
#299750000000
0!
1"
0'
1(
0/
10
#299760000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#299770000000
0!
0'
0/
#299780000000
1!
1'
1/
#299790000000
0!
0'
0/
#299800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#299810000000
0!
0'
0/
#299820000000
1!
1'
1/
#299830000000
0!
1"
0'
1(
0/
10
#299840000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#299850000000
0!
1$
0'
1+
0/
#299860000000
1!
1'
1/
#299870000000
0!
0'
0/
#299880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#299890000000
0!
0'
0/
#299900000000
1!
1'
1/
#299910000000
0!
0'
0/
#299920000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#299930000000
0!
0'
0/
#299940000000
1!
1'
1/
#299950000000
0!
0'
0/
#299960000000
1!
1'
1/
#299970000000
0!
0'
0/
#299980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#299990000000
0!
0'
0/
#300000000000
1!
1'
1/
#300010000000
0!
0'
0/
#300020000000
1!
1'
1/
#300030000000
0!
0'
0/
#300040000000
1!
1'
1/
#300050000000
0!
0'
0/
#300060000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#300070000000
0!
0'
0/
#300080000000
1!
1'
1/
#300090000000
0!
0'
0/
#300100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#300110000000
0!
0'
0/
#300120000000
1!
1'
1/
#300130000000
0!
0'
0/
#300140000000
#300150000000
1!
1'
1/
#300160000000
0!
0'
0/
#300170000000
1!
1'
1/
#300180000000
0!
1"
0'
1(
0/
10
#300190000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#300200000000
0!
0'
0/
#300210000000
1!
1'
1/
#300220000000
0!
0'
0/
#300230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#300240000000
0!
0'
0/
#300250000000
1!
1'
1/
#300260000000
0!
1"
0'
1(
0/
10
#300270000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#300280000000
0!
1$
0'
1+
0/
#300290000000
1!
1'
1/
#300300000000
0!
0'
0/
#300310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#300320000000
0!
0'
0/
#300330000000
1!
1'
1/
#300340000000
0!
0'
0/
#300350000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#300360000000
0!
0'
0/
#300370000000
1!
1'
1/
#300380000000
0!
0'
0/
#300390000000
1!
1'
1/
#300400000000
0!
0'
0/
#300410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#300420000000
0!
0'
0/
#300430000000
1!
1'
1/
#300440000000
0!
0'
0/
#300450000000
1!
1'
1/
#300460000000
0!
0'
0/
#300470000000
1!
1'
1/
#300480000000
0!
0'
0/
#300490000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#300500000000
0!
0'
0/
#300510000000
1!
1'
1/
#300520000000
0!
0'
0/
#300530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#300540000000
0!
0'
0/
#300550000000
1!
1'
1/
#300560000000
0!
0'
0/
#300570000000
#300580000000
1!
1'
1/
#300590000000
0!
0'
0/
#300600000000
1!
1'
1/
#300610000000
0!
1"
0'
1(
0/
10
#300620000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#300630000000
0!
0'
0/
#300640000000
1!
1'
1/
#300650000000
0!
0'
0/
#300660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#300670000000
0!
0'
0/
#300680000000
1!
1'
1/
#300690000000
0!
1"
0'
1(
0/
10
#300700000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#300710000000
0!
1$
0'
1+
0/
#300720000000
1!
1'
1/
#300730000000
0!
0'
0/
#300740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#300750000000
0!
0'
0/
#300760000000
1!
1'
1/
#300770000000
0!
0'
0/
#300780000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#300790000000
0!
0'
0/
#300800000000
1!
1'
1/
#300810000000
0!
0'
0/
#300820000000
1!
1'
1/
#300830000000
0!
0'
0/
#300840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#300850000000
0!
0'
0/
#300860000000
1!
1'
1/
#300870000000
0!
0'
0/
#300880000000
1!
1'
1/
#300890000000
0!
0'
0/
#300900000000
1!
1'
1/
#300910000000
0!
0'
0/
#300920000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#300930000000
0!
0'
0/
#300940000000
1!
1'
1/
#300950000000
0!
0'
0/
#300960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#300970000000
0!
0'
0/
#300980000000
1!
1'
1/
#300990000000
0!
0'
0/
#301000000000
#301010000000
1!
1'
1/
#301020000000
0!
0'
0/
#301030000000
1!
1'
1/
#301040000000
0!
1"
0'
1(
0/
10
#301050000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#301060000000
0!
0'
0/
#301070000000
1!
1'
1/
#301080000000
0!
0'
0/
#301090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#301100000000
0!
0'
0/
#301110000000
1!
1'
1/
#301120000000
0!
1"
0'
1(
0/
10
#301130000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#301140000000
0!
1$
0'
1+
0/
#301150000000
1!
1'
1/
#301160000000
0!
0'
0/
#301170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#301180000000
0!
0'
0/
#301190000000
1!
1'
1/
#301200000000
0!
0'
0/
#301210000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#301220000000
0!
0'
0/
#301230000000
1!
1'
1/
#301240000000
0!
0'
0/
#301250000000
1!
1'
1/
#301260000000
0!
0'
0/
#301270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#301280000000
0!
0'
0/
#301290000000
1!
1'
1/
#301300000000
0!
0'
0/
#301310000000
1!
1'
1/
#301320000000
0!
0'
0/
#301330000000
1!
1'
1/
#301340000000
0!
0'
0/
#301350000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#301360000000
0!
0'
0/
#301370000000
1!
1'
1/
#301380000000
0!
0'
0/
#301390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#301400000000
0!
0'
0/
#301410000000
1!
1'
1/
#301420000000
0!
0'
0/
#301430000000
#301440000000
1!
1'
1/
#301450000000
0!
0'
0/
#301460000000
1!
1'
1/
#301470000000
0!
1"
0'
1(
0/
10
#301480000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#301490000000
0!
0'
0/
#301500000000
1!
1'
1/
#301510000000
0!
0'
0/
#301520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#301530000000
0!
0'
0/
#301540000000
1!
1'
1/
#301550000000
0!
1"
0'
1(
0/
10
#301560000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#301570000000
0!
1$
0'
1+
0/
#301580000000
1!
1'
1/
#301590000000
0!
0'
0/
#301600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#301610000000
0!
0'
0/
#301620000000
1!
1'
1/
#301630000000
0!
0'
0/
#301640000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#301650000000
0!
0'
0/
#301660000000
1!
1'
1/
#301670000000
0!
0'
0/
#301680000000
1!
1'
1/
#301690000000
0!
0'
0/
#301700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#301710000000
0!
0'
0/
#301720000000
1!
1'
1/
#301730000000
0!
0'
0/
#301740000000
1!
1'
1/
#301750000000
0!
0'
0/
#301760000000
1!
1'
1/
#301770000000
0!
0'
0/
#301780000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#301790000000
0!
0'
0/
#301800000000
1!
1'
1/
#301810000000
0!
0'
0/
#301820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#301830000000
0!
0'
0/
#301840000000
1!
1'
1/
#301850000000
0!
0'
0/
#301860000000
#301870000000
1!
1'
1/
#301880000000
0!
0'
0/
#301890000000
1!
1'
1/
#301900000000
0!
1"
0'
1(
0/
10
#301910000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#301920000000
0!
0'
0/
#301930000000
1!
1'
1/
#301940000000
0!
0'
0/
#301950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#301960000000
0!
0'
0/
#301970000000
1!
1'
1/
#301980000000
0!
1"
0'
1(
0/
10
#301990000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#302000000000
0!
1$
0'
1+
0/
#302010000000
1!
1'
1/
#302020000000
0!
0'
0/
#302030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#302040000000
0!
0'
0/
#302050000000
1!
1'
1/
#302060000000
0!
0'
0/
#302070000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#302080000000
0!
0'
0/
#302090000000
1!
1'
1/
#302100000000
0!
0'
0/
#302110000000
1!
1'
1/
#302120000000
0!
0'
0/
#302130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#302140000000
0!
0'
0/
#302150000000
1!
1'
1/
#302160000000
0!
0'
0/
#302170000000
1!
1'
1/
#302180000000
0!
0'
0/
#302190000000
1!
1'
1/
#302200000000
0!
0'
0/
#302210000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#302220000000
0!
0'
0/
#302230000000
1!
1'
1/
#302240000000
0!
0'
0/
#302250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#302260000000
0!
0'
0/
#302270000000
1!
1'
1/
#302280000000
0!
0'
0/
#302290000000
#302300000000
1!
1'
1/
#302310000000
0!
0'
0/
#302320000000
1!
1'
1/
#302330000000
0!
1"
0'
1(
0/
10
#302340000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#302350000000
0!
0'
0/
#302360000000
1!
1'
1/
#302370000000
0!
0'
0/
#302380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#302390000000
0!
0'
0/
#302400000000
1!
1'
1/
#302410000000
0!
1"
0'
1(
0/
10
#302420000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#302430000000
0!
1$
0'
1+
0/
#302440000000
1!
1'
1/
#302450000000
0!
0'
0/
#302460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#302470000000
0!
0'
0/
#302480000000
1!
1'
1/
#302490000000
0!
0'
0/
#302500000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#302510000000
0!
0'
0/
#302520000000
1!
1'
1/
#302530000000
0!
0'
0/
#302540000000
1!
1'
1/
#302550000000
0!
0'
0/
#302560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#302570000000
0!
0'
0/
#302580000000
1!
1'
1/
#302590000000
0!
0'
0/
#302600000000
1!
1'
1/
#302610000000
0!
0'
0/
#302620000000
1!
1'
1/
#302630000000
0!
0'
0/
#302640000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#302650000000
0!
0'
0/
#302660000000
1!
1'
1/
#302670000000
0!
0'
0/
#302680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#302690000000
0!
0'
0/
#302700000000
1!
1'
1/
#302710000000
0!
0'
0/
#302720000000
#302730000000
1!
1'
1/
#302740000000
0!
0'
0/
#302750000000
1!
1'
1/
#302760000000
0!
1"
0'
1(
0/
10
#302770000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#302780000000
0!
0'
0/
#302790000000
1!
1'
1/
#302800000000
0!
0'
0/
#302810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#302820000000
0!
0'
0/
#302830000000
1!
1'
1/
#302840000000
0!
1"
0'
1(
0/
10
#302850000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#302860000000
0!
1$
0'
1+
0/
#302870000000
1!
1'
1/
#302880000000
0!
0'
0/
#302890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#302900000000
0!
0'
0/
#302910000000
1!
1'
1/
#302920000000
0!
0'
0/
#302930000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#302940000000
0!
0'
0/
#302950000000
1!
1'
1/
#302960000000
0!
0'
0/
#302970000000
1!
1'
1/
#302980000000
0!
0'
0/
#302990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#303000000000
0!
0'
0/
#303010000000
1!
1'
1/
#303020000000
0!
0'
0/
#303030000000
1!
1'
1/
#303040000000
0!
0'
0/
#303050000000
1!
1'
1/
#303060000000
0!
0'
0/
#303070000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#303080000000
0!
0'
0/
#303090000000
1!
1'
1/
#303100000000
0!
0'
0/
#303110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#303120000000
0!
0'
0/
#303130000000
1!
1'
1/
#303140000000
0!
0'
0/
#303150000000
#303160000000
1!
1'
1/
#303170000000
0!
0'
0/
#303180000000
1!
1'
1/
#303190000000
0!
1"
0'
1(
0/
10
#303200000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#303210000000
0!
0'
0/
#303220000000
1!
1'
1/
#303230000000
0!
0'
0/
#303240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#303250000000
0!
0'
0/
#303260000000
1!
1'
1/
#303270000000
0!
1"
0'
1(
0/
10
#303280000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#303290000000
0!
1$
0'
1+
0/
#303300000000
1!
1'
1/
#303310000000
0!
0'
0/
#303320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#303330000000
0!
0'
0/
#303340000000
1!
1'
1/
#303350000000
0!
0'
0/
#303360000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#303370000000
0!
0'
0/
#303380000000
1!
1'
1/
#303390000000
0!
0'
0/
#303400000000
1!
1'
1/
#303410000000
0!
0'
0/
#303420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#303430000000
0!
0'
0/
#303440000000
1!
1'
1/
#303450000000
0!
0'
0/
#303460000000
1!
1'
1/
#303470000000
0!
0'
0/
#303480000000
1!
1'
1/
#303490000000
0!
0'
0/
#303500000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#303510000000
0!
0'
0/
#303520000000
1!
1'
1/
#303530000000
0!
0'
0/
#303540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#303550000000
0!
0'
0/
#303560000000
1!
1'
1/
#303570000000
0!
0'
0/
#303580000000
#303590000000
1!
1'
1/
#303600000000
0!
0'
0/
#303610000000
1!
1'
1/
#303620000000
0!
1"
0'
1(
0/
10
#303630000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#303640000000
0!
0'
0/
#303650000000
1!
1'
1/
#303660000000
0!
0'
0/
#303670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#303680000000
0!
0'
0/
#303690000000
1!
1'
1/
#303700000000
0!
1"
0'
1(
0/
10
#303710000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#303720000000
0!
1$
0'
1+
0/
#303730000000
1!
1'
1/
#303740000000
0!
0'
0/
#303750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#303760000000
0!
0'
0/
#303770000000
1!
1'
1/
#303780000000
0!
0'
0/
#303790000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#303800000000
0!
0'
0/
#303810000000
1!
1'
1/
#303820000000
0!
0'
0/
#303830000000
1!
1'
1/
#303840000000
0!
0'
0/
#303850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#303860000000
0!
0'
0/
#303870000000
1!
1'
1/
#303880000000
0!
0'
0/
#303890000000
1!
1'
1/
#303900000000
0!
0'
0/
#303910000000
1!
1'
1/
#303920000000
0!
0'
0/
#303930000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#303940000000
0!
0'
0/
#303950000000
1!
1'
1/
#303960000000
0!
0'
0/
#303970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#303980000000
0!
0'
0/
#303990000000
1!
1'
1/
#304000000000
0!
0'
0/
#304010000000
#304020000000
1!
1'
1/
#304030000000
0!
0'
0/
#304040000000
1!
1'
1/
#304050000000
0!
1"
0'
1(
0/
10
#304060000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#304070000000
0!
0'
0/
#304080000000
1!
1'
1/
#304090000000
0!
0'
0/
#304100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#304110000000
0!
0'
0/
#304120000000
1!
1'
1/
#304130000000
0!
1"
0'
1(
0/
10
#304140000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#304150000000
0!
1$
0'
1+
0/
#304160000000
1!
1'
1/
#304170000000
0!
0'
0/
#304180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#304190000000
0!
0'
0/
#304200000000
1!
1'
1/
#304210000000
0!
0'
0/
#304220000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#304230000000
0!
0'
0/
#304240000000
1!
1'
1/
#304250000000
0!
0'
0/
#304260000000
1!
1'
1/
#304270000000
0!
0'
0/
#304280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#304290000000
0!
0'
0/
#304300000000
1!
1'
1/
#304310000000
0!
0'
0/
#304320000000
1!
1'
1/
#304330000000
0!
0'
0/
#304340000000
1!
1'
1/
#304350000000
0!
0'
0/
#304360000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#304370000000
0!
0'
0/
#304380000000
1!
1'
1/
#304390000000
0!
0'
0/
#304400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#304410000000
0!
0'
0/
#304420000000
1!
1'
1/
#304430000000
0!
0'
0/
#304440000000
#304450000000
1!
1'
1/
#304460000000
0!
0'
0/
#304470000000
1!
1'
1/
#304480000000
0!
1"
0'
1(
0/
10
#304490000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#304500000000
0!
0'
0/
#304510000000
1!
1'
1/
#304520000000
0!
0'
0/
#304530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#304540000000
0!
0'
0/
#304550000000
1!
1'
1/
#304560000000
0!
1"
0'
1(
0/
10
#304570000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#304580000000
0!
1$
0'
1+
0/
#304590000000
1!
1'
1/
#304600000000
0!
0'
0/
#304610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#304620000000
0!
0'
0/
#304630000000
1!
1'
1/
#304640000000
0!
0'
0/
#304650000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#304660000000
0!
0'
0/
#304670000000
1!
1'
1/
#304680000000
0!
0'
0/
#304690000000
1!
1'
1/
#304700000000
0!
0'
0/
#304710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#304720000000
0!
0'
0/
#304730000000
1!
1'
1/
#304740000000
0!
0'
0/
#304750000000
1!
1'
1/
#304760000000
0!
0'
0/
#304770000000
1!
1'
1/
#304780000000
0!
0'
0/
#304790000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#304800000000
0!
0'
0/
#304810000000
1!
1'
1/
#304820000000
0!
0'
0/
#304830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#304840000000
0!
0'
0/
#304850000000
1!
1'
1/
#304860000000
0!
0'
0/
#304870000000
#304880000000
1!
1'
1/
#304890000000
0!
0'
0/
#304900000000
1!
1'
1/
#304910000000
0!
1"
0'
1(
0/
10
#304920000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#304930000000
0!
0'
0/
#304940000000
1!
1'
1/
#304950000000
0!
0'
0/
#304960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#304970000000
0!
0'
0/
#304980000000
1!
1'
1/
#304990000000
0!
1"
0'
1(
0/
10
#305000000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#305010000000
0!
1$
0'
1+
0/
#305020000000
1!
1'
1/
#305030000000
0!
0'
0/
#305040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#305050000000
0!
0'
0/
#305060000000
1!
1'
1/
#305070000000
0!
0'
0/
#305080000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#305090000000
0!
0'
0/
#305100000000
1!
1'
1/
#305110000000
0!
0'
0/
#305120000000
1!
1'
1/
#305130000000
0!
0'
0/
#305140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#305150000000
0!
0'
0/
#305160000000
1!
1'
1/
#305170000000
0!
0'
0/
#305180000000
1!
1'
1/
#305190000000
0!
0'
0/
#305200000000
1!
1'
1/
#305210000000
0!
0'
0/
#305220000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#305230000000
0!
0'
0/
#305240000000
1!
1'
1/
#305250000000
0!
0'
0/
#305260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#305270000000
0!
0'
0/
#305280000000
1!
1'
1/
#305290000000
0!
0'
0/
#305300000000
#305310000000
1!
1'
1/
#305320000000
0!
0'
0/
#305330000000
1!
1'
1/
#305340000000
0!
1"
0'
1(
0/
10
#305350000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#305360000000
0!
0'
0/
#305370000000
1!
1'
1/
#305380000000
0!
0'
0/
#305390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#305400000000
0!
0'
0/
#305410000000
1!
1'
1/
#305420000000
0!
1"
0'
1(
0/
10
#305430000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#305440000000
0!
1$
0'
1+
0/
#305450000000
1!
1'
1/
#305460000000
0!
0'
0/
#305470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#305480000000
0!
0'
0/
#305490000000
1!
1'
1/
#305500000000
0!
0'
0/
#305510000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#305520000000
0!
0'
0/
#305530000000
1!
1'
1/
#305540000000
0!
0'
0/
#305550000000
1!
1'
1/
#305560000000
0!
0'
0/
#305570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#305580000000
0!
0'
0/
#305590000000
1!
1'
1/
#305600000000
0!
0'
0/
#305610000000
1!
1'
1/
#305620000000
0!
0'
0/
#305630000000
1!
1'
1/
#305640000000
0!
0'
0/
#305650000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#305660000000
0!
0'
0/
#305670000000
1!
1'
1/
#305680000000
0!
0'
0/
#305690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#305700000000
0!
0'
0/
#305710000000
1!
1'
1/
#305720000000
0!
0'
0/
#305730000000
#305740000000
1!
1'
1/
#305750000000
0!
0'
0/
#305760000000
1!
1'
1/
#305770000000
0!
1"
0'
1(
0/
10
#305780000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#305790000000
0!
0'
0/
#305800000000
1!
1'
1/
#305810000000
0!
0'
0/
#305820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#305830000000
0!
0'
0/
#305840000000
1!
1'
1/
#305850000000
0!
1"
0'
1(
0/
10
#305860000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#305870000000
0!
1$
0'
1+
0/
#305880000000
1!
1'
1/
#305890000000
0!
0'
0/
#305900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#305910000000
0!
0'
0/
#305920000000
1!
1'
1/
#305930000000
0!
0'
0/
#305940000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#305950000000
0!
0'
0/
#305960000000
1!
1'
1/
#305970000000
0!
0'
0/
#305980000000
1!
1'
1/
#305990000000
0!
0'
0/
#306000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#306010000000
0!
0'
0/
#306020000000
1!
1'
1/
#306030000000
0!
0'
0/
#306040000000
1!
1'
1/
#306050000000
0!
0'
0/
#306060000000
1!
1'
1/
#306070000000
0!
0'
0/
#306080000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#306090000000
0!
0'
0/
#306100000000
1!
1'
1/
#306110000000
0!
0'
0/
#306120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#306130000000
0!
0'
0/
#306140000000
1!
1'
1/
#306150000000
0!
0'
0/
#306160000000
#306170000000
1!
1'
1/
#306180000000
0!
0'
0/
#306190000000
1!
1'
1/
#306200000000
0!
1"
0'
1(
0/
10
#306210000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#306220000000
0!
0'
0/
#306230000000
1!
1'
1/
#306240000000
0!
0'
0/
#306250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#306260000000
0!
0'
0/
#306270000000
1!
1'
1/
#306280000000
0!
1"
0'
1(
0/
10
#306290000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#306300000000
0!
1$
0'
1+
0/
#306310000000
1!
1'
1/
#306320000000
0!
0'
0/
#306330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#306340000000
0!
0'
0/
#306350000000
1!
1'
1/
#306360000000
0!
0'
0/
#306370000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#306380000000
0!
0'
0/
#306390000000
1!
1'
1/
#306400000000
0!
0'
0/
#306410000000
1!
1'
1/
#306420000000
0!
0'
0/
#306430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#306440000000
0!
0'
0/
#306450000000
1!
1'
1/
#306460000000
0!
0'
0/
#306470000000
1!
1'
1/
#306480000000
0!
0'
0/
#306490000000
1!
1'
1/
#306500000000
0!
0'
0/
#306510000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#306520000000
0!
0'
0/
#306530000000
1!
1'
1/
#306540000000
0!
0'
0/
#306550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#306560000000
0!
0'
0/
#306570000000
1!
1'
1/
#306580000000
0!
0'
0/
#306590000000
#306600000000
1!
1'
1/
#306610000000
0!
0'
0/
#306620000000
1!
1'
1/
#306630000000
0!
1"
0'
1(
0/
10
#306640000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#306650000000
0!
0'
0/
#306660000000
1!
1'
1/
#306670000000
0!
0'
0/
#306680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#306690000000
0!
0'
0/
#306700000000
1!
1'
1/
#306710000000
0!
1"
0'
1(
0/
10
#306720000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#306730000000
0!
1$
0'
1+
0/
#306740000000
1!
1'
1/
#306750000000
0!
0'
0/
#306760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#306770000000
0!
0'
0/
#306780000000
1!
1'
1/
#306790000000
0!
0'
0/
#306800000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#306810000000
0!
0'
0/
#306820000000
1!
1'
1/
#306830000000
0!
0'
0/
#306840000000
1!
1'
1/
#306850000000
0!
0'
0/
#306860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#306870000000
0!
0'
0/
#306880000000
1!
1'
1/
#306890000000
0!
0'
0/
#306900000000
1!
1'
1/
#306910000000
0!
0'
0/
#306920000000
1!
1'
1/
#306930000000
0!
0'
0/
#306940000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#306950000000
0!
0'
0/
#306960000000
1!
1'
1/
#306970000000
0!
0'
0/
#306980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#306990000000
0!
0'
0/
#307000000000
1!
1'
1/
#307010000000
0!
0'
0/
#307020000000
#307030000000
1!
1'
1/
#307040000000
0!
0'
0/
#307050000000
1!
1'
1/
#307060000000
0!
1"
0'
1(
0/
10
#307070000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#307080000000
0!
0'
0/
#307090000000
1!
1'
1/
#307100000000
0!
0'
0/
#307110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#307120000000
0!
0'
0/
#307130000000
1!
1'
1/
#307140000000
0!
1"
0'
1(
0/
10
#307150000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#307160000000
0!
1$
0'
1+
0/
#307170000000
1!
1'
1/
#307180000000
0!
0'
0/
#307190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#307200000000
0!
0'
0/
#307210000000
1!
1'
1/
#307220000000
0!
0'
0/
#307230000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#307240000000
0!
0'
0/
#307250000000
1!
1'
1/
#307260000000
0!
0'
0/
#307270000000
1!
1'
1/
#307280000000
0!
0'
0/
#307290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#307300000000
0!
0'
0/
#307310000000
1!
1'
1/
#307320000000
0!
0'
0/
#307330000000
1!
1'
1/
#307340000000
0!
0'
0/
#307350000000
1!
1'
1/
#307360000000
0!
0'
0/
#307370000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#307380000000
0!
0'
0/
#307390000000
1!
1'
1/
#307400000000
0!
0'
0/
#307410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#307420000000
0!
0'
0/
#307430000000
1!
1'
1/
#307440000000
0!
0'
0/
#307450000000
#307460000000
1!
1'
1/
#307470000000
0!
0'
0/
#307480000000
1!
1'
1/
#307490000000
0!
1"
0'
1(
0/
10
#307500000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#307510000000
0!
0'
0/
#307520000000
1!
1'
1/
#307530000000
0!
0'
0/
#307540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#307550000000
0!
0'
0/
#307560000000
1!
1'
1/
#307570000000
0!
1"
0'
1(
0/
10
#307580000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#307590000000
0!
1$
0'
1+
0/
#307600000000
1!
1'
1/
#307610000000
0!
0'
0/
#307620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#307630000000
0!
0'
0/
#307640000000
1!
1'
1/
#307650000000
0!
0'
0/
#307660000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#307670000000
0!
0'
0/
#307680000000
1!
1'
1/
#307690000000
0!
0'
0/
#307700000000
1!
1'
1/
#307710000000
0!
0'
0/
#307720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#307730000000
0!
0'
0/
#307740000000
1!
1'
1/
#307750000000
0!
0'
0/
#307760000000
1!
1'
1/
#307770000000
0!
0'
0/
#307780000000
1!
1'
1/
#307790000000
0!
0'
0/
#307800000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#307810000000
0!
0'
0/
#307820000000
1!
1'
1/
#307830000000
0!
0'
0/
#307840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#307850000000
0!
0'
0/
#307860000000
1!
1'
1/
#307870000000
0!
0'
0/
#307880000000
#307890000000
1!
1'
1/
#307900000000
0!
0'
0/
#307910000000
1!
1'
1/
#307920000000
0!
1"
0'
1(
0/
10
#307930000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#307940000000
0!
0'
0/
#307950000000
1!
1'
1/
#307960000000
0!
0'
0/
#307970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#307980000000
0!
0'
0/
#307990000000
1!
1'
1/
#308000000000
0!
1"
0'
1(
0/
10
#308010000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#308020000000
0!
1$
0'
1+
0/
#308030000000
1!
1'
1/
#308040000000
0!
0'
0/
#308050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#308060000000
0!
0'
0/
#308070000000
1!
1'
1/
#308080000000
0!
0'
0/
#308090000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#308100000000
0!
0'
0/
#308110000000
1!
1'
1/
#308120000000
0!
0'
0/
#308130000000
1!
1'
1/
#308140000000
0!
0'
0/
#308150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#308160000000
0!
0'
0/
#308170000000
1!
1'
1/
#308180000000
0!
0'
0/
#308190000000
1!
1'
1/
#308200000000
0!
0'
0/
#308210000000
1!
1'
1/
#308220000000
0!
0'
0/
#308230000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#308240000000
0!
0'
0/
#308250000000
1!
1'
1/
#308260000000
0!
0'
0/
#308270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#308280000000
0!
0'
0/
#308290000000
1!
1'
1/
#308300000000
0!
0'
0/
#308310000000
#308320000000
1!
1'
1/
#308330000000
0!
0'
0/
#308340000000
1!
1'
1/
#308350000000
0!
1"
0'
1(
0/
10
#308360000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#308370000000
0!
0'
0/
#308380000000
1!
1'
1/
#308390000000
0!
0'
0/
#308400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#308410000000
0!
0'
0/
#308420000000
1!
1'
1/
#308430000000
0!
1"
0'
1(
0/
10
#308440000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#308450000000
0!
1$
0'
1+
0/
#308460000000
1!
1'
1/
#308470000000
0!
0'
0/
#308480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#308490000000
0!
0'
0/
#308500000000
1!
1'
1/
#308510000000
0!
0'
0/
#308520000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#308530000000
0!
0'
0/
#308540000000
1!
1'
1/
#308550000000
0!
0'
0/
#308560000000
1!
1'
1/
#308570000000
0!
0'
0/
#308580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#308590000000
0!
0'
0/
#308600000000
1!
1'
1/
#308610000000
0!
0'
0/
#308620000000
1!
1'
1/
#308630000000
0!
0'
0/
#308640000000
1!
1'
1/
#308650000000
0!
0'
0/
#308660000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#308670000000
0!
0'
0/
#308680000000
1!
1'
1/
#308690000000
0!
0'
0/
#308700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#308710000000
0!
0'
0/
#308720000000
1!
1'
1/
#308730000000
0!
0'
0/
#308740000000
#308750000000
1!
1'
1/
#308760000000
0!
0'
0/
#308770000000
1!
1'
1/
#308780000000
0!
1"
0'
1(
0/
10
#308790000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#308800000000
0!
0'
0/
#308810000000
1!
1'
1/
#308820000000
0!
0'
0/
#308830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#308840000000
0!
0'
0/
#308850000000
1!
1'
1/
#308860000000
0!
1"
0'
1(
0/
10
#308870000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#308880000000
0!
1$
0'
1+
0/
#308890000000
1!
1'
1/
#308900000000
0!
0'
0/
#308910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#308920000000
0!
0'
0/
#308930000000
1!
1'
1/
#308940000000
0!
0'
0/
#308950000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#308960000000
0!
0'
0/
#308970000000
1!
1'
1/
#308980000000
0!
0'
0/
#308990000000
1!
1'
1/
#309000000000
0!
0'
0/
#309010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#309020000000
0!
0'
0/
#309030000000
1!
1'
1/
#309040000000
0!
0'
0/
#309050000000
1!
1'
1/
#309060000000
0!
0'
0/
#309070000000
1!
1'
1/
#309080000000
0!
0'
0/
#309090000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#309100000000
0!
0'
0/
#309110000000
1!
1'
1/
#309120000000
0!
0'
0/
#309130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#309140000000
0!
0'
0/
#309150000000
1!
1'
1/
#309160000000
0!
0'
0/
#309170000000
#309180000000
1!
1'
1/
#309190000000
0!
0'
0/
#309200000000
1!
1'
1/
#309210000000
0!
1"
0'
1(
0/
10
#309220000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#309230000000
0!
0'
0/
#309240000000
1!
1'
1/
#309250000000
0!
0'
0/
#309260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#309270000000
0!
0'
0/
#309280000000
1!
1'
1/
#309290000000
0!
1"
0'
1(
0/
10
#309300000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#309310000000
0!
1$
0'
1+
0/
#309320000000
1!
1'
1/
#309330000000
0!
0'
0/
#309340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#309350000000
0!
0'
0/
#309360000000
1!
1'
1/
#309370000000
0!
0'
0/
#309380000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#309390000000
0!
0'
0/
#309400000000
1!
1'
1/
#309410000000
0!
0'
0/
#309420000000
1!
1'
1/
#309430000000
0!
0'
0/
#309440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#309450000000
0!
0'
0/
#309460000000
1!
1'
1/
#309470000000
0!
0'
0/
#309480000000
1!
1'
1/
#309490000000
0!
0'
0/
#309500000000
1!
1'
1/
#309510000000
0!
0'
0/
#309520000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#309530000000
0!
0'
0/
#309540000000
1!
1'
1/
#309550000000
0!
0'
0/
#309560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#309570000000
0!
0'
0/
#309580000000
1!
1'
1/
#309590000000
0!
0'
0/
#309600000000
#309610000000
1!
1'
1/
#309620000000
0!
0'
0/
#309630000000
1!
1'
1/
#309640000000
0!
1"
0'
1(
0/
10
#309650000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#309660000000
0!
0'
0/
#309670000000
1!
1'
1/
#309680000000
0!
0'
0/
#309690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#309700000000
0!
0'
0/
#309710000000
1!
1'
1/
#309720000000
0!
1"
0'
1(
0/
10
#309730000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#309740000000
0!
1$
0'
1+
0/
#309750000000
1!
1'
1/
#309760000000
0!
0'
0/
#309770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#309780000000
0!
0'
0/
#309790000000
1!
1'
1/
#309800000000
0!
0'
0/
#309810000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#309820000000
0!
0'
0/
#309830000000
1!
1'
1/
#309840000000
0!
0'
0/
#309850000000
1!
1'
1/
#309860000000
0!
0'
0/
#309870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#309880000000
0!
0'
0/
#309890000000
1!
1'
1/
#309900000000
0!
0'
0/
#309910000000
1!
1'
1/
#309920000000
0!
0'
0/
#309930000000
1!
1'
1/
#309940000000
0!
0'
0/
#309950000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#309960000000
0!
0'
0/
#309970000000
1!
1'
1/
#309980000000
0!
0'
0/
#309990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#310000000000
0!
0'
0/
#310010000000
1!
1'
1/
#310020000000
0!
0'
0/
#310030000000
#310040000000
1!
1'
1/
#310050000000
0!
0'
0/
#310060000000
1!
1'
1/
#310070000000
0!
1"
0'
1(
0/
10
#310080000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#310090000000
0!
0'
0/
#310100000000
1!
1'
1/
#310110000000
0!
0'
0/
#310120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#310130000000
0!
0'
0/
#310140000000
1!
1'
1/
#310150000000
0!
1"
0'
1(
0/
10
#310160000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#310170000000
0!
1$
0'
1+
0/
#310180000000
1!
1'
1/
#310190000000
0!
0'
0/
#310200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#310210000000
0!
0'
0/
#310220000000
1!
1'
1/
#310230000000
0!
0'
0/
#310240000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#310250000000
0!
0'
0/
#310260000000
1!
1'
1/
#310270000000
0!
0'
0/
#310280000000
1!
1'
1/
#310290000000
0!
0'
0/
#310300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#310310000000
0!
0'
0/
#310320000000
1!
1'
1/
#310330000000
0!
0'
0/
#310340000000
1!
1'
1/
#310350000000
0!
0'
0/
#310360000000
1!
1'
1/
#310370000000
0!
0'
0/
#310380000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#310390000000
0!
0'
0/
#310400000000
1!
1'
1/
#310410000000
0!
0'
0/
#310420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#310430000000
0!
0'
0/
#310440000000
1!
1'
1/
#310450000000
0!
0'
0/
#310460000000
#310470000000
1!
1'
1/
#310480000000
0!
0'
0/
#310490000000
1!
1'
1/
#310500000000
0!
1"
0'
1(
0/
10
#310510000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#310520000000
0!
0'
0/
#310530000000
1!
1'
1/
#310540000000
0!
0'
0/
#310550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#310560000000
0!
0'
0/
#310570000000
1!
1'
1/
#310580000000
0!
1"
0'
1(
0/
10
#310590000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#310600000000
0!
1$
0'
1+
0/
#310610000000
1!
1'
1/
#310620000000
0!
0'
0/
#310630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#310640000000
0!
0'
0/
#310650000000
1!
1'
1/
#310660000000
0!
0'
0/
#310670000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#310680000000
0!
0'
0/
#310690000000
1!
1'
1/
#310700000000
0!
0'
0/
#310710000000
1!
1'
1/
#310720000000
0!
0'
0/
#310730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#310740000000
0!
0'
0/
#310750000000
1!
1'
1/
#310760000000
0!
0'
0/
#310770000000
1!
1'
1/
#310780000000
0!
0'
0/
#310790000000
1!
1'
1/
#310800000000
0!
0'
0/
#310810000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#310820000000
0!
0'
0/
#310830000000
1!
1'
1/
#310840000000
0!
0'
0/
#310850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#310860000000
0!
0'
0/
#310870000000
1!
1'
1/
#310880000000
0!
0'
0/
#310890000000
#310900000000
1!
1'
1/
#310910000000
0!
0'
0/
#310920000000
1!
1'
1/
#310930000000
0!
1"
0'
1(
0/
10
#310940000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#310950000000
0!
0'
0/
#310960000000
1!
1'
1/
#310970000000
0!
0'
0/
#310980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#310990000000
0!
0'
0/
#311000000000
1!
1'
1/
#311010000000
0!
1"
0'
1(
0/
10
#311020000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#311030000000
0!
1$
0'
1+
0/
#311040000000
1!
1'
1/
#311050000000
0!
0'
0/
#311060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#311070000000
0!
0'
0/
#311080000000
1!
1'
1/
#311090000000
0!
0'
0/
#311100000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#311110000000
0!
0'
0/
#311120000000
1!
1'
1/
#311130000000
0!
0'
0/
#311140000000
1!
1'
1/
#311150000000
0!
0'
0/
#311160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#311170000000
0!
0'
0/
#311180000000
1!
1'
1/
#311190000000
0!
0'
0/
#311200000000
1!
1'
1/
#311210000000
0!
0'
0/
#311220000000
1!
1'
1/
#311230000000
0!
0'
0/
#311240000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#311250000000
0!
0'
0/
#311260000000
1!
1'
1/
#311270000000
0!
0'
0/
#311280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#311290000000
0!
0'
0/
#311300000000
1!
1'
1/
#311310000000
0!
0'
0/
#311320000000
#311330000000
1!
1'
1/
#311340000000
0!
0'
0/
#311350000000
1!
1'
1/
#311360000000
0!
1"
0'
1(
0/
10
#311370000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#311380000000
0!
0'
0/
#311390000000
1!
1'
1/
#311400000000
0!
0'
0/
#311410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#311420000000
0!
0'
0/
#311430000000
1!
1'
1/
#311440000000
0!
1"
0'
1(
0/
10
#311450000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#311460000000
0!
1$
0'
1+
0/
#311470000000
1!
1'
1/
#311480000000
0!
0'
0/
#311490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#311500000000
0!
0'
0/
#311510000000
1!
1'
1/
#311520000000
0!
0'
0/
#311530000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#311540000000
0!
0'
0/
#311550000000
1!
1'
1/
#311560000000
0!
0'
0/
#311570000000
1!
1'
1/
#311580000000
0!
0'
0/
#311590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#311600000000
0!
0'
0/
#311610000000
1!
1'
1/
#311620000000
0!
0'
0/
#311630000000
1!
1'
1/
#311640000000
0!
0'
0/
#311650000000
1!
1'
1/
#311660000000
0!
0'
0/
#311670000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#311680000000
0!
0'
0/
#311690000000
1!
1'
1/
#311700000000
0!
0'
0/
#311710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#311720000000
0!
0'
0/
#311730000000
1!
1'
1/
#311740000000
0!
0'
0/
#311750000000
#311760000000
1!
1'
1/
#311770000000
0!
0'
0/
#311780000000
1!
1'
1/
#311790000000
0!
1"
0'
1(
0/
10
#311800000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#311810000000
0!
0'
0/
#311820000000
1!
1'
1/
#311830000000
0!
0'
0/
#311840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#311850000000
0!
0'
0/
#311860000000
1!
1'
1/
#311870000000
0!
1"
0'
1(
0/
10
#311880000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#311890000000
0!
1$
0'
1+
0/
#311900000000
1!
1'
1/
#311910000000
0!
0'
0/
#311920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#311930000000
0!
0'
0/
#311940000000
1!
1'
1/
#311950000000
0!
0'
0/
#311960000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#311970000000
0!
0'
0/
#311980000000
1!
1'
1/
#311990000000
0!
0'
0/
#312000000000
1!
1'
1/
#312010000000
0!
0'
0/
#312020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#312030000000
0!
0'
0/
#312040000000
1!
1'
1/
#312050000000
0!
0'
0/
#312060000000
1!
1'
1/
#312070000000
0!
0'
0/
#312080000000
1!
1'
1/
#312090000000
0!
0'
0/
#312100000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#312110000000
0!
0'
0/
#312120000000
1!
1'
1/
#312130000000
0!
0'
0/
#312140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#312150000000
0!
0'
0/
#312160000000
1!
1'
1/
#312170000000
0!
0'
0/
#312180000000
#312190000000
1!
1'
1/
#312200000000
0!
0'
0/
#312210000000
1!
1'
1/
#312220000000
0!
1"
0'
1(
0/
10
#312230000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#312240000000
0!
0'
0/
#312250000000
1!
1'
1/
#312260000000
0!
0'
0/
#312270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#312280000000
0!
0'
0/
#312290000000
1!
1'
1/
#312300000000
0!
1"
0'
1(
0/
10
#312310000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#312320000000
0!
1$
0'
1+
0/
#312330000000
1!
1'
1/
#312340000000
0!
0'
0/
#312350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#312360000000
0!
0'
0/
#312370000000
1!
1'
1/
#312380000000
0!
0'
0/
#312390000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#312400000000
0!
0'
0/
#312410000000
1!
1'
1/
#312420000000
0!
0'
0/
#312430000000
1!
1'
1/
#312440000000
0!
0'
0/
#312450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#312460000000
0!
0'
0/
#312470000000
1!
1'
1/
#312480000000
0!
0'
0/
#312490000000
1!
1'
1/
#312500000000
0!
0'
0/
#312510000000
1!
1'
1/
#312520000000
0!
0'
0/
#312530000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#312540000000
0!
0'
0/
#312550000000
1!
1'
1/
#312560000000
0!
0'
0/
#312570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#312580000000
0!
0'
0/
#312590000000
1!
1'
1/
#312600000000
0!
0'
0/
#312610000000
#312620000000
1!
1'
1/
#312630000000
0!
0'
0/
#312640000000
1!
1'
1/
#312650000000
0!
1"
0'
1(
0/
10
#312660000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#312670000000
0!
0'
0/
#312680000000
1!
1'
1/
#312690000000
0!
0'
0/
#312700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#312710000000
0!
0'
0/
#312720000000
1!
1'
1/
#312730000000
0!
1"
0'
1(
0/
10
#312740000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#312750000000
0!
1$
0'
1+
0/
#312760000000
1!
1'
1/
#312770000000
0!
0'
0/
#312780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#312790000000
0!
0'
0/
#312800000000
1!
1'
1/
#312810000000
0!
0'
0/
#312820000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#312830000000
0!
0'
0/
#312840000000
1!
1'
1/
#312850000000
0!
0'
0/
#312860000000
1!
1'
1/
#312870000000
0!
0'
0/
#312880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#312890000000
0!
0'
0/
#312900000000
1!
1'
1/
#312910000000
0!
0'
0/
#312920000000
1!
1'
1/
#312930000000
0!
0'
0/
#312940000000
1!
1'
1/
#312950000000
0!
0'
0/
#312960000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#312970000000
0!
0'
0/
#312980000000
1!
1'
1/
#312990000000
0!
0'
0/
#313000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#313010000000
0!
0'
0/
#313020000000
1!
1'
1/
#313030000000
0!
0'
0/
#313040000000
#313050000000
1!
1'
1/
#313060000000
0!
0'
0/
#313070000000
1!
1'
1/
#313080000000
0!
1"
0'
1(
0/
10
#313090000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#313100000000
0!
0'
0/
#313110000000
1!
1'
1/
#313120000000
0!
0'
0/
#313130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#313140000000
0!
0'
0/
#313150000000
1!
1'
1/
#313160000000
0!
1"
0'
1(
0/
10
#313170000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#313180000000
0!
1$
0'
1+
0/
#313190000000
1!
1'
1/
#313200000000
0!
0'
0/
#313210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#313220000000
0!
0'
0/
#313230000000
1!
1'
1/
#313240000000
0!
0'
0/
#313250000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#313260000000
0!
0'
0/
#313270000000
1!
1'
1/
#313280000000
0!
0'
0/
#313290000000
1!
1'
1/
#313300000000
0!
0'
0/
#313310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#313320000000
0!
0'
0/
#313330000000
1!
1'
1/
#313340000000
0!
0'
0/
#313350000000
1!
1'
1/
#313360000000
0!
0'
0/
#313370000000
1!
1'
1/
#313380000000
0!
0'
0/
#313390000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#313400000000
0!
0'
0/
#313410000000
1!
1'
1/
#313420000000
0!
0'
0/
#313430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#313440000000
0!
0'
0/
#313450000000
1!
1'
1/
#313460000000
0!
0'
0/
#313470000000
#313480000000
1!
1'
1/
#313490000000
0!
0'
0/
#313500000000
1!
1'
1/
#313510000000
0!
1"
0'
1(
0/
10
#313520000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#313530000000
0!
0'
0/
#313540000000
1!
1'
1/
#313550000000
0!
0'
0/
#313560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#313570000000
0!
0'
0/
#313580000000
1!
1'
1/
#313590000000
0!
1"
0'
1(
0/
10
#313600000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#313610000000
0!
1$
0'
1+
0/
#313620000000
1!
1'
1/
#313630000000
0!
0'
0/
#313640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#313650000000
0!
0'
0/
#313660000000
1!
1'
1/
#313670000000
0!
0'
0/
#313680000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#313690000000
0!
0'
0/
#313700000000
1!
1'
1/
#313710000000
0!
0'
0/
#313720000000
1!
1'
1/
#313730000000
0!
0'
0/
#313740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#313750000000
0!
0'
0/
#313760000000
1!
1'
1/
#313770000000
0!
0'
0/
#313780000000
1!
1'
1/
#313790000000
0!
0'
0/
#313800000000
1!
1'
1/
#313810000000
0!
0'
0/
#313820000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#313830000000
0!
0'
0/
#313840000000
1!
1'
1/
#313850000000
0!
0'
0/
#313860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#313870000000
0!
0'
0/
#313880000000
1!
1'
1/
#313890000000
0!
0'
0/
#313900000000
#313910000000
1!
1'
1/
#313920000000
0!
0'
0/
#313930000000
1!
1'
1/
#313940000000
0!
1"
0'
1(
0/
10
#313950000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#313960000000
0!
0'
0/
#313970000000
1!
1'
1/
#313980000000
0!
0'
0/
#313990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#314000000000
0!
0'
0/
#314010000000
1!
1'
1/
#314020000000
0!
1"
0'
1(
0/
10
#314030000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#314040000000
0!
1$
0'
1+
0/
#314050000000
1!
1'
1/
#314060000000
0!
0'
0/
#314070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#314080000000
0!
0'
0/
#314090000000
1!
1'
1/
#314100000000
0!
0'
0/
#314110000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#314120000000
0!
0'
0/
#314130000000
1!
1'
1/
#314140000000
0!
0'
0/
#314150000000
1!
1'
1/
#314160000000
0!
0'
0/
#314170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#314180000000
0!
0'
0/
#314190000000
1!
1'
1/
#314200000000
0!
0'
0/
#314210000000
1!
1'
1/
#314220000000
0!
0'
0/
#314230000000
1!
1'
1/
#314240000000
0!
0'
0/
#314250000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#314260000000
0!
0'
0/
#314270000000
1!
1'
1/
#314280000000
0!
0'
0/
#314290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#314300000000
0!
0'
0/
#314310000000
1!
1'
1/
#314320000000
0!
0'
0/
#314330000000
#314340000000
1!
1'
1/
#314350000000
0!
0'
0/
#314360000000
1!
1'
1/
#314370000000
0!
1"
0'
1(
0/
10
#314380000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#314390000000
0!
0'
0/
#314400000000
1!
1'
1/
#314410000000
0!
0'
0/
#314420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#314430000000
0!
0'
0/
#314440000000
1!
1'
1/
#314450000000
0!
1"
0'
1(
0/
10
#314460000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#314470000000
0!
1$
0'
1+
0/
#314480000000
1!
1'
1/
#314490000000
0!
0'
0/
#314500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#314510000000
0!
0'
0/
#314520000000
1!
1'
1/
#314530000000
0!
0'
0/
#314540000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#314550000000
0!
0'
0/
#314560000000
1!
1'
1/
#314570000000
0!
0'
0/
#314580000000
1!
1'
1/
#314590000000
0!
0'
0/
#314600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#314610000000
0!
0'
0/
#314620000000
1!
1'
1/
#314630000000
0!
0'
0/
#314640000000
1!
1'
1/
#314650000000
0!
0'
0/
#314660000000
1!
1'
1/
#314670000000
0!
0'
0/
#314680000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#314690000000
0!
0'
0/
#314700000000
1!
1'
1/
#314710000000
0!
0'
0/
#314720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#314730000000
0!
0'
0/
#314740000000
1!
1'
1/
#314750000000
0!
0'
0/
#314760000000
#314770000000
1!
1'
1/
#314780000000
0!
0'
0/
#314790000000
1!
1'
1/
#314800000000
0!
1"
0'
1(
0/
10
#314810000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#314820000000
0!
0'
0/
#314830000000
1!
1'
1/
#314840000000
0!
0'
0/
#314850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#314860000000
0!
0'
0/
#314870000000
1!
1'
1/
#314880000000
0!
1"
0'
1(
0/
10
#314890000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#314900000000
0!
1$
0'
1+
0/
#314910000000
1!
1'
1/
#314920000000
0!
0'
0/
#314930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#314940000000
0!
0'
0/
#314950000000
1!
1'
1/
#314960000000
0!
0'
0/
#314970000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#314980000000
0!
0'
0/
#314990000000
1!
1'
1/
#315000000000
0!
0'
0/
#315010000000
1!
1'
1/
#315020000000
0!
0'
0/
#315030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#315040000000
0!
0'
0/
#315050000000
1!
1'
1/
#315060000000
0!
0'
0/
#315070000000
1!
1'
1/
#315080000000
0!
0'
0/
#315090000000
1!
1'
1/
#315100000000
0!
0'
0/
#315110000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#315120000000
0!
0'
0/
#315130000000
1!
1'
1/
#315140000000
0!
0'
0/
#315150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#315160000000
0!
0'
0/
#315170000000
1!
1'
1/
#315180000000
0!
0'
0/
#315190000000
#315200000000
1!
1'
1/
#315210000000
0!
0'
0/
#315220000000
1!
1'
1/
#315230000000
0!
1"
0'
1(
0/
10
#315240000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#315250000000
0!
0'
0/
#315260000000
1!
1'
1/
#315270000000
0!
0'
0/
#315280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#315290000000
0!
0'
0/
#315300000000
1!
1'
1/
#315310000000
0!
1"
0'
1(
0/
10
#315320000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#315330000000
0!
1$
0'
1+
0/
#315340000000
1!
1'
1/
#315350000000
0!
0'
0/
#315360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#315370000000
0!
0'
0/
#315380000000
1!
1'
1/
#315390000000
0!
0'
0/
#315400000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#315410000000
0!
0'
0/
#315420000000
1!
1'
1/
#315430000000
0!
0'
0/
#315440000000
1!
1'
1/
#315450000000
0!
0'
0/
#315460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#315470000000
0!
0'
0/
#315480000000
1!
1'
1/
#315490000000
0!
0'
0/
#315500000000
1!
1'
1/
#315510000000
0!
0'
0/
#315520000000
1!
1'
1/
#315530000000
0!
0'
0/
#315540000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#315550000000
0!
0'
0/
#315560000000
1!
1'
1/
#315570000000
0!
0'
0/
#315580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#315590000000
0!
0'
0/
#315600000000
1!
1'
1/
#315610000000
0!
0'
0/
#315620000000
#315630000000
1!
1'
1/
#315640000000
0!
0'
0/
#315650000000
1!
1'
1/
#315660000000
0!
1"
0'
1(
0/
10
#315670000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#315680000000
0!
0'
0/
#315690000000
1!
1'
1/
#315700000000
0!
0'
0/
#315710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#315720000000
0!
0'
0/
#315730000000
1!
1'
1/
#315740000000
0!
1"
0'
1(
0/
10
#315750000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#315760000000
0!
1$
0'
1+
0/
#315770000000
1!
1'
1/
#315780000000
0!
0'
0/
#315790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#315800000000
0!
0'
0/
#315810000000
1!
1'
1/
#315820000000
0!
0'
0/
#315830000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#315840000000
0!
0'
0/
#315850000000
1!
1'
1/
#315860000000
0!
0'
0/
#315870000000
1!
1'
1/
#315880000000
0!
0'
0/
#315890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#315900000000
0!
0'
0/
#315910000000
1!
1'
1/
#315920000000
0!
0'
0/
#315930000000
1!
1'
1/
#315940000000
0!
0'
0/
#315950000000
1!
1'
1/
#315960000000
0!
0'
0/
#315970000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#315980000000
0!
0'
0/
#315990000000
1!
1'
1/
#316000000000
0!
0'
0/
#316010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#316020000000
0!
0'
0/
#316030000000
1!
1'
1/
#316040000000
0!
0'
0/
#316050000000
#316060000000
1!
1'
1/
#316070000000
0!
0'
0/
#316080000000
1!
1'
1/
#316090000000
0!
1"
0'
1(
0/
10
#316100000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#316110000000
0!
0'
0/
#316120000000
1!
1'
1/
#316130000000
0!
0'
0/
#316140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#316150000000
0!
0'
0/
#316160000000
1!
1'
1/
#316170000000
0!
1"
0'
1(
0/
10
#316180000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#316190000000
0!
1$
0'
1+
0/
#316200000000
1!
1'
1/
#316210000000
0!
0'
0/
#316220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#316230000000
0!
0'
0/
#316240000000
1!
1'
1/
#316250000000
0!
0'
0/
#316260000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#316270000000
0!
0'
0/
#316280000000
1!
1'
1/
#316290000000
0!
0'
0/
#316300000000
1!
1'
1/
#316310000000
0!
0'
0/
#316320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#316330000000
0!
0'
0/
#316340000000
1!
1'
1/
#316350000000
0!
0'
0/
#316360000000
1!
1'
1/
#316370000000
0!
0'
0/
#316380000000
1!
1'
1/
#316390000000
0!
0'
0/
#316400000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#316410000000
0!
0'
0/
#316420000000
1!
1'
1/
#316430000000
0!
0'
0/
#316440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#316450000000
0!
0'
0/
#316460000000
1!
1'
1/
#316470000000
0!
0'
0/
#316480000000
#316490000000
1!
1'
1/
#316500000000
0!
0'
0/
#316510000000
1!
1'
1/
#316520000000
0!
1"
0'
1(
0/
10
#316530000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#316540000000
0!
0'
0/
#316550000000
1!
1'
1/
#316560000000
0!
0'
0/
#316570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#316580000000
0!
0'
0/
#316590000000
1!
1'
1/
#316600000000
0!
1"
0'
1(
0/
10
#316610000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#316620000000
0!
1$
0'
1+
0/
#316630000000
1!
1'
1/
#316640000000
0!
0'
0/
#316650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#316660000000
0!
0'
0/
#316670000000
1!
1'
1/
#316680000000
0!
0'
0/
#316690000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#316700000000
0!
0'
0/
#316710000000
1!
1'
1/
#316720000000
0!
0'
0/
#316730000000
1!
1'
1/
#316740000000
0!
0'
0/
#316750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#316760000000
0!
0'
0/
#316770000000
1!
1'
1/
#316780000000
0!
0'
0/
#316790000000
1!
1'
1/
#316800000000
0!
0'
0/
#316810000000
1!
1'
1/
#316820000000
0!
0'
0/
#316830000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#316840000000
0!
0'
0/
#316850000000
1!
1'
1/
#316860000000
0!
0'
0/
#316870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#316880000000
0!
0'
0/
#316890000000
1!
1'
1/
#316900000000
0!
0'
0/
#316910000000
#316920000000
1!
1'
1/
#316930000000
0!
0'
0/
#316940000000
1!
1'
1/
#316950000000
0!
1"
0'
1(
0/
10
#316960000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#316970000000
0!
0'
0/
#316980000000
1!
1'
1/
#316990000000
0!
0'
0/
#317000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#317010000000
0!
0'
0/
#317020000000
1!
1'
1/
#317030000000
0!
1"
0'
1(
0/
10
#317040000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#317050000000
0!
1$
0'
1+
0/
#317060000000
1!
1'
1/
#317070000000
0!
0'
0/
#317080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#317090000000
0!
0'
0/
#317100000000
1!
1'
1/
#317110000000
0!
0'
0/
#317120000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#317130000000
0!
0'
0/
#317140000000
1!
1'
1/
#317150000000
0!
0'
0/
#317160000000
1!
1'
1/
#317170000000
0!
0'
0/
#317180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#317190000000
0!
0'
0/
#317200000000
1!
1'
1/
#317210000000
0!
0'
0/
#317220000000
1!
1'
1/
#317230000000
0!
0'
0/
#317240000000
1!
1'
1/
#317250000000
0!
0'
0/
#317260000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#317270000000
0!
0'
0/
#317280000000
1!
1'
1/
#317290000000
0!
0'
0/
#317300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#317310000000
0!
0'
0/
#317320000000
1!
1'
1/
#317330000000
0!
0'
0/
#317340000000
#317350000000
1!
1'
1/
#317360000000
0!
0'
0/
#317370000000
1!
1'
1/
#317380000000
0!
1"
0'
1(
0/
10
#317390000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#317400000000
0!
0'
0/
#317410000000
1!
1'
1/
#317420000000
0!
0'
0/
#317430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#317440000000
0!
0'
0/
#317450000000
1!
1'
1/
#317460000000
0!
1"
0'
1(
0/
10
#317470000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#317480000000
0!
1$
0'
1+
0/
#317490000000
1!
1'
1/
#317500000000
0!
0'
0/
#317510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#317520000000
0!
0'
0/
#317530000000
1!
1'
1/
#317540000000
0!
0'
0/
#317550000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#317560000000
0!
0'
0/
#317570000000
1!
1'
1/
#317580000000
0!
0'
0/
#317590000000
1!
1'
1/
#317600000000
0!
0'
0/
#317610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#317620000000
0!
0'
0/
#317630000000
1!
1'
1/
#317640000000
0!
0'
0/
#317650000000
1!
1'
1/
#317660000000
0!
0'
0/
#317670000000
1!
1'
1/
#317680000000
0!
0'
0/
#317690000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#317700000000
0!
0'
0/
#317710000000
1!
1'
1/
#317720000000
0!
0'
0/
#317730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#317740000000
0!
0'
0/
#317750000000
1!
1'
1/
#317760000000
0!
0'
0/
#317770000000
#317780000000
1!
1'
1/
#317790000000
0!
0'
0/
#317800000000
1!
1'
1/
#317810000000
0!
1"
0'
1(
0/
10
#317820000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#317830000000
0!
0'
0/
#317840000000
1!
1'
1/
#317850000000
0!
0'
0/
#317860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#317870000000
0!
0'
0/
#317880000000
1!
1'
1/
#317890000000
0!
1"
0'
1(
0/
10
#317900000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#317910000000
0!
1$
0'
1+
0/
#317920000000
1!
1'
1/
#317930000000
0!
0'
0/
#317940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#317950000000
0!
0'
0/
#317960000000
1!
1'
1/
#317970000000
0!
0'
0/
#317980000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#317990000000
0!
0'
0/
#318000000000
1!
1'
1/
#318010000000
0!
0'
0/
#318020000000
1!
1'
1/
#318030000000
0!
0'
0/
#318040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#318050000000
0!
0'
0/
#318060000000
1!
1'
1/
#318070000000
0!
0'
0/
#318080000000
1!
1'
1/
#318090000000
0!
0'
0/
#318100000000
1!
1'
1/
#318110000000
0!
0'
0/
#318120000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#318130000000
0!
0'
0/
#318140000000
1!
1'
1/
#318150000000
0!
0'
0/
#318160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#318170000000
0!
0'
0/
#318180000000
1!
1'
1/
#318190000000
0!
0'
0/
#318200000000
#318210000000
1!
1'
1/
#318220000000
0!
0'
0/
#318230000000
1!
1'
1/
#318240000000
0!
1"
0'
1(
0/
10
#318250000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#318260000000
0!
0'
0/
#318270000000
1!
1'
1/
#318280000000
0!
0'
0/
#318290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#318300000000
0!
0'
0/
#318310000000
1!
1'
1/
#318320000000
0!
1"
0'
1(
0/
10
#318330000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#318340000000
0!
1$
0'
1+
0/
#318350000000
1!
1'
1/
#318360000000
0!
0'
0/
#318370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#318380000000
0!
0'
0/
#318390000000
1!
1'
1/
#318400000000
0!
0'
0/
#318410000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#318420000000
0!
0'
0/
#318430000000
1!
1'
1/
#318440000000
0!
0'
0/
#318450000000
1!
1'
1/
#318460000000
0!
0'
0/
#318470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#318480000000
0!
0'
0/
#318490000000
1!
1'
1/
#318500000000
0!
0'
0/
#318510000000
1!
1'
1/
#318520000000
0!
0'
0/
#318530000000
1!
1'
1/
#318540000000
0!
0'
0/
#318550000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#318560000000
0!
0'
0/
#318570000000
1!
1'
1/
#318580000000
0!
0'
0/
#318590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#318600000000
0!
0'
0/
#318610000000
1!
1'
1/
#318620000000
0!
0'
0/
#318630000000
#318640000000
1!
1'
1/
#318650000000
0!
0'
0/
#318660000000
1!
1'
1/
#318670000000
0!
1"
0'
1(
0/
10
#318680000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#318690000000
0!
0'
0/
#318700000000
1!
1'
1/
#318710000000
0!
0'
0/
#318720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#318730000000
0!
0'
0/
#318740000000
1!
1'
1/
#318750000000
0!
1"
0'
1(
0/
10
#318760000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#318770000000
0!
1$
0'
1+
0/
#318780000000
1!
1'
1/
#318790000000
0!
0'
0/
#318800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#318810000000
0!
0'
0/
#318820000000
1!
1'
1/
#318830000000
0!
0'
0/
#318840000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#318850000000
0!
0'
0/
#318860000000
1!
1'
1/
#318870000000
0!
0'
0/
#318880000000
1!
1'
1/
#318890000000
0!
0'
0/
#318900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#318910000000
0!
0'
0/
#318920000000
1!
1'
1/
#318930000000
0!
0'
0/
#318940000000
1!
1'
1/
#318950000000
0!
0'
0/
#318960000000
1!
1'
1/
#318970000000
0!
0'
0/
#318980000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#318990000000
0!
0'
0/
#319000000000
1!
1'
1/
#319010000000
0!
0'
0/
#319020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#319030000000
0!
0'
0/
#319040000000
1!
1'
1/
#319050000000
0!
0'
0/
#319060000000
#319070000000
1!
1'
1/
#319080000000
0!
0'
0/
#319090000000
1!
1'
1/
#319100000000
0!
1"
0'
1(
0/
10
#319110000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#319120000000
0!
0'
0/
#319130000000
1!
1'
1/
#319140000000
0!
0'
0/
#319150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#319160000000
0!
0'
0/
#319170000000
1!
1'
1/
#319180000000
0!
1"
0'
1(
0/
10
#319190000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#319200000000
0!
1$
0'
1+
0/
#319210000000
1!
1'
1/
#319220000000
0!
0'
0/
#319230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#319240000000
0!
0'
0/
#319250000000
1!
1'
1/
#319260000000
0!
0'
0/
#319270000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#319280000000
0!
0'
0/
#319290000000
1!
1'
1/
#319300000000
0!
0'
0/
#319310000000
1!
1'
1/
#319320000000
0!
0'
0/
#319330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#319340000000
0!
0'
0/
#319350000000
1!
1'
1/
#319360000000
0!
0'
0/
#319370000000
1!
1'
1/
#319380000000
0!
0'
0/
#319390000000
1!
1'
1/
#319400000000
0!
0'
0/
#319410000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#319420000000
0!
0'
0/
#319430000000
1!
1'
1/
#319440000000
0!
0'
0/
#319450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#319460000000
0!
0'
0/
#319470000000
1!
1'
1/
#319480000000
0!
0'
0/
#319490000000
#319500000000
1!
1'
1/
#319510000000
0!
0'
0/
#319520000000
1!
1'
1/
#319530000000
0!
1"
0'
1(
0/
10
#319540000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#319550000000
0!
0'
0/
#319560000000
1!
1'
1/
#319570000000
0!
0'
0/
#319580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#319590000000
0!
0'
0/
#319600000000
1!
1'
1/
#319610000000
0!
1"
0'
1(
0/
10
#319620000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#319630000000
0!
1$
0'
1+
0/
#319640000000
1!
1'
1/
#319650000000
0!
0'
0/
#319660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#319670000000
0!
0'
0/
#319680000000
1!
1'
1/
#319690000000
0!
0'
0/
#319700000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#319710000000
0!
0'
0/
#319720000000
1!
1'
1/
#319730000000
0!
0'
0/
#319740000000
1!
1'
1/
#319750000000
0!
0'
0/
#319760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#319770000000
0!
0'
0/
#319780000000
1!
1'
1/
#319790000000
0!
0'
0/
#319800000000
1!
1'
1/
#319810000000
0!
0'
0/
#319820000000
1!
1'
1/
#319830000000
0!
0'
0/
#319840000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#319850000000
0!
0'
0/
#319860000000
1!
1'
1/
#319870000000
0!
0'
0/
#319880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#319890000000
0!
0'
0/
#319900000000
1!
1'
1/
#319910000000
0!
0'
0/
#319920000000
#319930000000
1!
1'
1/
#319940000000
0!
0'
0/
#319950000000
1!
1'
1/
#319960000000
0!
1"
0'
1(
0/
10
#319970000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#319980000000
0!
0'
0/
#319990000000
1!
1'
1/
#320000000000
0!
0'
0/
#320010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#320020000000
0!
0'
0/
#320030000000
1!
1'
1/
#320040000000
0!
1"
0'
1(
0/
10
#320050000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#320060000000
0!
1$
0'
1+
0/
#320070000000
1!
1'
1/
#320080000000
0!
0'
0/
#320090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#320100000000
0!
0'
0/
#320110000000
1!
1'
1/
#320120000000
0!
0'
0/
#320130000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#320140000000
0!
0'
0/
#320150000000
1!
1'
1/
#320160000000
0!
0'
0/
#320170000000
1!
1'
1/
#320180000000
0!
0'
0/
#320190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#320200000000
0!
0'
0/
#320210000000
1!
1'
1/
#320220000000
0!
0'
0/
#320230000000
1!
1'
1/
#320240000000
0!
0'
0/
#320250000000
1!
1'
1/
#320260000000
0!
0'
0/
#320270000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#320280000000
0!
0'
0/
#320290000000
1!
1'
1/
#320300000000
0!
0'
0/
#320310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#320320000000
0!
0'
0/
#320330000000
1!
1'
1/
#320340000000
0!
0'
0/
#320350000000
#320360000000
1!
1'
1/
#320370000000
0!
0'
0/
#320380000000
1!
1'
1/
#320390000000
0!
1"
0'
1(
0/
10
#320400000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#320410000000
0!
0'
0/
#320420000000
1!
1'
1/
#320430000000
0!
0'
0/
#320440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#320450000000
0!
0'
0/
#320460000000
1!
1'
1/
#320470000000
0!
1"
0'
1(
0/
10
#320480000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#320490000000
0!
1$
0'
1+
0/
#320500000000
1!
1'
1/
#320510000000
0!
0'
0/
#320520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#320530000000
0!
0'
0/
#320540000000
1!
1'
1/
#320550000000
0!
0'
0/
#320560000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#320570000000
0!
0'
0/
#320580000000
1!
1'
1/
#320590000000
0!
0'
0/
#320600000000
1!
1'
1/
#320610000000
0!
0'
0/
#320620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#320630000000
0!
0'
0/
#320640000000
1!
1'
1/
#320650000000
0!
0'
0/
#320660000000
1!
1'
1/
#320670000000
0!
0'
0/
#320680000000
1!
1'
1/
#320690000000
0!
0'
0/
#320700000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#320710000000
0!
0'
0/
#320720000000
1!
1'
1/
#320730000000
0!
0'
0/
#320740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#320750000000
0!
0'
0/
#320760000000
1!
1'
1/
#320770000000
0!
0'
0/
#320780000000
#320790000000
1!
1'
1/
#320800000000
0!
0'
0/
#320810000000
1!
1'
1/
#320820000000
0!
1"
0'
1(
0/
10
#320830000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#320840000000
0!
0'
0/
#320850000000
1!
1'
1/
#320860000000
0!
0'
0/
#320870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#320880000000
0!
0'
0/
#320890000000
1!
1'
1/
#320900000000
0!
1"
0'
1(
0/
10
#320910000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#320920000000
0!
1$
0'
1+
0/
#320930000000
1!
1'
1/
#320940000000
0!
0'
0/
#320950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#320960000000
0!
0'
0/
#320970000000
1!
1'
1/
#320980000000
0!
0'
0/
#320990000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#321000000000
0!
0'
0/
#321010000000
1!
1'
1/
#321020000000
0!
0'
0/
#321030000000
1!
1'
1/
#321040000000
0!
0'
0/
#321050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#321060000000
0!
0'
0/
#321070000000
1!
1'
1/
#321080000000
0!
0'
0/
#321090000000
1!
1'
1/
#321100000000
0!
0'
0/
#321110000000
1!
1'
1/
#321120000000
0!
0'
0/
#321130000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#321140000000
0!
0'
0/
#321150000000
1!
1'
1/
#321160000000
0!
0'
0/
#321170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#321180000000
0!
0'
0/
#321190000000
1!
1'
1/
#321200000000
0!
0'
0/
#321210000000
#321220000000
1!
1'
1/
#321230000000
0!
0'
0/
#321240000000
1!
1'
1/
#321250000000
0!
1"
0'
1(
0/
10
#321260000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#321270000000
0!
0'
0/
#321280000000
1!
1'
1/
#321290000000
0!
0'
0/
#321300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#321310000000
0!
0'
0/
#321320000000
1!
1'
1/
#321330000000
0!
1"
0'
1(
0/
10
#321340000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#321350000000
0!
1$
0'
1+
0/
#321360000000
1!
1'
1/
#321370000000
0!
0'
0/
#321380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#321390000000
0!
0'
0/
#321400000000
1!
1'
1/
#321410000000
0!
0'
0/
#321420000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#321430000000
0!
0'
0/
#321440000000
1!
1'
1/
#321450000000
0!
0'
0/
#321460000000
1!
1'
1/
#321470000000
0!
0'
0/
#321480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#321490000000
0!
0'
0/
#321500000000
1!
1'
1/
#321510000000
0!
0'
0/
#321520000000
1!
1'
1/
#321530000000
0!
0'
0/
#321540000000
1!
1'
1/
#321550000000
0!
0'
0/
#321560000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#321570000000
0!
0'
0/
#321580000000
1!
1'
1/
#321590000000
0!
0'
0/
#321600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#321610000000
0!
0'
0/
#321620000000
1!
1'
1/
#321630000000
0!
0'
0/
#321640000000
#321650000000
1!
1'
1/
#321660000000
0!
0'
0/
#321670000000
1!
1'
1/
#321680000000
0!
1"
0'
1(
0/
10
#321690000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#321700000000
0!
0'
0/
#321710000000
1!
1'
1/
#321720000000
0!
0'
0/
#321730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#321740000000
0!
0'
0/
#321750000000
1!
1'
1/
#321760000000
0!
1"
0'
1(
0/
10
#321770000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#321780000000
0!
1$
0'
1+
0/
#321790000000
1!
1'
1/
#321800000000
0!
0'
0/
#321810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#321820000000
0!
0'
0/
#321830000000
1!
1'
1/
#321840000000
0!
0'
0/
#321850000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#321860000000
0!
0'
0/
#321870000000
1!
1'
1/
#321880000000
0!
0'
0/
#321890000000
1!
1'
1/
#321900000000
0!
0'
0/
#321910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#321920000000
0!
0'
0/
#321930000000
1!
1'
1/
#321940000000
0!
0'
0/
#321950000000
1!
1'
1/
#321960000000
0!
0'
0/
#321970000000
1!
1'
1/
#321980000000
0!
0'
0/
#321990000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#322000000000
0!
0'
0/
#322010000000
1!
1'
1/
#322020000000
0!
0'
0/
#322030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#322040000000
0!
0'
0/
#322050000000
1!
1'
1/
#322060000000
0!
0'
0/
#322070000000
#322080000000
1!
1'
1/
#322090000000
0!
0'
0/
#322100000000
1!
1'
1/
#322110000000
0!
1"
0'
1(
0/
10
#322120000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#322130000000
0!
0'
0/
#322140000000
1!
1'
1/
#322150000000
0!
0'
0/
#322160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#322170000000
0!
0'
0/
#322180000000
1!
1'
1/
#322190000000
0!
1"
0'
1(
0/
10
#322200000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#322210000000
0!
1$
0'
1+
0/
#322220000000
1!
1'
1/
#322230000000
0!
0'
0/
#322240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#322250000000
0!
0'
0/
#322260000000
1!
1'
1/
#322270000000
0!
0'
0/
#322280000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#322290000000
0!
0'
0/
#322300000000
1!
1'
1/
#322310000000
0!
0'
0/
#322320000000
1!
1'
1/
#322330000000
0!
0'
0/
#322340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#322350000000
0!
0'
0/
#322360000000
1!
1'
1/
#322370000000
0!
0'
0/
#322380000000
1!
1'
1/
#322390000000
0!
0'
0/
#322400000000
1!
1'
1/
#322410000000
0!
0'
0/
#322420000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#322430000000
0!
0'
0/
#322440000000
1!
1'
1/
#322450000000
0!
0'
0/
#322460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#322470000000
0!
0'
0/
#322480000000
1!
1'
1/
#322490000000
0!
0'
0/
#322500000000
#322510000000
1!
1'
1/
#322520000000
0!
0'
0/
#322530000000
1!
1'
1/
#322540000000
0!
1"
0'
1(
0/
10
#322550000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#322560000000
0!
0'
0/
#322570000000
1!
1'
1/
#322580000000
0!
0'
0/
#322590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#322600000000
0!
0'
0/
#322610000000
1!
1'
1/
#322620000000
0!
1"
0'
1(
0/
10
#322630000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#322640000000
0!
1$
0'
1+
0/
#322650000000
1!
1'
1/
#322660000000
0!
0'
0/
#322670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#322680000000
0!
0'
0/
#322690000000
1!
1'
1/
#322700000000
0!
0'
0/
#322710000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#322720000000
0!
0'
0/
#322730000000
1!
1'
1/
#322740000000
0!
0'
0/
#322750000000
1!
1'
1/
#322760000000
0!
0'
0/
#322770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#322780000000
0!
0'
0/
#322790000000
1!
1'
1/
#322800000000
0!
0'
0/
#322810000000
1!
1'
1/
#322820000000
0!
0'
0/
#322830000000
1!
1'
1/
#322840000000
0!
0'
0/
#322850000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#322860000000
0!
0'
0/
#322870000000
1!
1'
1/
#322880000000
0!
0'
0/
#322890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#322900000000
0!
0'
0/
#322910000000
1!
1'
1/
#322920000000
0!
0'
0/
#322930000000
#322940000000
1!
1'
1/
#322950000000
0!
0'
0/
#322960000000
1!
1'
1/
#322970000000
0!
1"
0'
1(
0/
10
#322980000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#322990000000
0!
0'
0/
#323000000000
1!
1'
1/
#323010000000
0!
0'
0/
#323020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#323030000000
0!
0'
0/
#323040000000
1!
1'
1/
#323050000000
0!
1"
0'
1(
0/
10
#323060000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#323070000000
0!
1$
0'
1+
0/
#323080000000
1!
1'
1/
#323090000000
0!
0'
0/
#323100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#323110000000
0!
0'
0/
#323120000000
1!
1'
1/
#323130000000
0!
0'
0/
#323140000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#323150000000
0!
0'
0/
#323160000000
1!
1'
1/
#323170000000
0!
0'
0/
#323180000000
1!
1'
1/
#323190000000
0!
0'
0/
#323200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#323210000000
0!
0'
0/
#323220000000
1!
1'
1/
#323230000000
0!
0'
0/
#323240000000
1!
1'
1/
#323250000000
0!
0'
0/
#323260000000
1!
1'
1/
#323270000000
0!
0'
0/
#323280000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#323290000000
0!
0'
0/
#323300000000
1!
1'
1/
#323310000000
0!
0'
0/
#323320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#323330000000
0!
0'
0/
#323340000000
1!
1'
1/
#323350000000
0!
0'
0/
#323360000000
#323370000000
1!
1'
1/
#323380000000
0!
0'
0/
#323390000000
1!
1'
1/
#323400000000
0!
1"
0'
1(
0/
10
#323410000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#323420000000
0!
0'
0/
#323430000000
1!
1'
1/
#323440000000
0!
0'
0/
#323450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#323460000000
0!
0'
0/
#323470000000
1!
1'
1/
#323480000000
0!
1"
0'
1(
0/
10
#323490000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#323500000000
0!
1$
0'
1+
0/
#323510000000
1!
1'
1/
#323520000000
0!
0'
0/
#323530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#323540000000
0!
0'
0/
#323550000000
1!
1'
1/
#323560000000
0!
0'
0/
#323570000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#323580000000
0!
0'
0/
#323590000000
1!
1'
1/
#323600000000
0!
0'
0/
#323610000000
1!
1'
1/
#323620000000
0!
0'
0/
#323630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#323640000000
0!
0'
0/
#323650000000
1!
1'
1/
#323660000000
0!
0'
0/
#323670000000
1!
1'
1/
#323680000000
0!
0'
0/
#323690000000
1!
1'
1/
#323700000000
0!
0'
0/
#323710000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#323720000000
0!
0'
0/
#323730000000
1!
1'
1/
#323740000000
0!
0'
0/
#323750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#323760000000
0!
0'
0/
#323770000000
1!
1'
1/
#323780000000
0!
0'
0/
#323790000000
#323800000000
1!
1'
1/
#323810000000
0!
0'
0/
#323820000000
1!
1'
1/
#323830000000
0!
1"
0'
1(
0/
10
#323840000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#323850000000
0!
0'
0/
#323860000000
1!
1'
1/
#323870000000
0!
0'
0/
#323880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#323890000000
0!
0'
0/
#323900000000
1!
1'
1/
#323910000000
0!
1"
0'
1(
0/
10
#323920000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#323930000000
0!
1$
0'
1+
0/
#323940000000
1!
1'
1/
#323950000000
0!
0'
0/
#323960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#323970000000
0!
0'
0/
#323980000000
1!
1'
1/
#323990000000
0!
0'
0/
#324000000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#324010000000
0!
0'
0/
#324020000000
1!
1'
1/
#324030000000
0!
0'
0/
#324040000000
1!
1'
1/
#324050000000
0!
0'
0/
#324060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#324070000000
0!
0'
0/
#324080000000
1!
1'
1/
#324090000000
0!
0'
0/
#324100000000
1!
1'
1/
#324110000000
0!
0'
0/
#324120000000
1!
1'
1/
#324130000000
0!
0'
0/
#324140000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#324150000000
0!
0'
0/
#324160000000
1!
1'
1/
#324170000000
0!
0'
0/
#324180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#324190000000
0!
0'
0/
#324200000000
1!
1'
1/
#324210000000
0!
0'
0/
#324220000000
#324230000000
1!
1'
1/
#324240000000
0!
0'
0/
#324250000000
1!
1'
1/
#324260000000
0!
1"
0'
1(
0/
10
#324270000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#324280000000
0!
0'
0/
#324290000000
1!
1'
1/
#324300000000
0!
0'
0/
#324310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#324320000000
0!
0'
0/
#324330000000
1!
1'
1/
#324340000000
0!
1"
0'
1(
0/
10
#324350000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#324360000000
0!
1$
0'
1+
0/
#324370000000
1!
1'
1/
#324380000000
0!
0'
0/
#324390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#324400000000
0!
0'
0/
#324410000000
1!
1'
1/
#324420000000
0!
0'
0/
#324430000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#324440000000
0!
0'
0/
#324450000000
1!
1'
1/
#324460000000
0!
0'
0/
#324470000000
1!
1'
1/
#324480000000
0!
0'
0/
#324490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#324500000000
0!
0'
0/
#324510000000
1!
1'
1/
#324520000000
0!
0'
0/
#324530000000
1!
1'
1/
#324540000000
0!
0'
0/
#324550000000
1!
1'
1/
#324560000000
0!
0'
0/
#324570000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#324580000000
0!
0'
0/
#324590000000
1!
1'
1/
#324600000000
0!
0'
0/
#324610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#324620000000
0!
0'
0/
#324630000000
1!
1'
1/
#324640000000
0!
0'
0/
#324650000000
#324660000000
1!
1'
1/
#324670000000
0!
0'
0/
#324680000000
1!
1'
1/
#324690000000
0!
1"
0'
1(
0/
10
#324700000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#324710000000
0!
0'
0/
#324720000000
1!
1'
1/
#324730000000
0!
0'
0/
#324740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#324750000000
0!
0'
0/
#324760000000
1!
1'
1/
#324770000000
0!
1"
0'
1(
0/
10
#324780000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#324790000000
0!
1$
0'
1+
0/
#324800000000
1!
1'
1/
#324810000000
0!
0'
0/
#324820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#324830000000
0!
0'
0/
#324840000000
1!
1'
1/
#324850000000
0!
0'
0/
#324860000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#324870000000
0!
0'
0/
#324880000000
1!
1'
1/
#324890000000
0!
0'
0/
#324900000000
1!
1'
1/
#324910000000
0!
0'
0/
#324920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#324930000000
0!
0'
0/
#324940000000
1!
1'
1/
#324950000000
0!
0'
0/
#324960000000
1!
1'
1/
#324970000000
0!
0'
0/
#324980000000
1!
1'
1/
#324990000000
0!
0'
0/
#325000000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#325010000000
0!
0'
0/
#325020000000
1!
1'
1/
#325030000000
0!
0'
0/
#325040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#325050000000
0!
0'
0/
#325060000000
1!
1'
1/
#325070000000
0!
0'
0/
#325080000000
#325090000000
1!
1'
1/
#325100000000
0!
0'
0/
#325110000000
1!
1'
1/
#325120000000
0!
1"
0'
1(
0/
10
#325130000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#325140000000
0!
0'
0/
#325150000000
1!
1'
1/
#325160000000
0!
0'
0/
#325170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#325180000000
0!
0'
0/
#325190000000
1!
1'
1/
#325200000000
0!
1"
0'
1(
0/
10
#325210000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#325220000000
0!
1$
0'
1+
0/
#325230000000
1!
1'
1/
#325240000000
0!
0'
0/
#325250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#325260000000
0!
0'
0/
#325270000000
1!
1'
1/
#325280000000
0!
0'
0/
#325290000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#325300000000
0!
0'
0/
#325310000000
1!
1'
1/
#325320000000
0!
0'
0/
#325330000000
1!
1'
1/
#325340000000
0!
0'
0/
#325350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#325360000000
0!
0'
0/
#325370000000
1!
1'
1/
#325380000000
0!
0'
0/
#325390000000
1!
1'
1/
#325400000000
0!
0'
0/
#325410000000
1!
1'
1/
#325420000000
0!
0'
0/
#325430000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#325440000000
0!
0'
0/
#325450000000
1!
1'
1/
#325460000000
0!
0'
0/
#325470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#325480000000
0!
0'
0/
#325490000000
1!
1'
1/
#325500000000
0!
0'
0/
#325510000000
#325520000000
1!
1'
1/
#325530000000
0!
0'
0/
#325540000000
1!
1'
1/
#325550000000
0!
1"
0'
1(
0/
10
#325560000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#325570000000
0!
0'
0/
#325580000000
1!
1'
1/
#325590000000
0!
0'
0/
#325600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#325610000000
0!
0'
0/
#325620000000
1!
1'
1/
#325630000000
0!
1"
0'
1(
0/
10
#325640000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#325650000000
0!
1$
0'
1+
0/
#325660000000
1!
1'
1/
#325670000000
0!
0'
0/
#325680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#325690000000
0!
0'
0/
#325700000000
1!
1'
1/
#325710000000
0!
0'
0/
#325720000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#325730000000
0!
0'
0/
#325740000000
1!
1'
1/
#325750000000
0!
0'
0/
#325760000000
1!
1'
1/
#325770000000
0!
0'
0/
#325780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#325790000000
0!
0'
0/
#325800000000
1!
1'
1/
#325810000000
0!
0'
0/
#325820000000
1!
1'
1/
#325830000000
0!
0'
0/
#325840000000
1!
1'
1/
#325850000000
0!
0'
0/
#325860000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#325870000000
0!
0'
0/
#325880000000
1!
1'
1/
#325890000000
0!
0'
0/
#325900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#325910000000
0!
0'
0/
#325920000000
1!
1'
1/
#325930000000
0!
0'
0/
#325940000000
#325950000000
1!
1'
1/
#325960000000
0!
0'
0/
#325970000000
1!
1'
1/
#325980000000
0!
1"
0'
1(
0/
10
#325990000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#326000000000
0!
0'
0/
#326010000000
1!
1'
1/
#326020000000
0!
0'
0/
#326030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#326040000000
0!
0'
0/
#326050000000
1!
1'
1/
#326060000000
0!
1"
0'
1(
0/
10
#326070000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#326080000000
0!
1$
0'
1+
0/
#326090000000
1!
1'
1/
#326100000000
0!
0'
0/
#326110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#326120000000
0!
0'
0/
#326130000000
1!
1'
1/
#326140000000
0!
0'
0/
#326150000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#326160000000
0!
0'
0/
#326170000000
1!
1'
1/
#326180000000
0!
0'
0/
#326190000000
1!
1'
1/
#326200000000
0!
0'
0/
#326210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#326220000000
0!
0'
0/
#326230000000
1!
1'
1/
#326240000000
0!
0'
0/
#326250000000
1!
1'
1/
#326260000000
0!
0'
0/
#326270000000
1!
1'
1/
#326280000000
0!
0'
0/
#326290000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#326300000000
0!
0'
0/
#326310000000
1!
1'
1/
#326320000000
0!
0'
0/
#326330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#326340000000
0!
0'
0/
#326350000000
1!
1'
1/
#326360000000
0!
0'
0/
#326370000000
#326380000000
1!
1'
1/
#326390000000
0!
0'
0/
#326400000000
1!
1'
1/
#326410000000
0!
1"
0'
1(
0/
10
#326420000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#326430000000
0!
0'
0/
#326440000000
1!
1'
1/
#326450000000
0!
0'
0/
#326460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#326470000000
0!
0'
0/
#326480000000
1!
1'
1/
#326490000000
0!
1"
0'
1(
0/
10
#326500000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#326510000000
0!
1$
0'
1+
0/
#326520000000
1!
1'
1/
#326530000000
0!
0'
0/
#326540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#326550000000
0!
0'
0/
#326560000000
1!
1'
1/
#326570000000
0!
0'
0/
#326580000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#326590000000
0!
0'
0/
#326600000000
1!
1'
1/
#326610000000
0!
0'
0/
#326620000000
1!
1'
1/
#326630000000
0!
0'
0/
#326640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#326650000000
0!
0'
0/
#326660000000
1!
1'
1/
#326670000000
0!
0'
0/
#326680000000
1!
1'
1/
#326690000000
0!
0'
0/
#326700000000
1!
1'
1/
#326710000000
0!
0'
0/
#326720000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#326730000000
0!
0'
0/
#326740000000
1!
1'
1/
#326750000000
0!
0'
0/
#326760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#326770000000
0!
0'
0/
#326780000000
1!
1'
1/
#326790000000
0!
0'
0/
#326800000000
#326810000000
1!
1'
1/
#326820000000
0!
0'
0/
#326830000000
1!
1'
1/
#326840000000
0!
1"
0'
1(
0/
10
#326850000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#326860000000
0!
0'
0/
#326870000000
1!
1'
1/
#326880000000
0!
0'
0/
#326890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#326900000000
0!
0'
0/
#326910000000
1!
1'
1/
#326920000000
0!
1"
0'
1(
0/
10
#326930000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#326940000000
0!
1$
0'
1+
0/
#326950000000
1!
1'
1/
#326960000000
0!
0'
0/
#326970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#326980000000
0!
0'
0/
#326990000000
1!
1'
1/
#327000000000
0!
0'
0/
#327010000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#327020000000
0!
0'
0/
#327030000000
1!
1'
1/
#327040000000
0!
0'
0/
#327050000000
1!
1'
1/
#327060000000
0!
0'
0/
#327070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#327080000000
0!
0'
0/
#327090000000
1!
1'
1/
#327100000000
0!
0'
0/
#327110000000
1!
1'
1/
#327120000000
0!
0'
0/
#327130000000
1!
1'
1/
#327140000000
0!
0'
0/
#327150000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#327160000000
0!
0'
0/
#327170000000
1!
1'
1/
#327180000000
0!
0'
0/
#327190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#327200000000
0!
0'
0/
#327210000000
1!
1'
1/
#327220000000
0!
0'
0/
#327230000000
#327240000000
1!
1'
1/
#327250000000
0!
0'
0/
#327260000000
1!
1'
1/
#327270000000
0!
1"
0'
1(
0/
10
#327280000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#327290000000
0!
0'
0/
#327300000000
1!
1'
1/
#327310000000
0!
0'
0/
#327320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#327330000000
0!
0'
0/
#327340000000
1!
1'
1/
#327350000000
0!
1"
0'
1(
0/
10
#327360000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#327370000000
0!
1$
0'
1+
0/
#327380000000
1!
1'
1/
#327390000000
0!
0'
0/
#327400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#327410000000
0!
0'
0/
#327420000000
1!
1'
1/
#327430000000
0!
0'
0/
#327440000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#327450000000
0!
0'
0/
#327460000000
1!
1'
1/
#327470000000
0!
0'
0/
#327480000000
1!
1'
1/
#327490000000
0!
0'
0/
#327500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#327510000000
0!
0'
0/
#327520000000
1!
1'
1/
#327530000000
0!
0'
0/
#327540000000
1!
1'
1/
#327550000000
0!
0'
0/
#327560000000
1!
1'
1/
#327570000000
0!
0'
0/
#327580000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#327590000000
0!
0'
0/
#327600000000
1!
1'
1/
#327610000000
0!
0'
0/
#327620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#327630000000
0!
0'
0/
#327640000000
1!
1'
1/
#327650000000
0!
0'
0/
#327660000000
#327670000000
1!
1'
1/
#327680000000
0!
0'
0/
#327690000000
1!
1'
1/
#327700000000
0!
1"
0'
1(
0/
10
#327710000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#327720000000
0!
0'
0/
#327730000000
1!
1'
1/
#327740000000
0!
0'
0/
#327750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#327760000000
0!
0'
0/
#327770000000
1!
1'
1/
#327780000000
0!
1"
0'
1(
0/
10
#327790000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#327800000000
0!
1$
0'
1+
0/
#327810000000
1!
1'
1/
#327820000000
0!
0'
0/
#327830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#327840000000
0!
0'
0/
#327850000000
1!
1'
1/
#327860000000
0!
0'
0/
#327870000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#327880000000
0!
0'
0/
#327890000000
1!
1'
1/
#327900000000
0!
0'
0/
#327910000000
1!
1'
1/
#327920000000
0!
0'
0/
#327930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#327940000000
0!
0'
0/
#327950000000
1!
1'
1/
#327960000000
0!
0'
0/
#327970000000
1!
1'
1/
#327980000000
0!
0'
0/
#327990000000
1!
1'
1/
#328000000000
0!
0'
0/
#328010000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#328020000000
0!
0'
0/
#328030000000
1!
1'
1/
#328040000000
0!
0'
0/
#328050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#328060000000
0!
0'
0/
#328070000000
1!
1'
1/
#328080000000
0!
0'
0/
#328090000000
#328100000000
1!
1'
1/
#328110000000
0!
0'
0/
#328120000000
1!
1'
1/
#328130000000
0!
1"
0'
1(
0/
10
#328140000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#328150000000
0!
0'
0/
#328160000000
1!
1'
1/
#328170000000
0!
0'
0/
#328180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#328190000000
0!
0'
0/
#328200000000
1!
1'
1/
#328210000000
0!
1"
0'
1(
0/
10
#328220000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#328230000000
0!
1$
0'
1+
0/
#328240000000
1!
1'
1/
#328250000000
0!
0'
0/
#328260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#328270000000
0!
0'
0/
#328280000000
1!
1'
1/
#328290000000
0!
0'
0/
#328300000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#328310000000
0!
0'
0/
#328320000000
1!
1'
1/
#328330000000
0!
0'
0/
#328340000000
1!
1'
1/
#328350000000
0!
0'
0/
#328360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#328370000000
0!
0'
0/
#328380000000
1!
1'
1/
#328390000000
0!
0'
0/
#328400000000
1!
1'
1/
#328410000000
0!
0'
0/
#328420000000
1!
1'
1/
#328430000000
0!
0'
0/
#328440000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#328450000000
0!
0'
0/
#328460000000
1!
1'
1/
#328470000000
0!
0'
0/
#328480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#328490000000
0!
0'
0/
#328500000000
1!
1'
1/
#328510000000
0!
0'
0/
#328520000000
#328530000000
1!
1'
1/
#328540000000
0!
0'
0/
#328550000000
1!
1'
1/
#328560000000
0!
1"
0'
1(
0/
10
#328570000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#328580000000
0!
0'
0/
#328590000000
1!
1'
1/
#328600000000
0!
0'
0/
#328610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#328620000000
0!
0'
0/
#328630000000
1!
1'
1/
#328640000000
0!
1"
0'
1(
0/
10
#328650000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#328660000000
0!
1$
0'
1+
0/
#328670000000
1!
1'
1/
#328680000000
0!
0'
0/
#328690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#328700000000
0!
0'
0/
#328710000000
1!
1'
1/
#328720000000
0!
0'
0/
#328730000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#328740000000
0!
0'
0/
#328750000000
1!
1'
1/
#328760000000
0!
0'
0/
#328770000000
1!
1'
1/
#328780000000
0!
0'
0/
#328790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#328800000000
0!
0'
0/
#328810000000
1!
1'
1/
#328820000000
0!
0'
0/
#328830000000
1!
1'
1/
#328840000000
0!
0'
0/
#328850000000
1!
1'
1/
#328860000000
0!
0'
0/
#328870000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#328880000000
0!
0'
0/
#328890000000
1!
1'
1/
#328900000000
0!
0'
0/
#328910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#328920000000
0!
0'
0/
#328930000000
1!
1'
1/
#328940000000
0!
0'
0/
#328950000000
#328960000000
1!
1'
1/
#328970000000
0!
0'
0/
#328980000000
1!
1'
1/
#328990000000
0!
1"
0'
1(
0/
10
#329000000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#329010000000
0!
0'
0/
#329020000000
1!
1'
1/
#329030000000
0!
0'
0/
#329040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#329050000000
0!
0'
0/
#329060000000
1!
1'
1/
#329070000000
0!
1"
0'
1(
0/
10
#329080000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#329090000000
0!
1$
0'
1+
0/
#329100000000
1!
1'
1/
#329110000000
0!
0'
0/
#329120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#329130000000
0!
0'
0/
#329140000000
1!
1'
1/
#329150000000
0!
0'
0/
#329160000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#329170000000
0!
0'
0/
#329180000000
1!
1'
1/
#329190000000
0!
0'
0/
#329200000000
1!
1'
1/
#329210000000
0!
0'
0/
#329220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#329230000000
0!
0'
0/
#329240000000
1!
1'
1/
#329250000000
0!
0'
0/
#329260000000
1!
1'
1/
#329270000000
0!
0'
0/
#329280000000
1!
1'
1/
#329290000000
0!
0'
0/
#329300000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#329310000000
0!
0'
0/
#329320000000
1!
1'
1/
#329330000000
0!
0'
0/
#329340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#329350000000
0!
0'
0/
#329360000000
1!
1'
1/
#329370000000
0!
0'
0/
#329380000000
#329390000000
1!
1'
1/
#329400000000
0!
0'
0/
#329410000000
1!
1'
1/
#329420000000
0!
1"
0'
1(
0/
10
#329430000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#329440000000
0!
0'
0/
#329450000000
1!
1'
1/
#329460000000
0!
0'
0/
#329470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#329480000000
0!
0'
0/
#329490000000
1!
1'
1/
#329500000000
0!
1"
0'
1(
0/
10
#329510000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#329520000000
0!
1$
0'
1+
0/
#329530000000
1!
1'
1/
#329540000000
0!
0'
0/
#329550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#329560000000
0!
0'
0/
#329570000000
1!
1'
1/
#329580000000
0!
0'
0/
#329590000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#329600000000
0!
0'
0/
#329610000000
1!
1'
1/
#329620000000
0!
0'
0/
#329630000000
1!
1'
1/
#329640000000
0!
0'
0/
#329650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#329660000000
0!
0'
0/
#329670000000
1!
1'
1/
#329680000000
0!
0'
0/
#329690000000
1!
1'
1/
#329700000000
0!
0'
0/
#329710000000
1!
1'
1/
#329720000000
0!
0'
0/
#329730000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#329740000000
0!
0'
0/
#329750000000
1!
1'
1/
#329760000000
0!
0'
0/
#329770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#329780000000
0!
0'
0/
#329790000000
1!
1'
1/
#329800000000
0!
0'
0/
#329810000000
#329820000000
1!
1'
1/
#329830000000
0!
0'
0/
#329840000000
1!
1'
1/
#329850000000
0!
1"
0'
1(
0/
10
#329860000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#329870000000
0!
0'
0/
#329880000000
1!
1'
1/
#329890000000
0!
0'
0/
#329900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#329910000000
0!
0'
0/
#329920000000
1!
1'
1/
#329930000000
0!
1"
0'
1(
0/
10
#329940000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#329950000000
0!
1$
0'
1+
0/
#329960000000
1!
1'
1/
#329970000000
0!
0'
0/
#329980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#329990000000
0!
0'
0/
#330000000000
1!
1'
1/
#330010000000
0!
0'
0/
#330020000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#330030000000
0!
0'
0/
#330040000000
1!
1'
1/
#330050000000
0!
0'
0/
#330060000000
1!
1'
1/
#330070000000
0!
0'
0/
#330080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#330090000000
0!
0'
0/
#330100000000
1!
1'
1/
#330110000000
0!
0'
0/
#330120000000
1!
1'
1/
#330130000000
0!
0'
0/
#330140000000
1!
1'
1/
#330150000000
0!
0'
0/
#330160000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#330170000000
0!
0'
0/
#330180000000
1!
1'
1/
#330190000000
0!
0'
0/
#330200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#330210000000
0!
0'
0/
#330220000000
1!
1'
1/
#330230000000
0!
0'
0/
#330240000000
#330250000000
1!
1'
1/
#330260000000
0!
0'
0/
#330270000000
1!
1'
1/
#330280000000
0!
1"
0'
1(
0/
10
#330290000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#330300000000
0!
0'
0/
#330310000000
1!
1'
1/
#330320000000
0!
0'
0/
#330330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#330340000000
0!
0'
0/
#330350000000
1!
1'
1/
#330360000000
0!
1"
0'
1(
0/
10
#330370000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#330380000000
0!
1$
0'
1+
0/
#330390000000
1!
1'
1/
#330400000000
0!
0'
0/
#330410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#330420000000
0!
0'
0/
#330430000000
1!
1'
1/
#330440000000
0!
0'
0/
#330450000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#330460000000
0!
0'
0/
#330470000000
1!
1'
1/
#330480000000
0!
0'
0/
#330490000000
1!
1'
1/
#330500000000
0!
0'
0/
#330510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#330520000000
0!
0'
0/
#330530000000
1!
1'
1/
#330540000000
0!
0'
0/
#330550000000
1!
1'
1/
#330560000000
0!
0'
0/
#330570000000
1!
1'
1/
#330580000000
0!
0'
0/
#330590000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#330600000000
0!
0'
0/
#330610000000
1!
1'
1/
#330620000000
0!
0'
0/
#330630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#330640000000
0!
0'
0/
#330650000000
1!
1'
1/
#330660000000
0!
0'
0/
#330670000000
#330680000000
1!
1'
1/
#330690000000
0!
0'
0/
#330700000000
1!
1'
1/
#330710000000
0!
1"
0'
1(
0/
10
#330720000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#330730000000
0!
0'
0/
#330740000000
1!
1'
1/
#330750000000
0!
0'
0/
#330760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#330770000000
0!
0'
0/
#330780000000
1!
1'
1/
#330790000000
0!
1"
0'
1(
0/
10
#330800000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#330810000000
0!
1$
0'
1+
0/
#330820000000
1!
1'
1/
#330830000000
0!
0'
0/
#330840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#330850000000
0!
0'
0/
#330860000000
1!
1'
1/
#330870000000
0!
0'
0/
#330880000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#330890000000
0!
0'
0/
#330900000000
1!
1'
1/
#330910000000
0!
0'
0/
#330920000000
1!
1'
1/
#330930000000
0!
0'
0/
#330940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#330950000000
0!
0'
0/
#330960000000
1!
1'
1/
#330970000000
0!
0'
0/
#330980000000
1!
1'
1/
#330990000000
0!
0'
0/
#331000000000
1!
1'
1/
#331010000000
0!
0'
0/
#331020000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#331030000000
0!
0'
0/
#331040000000
1!
1'
1/
#331050000000
0!
0'
0/
#331060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#331070000000
0!
0'
0/
#331080000000
1!
1'
1/
#331090000000
0!
0'
0/
#331100000000
#331110000000
1!
1'
1/
#331120000000
0!
0'
0/
#331130000000
1!
1'
1/
#331140000000
0!
1"
0'
1(
0/
10
#331150000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#331160000000
0!
0'
0/
#331170000000
1!
1'
1/
#331180000000
0!
0'
0/
#331190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#331200000000
0!
0'
0/
#331210000000
1!
1'
1/
#331220000000
0!
1"
0'
1(
0/
10
#331230000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#331240000000
0!
1$
0'
1+
0/
#331250000000
1!
1'
1/
#331260000000
0!
0'
0/
#331270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#331280000000
0!
0'
0/
#331290000000
1!
1'
1/
#331300000000
0!
0'
0/
#331310000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#331320000000
0!
0'
0/
#331330000000
1!
1'
1/
#331340000000
0!
0'
0/
#331350000000
1!
1'
1/
#331360000000
0!
0'
0/
#331370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#331380000000
0!
0'
0/
#331390000000
1!
1'
1/
#331400000000
0!
0'
0/
#331410000000
1!
1'
1/
#331420000000
0!
0'
0/
#331430000000
1!
1'
1/
#331440000000
0!
0'
0/
#331450000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#331460000000
0!
0'
0/
#331470000000
1!
1'
1/
#331480000000
0!
0'
0/
#331490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#331500000000
0!
0'
0/
#331510000000
1!
1'
1/
#331520000000
0!
0'
0/
#331530000000
#331540000000
1!
1'
1/
#331550000000
0!
0'
0/
#331560000000
1!
1'
1/
#331570000000
0!
1"
0'
1(
0/
10
#331580000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#331590000000
0!
0'
0/
#331600000000
1!
1'
1/
#331610000000
0!
0'
0/
#331620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#331630000000
0!
0'
0/
#331640000000
1!
1'
1/
#331650000000
0!
1"
0'
1(
0/
10
#331660000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#331670000000
0!
1$
0'
1+
0/
#331680000000
1!
1'
1/
#331690000000
0!
0'
0/
#331700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#331710000000
0!
0'
0/
#331720000000
1!
1'
1/
#331730000000
0!
0'
0/
#331740000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#331750000000
0!
0'
0/
#331760000000
1!
1'
1/
#331770000000
0!
0'
0/
#331780000000
1!
1'
1/
#331790000000
0!
0'
0/
#331800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#331810000000
0!
0'
0/
#331820000000
1!
1'
1/
#331830000000
0!
0'
0/
#331840000000
1!
1'
1/
#331850000000
0!
0'
0/
#331860000000
1!
1'
1/
#331870000000
0!
0'
0/
#331880000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#331890000000
0!
0'
0/
#331900000000
1!
1'
1/
#331910000000
0!
0'
0/
#331920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#331930000000
0!
0'
0/
#331940000000
1!
1'
1/
#331950000000
0!
0'
0/
#331960000000
#331970000000
1!
1'
1/
#331980000000
0!
0'
0/
#331990000000
1!
1'
1/
#332000000000
0!
1"
0'
1(
0/
10
#332010000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#332020000000
0!
0'
0/
#332030000000
1!
1'
1/
#332040000000
0!
0'
0/
#332050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#332060000000
0!
0'
0/
#332070000000
1!
1'
1/
#332080000000
0!
1"
0'
1(
0/
10
#332090000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#332100000000
0!
1$
0'
1+
0/
#332110000000
1!
1'
1/
#332120000000
0!
0'
0/
#332130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#332140000000
0!
0'
0/
#332150000000
1!
1'
1/
#332160000000
0!
0'
0/
#332170000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#332180000000
0!
0'
0/
#332190000000
1!
1'
1/
#332200000000
0!
0'
0/
#332210000000
1!
1'
1/
#332220000000
0!
0'
0/
#332230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#332240000000
0!
0'
0/
#332250000000
1!
1'
1/
#332260000000
0!
0'
0/
#332270000000
1!
1'
1/
#332280000000
0!
0'
0/
#332290000000
1!
1'
1/
#332300000000
0!
0'
0/
#332310000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#332320000000
0!
0'
0/
#332330000000
1!
1'
1/
#332340000000
0!
0'
0/
#332350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#332360000000
0!
0'
0/
#332370000000
1!
1'
1/
#332380000000
0!
0'
0/
#332390000000
#332400000000
1!
1'
1/
#332410000000
0!
0'
0/
#332420000000
1!
1'
1/
#332430000000
0!
1"
0'
1(
0/
10
#332440000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#332450000000
0!
0'
0/
#332460000000
1!
1'
1/
#332470000000
0!
0'
0/
#332480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#332490000000
0!
0'
0/
#332500000000
1!
1'
1/
#332510000000
0!
1"
0'
1(
0/
10
#332520000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#332530000000
0!
1$
0'
1+
0/
#332540000000
1!
1'
1/
#332550000000
0!
0'
0/
#332560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#332570000000
0!
0'
0/
#332580000000
1!
1'
1/
#332590000000
0!
0'
0/
#332600000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#332610000000
0!
0'
0/
#332620000000
1!
1'
1/
#332630000000
0!
0'
0/
#332640000000
1!
1'
1/
#332650000000
0!
0'
0/
#332660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#332670000000
0!
0'
0/
#332680000000
1!
1'
1/
#332690000000
0!
0'
0/
#332700000000
1!
1'
1/
#332710000000
0!
0'
0/
#332720000000
1!
1'
1/
#332730000000
0!
0'
0/
#332740000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#332750000000
0!
0'
0/
#332760000000
1!
1'
1/
#332770000000
0!
0'
0/
#332780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#332790000000
0!
0'
0/
#332800000000
1!
1'
1/
#332810000000
0!
0'
0/
#332820000000
#332830000000
1!
1'
1/
#332840000000
0!
0'
0/
#332850000000
1!
1'
1/
#332860000000
0!
1"
0'
1(
0/
10
#332870000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#332880000000
0!
0'
0/
#332890000000
1!
1'
1/
#332900000000
0!
0'
0/
#332910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#332920000000
0!
0'
0/
#332930000000
1!
1'
1/
#332940000000
0!
1"
0'
1(
0/
10
#332950000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#332960000000
0!
1$
0'
1+
0/
#332970000000
1!
1'
1/
#332980000000
0!
0'
0/
#332990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#333000000000
0!
0'
0/
#333010000000
1!
1'
1/
#333020000000
0!
0'
0/
#333030000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#333040000000
0!
0'
0/
#333050000000
1!
1'
1/
#333060000000
0!
0'
0/
#333070000000
1!
1'
1/
#333080000000
0!
0'
0/
#333090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#333100000000
0!
0'
0/
#333110000000
1!
1'
1/
#333120000000
0!
0'
0/
#333130000000
1!
1'
1/
#333140000000
0!
0'
0/
#333150000000
1!
1'
1/
#333160000000
0!
0'
0/
#333170000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#333180000000
0!
0'
0/
#333190000000
1!
1'
1/
#333200000000
0!
0'
0/
#333210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#333220000000
0!
0'
0/
#333230000000
1!
1'
1/
#333240000000
0!
0'
0/
#333250000000
#333260000000
1!
1'
1/
#333270000000
0!
0'
0/
#333280000000
1!
1'
1/
#333290000000
0!
1"
0'
1(
0/
10
#333300000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#333310000000
0!
0'
0/
#333320000000
1!
1'
1/
#333330000000
0!
0'
0/
#333340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#333350000000
0!
0'
0/
#333360000000
1!
1'
1/
#333370000000
0!
1"
0'
1(
0/
10
#333380000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#333390000000
0!
1$
0'
1+
0/
#333400000000
1!
1'
1/
#333410000000
0!
0'
0/
#333420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#333430000000
0!
0'
0/
#333440000000
1!
1'
1/
#333450000000
0!
0'
0/
#333460000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#333470000000
0!
0'
0/
#333480000000
1!
1'
1/
#333490000000
0!
0'
0/
#333500000000
1!
1'
1/
#333510000000
0!
0'
0/
#333520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#333530000000
0!
0'
0/
#333540000000
1!
1'
1/
#333550000000
0!
0'
0/
#333560000000
1!
1'
1/
#333570000000
0!
0'
0/
#333580000000
1!
1'
1/
#333590000000
0!
0'
0/
#333600000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#333610000000
0!
0'
0/
#333620000000
1!
1'
1/
#333630000000
0!
0'
0/
#333640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#333650000000
0!
0'
0/
#333660000000
1!
1'
1/
#333670000000
0!
0'
0/
#333680000000
#333690000000
1!
1'
1/
#333700000000
0!
0'
0/
#333710000000
1!
1'
1/
#333720000000
0!
1"
0'
1(
0/
10
#333730000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#333740000000
0!
0'
0/
#333750000000
1!
1'
1/
#333760000000
0!
0'
0/
#333770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#333780000000
0!
0'
0/
#333790000000
1!
1'
1/
#333800000000
0!
1"
0'
1(
0/
10
#333810000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#333820000000
0!
1$
0'
1+
0/
#333830000000
1!
1'
1/
#333840000000
0!
0'
0/
#333850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#333860000000
0!
0'
0/
#333870000000
1!
1'
1/
#333880000000
0!
0'
0/
#333890000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#333900000000
0!
0'
0/
#333910000000
1!
1'
1/
#333920000000
0!
0'
0/
#333930000000
1!
1'
1/
#333940000000
0!
0'
0/
#333950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#333960000000
0!
0'
0/
#333970000000
1!
1'
1/
#333980000000
0!
0'
0/
#333990000000
1!
1'
1/
#334000000000
0!
0'
0/
#334010000000
1!
1'
1/
#334020000000
0!
0'
0/
#334030000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#334040000000
0!
0'
0/
#334050000000
1!
1'
1/
#334060000000
0!
0'
0/
#334070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#334080000000
0!
0'
0/
#334090000000
1!
1'
1/
#334100000000
0!
0'
0/
#334110000000
#334120000000
1!
1'
1/
#334130000000
0!
0'
0/
#334140000000
1!
1'
1/
#334150000000
0!
1"
0'
1(
0/
10
#334160000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#334170000000
0!
0'
0/
#334180000000
1!
1'
1/
#334190000000
0!
0'
0/
#334200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#334210000000
0!
0'
0/
#334220000000
1!
1'
1/
#334230000000
0!
1"
0'
1(
0/
10
#334240000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#334250000000
0!
1$
0'
1+
0/
#334260000000
1!
1'
1/
#334270000000
0!
0'
0/
#334280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#334290000000
0!
0'
0/
#334300000000
1!
1'
1/
#334310000000
0!
0'
0/
#334320000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#334330000000
0!
0'
0/
#334340000000
1!
1'
1/
#334350000000
0!
0'
0/
#334360000000
1!
1'
1/
#334370000000
0!
0'
0/
#334380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#334390000000
0!
0'
0/
#334400000000
1!
1'
1/
#334410000000
0!
0'
0/
#334420000000
1!
1'
1/
#334430000000
0!
0'
0/
#334440000000
1!
1'
1/
#334450000000
0!
0'
0/
#334460000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#334470000000
0!
0'
0/
#334480000000
1!
1'
1/
#334490000000
0!
0'
0/
#334500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#334510000000
0!
0'
0/
#334520000000
1!
1'
1/
#334530000000
0!
0'
0/
#334540000000
#334550000000
1!
1'
1/
#334560000000
0!
0'
0/
#334570000000
1!
1'
1/
#334580000000
0!
1"
0'
1(
0/
10
#334590000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#334600000000
0!
0'
0/
#334610000000
1!
1'
1/
#334620000000
0!
0'
0/
#334630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#334640000000
0!
0'
0/
#334650000000
1!
1'
1/
#334660000000
0!
1"
0'
1(
0/
10
#334670000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#334680000000
0!
1$
0'
1+
0/
#334690000000
1!
1'
1/
#334700000000
0!
0'
0/
#334710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#334720000000
0!
0'
0/
#334730000000
1!
1'
1/
#334740000000
0!
0'
0/
#334750000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#334760000000
0!
0'
0/
#334770000000
1!
1'
1/
#334780000000
0!
0'
0/
#334790000000
1!
1'
1/
#334800000000
0!
0'
0/
#334810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#334820000000
0!
0'
0/
#334830000000
1!
1'
1/
#334840000000
0!
0'
0/
#334850000000
1!
1'
1/
#334860000000
0!
0'
0/
#334870000000
1!
1'
1/
#334880000000
0!
0'
0/
#334890000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#334900000000
0!
0'
0/
#334910000000
1!
1'
1/
#334920000000
0!
0'
0/
#334930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#334940000000
0!
0'
0/
#334950000000
1!
1'
1/
#334960000000
0!
0'
0/
#334970000000
#334980000000
1!
1'
1/
#334990000000
0!
0'
0/
#335000000000
1!
1'
1/
#335010000000
0!
1"
0'
1(
0/
10
#335020000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#335030000000
0!
0'
0/
#335040000000
1!
1'
1/
#335050000000
0!
0'
0/
#335060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#335070000000
0!
0'
0/
#335080000000
1!
1'
1/
#335090000000
0!
1"
0'
1(
0/
10
#335100000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#335110000000
0!
1$
0'
1+
0/
#335120000000
1!
1'
1/
#335130000000
0!
0'
0/
#335140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#335150000000
0!
0'
0/
#335160000000
1!
1'
1/
#335170000000
0!
0'
0/
#335180000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#335190000000
0!
0'
0/
#335200000000
1!
1'
1/
#335210000000
0!
0'
0/
#335220000000
1!
1'
1/
#335230000000
0!
0'
0/
#335240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#335250000000
0!
0'
0/
#335260000000
1!
1'
1/
#335270000000
0!
0'
0/
#335280000000
1!
1'
1/
#335290000000
0!
0'
0/
#335300000000
1!
1'
1/
#335310000000
0!
0'
0/
#335320000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#335330000000
0!
0'
0/
#335340000000
1!
1'
1/
#335350000000
0!
0'
0/
#335360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#335370000000
0!
0'
0/
#335380000000
1!
1'
1/
#335390000000
0!
0'
0/
#335400000000
#335410000000
1!
1'
1/
#335420000000
0!
0'
0/
#335430000000
1!
1'
1/
#335440000000
0!
1"
0'
1(
0/
10
#335450000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#335460000000
0!
0'
0/
#335470000000
1!
1'
1/
#335480000000
0!
0'
0/
#335490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#335500000000
0!
0'
0/
#335510000000
1!
1'
1/
#335520000000
0!
1"
0'
1(
0/
10
#335530000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#335540000000
0!
1$
0'
1+
0/
#335550000000
1!
1'
1/
#335560000000
0!
0'
0/
#335570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#335580000000
0!
0'
0/
#335590000000
1!
1'
1/
#335600000000
0!
0'
0/
#335610000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#335620000000
0!
0'
0/
#335630000000
1!
1'
1/
#335640000000
0!
0'
0/
#335650000000
1!
1'
1/
#335660000000
0!
0'
0/
#335670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#335680000000
0!
0'
0/
#335690000000
1!
1'
1/
#335700000000
0!
0'
0/
#335710000000
1!
1'
1/
#335720000000
0!
0'
0/
#335730000000
1!
1'
1/
#335740000000
0!
0'
0/
#335750000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#335760000000
0!
0'
0/
#335770000000
1!
1'
1/
#335780000000
0!
0'
0/
#335790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#335800000000
0!
0'
0/
#335810000000
1!
1'
1/
#335820000000
0!
0'
0/
#335830000000
#335840000000
1!
1'
1/
#335850000000
0!
0'
0/
#335860000000
1!
1'
1/
#335870000000
0!
1"
0'
1(
0/
10
#335880000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#335890000000
0!
0'
0/
#335900000000
1!
1'
1/
#335910000000
0!
0'
0/
#335920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#335930000000
0!
0'
0/
#335940000000
1!
1'
1/
#335950000000
0!
1"
0'
1(
0/
10
#335960000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#335970000000
0!
1$
0'
1+
0/
#335980000000
1!
1'
1/
#335990000000
0!
0'
0/
#336000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#336010000000
0!
0'
0/
#336020000000
1!
1'
1/
#336030000000
0!
0'
0/
#336040000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#336050000000
0!
0'
0/
#336060000000
1!
1'
1/
#336070000000
0!
0'
0/
#336080000000
1!
1'
1/
#336090000000
0!
0'
0/
#336100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#336110000000
0!
0'
0/
#336120000000
1!
1'
1/
#336130000000
0!
0'
0/
#336140000000
1!
1'
1/
#336150000000
0!
0'
0/
#336160000000
1!
1'
1/
#336170000000
0!
0'
0/
#336180000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#336190000000
0!
0'
0/
#336200000000
1!
1'
1/
#336210000000
0!
0'
0/
#336220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#336230000000
0!
0'
0/
#336240000000
1!
1'
1/
#336250000000
0!
0'
0/
#336260000000
#336270000000
1!
1'
1/
#336280000000
0!
0'
0/
#336290000000
1!
1'
1/
#336300000000
0!
1"
0'
1(
0/
10
#336310000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#336320000000
0!
0'
0/
#336330000000
1!
1'
1/
#336340000000
0!
0'
0/
#336350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#336360000000
0!
0'
0/
#336370000000
1!
1'
1/
#336380000000
0!
1"
0'
1(
0/
10
#336390000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#336400000000
0!
1$
0'
1+
0/
#336410000000
1!
1'
1/
#336420000000
0!
0'
0/
#336430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#336440000000
0!
0'
0/
#336450000000
1!
1'
1/
#336460000000
0!
0'
0/
#336470000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#336480000000
0!
0'
0/
#336490000000
1!
1'
1/
#336500000000
0!
0'
0/
#336510000000
1!
1'
1/
#336520000000
0!
0'
0/
#336530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#336540000000
0!
0'
0/
#336550000000
1!
1'
1/
#336560000000
0!
0'
0/
#336570000000
1!
1'
1/
#336580000000
0!
0'
0/
#336590000000
1!
1'
1/
#336600000000
0!
0'
0/
#336610000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#336620000000
0!
0'
0/
#336630000000
1!
1'
1/
#336640000000
0!
0'
0/
#336650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#336660000000
0!
0'
0/
#336670000000
1!
1'
1/
#336680000000
0!
0'
0/
#336690000000
#336700000000
1!
1'
1/
#336710000000
0!
0'
0/
#336720000000
1!
1'
1/
#336730000000
0!
1"
0'
1(
0/
10
#336740000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#336750000000
0!
0'
0/
#336760000000
1!
1'
1/
#336770000000
0!
0'
0/
#336780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#336790000000
0!
0'
0/
#336800000000
1!
1'
1/
#336810000000
0!
1"
0'
1(
0/
10
#336820000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#336830000000
0!
1$
0'
1+
0/
#336840000000
1!
1'
1/
#336850000000
0!
0'
0/
#336860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#336870000000
0!
0'
0/
#336880000000
1!
1'
1/
#336890000000
0!
0'
0/
#336900000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#336910000000
0!
0'
0/
#336920000000
1!
1'
1/
#336930000000
0!
0'
0/
#336940000000
1!
1'
1/
#336950000000
0!
0'
0/
#336960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#336970000000
0!
0'
0/
#336980000000
1!
1'
1/
#336990000000
0!
0'
0/
#337000000000
1!
1'
1/
#337010000000
0!
0'
0/
#337020000000
1!
1'
1/
#337030000000
0!
0'
0/
#337040000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#337050000000
0!
0'
0/
#337060000000
1!
1'
1/
#337070000000
0!
0'
0/
#337080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#337090000000
0!
0'
0/
#337100000000
1!
1'
1/
#337110000000
0!
0'
0/
#337120000000
#337130000000
1!
1'
1/
#337140000000
0!
0'
0/
#337150000000
1!
1'
1/
#337160000000
0!
1"
0'
1(
0/
10
#337170000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#337180000000
0!
0'
0/
#337190000000
1!
1'
1/
#337200000000
0!
0'
0/
#337210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#337220000000
0!
0'
0/
#337230000000
1!
1'
1/
#337240000000
0!
1"
0'
1(
0/
10
#337250000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#337260000000
0!
1$
0'
1+
0/
#337270000000
1!
1'
1/
#337280000000
0!
0'
0/
#337290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#337300000000
0!
0'
0/
#337310000000
1!
1'
1/
#337320000000
0!
0'
0/
#337330000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#337340000000
0!
0'
0/
#337350000000
1!
1'
1/
#337360000000
0!
0'
0/
#337370000000
1!
1'
1/
#337380000000
0!
0'
0/
#337390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#337400000000
0!
0'
0/
#337410000000
1!
1'
1/
#337420000000
0!
0'
0/
#337430000000
1!
1'
1/
#337440000000
0!
0'
0/
#337450000000
1!
1'
1/
#337460000000
0!
0'
0/
#337470000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#337480000000
0!
0'
0/
#337490000000
1!
1'
1/
#337500000000
0!
0'
0/
#337510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#337520000000
0!
0'
0/
#337530000000
1!
1'
1/
#337540000000
0!
0'
0/
#337550000000
#337560000000
1!
1'
1/
#337570000000
0!
0'
0/
#337580000000
1!
1'
1/
#337590000000
0!
1"
0'
1(
0/
10
#337600000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#337610000000
0!
0'
0/
#337620000000
1!
1'
1/
#337630000000
0!
0'
0/
#337640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#337650000000
0!
0'
0/
#337660000000
1!
1'
1/
#337670000000
0!
1"
0'
1(
0/
10
#337680000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#337690000000
0!
1$
0'
1+
0/
#337700000000
1!
1'
1/
#337710000000
0!
0'
0/
#337720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#337730000000
0!
0'
0/
#337740000000
1!
1'
1/
#337750000000
0!
0'
0/
#337760000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#337770000000
0!
0'
0/
#337780000000
1!
1'
1/
#337790000000
0!
0'
0/
#337800000000
1!
1'
1/
#337810000000
0!
0'
0/
#337820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#337830000000
0!
0'
0/
#337840000000
1!
1'
1/
#337850000000
0!
0'
0/
#337860000000
1!
1'
1/
#337870000000
0!
0'
0/
#337880000000
1!
1'
1/
#337890000000
0!
0'
0/
#337900000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#337910000000
0!
0'
0/
#337920000000
1!
1'
1/
#337930000000
0!
0'
0/
#337940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#337950000000
0!
0'
0/
#337960000000
1!
1'
1/
#337970000000
0!
0'
0/
#337980000000
#337990000000
1!
1'
1/
#338000000000
0!
0'
0/
#338010000000
1!
1'
1/
#338020000000
0!
1"
0'
1(
0/
10
#338030000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#338040000000
0!
0'
0/
#338050000000
1!
1'
1/
#338060000000
0!
0'
0/
#338070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#338080000000
0!
0'
0/
#338090000000
1!
1'
1/
#338100000000
0!
1"
0'
1(
0/
10
#338110000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#338120000000
0!
1$
0'
1+
0/
#338130000000
1!
1'
1/
#338140000000
0!
0'
0/
#338150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#338160000000
0!
0'
0/
#338170000000
1!
1'
1/
#338180000000
0!
0'
0/
#338190000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#338200000000
0!
0'
0/
#338210000000
1!
1'
1/
#338220000000
0!
0'
0/
#338230000000
1!
1'
1/
#338240000000
0!
0'
0/
#338250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#338260000000
0!
0'
0/
#338270000000
1!
1'
1/
#338280000000
0!
0'
0/
#338290000000
1!
1'
1/
#338300000000
0!
0'
0/
#338310000000
1!
1'
1/
#338320000000
0!
0'
0/
#338330000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#338340000000
0!
0'
0/
#338350000000
1!
1'
1/
#338360000000
0!
0'
0/
#338370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#338380000000
0!
0'
0/
#338390000000
1!
1'
1/
#338400000000
0!
0'
0/
#338410000000
#338420000000
1!
1'
1/
#338430000000
0!
0'
0/
#338440000000
1!
1'
1/
#338450000000
0!
1"
0'
1(
0/
10
#338460000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#338470000000
0!
0'
0/
#338480000000
1!
1'
1/
#338490000000
0!
0'
0/
#338500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#338510000000
0!
0'
0/
#338520000000
1!
1'
1/
#338530000000
0!
1"
0'
1(
0/
10
#338540000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#338550000000
0!
1$
0'
1+
0/
#338560000000
1!
1'
1/
#338570000000
0!
0'
0/
#338580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#338590000000
0!
0'
0/
#338600000000
1!
1'
1/
#338610000000
0!
0'
0/
#338620000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#338630000000
0!
0'
0/
#338640000000
1!
1'
1/
#338650000000
0!
0'
0/
#338660000000
1!
1'
1/
#338670000000
0!
0'
0/
#338680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#338690000000
0!
0'
0/
#338700000000
1!
1'
1/
#338710000000
0!
0'
0/
#338720000000
1!
1'
1/
#338730000000
0!
0'
0/
#338740000000
1!
1'
1/
#338750000000
0!
0'
0/
#338760000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#338770000000
0!
0'
0/
#338780000000
1!
1'
1/
#338790000000
0!
0'
0/
#338800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#338810000000
0!
0'
0/
#338820000000
1!
1'
1/
#338830000000
0!
0'
0/
#338840000000
#338850000000
1!
1'
1/
#338860000000
0!
0'
0/
#338870000000
1!
1'
1/
#338880000000
0!
1"
0'
1(
0/
10
#338890000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#338900000000
0!
0'
0/
#338910000000
1!
1'
1/
#338920000000
0!
0'
0/
#338930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#338940000000
0!
0'
0/
#338950000000
1!
1'
1/
#338960000000
0!
1"
0'
1(
0/
10
#338970000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#338980000000
0!
1$
0'
1+
0/
#338990000000
1!
1'
1/
#339000000000
0!
0'
0/
#339010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#339020000000
0!
0'
0/
#339030000000
1!
1'
1/
#339040000000
0!
0'
0/
#339050000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#339060000000
0!
0'
0/
#339070000000
1!
1'
1/
#339080000000
0!
0'
0/
#339090000000
1!
1'
1/
#339100000000
0!
0'
0/
#339110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#339120000000
0!
0'
0/
#339130000000
1!
1'
1/
#339140000000
0!
0'
0/
#339150000000
1!
1'
1/
#339160000000
0!
0'
0/
#339170000000
1!
1'
1/
#339180000000
0!
0'
0/
#339190000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#339200000000
0!
0'
0/
#339210000000
1!
1'
1/
#339220000000
0!
0'
0/
#339230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#339240000000
0!
0'
0/
#339250000000
1!
1'
1/
#339260000000
0!
0'
0/
#339270000000
#339280000000
1!
1'
1/
#339290000000
0!
0'
0/
#339300000000
1!
1'
1/
#339310000000
0!
1"
0'
1(
0/
10
#339320000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#339330000000
0!
0'
0/
#339340000000
1!
1'
1/
#339350000000
0!
0'
0/
#339360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#339370000000
0!
0'
0/
#339380000000
1!
1'
1/
#339390000000
0!
1"
0'
1(
0/
10
#339400000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#339410000000
0!
1$
0'
1+
0/
#339420000000
1!
1'
1/
#339430000000
0!
0'
0/
#339440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#339450000000
0!
0'
0/
#339460000000
1!
1'
1/
#339470000000
0!
0'
0/
#339480000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#339490000000
0!
0'
0/
#339500000000
1!
1'
1/
#339510000000
0!
0'
0/
#339520000000
1!
1'
1/
#339530000000
0!
0'
0/
#339540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#339550000000
0!
0'
0/
#339560000000
1!
1'
1/
#339570000000
0!
0'
0/
#339580000000
1!
1'
1/
#339590000000
0!
0'
0/
#339600000000
1!
1'
1/
#339610000000
0!
0'
0/
#339620000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#339630000000
0!
0'
0/
#339640000000
1!
1'
1/
#339650000000
0!
0'
0/
#339660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#339670000000
0!
0'
0/
#339680000000
1!
1'
1/
#339690000000
0!
0'
0/
#339700000000
#339710000000
1!
1'
1/
#339720000000
0!
0'
0/
#339730000000
1!
1'
1/
#339740000000
0!
1"
0'
1(
0/
10
#339750000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#339760000000
0!
0'
0/
#339770000000
1!
1'
1/
#339780000000
0!
0'
0/
#339790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#339800000000
0!
0'
0/
#339810000000
1!
1'
1/
#339820000000
0!
1"
0'
1(
0/
10
#339830000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#339840000000
0!
1$
0'
1+
0/
#339850000000
1!
1'
1/
#339860000000
0!
0'
0/
#339870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#339880000000
0!
0'
0/
#339890000000
1!
1'
1/
#339900000000
0!
0'
0/
#339910000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#339920000000
0!
0'
0/
#339930000000
1!
1'
1/
#339940000000
0!
0'
0/
#339950000000
1!
1'
1/
#339960000000
0!
0'
0/
#339970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#339980000000
0!
0'
0/
#339990000000
1!
1'
1/
#340000000000
0!
0'
0/
#340010000000
1!
1'
1/
#340020000000
0!
0'
0/
#340030000000
1!
1'
1/
#340040000000
0!
0'
0/
#340050000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#340060000000
0!
0'
0/
#340070000000
1!
1'
1/
#340080000000
0!
0'
0/
#340090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#340100000000
0!
0'
0/
#340110000000
1!
1'
1/
#340120000000
0!
0'
0/
#340130000000
#340140000000
1!
1'
1/
#340150000000
0!
0'
0/
#340160000000
1!
1'
1/
#340170000000
0!
1"
0'
1(
0/
10
#340180000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#340190000000
0!
0'
0/
#340200000000
1!
1'
1/
#340210000000
0!
0'
0/
#340220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#340230000000
0!
0'
0/
#340240000000
1!
1'
1/
#340250000000
0!
1"
0'
1(
0/
10
#340260000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#340270000000
0!
1$
0'
1+
0/
#340280000000
1!
1'
1/
#340290000000
0!
0'
0/
#340300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#340310000000
0!
0'
0/
#340320000000
1!
1'
1/
#340330000000
0!
0'
0/
#340340000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#340350000000
0!
0'
0/
#340360000000
1!
1'
1/
#340370000000
0!
0'
0/
#340380000000
1!
1'
1/
#340390000000
0!
0'
0/
#340400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#340410000000
0!
0'
0/
#340420000000
1!
1'
1/
#340430000000
0!
0'
0/
#340440000000
1!
1'
1/
#340450000000
0!
0'
0/
#340460000000
1!
1'
1/
#340470000000
0!
0'
0/
#340480000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#340490000000
0!
0'
0/
#340500000000
1!
1'
1/
#340510000000
0!
0'
0/
#340520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#340530000000
0!
0'
0/
#340540000000
1!
1'
1/
#340550000000
0!
0'
0/
#340560000000
#340570000000
1!
1'
1/
#340580000000
0!
0'
0/
#340590000000
1!
1'
1/
#340600000000
0!
1"
0'
1(
0/
10
#340610000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#340620000000
0!
0'
0/
#340630000000
1!
1'
1/
#340640000000
0!
0'
0/
#340650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#340660000000
0!
0'
0/
#340670000000
1!
1'
1/
#340680000000
0!
1"
0'
1(
0/
10
#340690000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#340700000000
0!
1$
0'
1+
0/
#340710000000
1!
1'
1/
#340720000000
0!
0'
0/
#340730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#340740000000
0!
0'
0/
#340750000000
1!
1'
1/
#340760000000
0!
0'
0/
#340770000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#340780000000
0!
0'
0/
#340790000000
1!
1'
1/
#340800000000
0!
0'
0/
#340810000000
1!
1'
1/
#340820000000
0!
0'
0/
#340830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#340840000000
0!
0'
0/
#340850000000
1!
1'
1/
#340860000000
0!
0'
0/
#340870000000
1!
1'
1/
#340880000000
0!
0'
0/
#340890000000
1!
1'
1/
#340900000000
0!
0'
0/
#340910000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#340920000000
0!
0'
0/
#340930000000
1!
1'
1/
#340940000000
0!
0'
0/
#340950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#340960000000
0!
0'
0/
#340970000000
1!
1'
1/
#340980000000
0!
0'
0/
#340990000000
#341000000000
1!
1'
1/
#341010000000
0!
0'
0/
#341020000000
1!
1'
1/
#341030000000
0!
1"
0'
1(
0/
10
#341040000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#341050000000
0!
0'
0/
#341060000000
1!
1'
1/
#341070000000
0!
0'
0/
#341080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#341090000000
0!
0'
0/
#341100000000
1!
1'
1/
#341110000000
0!
1"
0'
1(
0/
10
#341120000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#341130000000
0!
1$
0'
1+
0/
#341140000000
1!
1'
1/
#341150000000
0!
0'
0/
#341160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#341170000000
0!
0'
0/
#341180000000
1!
1'
1/
#341190000000
0!
0'
0/
#341200000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#341210000000
0!
0'
0/
#341220000000
1!
1'
1/
#341230000000
0!
0'
0/
#341240000000
1!
1'
1/
#341250000000
0!
0'
0/
#341260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#341270000000
0!
0'
0/
#341280000000
1!
1'
1/
#341290000000
0!
0'
0/
#341300000000
1!
1'
1/
#341310000000
0!
0'
0/
#341320000000
1!
1'
1/
#341330000000
0!
0'
0/
#341340000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#341350000000
0!
0'
0/
#341360000000
1!
1'
1/
#341370000000
0!
0'
0/
#341380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#341390000000
0!
0'
0/
#341400000000
1!
1'
1/
#341410000000
0!
0'
0/
#341420000000
#341430000000
1!
1'
1/
#341440000000
0!
0'
0/
#341450000000
1!
1'
1/
#341460000000
0!
1"
0'
1(
0/
10
#341470000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#341480000000
0!
0'
0/
#341490000000
1!
1'
1/
#341500000000
0!
0'
0/
#341510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#341520000000
0!
0'
0/
#341530000000
1!
1'
1/
#341540000000
0!
1"
0'
1(
0/
10
#341550000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#341560000000
0!
1$
0'
1+
0/
#341570000000
1!
1'
1/
#341580000000
0!
0'
0/
#341590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#341600000000
0!
0'
0/
#341610000000
1!
1'
1/
#341620000000
0!
0'
0/
#341630000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#341640000000
0!
0'
0/
#341650000000
1!
1'
1/
#341660000000
0!
0'
0/
#341670000000
1!
1'
1/
#341680000000
0!
0'
0/
#341690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#341700000000
0!
0'
0/
#341710000000
1!
1'
1/
#341720000000
0!
0'
0/
#341730000000
1!
1'
1/
#341740000000
0!
0'
0/
#341750000000
1!
1'
1/
#341760000000
0!
0'
0/
#341770000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#341780000000
0!
0'
0/
#341790000000
1!
1'
1/
#341800000000
0!
0'
0/
#341810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#341820000000
0!
0'
0/
#341830000000
1!
1'
1/
#341840000000
0!
0'
0/
#341850000000
#341860000000
1!
1'
1/
#341870000000
0!
0'
0/
#341880000000
1!
1'
1/
#341890000000
0!
1"
0'
1(
0/
10
#341900000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#341910000000
0!
0'
0/
#341920000000
1!
1'
1/
#341930000000
0!
0'
0/
#341940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#341950000000
0!
0'
0/
#341960000000
1!
1'
1/
#341970000000
0!
1"
0'
1(
0/
10
#341980000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#341990000000
0!
1$
0'
1+
0/
#342000000000
1!
1'
1/
#342010000000
0!
0'
0/
#342020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#342030000000
0!
0'
0/
#342040000000
1!
1'
1/
#342050000000
0!
0'
0/
#342060000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#342070000000
0!
0'
0/
#342080000000
1!
1'
1/
#342090000000
0!
0'
0/
#342100000000
1!
1'
1/
#342110000000
0!
0'
0/
#342120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#342130000000
0!
0'
0/
#342140000000
1!
1'
1/
#342150000000
0!
0'
0/
#342160000000
1!
1'
1/
#342170000000
0!
0'
0/
#342180000000
1!
1'
1/
#342190000000
0!
0'
0/
#342200000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#342210000000
0!
0'
0/
#342220000000
1!
1'
1/
#342230000000
0!
0'
0/
#342240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#342250000000
0!
0'
0/
#342260000000
1!
1'
1/
#342270000000
0!
0'
0/
#342280000000
#342290000000
1!
1'
1/
#342300000000
0!
0'
0/
#342310000000
1!
1'
1/
#342320000000
0!
1"
0'
1(
0/
10
#342330000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#342340000000
0!
0'
0/
#342350000000
1!
1'
1/
#342360000000
0!
0'
0/
#342370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#342380000000
0!
0'
0/
#342390000000
1!
1'
1/
#342400000000
0!
1"
0'
1(
0/
10
#342410000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#342420000000
0!
1$
0'
1+
0/
#342430000000
1!
1'
1/
#342440000000
0!
0'
0/
#342450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#342460000000
0!
0'
0/
#342470000000
1!
1'
1/
#342480000000
0!
0'
0/
#342490000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#342500000000
0!
0'
0/
#342510000000
1!
1'
1/
#342520000000
0!
0'
0/
#342530000000
1!
1'
1/
#342540000000
0!
0'
0/
#342550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#342560000000
0!
0'
0/
#342570000000
1!
1'
1/
#342580000000
0!
0'
0/
#342590000000
1!
1'
1/
#342600000000
0!
0'
0/
#342610000000
1!
1'
1/
#342620000000
0!
0'
0/
#342630000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#342640000000
0!
0'
0/
#342650000000
1!
1'
1/
#342660000000
0!
0'
0/
#342670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#342680000000
0!
0'
0/
#342690000000
1!
1'
1/
#342700000000
0!
0'
0/
#342710000000
#342720000000
1!
1'
1/
#342730000000
0!
0'
0/
#342740000000
1!
1'
1/
#342750000000
0!
1"
0'
1(
0/
10
#342760000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#342770000000
0!
0'
0/
#342780000000
1!
1'
1/
#342790000000
0!
0'
0/
#342800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#342810000000
0!
0'
0/
#342820000000
1!
1'
1/
#342830000000
0!
1"
0'
1(
0/
10
#342840000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#342850000000
0!
1$
0'
1+
0/
#342860000000
1!
1'
1/
#342870000000
0!
0'
0/
#342880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#342890000000
0!
0'
0/
#342900000000
1!
1'
1/
#342910000000
0!
0'
0/
#342920000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#342930000000
0!
0'
0/
#342940000000
1!
1'
1/
#342950000000
0!
0'
0/
#342960000000
1!
1'
1/
#342970000000
0!
0'
0/
#342980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#342990000000
0!
0'
0/
#343000000000
1!
1'
1/
#343010000000
0!
0'
0/
#343020000000
1!
1'
1/
#343030000000
0!
0'
0/
#343040000000
1!
1'
1/
#343050000000
0!
0'
0/
#343060000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#343070000000
0!
0'
0/
#343080000000
1!
1'
1/
#343090000000
0!
0'
0/
#343100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#343110000000
0!
0'
0/
#343120000000
1!
1'
1/
#343130000000
0!
0'
0/
#343140000000
#343150000000
1!
1'
1/
#343160000000
0!
0'
0/
#343170000000
1!
1'
1/
#343180000000
0!
1"
0'
1(
0/
10
#343190000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#343200000000
0!
0'
0/
#343210000000
1!
1'
1/
#343220000000
0!
0'
0/
#343230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#343240000000
0!
0'
0/
#343250000000
1!
1'
1/
#343260000000
0!
1"
0'
1(
0/
10
#343270000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#343280000000
0!
1$
0'
1+
0/
#343290000000
1!
1'
1/
#343300000000
0!
0'
0/
#343310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#343320000000
0!
0'
0/
#343330000000
1!
1'
1/
#343340000000
0!
0'
0/
#343350000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#343360000000
0!
0'
0/
#343370000000
1!
1'
1/
#343380000000
0!
0'
0/
#343390000000
1!
1'
1/
#343400000000
0!
0'
0/
#343410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#343420000000
0!
0'
0/
#343430000000
1!
1'
1/
#343440000000
0!
0'
0/
#343450000000
1!
1'
1/
#343460000000
0!
0'
0/
#343470000000
1!
1'
1/
#343480000000
0!
0'
0/
#343490000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#343500000000
0!
0'
0/
#343510000000
1!
1'
1/
#343520000000
0!
0'
0/
#343530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#343540000000
0!
0'
0/
#343550000000
1!
1'
1/
#343560000000
0!
0'
0/
#343570000000
#343580000000
1!
1'
1/
#343590000000
0!
0'
0/
#343600000000
1!
1'
1/
#343610000000
0!
1"
0'
1(
0/
10
#343620000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#343630000000
0!
0'
0/
#343640000000
1!
1'
1/
#343650000000
0!
0'
0/
#343660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#343670000000
0!
0'
0/
#343680000000
1!
1'
1/
#343690000000
0!
1"
0'
1(
0/
10
#343700000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#343710000000
0!
1$
0'
1+
0/
#343720000000
1!
1'
1/
#343730000000
0!
0'
0/
#343740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#343750000000
0!
0'
0/
#343760000000
1!
1'
1/
#343770000000
0!
0'
0/
#343780000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#343790000000
0!
0'
0/
#343800000000
1!
1'
1/
#343810000000
0!
0'
0/
#343820000000
1!
1'
1/
#343830000000
0!
0'
0/
#343840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#343850000000
0!
0'
0/
#343860000000
1!
1'
1/
#343870000000
0!
0'
0/
#343880000000
1!
1'
1/
#343890000000
0!
0'
0/
#343900000000
1!
1'
1/
#343910000000
0!
0'
0/
#343920000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#343930000000
0!
0'
0/
#343940000000
1!
1'
1/
#343950000000
0!
0'
0/
#343960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#343970000000
0!
0'
0/
#343980000000
1!
1'
1/
#343990000000
0!
0'
0/
#344000000000
#344010000000
1!
1'
1/
#344020000000
0!
0'
0/
#344030000000
1!
1'
1/
#344040000000
0!
1"
0'
1(
0/
10
#344050000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#344060000000
0!
0'
0/
#344070000000
1!
1'
1/
#344080000000
0!
0'
0/
#344090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#344100000000
0!
0'
0/
#344110000000
1!
1'
1/
#344120000000
0!
1"
0'
1(
0/
10
#344130000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#344140000000
0!
1$
0'
1+
0/
#344150000000
1!
1'
1/
#344160000000
0!
0'
0/
#344170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#344180000000
0!
0'
0/
#344190000000
1!
1'
1/
#344200000000
0!
0'
0/
#344210000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#344220000000
0!
0'
0/
#344230000000
1!
1'
1/
#344240000000
0!
0'
0/
#344250000000
1!
1'
1/
#344260000000
0!
0'
0/
#344270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#344280000000
0!
0'
0/
#344290000000
1!
1'
1/
#344300000000
0!
0'
0/
#344310000000
1!
1'
1/
#344320000000
0!
0'
0/
#344330000000
1!
1'
1/
#344340000000
0!
0'
0/
#344350000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#344360000000
0!
0'
0/
#344370000000
1!
1'
1/
#344380000000
0!
0'
0/
#344390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#344400000000
0!
0'
0/
#344410000000
1!
1'
1/
#344420000000
0!
0'
0/
#344430000000
#344440000000
1!
1'
1/
#344450000000
0!
0'
0/
#344460000000
1!
1'
1/
#344470000000
0!
1"
0'
1(
0/
10
#344480000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#344490000000
0!
0'
0/
#344500000000
1!
1'
1/
#344510000000
0!
0'
0/
#344520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#344530000000
0!
0'
0/
#344540000000
1!
1'
1/
#344550000000
0!
1"
0'
1(
0/
10
#344560000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#344570000000
0!
1$
0'
1+
0/
#344580000000
1!
1'
1/
#344590000000
0!
0'
0/
#344600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#344610000000
0!
0'
0/
#344620000000
1!
1'
1/
#344630000000
0!
0'
0/
#344640000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#344650000000
0!
0'
0/
#344660000000
1!
1'
1/
#344670000000
0!
0'
0/
#344680000000
1!
1'
1/
#344690000000
0!
0'
0/
#344700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#344710000000
0!
0'
0/
#344720000000
1!
1'
1/
#344730000000
0!
0'
0/
#344740000000
1!
1'
1/
#344750000000
0!
0'
0/
#344760000000
1!
1'
1/
#344770000000
0!
0'
0/
#344780000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#344790000000
0!
0'
0/
#344800000000
1!
1'
1/
#344810000000
0!
0'
0/
#344820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#344830000000
0!
0'
0/
#344840000000
1!
1'
1/
#344850000000
0!
0'
0/
#344860000000
#344870000000
1!
1'
1/
#344880000000
0!
0'
0/
#344890000000
1!
1'
1/
#344900000000
0!
1"
0'
1(
0/
10
#344910000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#344920000000
0!
0'
0/
#344930000000
1!
1'
1/
#344940000000
0!
0'
0/
#344950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#344960000000
0!
0'
0/
#344970000000
1!
1'
1/
#344980000000
0!
1"
0'
1(
0/
10
#344990000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#345000000000
0!
1$
0'
1+
0/
#345010000000
1!
1'
1/
#345020000000
0!
0'
0/
#345030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#345040000000
0!
0'
0/
#345050000000
1!
1'
1/
#345060000000
0!
0'
0/
#345070000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#345080000000
0!
0'
0/
#345090000000
1!
1'
1/
#345100000000
0!
0'
0/
#345110000000
1!
1'
1/
#345120000000
0!
0'
0/
#345130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#345140000000
0!
0'
0/
#345150000000
1!
1'
1/
#345160000000
0!
0'
0/
#345170000000
1!
1'
1/
#345180000000
0!
0'
0/
#345190000000
1!
1'
1/
#345200000000
0!
0'
0/
#345210000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#345220000000
0!
0'
0/
#345230000000
1!
1'
1/
#345240000000
0!
0'
0/
#345250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#345260000000
0!
0'
0/
#345270000000
1!
1'
1/
#345280000000
0!
0'
0/
#345290000000
#345300000000
1!
1'
1/
#345310000000
0!
0'
0/
#345320000000
1!
1'
1/
#345330000000
0!
1"
0'
1(
0/
10
#345340000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#345350000000
0!
0'
0/
#345360000000
1!
1'
1/
#345370000000
0!
0'
0/
#345380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#345390000000
0!
0'
0/
#345400000000
1!
1'
1/
#345410000000
0!
1"
0'
1(
0/
10
#345420000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#345430000000
0!
1$
0'
1+
0/
#345440000000
1!
1'
1/
#345450000000
0!
0'
0/
#345460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#345470000000
0!
0'
0/
#345480000000
1!
1'
1/
#345490000000
0!
0'
0/
#345500000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#345510000000
0!
0'
0/
#345520000000
1!
1'
1/
#345530000000
0!
0'
0/
#345540000000
1!
1'
1/
#345550000000
0!
0'
0/
#345560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#345570000000
0!
0'
0/
#345580000000
1!
1'
1/
#345590000000
0!
0'
0/
#345600000000
1!
1'
1/
#345610000000
0!
0'
0/
#345620000000
1!
1'
1/
#345630000000
0!
0'
0/
#345640000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#345650000000
0!
0'
0/
#345660000000
1!
1'
1/
#345670000000
0!
0'
0/
#345680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#345690000000
0!
0'
0/
#345700000000
1!
1'
1/
#345710000000
0!
0'
0/
#345720000000
#345730000000
1!
1'
1/
#345740000000
0!
0'
0/
#345750000000
1!
1'
1/
#345760000000
0!
1"
0'
1(
0/
10
#345770000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#345780000000
0!
0'
0/
#345790000000
1!
1'
1/
#345800000000
0!
0'
0/
#345810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#345820000000
0!
0'
0/
#345830000000
1!
1'
1/
#345840000000
0!
1"
0'
1(
0/
10
#345850000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#345860000000
0!
1$
0'
1+
0/
#345870000000
1!
1'
1/
#345880000000
0!
0'
0/
#345890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#345900000000
0!
0'
0/
#345910000000
1!
1'
1/
#345920000000
0!
0'
0/
#345930000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#345940000000
0!
0'
0/
#345950000000
1!
1'
1/
#345960000000
0!
0'
0/
#345970000000
1!
1'
1/
#345980000000
0!
0'
0/
#345990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#346000000000
0!
0'
0/
#346010000000
1!
1'
1/
#346020000000
0!
0'
0/
#346030000000
1!
1'
1/
#346040000000
0!
0'
0/
#346050000000
1!
1'
1/
#346060000000
0!
0'
0/
#346070000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#346080000000
0!
0'
0/
#346090000000
1!
1'
1/
#346100000000
0!
0'
0/
#346110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#346120000000
0!
0'
0/
#346130000000
1!
1'
1/
#346140000000
0!
0'
0/
#346150000000
#346160000000
1!
1'
1/
#346170000000
0!
0'
0/
#346180000000
1!
1'
1/
#346190000000
0!
1"
0'
1(
0/
10
#346200000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#346210000000
0!
0'
0/
#346220000000
1!
1'
1/
#346230000000
0!
0'
0/
#346240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#346250000000
0!
0'
0/
#346260000000
1!
1'
1/
#346270000000
0!
1"
0'
1(
0/
10
#346280000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#346290000000
0!
1$
0'
1+
0/
#346300000000
1!
1'
1/
#346310000000
0!
0'
0/
#346320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#346330000000
0!
0'
0/
#346340000000
1!
1'
1/
#346350000000
0!
0'
0/
#346360000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#346370000000
0!
0'
0/
#346380000000
1!
1'
1/
#346390000000
0!
0'
0/
#346400000000
1!
1'
1/
#346410000000
0!
0'
0/
#346420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#346430000000
0!
0'
0/
#346440000000
1!
1'
1/
#346450000000
0!
0'
0/
#346460000000
1!
1'
1/
#346470000000
0!
0'
0/
#346480000000
1!
1'
1/
#346490000000
0!
0'
0/
#346500000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#346510000000
0!
0'
0/
#346520000000
1!
1'
1/
#346530000000
0!
0'
0/
#346540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#346550000000
0!
0'
0/
#346560000000
1!
1'
1/
#346570000000
0!
0'
0/
#346580000000
#346590000000
1!
1'
1/
#346600000000
0!
0'
0/
#346610000000
1!
1'
1/
#346620000000
0!
1"
0'
1(
0/
10
#346630000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#346640000000
0!
0'
0/
#346650000000
1!
1'
1/
#346660000000
0!
0'
0/
#346670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#346680000000
0!
0'
0/
#346690000000
1!
1'
1/
#346700000000
0!
1"
0'
1(
0/
10
#346710000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#346720000000
0!
1$
0'
1+
0/
#346730000000
1!
1'
1/
#346740000000
0!
0'
0/
#346750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#346760000000
0!
0'
0/
#346770000000
1!
1'
1/
#346780000000
0!
0'
0/
#346790000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#346800000000
0!
0'
0/
#346810000000
1!
1'
1/
#346820000000
0!
0'
0/
#346830000000
1!
1'
1/
#346840000000
0!
0'
0/
#346850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#346860000000
0!
0'
0/
#346870000000
1!
1'
1/
#346880000000
0!
0'
0/
#346890000000
1!
1'
1/
#346900000000
0!
0'
0/
#346910000000
1!
1'
1/
#346920000000
0!
0'
0/
#346930000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#346940000000
0!
0'
0/
#346950000000
1!
1'
1/
#346960000000
0!
0'
0/
#346970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#346980000000
0!
0'
0/
#346990000000
1!
1'
1/
#347000000000
0!
0'
0/
#347010000000
#347020000000
1!
1'
1/
#347030000000
0!
0'
0/
#347040000000
1!
1'
1/
#347050000000
0!
1"
0'
1(
0/
10
#347060000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#347070000000
0!
0'
0/
#347080000000
1!
1'
1/
#347090000000
0!
0'
0/
#347100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#347110000000
0!
0'
0/
#347120000000
1!
1'
1/
#347130000000
0!
1"
0'
1(
0/
10
#347140000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#347150000000
0!
1$
0'
1+
0/
#347160000000
1!
1'
1/
#347170000000
0!
0'
0/
#347180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#347190000000
0!
0'
0/
#347200000000
1!
1'
1/
#347210000000
0!
0'
0/
#347220000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#347230000000
0!
0'
0/
#347240000000
1!
1'
1/
#347250000000
0!
0'
0/
#347260000000
1!
1'
1/
#347270000000
0!
0'
0/
#347280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#347290000000
0!
0'
0/
#347300000000
1!
1'
1/
#347310000000
0!
0'
0/
#347320000000
1!
1'
1/
#347330000000
0!
0'
0/
#347340000000
1!
1'
1/
#347350000000
0!
0'
0/
#347360000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#347370000000
0!
0'
0/
#347380000000
1!
1'
1/
#347390000000
0!
0'
0/
#347400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#347410000000
0!
0'
0/
#347420000000
1!
1'
1/
#347430000000
0!
0'
0/
#347440000000
#347450000000
1!
1'
1/
#347460000000
0!
0'
0/
#347470000000
1!
1'
1/
#347480000000
0!
1"
0'
1(
0/
10
#347490000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#347500000000
0!
0'
0/
#347510000000
1!
1'
1/
#347520000000
0!
0'
0/
#347530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#347540000000
0!
0'
0/
#347550000000
1!
1'
1/
#347560000000
0!
1"
0'
1(
0/
10
#347570000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#347580000000
0!
1$
0'
1+
0/
#347590000000
1!
1'
1/
#347600000000
0!
0'
0/
#347610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#347620000000
0!
0'
0/
#347630000000
1!
1'
1/
#347640000000
0!
0'
0/
#347650000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#347660000000
0!
0'
0/
#347670000000
1!
1'
1/
#347680000000
0!
0'
0/
#347690000000
1!
1'
1/
#347700000000
0!
0'
0/
#347710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#347720000000
0!
0'
0/
#347730000000
1!
1'
1/
#347740000000
0!
0'
0/
#347750000000
1!
1'
1/
#347760000000
0!
0'
0/
#347770000000
1!
1'
1/
#347780000000
0!
0'
0/
#347790000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#347800000000
0!
0'
0/
#347810000000
1!
1'
1/
#347820000000
0!
0'
0/
#347830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#347840000000
0!
0'
0/
#347850000000
1!
1'
1/
#347860000000
0!
0'
0/
#347870000000
#347880000000
1!
1'
1/
#347890000000
0!
0'
0/
#347900000000
1!
1'
1/
#347910000000
0!
1"
0'
1(
0/
10
#347920000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#347930000000
0!
0'
0/
#347940000000
1!
1'
1/
#347950000000
0!
0'
0/
#347960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#347970000000
0!
0'
0/
#347980000000
1!
1'
1/
#347990000000
0!
1"
0'
1(
0/
10
#348000000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#348010000000
0!
1$
0'
1+
0/
#348020000000
1!
1'
1/
#348030000000
0!
0'
0/
#348040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#348050000000
0!
0'
0/
#348060000000
1!
1'
1/
#348070000000
0!
0'
0/
#348080000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#348090000000
0!
0'
0/
#348100000000
1!
1'
1/
#348110000000
0!
0'
0/
#348120000000
1!
1'
1/
#348130000000
0!
0'
0/
#348140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#348150000000
0!
0'
0/
#348160000000
1!
1'
1/
#348170000000
0!
0'
0/
#348180000000
1!
1'
1/
#348190000000
0!
0'
0/
#348200000000
1!
1'
1/
#348210000000
0!
0'
0/
#348220000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#348230000000
0!
0'
0/
#348240000000
1!
1'
1/
#348250000000
0!
0'
0/
#348260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#348270000000
0!
0'
0/
#348280000000
1!
1'
1/
#348290000000
0!
0'
0/
#348300000000
#348310000000
1!
1'
1/
#348320000000
0!
0'
0/
#348330000000
1!
1'
1/
#348340000000
0!
1"
0'
1(
0/
10
#348350000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#348360000000
0!
0'
0/
#348370000000
1!
1'
1/
#348380000000
0!
0'
0/
#348390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#348400000000
0!
0'
0/
#348410000000
1!
1'
1/
#348420000000
0!
1"
0'
1(
0/
10
#348430000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#348440000000
0!
1$
0'
1+
0/
#348450000000
1!
1'
1/
#348460000000
0!
0'
0/
#348470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#348480000000
0!
0'
0/
#348490000000
1!
1'
1/
#348500000000
0!
0'
0/
#348510000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#348520000000
0!
0'
0/
#348530000000
1!
1'
1/
#348540000000
0!
0'
0/
#348550000000
1!
1'
1/
#348560000000
0!
0'
0/
#348570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#348580000000
0!
0'
0/
#348590000000
1!
1'
1/
#348600000000
0!
0'
0/
#348610000000
1!
1'
1/
#348620000000
0!
0'
0/
#348630000000
1!
1'
1/
#348640000000
0!
0'
0/
#348650000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#348660000000
0!
0'
0/
#348670000000
1!
1'
1/
#348680000000
0!
0'
0/
#348690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#348700000000
0!
0'
0/
#348710000000
1!
1'
1/
#348720000000
0!
0'
0/
#348730000000
#348740000000
1!
1'
1/
#348750000000
0!
0'
0/
#348760000000
1!
1'
1/
#348770000000
0!
1"
0'
1(
0/
10
#348780000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#348790000000
0!
0'
0/
#348800000000
1!
1'
1/
#348810000000
0!
0'
0/
#348820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#348830000000
0!
0'
0/
#348840000000
1!
1'
1/
#348850000000
0!
1"
0'
1(
0/
10
#348860000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#348870000000
0!
1$
0'
1+
0/
#348880000000
1!
1'
1/
#348890000000
0!
0'
0/
#348900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#348910000000
0!
0'
0/
#348920000000
1!
1'
1/
#348930000000
0!
0'
0/
#348940000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#348950000000
0!
0'
0/
#348960000000
1!
1'
1/
#348970000000
0!
0'
0/
#348980000000
1!
1'
1/
#348990000000
0!
0'
0/
#349000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#349010000000
0!
0'
0/
#349020000000
1!
1'
1/
#349030000000
0!
0'
0/
#349040000000
1!
1'
1/
#349050000000
0!
0'
0/
#349060000000
1!
1'
1/
#349070000000
0!
0'
0/
#349080000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#349090000000
0!
0'
0/
#349100000000
1!
1'
1/
#349110000000
0!
0'
0/
#349120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#349130000000
0!
0'
0/
#349140000000
1!
1'
1/
#349150000000
0!
0'
0/
#349160000000
#349170000000
1!
1'
1/
#349180000000
0!
0'
0/
#349190000000
1!
1'
1/
#349200000000
0!
1"
0'
1(
0/
10
#349210000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#349220000000
0!
0'
0/
#349230000000
1!
1'
1/
#349240000000
0!
0'
0/
#349250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#349260000000
0!
0'
0/
#349270000000
1!
1'
1/
#349280000000
0!
1"
0'
1(
0/
10
#349290000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#349300000000
0!
1$
0'
1+
0/
#349310000000
1!
1'
1/
#349320000000
0!
0'
0/
#349330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#349340000000
0!
0'
0/
#349350000000
1!
1'
1/
#349360000000
0!
0'
0/
#349370000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#349380000000
0!
0'
0/
#349390000000
1!
1'
1/
#349400000000
0!
0'
0/
#349410000000
1!
1'
1/
#349420000000
0!
0'
0/
#349430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#349440000000
0!
0'
0/
#349450000000
1!
1'
1/
#349460000000
0!
0'
0/
#349470000000
1!
1'
1/
#349480000000
0!
0'
0/
#349490000000
1!
1'
1/
#349500000000
0!
0'
0/
#349510000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#349520000000
0!
0'
0/
#349530000000
1!
1'
1/
#349540000000
0!
0'
0/
#349550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#349560000000
0!
0'
0/
#349570000000
1!
1'
1/
#349580000000
0!
0'
0/
#349590000000
#349600000000
1!
1'
1/
#349610000000
0!
0'
0/
#349620000000
1!
1'
1/
#349630000000
0!
1"
0'
1(
0/
10
#349640000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#349650000000
0!
0'
0/
#349660000000
1!
1'
1/
#349670000000
0!
0'
0/
#349680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#349690000000
0!
0'
0/
#349700000000
1!
1'
1/
#349710000000
0!
1"
0'
1(
0/
10
#349720000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#349730000000
0!
1$
0'
1+
0/
#349740000000
1!
1'
1/
#349750000000
0!
0'
0/
#349760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#349770000000
0!
0'
0/
#349780000000
1!
1'
1/
#349790000000
0!
0'
0/
#349800000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#349810000000
0!
0'
0/
#349820000000
1!
1'
1/
#349830000000
0!
0'
0/
#349840000000
1!
1'
1/
#349850000000
0!
0'
0/
#349860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#349870000000
0!
0'
0/
#349880000000
1!
1'
1/
#349890000000
0!
0'
0/
#349900000000
1!
1'
1/
#349910000000
0!
0'
0/
#349920000000
1!
1'
1/
#349930000000
0!
0'
0/
#349940000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#349950000000
0!
0'
0/
#349960000000
1!
1'
1/
#349970000000
0!
0'
0/
#349980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#349990000000
0!
0'
0/
#350000000000
1!
1'
1/
#350010000000
0!
0'
0/
#350020000000
#350030000000
1!
1'
1/
#350040000000
0!
0'
0/
#350050000000
1!
1'
1/
#350060000000
0!
1"
0'
1(
0/
10
#350070000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#350080000000
0!
0'
0/
#350090000000
1!
1'
1/
#350100000000
0!
0'
0/
#350110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#350120000000
0!
0'
0/
#350130000000
1!
1'
1/
#350140000000
0!
1"
0'
1(
0/
10
#350150000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#350160000000
0!
1$
0'
1+
0/
#350170000000
1!
1'
1/
#350180000000
0!
0'
0/
#350190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#350200000000
0!
0'
0/
#350210000000
1!
1'
1/
#350220000000
0!
0'
0/
#350230000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#350240000000
0!
0'
0/
#350250000000
1!
1'
1/
#350260000000
0!
0'
0/
#350270000000
1!
1'
1/
#350280000000
0!
0'
0/
#350290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#350300000000
0!
0'
0/
#350310000000
1!
1'
1/
#350320000000
0!
0'
0/
#350330000000
1!
1'
1/
#350340000000
0!
0'
0/
#350350000000
1!
1'
1/
#350360000000
0!
0'
0/
#350370000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#350380000000
0!
0'
0/
#350390000000
1!
1'
1/
#350400000000
0!
0'
0/
#350410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#350420000000
0!
0'
0/
#350430000000
1!
1'
1/
#350440000000
0!
0'
0/
#350450000000
#350460000000
1!
1'
1/
#350470000000
0!
0'
0/
#350480000000
1!
1'
1/
#350490000000
0!
1"
0'
1(
0/
10
#350500000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#350510000000
0!
0'
0/
#350520000000
1!
1'
1/
#350530000000
0!
0'
0/
#350540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#350550000000
0!
0'
0/
#350560000000
1!
1'
1/
#350570000000
0!
1"
0'
1(
0/
10
#350580000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#350590000000
0!
1$
0'
1+
0/
#350600000000
1!
1'
1/
#350610000000
0!
0'
0/
#350620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#350630000000
0!
0'
0/
#350640000000
1!
1'
1/
#350650000000
0!
0'
0/
#350660000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#350670000000
0!
0'
0/
#350680000000
1!
1'
1/
#350690000000
0!
0'
0/
#350700000000
1!
1'
1/
#350710000000
0!
0'
0/
#350720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#350730000000
0!
0'
0/
#350740000000
1!
1'
1/
#350750000000
0!
0'
0/
#350760000000
1!
1'
1/
#350770000000
0!
0'
0/
#350780000000
1!
1'
1/
#350790000000
0!
0'
0/
#350800000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#350810000000
0!
0'
0/
#350820000000
1!
1'
1/
#350830000000
0!
0'
0/
#350840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#350850000000
0!
0'
0/
#350860000000
1!
1'
1/
#350870000000
0!
0'
0/
#350880000000
#350890000000
1!
1'
1/
#350900000000
0!
0'
0/
#350910000000
1!
1'
1/
#350920000000
0!
1"
0'
1(
0/
10
#350930000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#350940000000
0!
0'
0/
#350950000000
1!
1'
1/
#350960000000
0!
0'
0/
#350970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#350980000000
0!
0'
0/
#350990000000
1!
1'
1/
#351000000000
0!
1"
0'
1(
0/
10
#351010000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#351020000000
0!
1$
0'
1+
0/
#351030000000
1!
1'
1/
#351040000000
0!
0'
0/
#351050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#351060000000
0!
0'
0/
#351070000000
1!
1'
1/
#351080000000
0!
0'
0/
#351090000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#351100000000
0!
0'
0/
#351110000000
1!
1'
1/
#351120000000
0!
0'
0/
#351130000000
1!
1'
1/
#351140000000
0!
0'
0/
#351150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#351160000000
0!
0'
0/
#351170000000
1!
1'
1/
#351180000000
0!
0'
0/
#351190000000
1!
1'
1/
#351200000000
0!
0'
0/
#351210000000
1!
1'
1/
#351220000000
0!
0'
0/
#351230000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#351240000000
0!
0'
0/
#351250000000
1!
1'
1/
#351260000000
0!
0'
0/
#351270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#351280000000
0!
0'
0/
#351290000000
1!
1'
1/
#351300000000
0!
0'
0/
#351310000000
#351320000000
1!
1'
1/
#351330000000
0!
0'
0/
#351340000000
1!
1'
1/
#351350000000
0!
1"
0'
1(
0/
10
#351360000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#351370000000
0!
0'
0/
#351380000000
1!
1'
1/
#351390000000
0!
0'
0/
#351400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#351410000000
0!
0'
0/
#351420000000
1!
1'
1/
#351430000000
0!
1"
0'
1(
0/
10
#351440000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#351450000000
0!
1$
0'
1+
0/
#351460000000
1!
1'
1/
#351470000000
0!
0'
0/
#351480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#351490000000
0!
0'
0/
#351500000000
1!
1'
1/
#351510000000
0!
0'
0/
#351520000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#351530000000
0!
0'
0/
#351540000000
1!
1'
1/
#351550000000
0!
0'
0/
#351560000000
1!
1'
1/
#351570000000
0!
0'
0/
#351580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#351590000000
0!
0'
0/
#351600000000
1!
1'
1/
#351610000000
0!
0'
0/
#351620000000
1!
1'
1/
#351630000000
0!
0'
0/
#351640000000
1!
1'
1/
#351650000000
0!
0'
0/
#351660000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#351670000000
0!
0'
0/
#351680000000
1!
1'
1/
#351690000000
0!
0'
0/
#351700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#351710000000
0!
0'
0/
#351720000000
1!
1'
1/
#351730000000
0!
0'
0/
#351740000000
#351750000000
1!
1'
1/
#351760000000
0!
0'
0/
#351770000000
1!
1'
1/
#351780000000
0!
1"
0'
1(
0/
10
#351790000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#351800000000
0!
0'
0/
#351810000000
1!
1'
1/
#351820000000
0!
0'
0/
#351830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#351840000000
0!
0'
0/
#351850000000
1!
1'
1/
#351860000000
0!
1"
0'
1(
0/
10
#351870000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#351880000000
0!
1$
0'
1+
0/
#351890000000
1!
1'
1/
#351900000000
0!
0'
0/
#351910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#351920000000
0!
0'
0/
#351930000000
1!
1'
1/
#351940000000
0!
0'
0/
#351950000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#351960000000
0!
0'
0/
#351970000000
1!
1'
1/
#351980000000
0!
0'
0/
#351990000000
1!
1'
1/
#352000000000
0!
0'
0/
#352010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#352020000000
0!
0'
0/
#352030000000
1!
1'
1/
#352040000000
0!
0'
0/
#352050000000
1!
1'
1/
#352060000000
0!
0'
0/
#352070000000
1!
1'
1/
#352080000000
0!
0'
0/
#352090000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#352100000000
0!
0'
0/
#352110000000
1!
1'
1/
#352120000000
0!
0'
0/
#352130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#352140000000
0!
0'
0/
#352150000000
1!
1'
1/
#352160000000
0!
0'
0/
#352170000000
#352180000000
1!
1'
1/
#352190000000
0!
0'
0/
#352200000000
1!
1'
1/
#352210000000
0!
1"
0'
1(
0/
10
#352220000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#352230000000
0!
0'
0/
#352240000000
1!
1'
1/
#352250000000
0!
0'
0/
#352260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#352270000000
0!
0'
0/
#352280000000
1!
1'
1/
#352290000000
0!
1"
0'
1(
0/
10
#352300000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#352310000000
0!
1$
0'
1+
0/
#352320000000
1!
1'
1/
#352330000000
0!
0'
0/
#352340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#352350000000
0!
0'
0/
#352360000000
1!
1'
1/
#352370000000
0!
0'
0/
#352380000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#352390000000
0!
0'
0/
#352400000000
1!
1'
1/
#352410000000
0!
0'
0/
#352420000000
1!
1'
1/
#352430000000
0!
0'
0/
#352440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#352450000000
0!
0'
0/
#352460000000
1!
1'
1/
#352470000000
0!
0'
0/
#352480000000
1!
1'
1/
#352490000000
0!
0'
0/
#352500000000
1!
1'
1/
#352510000000
0!
0'
0/
#352520000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#352530000000
0!
0'
0/
#352540000000
1!
1'
1/
#352550000000
0!
0'
0/
#352560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#352570000000
0!
0'
0/
#352580000000
1!
1'
1/
#352590000000
0!
0'
0/
#352600000000
#352610000000
1!
1'
1/
#352620000000
0!
0'
0/
#352630000000
1!
1'
1/
#352640000000
0!
1"
0'
1(
0/
10
#352650000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#352660000000
0!
0'
0/
#352670000000
1!
1'
1/
#352680000000
0!
0'
0/
#352690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#352700000000
0!
0'
0/
#352710000000
1!
1'
1/
#352720000000
0!
1"
0'
1(
0/
10
#352730000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#352740000000
0!
1$
0'
1+
0/
#352750000000
1!
1'
1/
#352760000000
0!
0'
0/
#352770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#352780000000
0!
0'
0/
#352790000000
1!
1'
1/
#352800000000
0!
0'
0/
#352810000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#352820000000
0!
0'
0/
#352830000000
1!
1'
1/
#352840000000
0!
0'
0/
#352850000000
1!
1'
1/
#352860000000
0!
0'
0/
#352870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#352880000000
0!
0'
0/
#352890000000
1!
1'
1/
#352900000000
0!
0'
0/
#352910000000
1!
1'
1/
#352920000000
0!
0'
0/
#352930000000
1!
1'
1/
#352940000000
0!
0'
0/
#352950000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#352960000000
0!
0'
0/
#352970000000
1!
1'
1/
#352980000000
0!
0'
0/
#352990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#353000000000
0!
0'
0/
#353010000000
1!
1'
1/
#353020000000
0!
0'
0/
#353030000000
#353040000000
1!
1'
1/
#353050000000
0!
0'
0/
#353060000000
1!
1'
1/
#353070000000
0!
1"
0'
1(
0/
10
#353080000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#353090000000
0!
0'
0/
#353100000000
1!
1'
1/
#353110000000
0!
0'
0/
#353120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#353130000000
0!
0'
0/
#353140000000
1!
1'
1/
#353150000000
0!
1"
0'
1(
0/
10
#353160000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#353170000000
0!
1$
0'
1+
0/
#353180000000
1!
1'
1/
#353190000000
0!
0'
0/
#353200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#353210000000
0!
0'
0/
#353220000000
1!
1'
1/
#353230000000
0!
0'
0/
#353240000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#353250000000
0!
0'
0/
#353260000000
1!
1'
1/
#353270000000
0!
0'
0/
#353280000000
1!
1'
1/
#353290000000
0!
0'
0/
#353300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#353310000000
0!
0'
0/
#353320000000
1!
1'
1/
#353330000000
0!
0'
0/
#353340000000
1!
1'
1/
#353350000000
0!
0'
0/
#353360000000
1!
1'
1/
#353370000000
0!
0'
0/
#353380000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#353390000000
0!
0'
0/
#353400000000
1!
1'
1/
#353410000000
0!
0'
0/
#353420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#353430000000
0!
0'
0/
#353440000000
1!
1'
1/
#353450000000
0!
0'
0/
#353460000000
#353470000000
1!
1'
1/
#353480000000
0!
0'
0/
#353490000000
1!
1'
1/
#353500000000
0!
1"
0'
1(
0/
10
#353510000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#353520000000
0!
0'
0/
#353530000000
1!
1'
1/
#353540000000
0!
0'
0/
#353550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#353560000000
0!
0'
0/
#353570000000
1!
1'
1/
#353580000000
0!
1"
0'
1(
0/
10
#353590000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#353600000000
0!
1$
0'
1+
0/
#353610000000
1!
1'
1/
#353620000000
0!
0'
0/
#353630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#353640000000
0!
0'
0/
#353650000000
1!
1'
1/
#353660000000
0!
0'
0/
#353670000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#353680000000
0!
0'
0/
#353690000000
1!
1'
1/
#353700000000
0!
0'
0/
#353710000000
1!
1'
1/
#353720000000
0!
0'
0/
#353730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#353740000000
0!
0'
0/
#353750000000
1!
1'
1/
#353760000000
0!
0'
0/
#353770000000
1!
1'
1/
#353780000000
0!
0'
0/
#353790000000
1!
1'
1/
#353800000000
0!
0'
0/
#353810000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#353820000000
0!
0'
0/
#353830000000
1!
1'
1/
#353840000000
0!
0'
0/
#353850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#353860000000
0!
0'
0/
#353870000000
1!
1'
1/
#353880000000
0!
0'
0/
#353890000000
#353900000000
1!
1'
1/
#353910000000
0!
0'
0/
#353920000000
1!
1'
1/
#353930000000
0!
1"
0'
1(
0/
10
#353940000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#353950000000
0!
0'
0/
#353960000000
1!
1'
1/
#353970000000
0!
0'
0/
#353980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#353990000000
0!
0'
0/
#354000000000
1!
1'
1/
#354010000000
0!
1"
0'
1(
0/
10
#354020000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#354030000000
0!
1$
0'
1+
0/
#354040000000
1!
1'
1/
#354050000000
0!
0'
0/
#354060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#354070000000
0!
0'
0/
#354080000000
1!
1'
1/
#354090000000
0!
0'
0/
#354100000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#354110000000
0!
0'
0/
#354120000000
1!
1'
1/
#354130000000
0!
0'
0/
#354140000000
1!
1'
1/
#354150000000
0!
0'
0/
#354160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#354170000000
0!
0'
0/
#354180000000
1!
1'
1/
#354190000000
0!
0'
0/
#354200000000
1!
1'
1/
#354210000000
0!
0'
0/
#354220000000
1!
1'
1/
#354230000000
0!
0'
0/
#354240000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#354250000000
0!
0'
0/
#354260000000
1!
1'
1/
#354270000000
0!
0'
0/
#354280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#354290000000
0!
0'
0/
#354300000000
1!
1'
1/
#354310000000
0!
0'
0/
#354320000000
#354330000000
1!
1'
1/
#354340000000
0!
0'
0/
#354350000000
1!
1'
1/
#354360000000
0!
1"
0'
1(
0/
10
#354370000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#354380000000
0!
0'
0/
#354390000000
1!
1'
1/
#354400000000
0!
0'
0/
#354410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#354420000000
0!
0'
0/
#354430000000
1!
1'
1/
#354440000000
0!
1"
0'
1(
0/
10
#354450000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#354460000000
0!
1$
0'
1+
0/
#354470000000
1!
1'
1/
#354480000000
0!
0'
0/
#354490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#354500000000
0!
0'
0/
#354510000000
1!
1'
1/
#354520000000
0!
0'
0/
#354530000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#354540000000
0!
0'
0/
#354550000000
1!
1'
1/
#354560000000
0!
0'
0/
#354570000000
1!
1'
1/
#354580000000
0!
0'
0/
#354590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#354600000000
0!
0'
0/
#354610000000
1!
1'
1/
#354620000000
0!
0'
0/
#354630000000
1!
1'
1/
#354640000000
0!
0'
0/
#354650000000
1!
1'
1/
#354660000000
0!
0'
0/
#354670000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#354680000000
0!
0'
0/
#354690000000
1!
1'
1/
#354700000000
0!
0'
0/
#354710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#354720000000
0!
0'
0/
#354730000000
1!
1'
1/
#354740000000
0!
0'
0/
#354750000000
#354760000000
1!
1'
1/
#354770000000
0!
0'
0/
#354780000000
1!
1'
1/
#354790000000
0!
1"
0'
1(
0/
10
#354800000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#354810000000
0!
0'
0/
#354820000000
1!
1'
1/
#354830000000
0!
0'
0/
#354840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#354850000000
0!
0'
0/
#354860000000
1!
1'
1/
#354870000000
0!
1"
0'
1(
0/
10
#354880000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#354890000000
0!
1$
0'
1+
0/
#354900000000
1!
1'
1/
#354910000000
0!
0'
0/
#354920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#354930000000
0!
0'
0/
#354940000000
1!
1'
1/
#354950000000
0!
0'
0/
#354960000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#354970000000
0!
0'
0/
#354980000000
1!
1'
1/
#354990000000
0!
0'
0/
#355000000000
1!
1'
1/
#355010000000
0!
0'
0/
#355020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#355030000000
0!
0'
0/
#355040000000
1!
1'
1/
#355050000000
0!
0'
0/
#355060000000
1!
1'
1/
#355070000000
0!
0'
0/
#355080000000
1!
1'
1/
#355090000000
0!
0'
0/
#355100000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#355110000000
0!
0'
0/
#355120000000
1!
1'
1/
#355130000000
0!
0'
0/
#355140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#355150000000
0!
0'
0/
#355160000000
1!
1'
1/
#355170000000
0!
0'
0/
#355180000000
#355190000000
1!
1'
1/
#355200000000
0!
0'
0/
#355210000000
1!
1'
1/
#355220000000
0!
1"
0'
1(
0/
10
#355230000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#355240000000
0!
0'
0/
#355250000000
1!
1'
1/
#355260000000
0!
0'
0/
#355270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#355280000000
0!
0'
0/
#355290000000
1!
1'
1/
#355300000000
0!
1"
0'
1(
0/
10
#355310000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#355320000000
0!
1$
0'
1+
0/
#355330000000
1!
1'
1/
#355340000000
0!
0'
0/
#355350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#355360000000
0!
0'
0/
#355370000000
1!
1'
1/
#355380000000
0!
0'
0/
#355390000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#355400000000
0!
0'
0/
#355410000000
1!
1'
1/
#355420000000
0!
0'
0/
#355430000000
1!
1'
1/
#355440000000
0!
0'
0/
#355450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#355460000000
0!
0'
0/
#355470000000
1!
1'
1/
#355480000000
0!
0'
0/
#355490000000
1!
1'
1/
#355500000000
0!
0'
0/
#355510000000
1!
1'
1/
#355520000000
0!
0'
0/
#355530000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#355540000000
0!
0'
0/
#355550000000
1!
1'
1/
#355560000000
0!
0'
0/
#355570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#355580000000
0!
0'
0/
#355590000000
1!
1'
1/
#355600000000
0!
0'
0/
#355610000000
#355620000000
1!
1'
1/
#355630000000
0!
0'
0/
#355640000000
1!
1'
1/
#355650000000
0!
1"
0'
1(
0/
10
#355660000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#355670000000
0!
0'
0/
#355680000000
1!
1'
1/
#355690000000
0!
0'
0/
#355700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#355710000000
0!
0'
0/
#355720000000
1!
1'
1/
#355730000000
0!
1"
0'
1(
0/
10
#355740000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#355750000000
0!
1$
0'
1+
0/
#355760000000
1!
1'
1/
#355770000000
0!
0'
0/
#355780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#355790000000
0!
0'
0/
#355800000000
1!
1'
1/
#355810000000
0!
0'
0/
#355820000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#355830000000
0!
0'
0/
#355840000000
1!
1'
1/
#355850000000
0!
0'
0/
#355860000000
1!
1'
1/
#355870000000
0!
0'
0/
#355880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#355890000000
0!
0'
0/
#355900000000
1!
1'
1/
#355910000000
0!
0'
0/
#355920000000
1!
1'
1/
#355930000000
0!
0'
0/
#355940000000
1!
1'
1/
#355950000000
0!
0'
0/
#355960000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#355970000000
0!
0'
0/
#355980000000
1!
1'
1/
#355990000000
0!
0'
0/
#356000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#356010000000
0!
0'
0/
#356020000000
1!
1'
1/
#356030000000
0!
0'
0/
#356040000000
#356050000000
1!
1'
1/
#356060000000
0!
0'
0/
#356070000000
1!
1'
1/
#356080000000
0!
1"
0'
1(
0/
10
#356090000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#356100000000
0!
0'
0/
#356110000000
1!
1'
1/
#356120000000
0!
0'
0/
#356130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#356140000000
0!
0'
0/
#356150000000
1!
1'
1/
#356160000000
0!
1"
0'
1(
0/
10
#356170000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#356180000000
0!
1$
0'
1+
0/
#356190000000
1!
1'
1/
#356200000000
0!
0'
0/
#356210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#356220000000
0!
0'
0/
#356230000000
1!
1'
1/
#356240000000
0!
0'
0/
#356250000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#356260000000
0!
0'
0/
#356270000000
1!
1'
1/
#356280000000
0!
0'
0/
#356290000000
1!
1'
1/
#356300000000
0!
0'
0/
#356310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#356320000000
0!
0'
0/
#356330000000
1!
1'
1/
#356340000000
0!
0'
0/
#356350000000
1!
1'
1/
#356360000000
0!
0'
0/
#356370000000
1!
1'
1/
#356380000000
0!
0'
0/
#356390000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#356400000000
0!
0'
0/
#356410000000
1!
1'
1/
#356420000000
0!
0'
0/
#356430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#356440000000
0!
0'
0/
#356450000000
1!
1'
1/
#356460000000
0!
0'
0/
#356470000000
#356480000000
1!
1'
1/
#356490000000
0!
0'
0/
#356500000000
1!
1'
1/
#356510000000
0!
1"
0'
1(
0/
10
#356520000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#356530000000
0!
0'
0/
#356540000000
1!
1'
1/
#356550000000
0!
0'
0/
#356560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#356570000000
0!
0'
0/
#356580000000
1!
1'
1/
#356590000000
0!
1"
0'
1(
0/
10
#356600000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#356610000000
0!
1$
0'
1+
0/
#356620000000
1!
1'
1/
#356630000000
0!
0'
0/
#356640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#356650000000
0!
0'
0/
#356660000000
1!
1'
1/
#356670000000
0!
0'
0/
#356680000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#356690000000
0!
0'
0/
#356700000000
1!
1'
1/
#356710000000
0!
0'
0/
#356720000000
1!
1'
1/
#356730000000
0!
0'
0/
#356740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#356750000000
0!
0'
0/
#356760000000
1!
1'
1/
#356770000000
0!
0'
0/
#356780000000
1!
1'
1/
#356790000000
0!
0'
0/
#356800000000
1!
1'
1/
#356810000000
0!
0'
0/
#356820000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#356830000000
0!
0'
0/
#356840000000
1!
1'
1/
#356850000000
0!
0'
0/
#356860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#356870000000
0!
0'
0/
#356880000000
1!
1'
1/
#356890000000
0!
0'
0/
#356900000000
#356910000000
1!
1'
1/
#356920000000
0!
0'
0/
#356930000000
1!
1'
1/
#356940000000
0!
1"
0'
1(
0/
10
#356950000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#356960000000
0!
0'
0/
#356970000000
1!
1'
1/
#356980000000
0!
0'
0/
#356990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#357000000000
0!
0'
0/
#357010000000
1!
1'
1/
#357020000000
0!
1"
0'
1(
0/
10
#357030000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#357040000000
0!
1$
0'
1+
0/
#357050000000
1!
1'
1/
#357060000000
0!
0'
0/
#357070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#357080000000
0!
0'
0/
#357090000000
1!
1'
1/
#357100000000
0!
0'
0/
#357110000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#357120000000
0!
0'
0/
#357130000000
1!
1'
1/
#357140000000
0!
0'
0/
#357150000000
1!
1'
1/
#357160000000
0!
0'
0/
#357170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#357180000000
0!
0'
0/
#357190000000
1!
1'
1/
#357200000000
0!
0'
0/
#357210000000
1!
1'
1/
#357220000000
0!
0'
0/
#357230000000
1!
1'
1/
#357240000000
0!
0'
0/
#357250000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#357260000000
0!
0'
0/
#357270000000
1!
1'
1/
#357280000000
0!
0'
0/
#357290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#357300000000
0!
0'
0/
#357310000000
1!
1'
1/
#357320000000
0!
0'
0/
#357330000000
#357340000000
1!
1'
1/
#357350000000
0!
0'
0/
#357360000000
1!
1'
1/
#357370000000
0!
1"
0'
1(
0/
10
#357380000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#357390000000
0!
0'
0/
#357400000000
1!
1'
1/
#357410000000
0!
0'
0/
#357420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#357430000000
0!
0'
0/
#357440000000
1!
1'
1/
#357450000000
0!
1"
0'
1(
0/
10
#357460000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#357470000000
0!
1$
0'
1+
0/
#357480000000
1!
1'
1/
#357490000000
0!
0'
0/
#357500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#357510000000
0!
0'
0/
#357520000000
1!
1'
1/
#357530000000
0!
0'
0/
#357540000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#357550000000
0!
0'
0/
#357560000000
1!
1'
1/
#357570000000
0!
0'
0/
#357580000000
1!
1'
1/
#357590000000
0!
0'
0/
#357600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#357610000000
0!
0'
0/
#357620000000
1!
1'
1/
#357630000000
0!
0'
0/
#357640000000
1!
1'
1/
#357650000000
0!
0'
0/
#357660000000
1!
1'
1/
#357670000000
0!
0'
0/
#357680000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#357690000000
0!
0'
0/
#357700000000
1!
1'
1/
#357710000000
0!
0'
0/
#357720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#357730000000
0!
0'
0/
#357740000000
1!
1'
1/
#357750000000
0!
0'
0/
#357760000000
#357770000000
1!
1'
1/
#357780000000
0!
0'
0/
#357790000000
1!
1'
1/
#357800000000
0!
1"
0'
1(
0/
10
#357810000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#357820000000
0!
0'
0/
#357830000000
1!
1'
1/
#357840000000
0!
0'
0/
#357850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#357860000000
0!
0'
0/
#357870000000
1!
1'
1/
#357880000000
0!
1"
0'
1(
0/
10
#357890000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#357900000000
0!
1$
0'
1+
0/
#357910000000
1!
1'
1/
#357920000000
0!
0'
0/
#357930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#357940000000
0!
0'
0/
#357950000000
1!
1'
1/
#357960000000
0!
0'
0/
#357970000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#357980000000
0!
0'
0/
#357990000000
1!
1'
1/
#358000000000
0!
0'
0/
#358010000000
1!
1'
1/
#358020000000
0!
0'
0/
#358030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#358040000000
0!
0'
0/
#358050000000
1!
1'
1/
#358060000000
0!
0'
0/
#358070000000
1!
1'
1/
#358080000000
0!
0'
0/
#358090000000
1!
1'
1/
#358100000000
0!
0'
0/
#358110000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#358120000000
0!
0'
0/
#358130000000
1!
1'
1/
#358140000000
0!
0'
0/
#358150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#358160000000
0!
0'
0/
#358170000000
1!
1'
1/
#358180000000
0!
0'
0/
#358190000000
#358200000000
1!
1'
1/
#358210000000
0!
0'
0/
#358220000000
1!
1'
1/
#358230000000
0!
1"
0'
1(
0/
10
#358240000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#358250000000
0!
0'
0/
#358260000000
1!
1'
1/
#358270000000
0!
0'
0/
#358280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#358290000000
0!
0'
0/
#358300000000
1!
1'
1/
#358310000000
0!
1"
0'
1(
0/
10
#358320000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#358330000000
0!
1$
0'
1+
0/
#358340000000
1!
1'
1/
#358350000000
0!
0'
0/
#358360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#358370000000
0!
0'
0/
#358380000000
1!
1'
1/
#358390000000
0!
0'
0/
#358400000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#358410000000
0!
0'
0/
#358420000000
1!
1'
1/
#358430000000
0!
0'
0/
#358440000000
1!
1'
1/
#358450000000
0!
0'
0/
#358460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#358470000000
0!
0'
0/
#358480000000
1!
1'
1/
#358490000000
0!
0'
0/
#358500000000
1!
1'
1/
#358510000000
0!
0'
0/
#358520000000
1!
1'
1/
#358530000000
0!
0'
0/
#358540000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#358550000000
0!
0'
0/
#358560000000
1!
1'
1/
#358570000000
0!
0'
0/
#358580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#358590000000
0!
0'
0/
#358600000000
1!
1'
1/
#358610000000
0!
0'
0/
#358620000000
#358630000000
1!
1'
1/
#358640000000
0!
0'
0/
#358650000000
1!
1'
1/
#358660000000
0!
1"
0'
1(
0/
10
#358670000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#358680000000
0!
0'
0/
#358690000000
1!
1'
1/
#358700000000
0!
0'
0/
#358710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#358720000000
0!
0'
0/
#358730000000
1!
1'
1/
#358740000000
0!
1"
0'
1(
0/
10
#358750000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#358760000000
0!
1$
0'
1+
0/
#358770000000
1!
1'
1/
#358780000000
0!
0'
0/
#358790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#358800000000
0!
0'
0/
#358810000000
1!
1'
1/
#358820000000
0!
0'
0/
#358830000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#358840000000
0!
0'
0/
#358850000000
1!
1'
1/
#358860000000
0!
0'
0/
#358870000000
1!
1'
1/
#358880000000
0!
0'
0/
#358890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#358900000000
0!
0'
0/
#358910000000
1!
1'
1/
#358920000000
0!
0'
0/
#358930000000
1!
1'
1/
#358940000000
0!
0'
0/
#358950000000
1!
1'
1/
#358960000000
0!
0'
0/
#358970000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#358980000000
0!
0'
0/
#358990000000
1!
1'
1/
#359000000000
0!
0'
0/
#359010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#359020000000
0!
0'
0/
#359030000000
1!
1'
1/
#359040000000
0!
0'
0/
#359050000000
#359060000000
1!
1'
1/
#359070000000
0!
0'
0/
#359080000000
1!
1'
1/
#359090000000
0!
1"
0'
1(
0/
10
#359100000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#359110000000
0!
0'
0/
#359120000000
1!
1'
1/
#359130000000
0!
0'
0/
#359140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#359150000000
0!
0'
0/
#359160000000
1!
1'
1/
#359170000000
0!
1"
0'
1(
0/
10
#359180000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#359190000000
0!
1$
0'
1+
0/
#359200000000
1!
1'
1/
#359210000000
0!
0'
0/
#359220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#359230000000
0!
0'
0/
#359240000000
1!
1'
1/
#359250000000
0!
0'
0/
#359260000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#359270000000
0!
0'
0/
#359280000000
1!
1'
1/
#359290000000
0!
0'
0/
#359300000000
1!
1'
1/
#359310000000
0!
0'
0/
#359320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#359330000000
0!
0'
0/
#359340000000
1!
1'
1/
#359350000000
0!
0'
0/
#359360000000
1!
1'
1/
#359370000000
0!
0'
0/
#359380000000
1!
1'
1/
#359390000000
0!
0'
0/
#359400000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#359410000000
0!
0'
0/
#359420000000
1!
1'
1/
#359430000000
0!
0'
0/
#359440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#359450000000
0!
0'
0/
#359460000000
1!
1'
1/
#359470000000
0!
0'
0/
#359480000000
#359490000000
1!
1'
1/
#359500000000
0!
0'
0/
#359510000000
1!
1'
1/
#359520000000
0!
1"
0'
1(
0/
10
#359530000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#359540000000
0!
0'
0/
#359550000000
1!
1'
1/
#359560000000
0!
0'
0/
#359570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#359580000000
0!
0'
0/
#359590000000
1!
1'
1/
#359600000000
0!
1"
0'
1(
0/
10
#359610000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#359620000000
0!
1$
0'
1+
0/
#359630000000
1!
1'
1/
#359640000000
0!
0'
0/
#359650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#359660000000
0!
0'
0/
#359670000000
1!
1'
1/
#359680000000
0!
0'
0/
#359690000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#359700000000
0!
0'
0/
#359710000000
1!
1'
1/
#359720000000
0!
0'
0/
#359730000000
1!
1'
1/
#359740000000
0!
0'
0/
#359750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#359760000000
0!
0'
0/
#359770000000
1!
1'
1/
#359780000000
0!
0'
0/
#359790000000
1!
1'
1/
#359800000000
0!
0'
0/
#359810000000
1!
1'
1/
#359820000000
0!
0'
0/
#359830000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#359840000000
0!
0'
0/
#359850000000
1!
1'
1/
#359860000000
0!
0'
0/
#359870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#359880000000
0!
0'
0/
#359890000000
1!
1'
1/
#359900000000
0!
0'
0/
#359910000000
#359920000000
1!
1'
1/
#359930000000
0!
0'
0/
#359940000000
1!
1'
1/
#359950000000
0!
1"
0'
1(
0/
10
#359960000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#359970000000
0!
0'
0/
#359980000000
1!
1'
1/
#359990000000
0!
0'
0/
#360000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#360010000000
0!
0'
0/
#360020000000
1!
1'
1/
#360030000000
0!
1"
0'
1(
0/
10
#360040000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#360050000000
0!
1$
0'
1+
0/
#360060000000
1!
1'
1/
#360070000000
0!
0'
0/
#360080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#360090000000
0!
0'
0/
#360100000000
1!
1'
1/
#360110000000
0!
0'
0/
#360120000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#360130000000
0!
0'
0/
#360140000000
1!
1'
1/
#360150000000
0!
0'
0/
#360160000000
1!
1'
1/
#360170000000
0!
0'
0/
#360180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#360190000000
0!
0'
0/
#360200000000
1!
1'
1/
#360210000000
0!
0'
0/
#360220000000
1!
1'
1/
#360230000000
0!
0'
0/
#360240000000
1!
1'
1/
#360250000000
0!
0'
0/
#360260000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#360270000000
0!
0'
0/
#360280000000
1!
1'
1/
#360290000000
0!
0'
0/
#360300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#360310000000
0!
0'
0/
#360320000000
1!
1'
1/
#360330000000
0!
0'
0/
#360340000000
#360350000000
1!
1'
1/
#360360000000
0!
0'
0/
#360370000000
1!
1'
1/
#360380000000
0!
1"
0'
1(
0/
10
#360390000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#360400000000
0!
0'
0/
#360410000000
1!
1'
1/
#360420000000
0!
0'
0/
#360430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#360440000000
0!
0'
0/
#360450000000
1!
1'
1/
#360460000000
0!
1"
0'
1(
0/
10
#360470000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#360480000000
0!
1$
0'
1+
0/
#360490000000
1!
1'
1/
#360500000000
0!
0'
0/
#360510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#360520000000
0!
0'
0/
#360530000000
1!
1'
1/
#360540000000
0!
0'
0/
#360550000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#360560000000
0!
0'
0/
#360570000000
1!
1'
1/
#360580000000
0!
0'
0/
#360590000000
1!
1'
1/
#360600000000
0!
0'
0/
#360610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#360620000000
0!
0'
0/
#360630000000
1!
1'
1/
#360640000000
0!
0'
0/
#360650000000
1!
1'
1/
#360660000000
0!
0'
0/
#360670000000
1!
1'
1/
#360680000000
0!
0'
0/
#360690000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#360700000000
0!
0'
0/
#360710000000
1!
1'
1/
#360720000000
0!
0'
0/
#360730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#360740000000
0!
0'
0/
#360750000000
1!
1'
1/
#360760000000
0!
0'
0/
#360770000000
#360780000000
1!
1'
1/
#360790000000
0!
0'
0/
#360800000000
1!
1'
1/
#360810000000
0!
1"
0'
1(
0/
10
#360820000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#360830000000
0!
0'
0/
#360840000000
1!
1'
1/
#360850000000
0!
0'
0/
#360860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#360870000000
0!
0'
0/
#360880000000
1!
1'
1/
#360890000000
0!
1"
0'
1(
0/
10
#360900000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#360910000000
0!
1$
0'
1+
0/
#360920000000
1!
1'
1/
#360930000000
0!
0'
0/
#360940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#360950000000
0!
0'
0/
#360960000000
1!
1'
1/
#360970000000
0!
0'
0/
#360980000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#360990000000
0!
0'
0/
#361000000000
1!
1'
1/
#361010000000
0!
0'
0/
#361020000000
1!
1'
1/
#361030000000
0!
0'
0/
#361040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#361050000000
0!
0'
0/
#361060000000
1!
1'
1/
#361070000000
0!
0'
0/
#361080000000
1!
1'
1/
#361090000000
0!
0'
0/
#361100000000
1!
1'
1/
#361110000000
0!
0'
0/
#361120000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#361130000000
0!
0'
0/
#361140000000
1!
1'
1/
#361150000000
0!
0'
0/
#361160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#361170000000
0!
0'
0/
#361180000000
1!
1'
1/
#361190000000
0!
0'
0/
#361200000000
#361210000000
1!
1'
1/
#361220000000
0!
0'
0/
#361230000000
1!
1'
1/
#361240000000
0!
1"
0'
1(
0/
10
#361250000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#361260000000
0!
0'
0/
#361270000000
1!
1'
1/
#361280000000
0!
0'
0/
#361290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#361300000000
0!
0'
0/
#361310000000
1!
1'
1/
#361320000000
0!
1"
0'
1(
0/
10
#361330000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#361340000000
0!
1$
0'
1+
0/
#361350000000
1!
1'
1/
#361360000000
0!
0'
0/
#361370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#361380000000
0!
0'
0/
#361390000000
1!
1'
1/
#361400000000
0!
0'
0/
#361410000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#361420000000
0!
0'
0/
#361430000000
1!
1'
1/
#361440000000
0!
0'
0/
#361450000000
1!
1'
1/
#361460000000
0!
0'
0/
#361470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#361480000000
0!
0'
0/
#361490000000
1!
1'
1/
#361500000000
0!
0'
0/
#361510000000
1!
1'
1/
#361520000000
0!
0'
0/
#361530000000
1!
1'
1/
#361540000000
0!
0'
0/
#361550000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#361560000000
0!
0'
0/
#361570000000
1!
1'
1/
#361580000000
0!
0'
0/
#361590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#361600000000
0!
0'
0/
#361610000000
1!
1'
1/
#361620000000
0!
0'
0/
#361630000000
#361640000000
1!
1'
1/
#361650000000
0!
0'
0/
#361660000000
1!
1'
1/
#361670000000
0!
1"
0'
1(
0/
10
#361680000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#361690000000
0!
0'
0/
#361700000000
1!
1'
1/
#361710000000
0!
0'
0/
#361720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#361730000000
0!
0'
0/
#361740000000
1!
1'
1/
#361750000000
0!
1"
0'
1(
0/
10
#361760000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#361770000000
0!
1$
0'
1+
0/
#361780000000
1!
1'
1/
#361790000000
0!
0'
0/
#361800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#361810000000
0!
0'
0/
#361820000000
1!
1'
1/
#361830000000
0!
0'
0/
#361840000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#361850000000
0!
0'
0/
#361860000000
1!
1'
1/
#361870000000
0!
0'
0/
#361880000000
1!
1'
1/
#361890000000
0!
0'
0/
#361900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#361910000000
0!
0'
0/
#361920000000
1!
1'
1/
#361930000000
0!
0'
0/
#361940000000
1!
1'
1/
#361950000000
0!
0'
0/
#361960000000
1!
1'
1/
#361970000000
0!
0'
0/
#361980000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#361990000000
0!
0'
0/
#362000000000
1!
1'
1/
#362010000000
0!
0'
0/
#362020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#362030000000
0!
0'
0/
#362040000000
1!
1'
1/
#362050000000
0!
0'
0/
#362060000000
#362070000000
1!
1'
1/
#362080000000
0!
0'
0/
#362090000000
1!
1'
1/
#362100000000
0!
1"
0'
1(
0/
10
#362110000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#362120000000
0!
0'
0/
#362130000000
1!
1'
1/
#362140000000
0!
0'
0/
#362150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#362160000000
0!
0'
0/
#362170000000
1!
1'
1/
#362180000000
0!
1"
0'
1(
0/
10
#362190000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#362200000000
0!
1$
0'
1+
0/
#362210000000
1!
1'
1/
#362220000000
0!
0'
0/
#362230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#362240000000
0!
0'
0/
#362250000000
1!
1'
1/
#362260000000
0!
0'
0/
#362270000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#362280000000
0!
0'
0/
#362290000000
1!
1'
1/
#362300000000
0!
0'
0/
#362310000000
1!
1'
1/
#362320000000
0!
0'
0/
#362330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#362340000000
0!
0'
0/
#362350000000
1!
1'
1/
#362360000000
0!
0'
0/
#362370000000
1!
1'
1/
#362380000000
0!
0'
0/
#362390000000
1!
1'
1/
#362400000000
0!
0'
0/
#362410000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#362420000000
0!
0'
0/
#362430000000
1!
1'
1/
#362440000000
0!
0'
0/
#362450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#362460000000
0!
0'
0/
#362470000000
1!
1'
1/
#362480000000
0!
0'
0/
#362490000000
#362500000000
1!
1'
1/
#362510000000
0!
0'
0/
#362520000000
1!
1'
1/
#362530000000
0!
1"
0'
1(
0/
10
#362540000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#362550000000
0!
0'
0/
#362560000000
1!
1'
1/
#362570000000
0!
0'
0/
#362580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#362590000000
0!
0'
0/
#362600000000
1!
1'
1/
#362610000000
0!
1"
0'
1(
0/
10
#362620000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#362630000000
0!
1$
0'
1+
0/
#362640000000
1!
1'
1/
#362650000000
0!
0'
0/
#362660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#362670000000
0!
0'
0/
#362680000000
1!
1'
1/
#362690000000
0!
0'
0/
#362700000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#362710000000
0!
0'
0/
#362720000000
1!
1'
1/
#362730000000
0!
0'
0/
#362740000000
1!
1'
1/
#362750000000
0!
0'
0/
#362760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#362770000000
0!
0'
0/
#362780000000
1!
1'
1/
#362790000000
0!
0'
0/
#362800000000
1!
1'
1/
#362810000000
0!
0'
0/
#362820000000
1!
1'
1/
#362830000000
0!
0'
0/
#362840000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#362850000000
0!
0'
0/
#362860000000
1!
1'
1/
#362870000000
0!
0'
0/
#362880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#362890000000
0!
0'
0/
#362900000000
1!
1'
1/
#362910000000
0!
0'
0/
#362920000000
#362930000000
1!
1'
1/
#362940000000
0!
0'
0/
#362950000000
1!
1'
1/
#362960000000
0!
1"
0'
1(
0/
10
#362970000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#362980000000
0!
0'
0/
#362990000000
1!
1'
1/
#363000000000
0!
0'
0/
#363010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#363020000000
0!
0'
0/
#363030000000
1!
1'
1/
#363040000000
0!
1"
0'
1(
0/
10
#363050000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#363060000000
0!
1$
0'
1+
0/
#363070000000
1!
1'
1/
#363080000000
0!
0'
0/
#363090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#363100000000
0!
0'
0/
#363110000000
1!
1'
1/
#363120000000
0!
0'
0/
#363130000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#363140000000
0!
0'
0/
#363150000000
1!
1'
1/
#363160000000
0!
0'
0/
#363170000000
1!
1'
1/
#363180000000
0!
0'
0/
#363190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#363200000000
0!
0'
0/
#363210000000
1!
1'
1/
#363220000000
0!
0'
0/
#363230000000
1!
1'
1/
#363240000000
0!
0'
0/
#363250000000
1!
1'
1/
#363260000000
0!
0'
0/
#363270000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#363280000000
0!
0'
0/
#363290000000
1!
1'
1/
#363300000000
0!
0'
0/
#363310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#363320000000
0!
0'
0/
#363330000000
1!
1'
1/
#363340000000
0!
0'
0/
#363350000000
#363360000000
1!
1'
1/
#363370000000
0!
0'
0/
#363380000000
1!
1'
1/
#363390000000
0!
1"
0'
1(
0/
10
#363400000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#363410000000
0!
0'
0/
#363420000000
1!
1'
1/
#363430000000
0!
0'
0/
#363440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#363450000000
0!
0'
0/
#363460000000
1!
1'
1/
#363470000000
0!
1"
0'
1(
0/
10
#363480000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#363490000000
0!
1$
0'
1+
0/
#363500000000
1!
1'
1/
#363510000000
0!
0'
0/
#363520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#363530000000
0!
0'
0/
#363540000000
1!
1'
1/
#363550000000
0!
0'
0/
#363560000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#363570000000
0!
0'
0/
#363580000000
1!
1'
1/
#363590000000
0!
0'
0/
#363600000000
1!
1'
1/
#363610000000
0!
0'
0/
#363620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#363630000000
0!
0'
0/
#363640000000
1!
1'
1/
#363650000000
0!
0'
0/
#363660000000
1!
1'
1/
#363670000000
0!
0'
0/
#363680000000
1!
1'
1/
#363690000000
0!
0'
0/
#363700000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#363710000000
0!
0'
0/
#363720000000
1!
1'
1/
#363730000000
0!
0'
0/
#363740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#363750000000
0!
0'
0/
#363760000000
1!
1'
1/
#363770000000
0!
0'
0/
#363780000000
#363790000000
1!
1'
1/
#363800000000
0!
0'
0/
#363810000000
1!
1'
1/
#363820000000
0!
1"
0'
1(
0/
10
#363830000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#363840000000
0!
0'
0/
#363850000000
1!
1'
1/
#363860000000
0!
0'
0/
#363870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#363880000000
0!
0'
0/
#363890000000
1!
1'
1/
#363900000000
0!
1"
0'
1(
0/
10
#363910000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#363920000000
0!
1$
0'
1+
0/
#363930000000
1!
1'
1/
#363940000000
0!
0'
0/
#363950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#363960000000
0!
0'
0/
#363970000000
1!
1'
1/
#363980000000
0!
0'
0/
#363990000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#364000000000
0!
0'
0/
#364010000000
1!
1'
1/
#364020000000
0!
0'
0/
#364030000000
1!
1'
1/
#364040000000
0!
0'
0/
#364050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#364060000000
0!
0'
0/
#364070000000
1!
1'
1/
#364080000000
0!
0'
0/
#364090000000
1!
1'
1/
#364100000000
0!
0'
0/
#364110000000
1!
1'
1/
#364120000000
0!
0'
0/
#364130000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#364140000000
0!
0'
0/
#364150000000
1!
1'
1/
#364160000000
0!
0'
0/
#364170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#364180000000
0!
0'
0/
#364190000000
1!
1'
1/
#364200000000
0!
0'
0/
#364210000000
#364220000000
1!
1'
1/
#364230000000
0!
0'
0/
#364240000000
1!
1'
1/
#364250000000
0!
1"
0'
1(
0/
10
#364260000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#364270000000
0!
0'
0/
#364280000000
1!
1'
1/
#364290000000
0!
0'
0/
#364300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#364310000000
0!
0'
0/
#364320000000
1!
1'
1/
#364330000000
0!
1"
0'
1(
0/
10
#364340000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#364350000000
0!
1$
0'
1+
0/
#364360000000
1!
1'
1/
#364370000000
0!
0'
0/
#364380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#364390000000
0!
0'
0/
#364400000000
1!
1'
1/
#364410000000
0!
0'
0/
#364420000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#364430000000
0!
0'
0/
#364440000000
1!
1'
1/
#364450000000
0!
0'
0/
#364460000000
1!
1'
1/
#364470000000
0!
0'
0/
#364480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#364490000000
0!
0'
0/
#364500000000
1!
1'
1/
#364510000000
0!
0'
0/
#364520000000
1!
1'
1/
#364530000000
0!
0'
0/
#364540000000
1!
1'
1/
#364550000000
0!
0'
0/
#364560000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#364570000000
0!
0'
0/
#364580000000
1!
1'
1/
#364590000000
0!
0'
0/
#364600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#364610000000
0!
0'
0/
#364620000000
1!
1'
1/
#364630000000
0!
0'
0/
#364640000000
#364650000000
1!
1'
1/
#364660000000
0!
0'
0/
#364670000000
1!
1'
1/
#364680000000
0!
1"
0'
1(
0/
10
#364690000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#364700000000
0!
0'
0/
#364710000000
1!
1'
1/
#364720000000
0!
0'
0/
#364730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#364740000000
0!
0'
0/
#364750000000
1!
1'
1/
#364760000000
0!
1"
0'
1(
0/
10
#364770000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#364780000000
0!
1$
0'
1+
0/
#364790000000
1!
1'
1/
#364800000000
0!
0'
0/
#364810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#364820000000
0!
0'
0/
#364830000000
1!
1'
1/
#364840000000
0!
0'
0/
#364850000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#364860000000
0!
0'
0/
#364870000000
1!
1'
1/
#364880000000
0!
0'
0/
#364890000000
1!
1'
1/
#364900000000
0!
0'
0/
#364910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#364920000000
0!
0'
0/
#364930000000
1!
1'
1/
#364940000000
0!
0'
0/
#364950000000
1!
1'
1/
#364960000000
0!
0'
0/
#364970000000
1!
1'
1/
#364980000000
0!
0'
0/
#364990000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#365000000000
0!
0'
0/
#365010000000
1!
1'
1/
#365020000000
0!
0'
0/
#365030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#365040000000
0!
0'
0/
#365050000000
1!
1'
1/
#365060000000
0!
0'
0/
#365070000000
#365080000000
1!
1'
1/
#365090000000
0!
0'
0/
#365100000000
1!
1'
1/
#365110000000
0!
1"
0'
1(
0/
10
#365120000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#365130000000
0!
0'
0/
#365140000000
1!
1'
1/
#365150000000
0!
0'
0/
#365160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#365170000000
0!
0'
0/
#365180000000
1!
1'
1/
#365190000000
0!
1"
0'
1(
0/
10
#365200000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#365210000000
0!
1$
0'
1+
0/
#365220000000
1!
1'
1/
#365230000000
0!
0'
0/
#365240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#365250000000
0!
0'
0/
#365260000000
1!
1'
1/
#365270000000
0!
0'
0/
#365280000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#365290000000
0!
0'
0/
#365300000000
1!
1'
1/
#365310000000
0!
0'
0/
#365320000000
1!
1'
1/
#365330000000
0!
0'
0/
#365340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#365350000000
0!
0'
0/
#365360000000
1!
1'
1/
#365370000000
0!
0'
0/
#365380000000
1!
1'
1/
#365390000000
0!
0'
0/
#365400000000
1!
1'
1/
#365410000000
0!
0'
0/
#365420000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#365430000000
0!
0'
0/
#365440000000
1!
1'
1/
#365450000000
0!
0'
0/
#365460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#365470000000
0!
0'
0/
#365480000000
1!
1'
1/
#365490000000
0!
0'
0/
#365500000000
#365510000000
1!
1'
1/
#365520000000
0!
0'
0/
#365530000000
1!
1'
1/
#365540000000
0!
1"
0'
1(
0/
10
#365550000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#365560000000
0!
0'
0/
#365570000000
1!
1'
1/
#365580000000
0!
0'
0/
#365590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#365600000000
0!
0'
0/
#365610000000
1!
1'
1/
#365620000000
0!
1"
0'
1(
0/
10
#365630000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#365640000000
0!
1$
0'
1+
0/
#365650000000
1!
1'
1/
#365660000000
0!
0'
0/
#365670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#365680000000
0!
0'
0/
#365690000000
1!
1'
1/
#365700000000
0!
0'
0/
#365710000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#365720000000
0!
0'
0/
#365730000000
1!
1'
1/
#365740000000
0!
0'
0/
#365750000000
1!
1'
1/
#365760000000
0!
0'
0/
#365770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#365780000000
0!
0'
0/
#365790000000
1!
1'
1/
#365800000000
0!
0'
0/
#365810000000
1!
1'
1/
#365820000000
0!
0'
0/
#365830000000
1!
1'
1/
#365840000000
0!
0'
0/
#365850000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#365860000000
0!
0'
0/
#365870000000
1!
1'
1/
#365880000000
0!
0'
0/
#365890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#365900000000
0!
0'
0/
#365910000000
1!
1'
1/
#365920000000
0!
0'
0/
#365930000000
#365940000000
1!
1'
1/
#365950000000
0!
0'
0/
#365960000000
1!
1'
1/
#365970000000
0!
1"
0'
1(
0/
10
#365980000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#365990000000
0!
0'
0/
#366000000000
1!
1'
1/
#366010000000
0!
0'
0/
#366020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#366030000000
0!
0'
0/
#366040000000
1!
1'
1/
#366050000000
0!
1"
0'
1(
0/
10
#366060000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#366070000000
0!
1$
0'
1+
0/
#366080000000
1!
1'
1/
#366090000000
0!
0'
0/
#366100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#366110000000
0!
0'
0/
#366120000000
1!
1'
1/
#366130000000
0!
0'
0/
#366140000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#366150000000
0!
0'
0/
#366160000000
1!
1'
1/
#366170000000
0!
0'
0/
#366180000000
1!
1'
1/
#366190000000
0!
0'
0/
#366200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#366210000000
0!
0'
0/
#366220000000
1!
1'
1/
#366230000000
0!
0'
0/
#366240000000
1!
1'
1/
#366250000000
0!
0'
0/
#366260000000
1!
1'
1/
#366270000000
0!
0'
0/
#366280000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#366290000000
0!
0'
0/
#366300000000
1!
1'
1/
#366310000000
0!
0'
0/
#366320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#366330000000
0!
0'
0/
#366340000000
1!
1'
1/
#366350000000
0!
0'
0/
#366360000000
#366370000000
1!
1'
1/
#366380000000
0!
0'
0/
#366390000000
1!
1'
1/
#366400000000
0!
1"
0'
1(
0/
10
#366410000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#366420000000
0!
0'
0/
#366430000000
1!
1'
1/
#366440000000
0!
0'
0/
#366450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#366460000000
0!
0'
0/
#366470000000
1!
1'
1/
#366480000000
0!
1"
0'
1(
0/
10
#366490000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#366500000000
0!
1$
0'
1+
0/
#366510000000
1!
1'
1/
#366520000000
0!
0'
0/
#366530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#366540000000
0!
0'
0/
#366550000000
1!
1'
1/
#366560000000
0!
0'
0/
#366570000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#366580000000
0!
0'
0/
#366590000000
1!
1'
1/
#366600000000
0!
0'
0/
#366610000000
1!
1'
1/
#366620000000
0!
0'
0/
#366630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#366640000000
0!
0'
0/
#366650000000
1!
1'
1/
#366660000000
0!
0'
0/
#366670000000
1!
1'
1/
#366680000000
0!
0'
0/
#366690000000
1!
1'
1/
#366700000000
0!
0'
0/
#366710000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#366720000000
0!
0'
0/
#366730000000
1!
1'
1/
#366740000000
0!
0'
0/
#366750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#366760000000
0!
0'
0/
#366770000000
1!
1'
1/
#366780000000
0!
0'
0/
#366790000000
#366800000000
1!
1'
1/
#366810000000
0!
0'
0/
#366820000000
1!
1'
1/
#366830000000
0!
1"
0'
1(
0/
10
#366840000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#366850000000
0!
0'
0/
#366860000000
1!
1'
1/
#366870000000
0!
0'
0/
#366880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#366890000000
0!
0'
0/
#366900000000
1!
1'
1/
#366910000000
0!
1"
0'
1(
0/
10
#366920000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#366930000000
0!
1$
0'
1+
0/
#366940000000
1!
1'
1/
#366950000000
0!
0'
0/
#366960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#366970000000
0!
0'
0/
#366980000000
1!
1'
1/
#366990000000
0!
0'
0/
#367000000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#367010000000
0!
0'
0/
#367020000000
1!
1'
1/
#367030000000
0!
0'
0/
#367040000000
1!
1'
1/
#367050000000
0!
0'
0/
#367060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#367070000000
0!
0'
0/
#367080000000
1!
1'
1/
#367090000000
0!
0'
0/
#367100000000
1!
1'
1/
#367110000000
0!
0'
0/
#367120000000
1!
1'
1/
#367130000000
0!
0'
0/
#367140000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#367150000000
0!
0'
0/
#367160000000
1!
1'
1/
#367170000000
0!
0'
0/
#367180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#367190000000
0!
0'
0/
#367200000000
1!
1'
1/
#367210000000
0!
0'
0/
#367220000000
#367230000000
1!
1'
1/
#367240000000
0!
0'
0/
#367250000000
1!
1'
1/
#367260000000
0!
1"
0'
1(
0/
10
#367270000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#367280000000
0!
0'
0/
#367290000000
1!
1'
1/
#367300000000
0!
0'
0/
#367310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#367320000000
0!
0'
0/
#367330000000
1!
1'
1/
#367340000000
0!
1"
0'
1(
0/
10
#367350000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#367360000000
0!
1$
0'
1+
0/
#367370000000
1!
1'
1/
#367380000000
0!
0'
0/
#367390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#367400000000
0!
0'
0/
#367410000000
1!
1'
1/
#367420000000
0!
0'
0/
#367430000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#367440000000
0!
0'
0/
#367450000000
1!
1'
1/
#367460000000
0!
0'
0/
#367470000000
1!
1'
1/
#367480000000
0!
0'
0/
#367490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#367500000000
0!
0'
0/
#367510000000
1!
1'
1/
#367520000000
0!
0'
0/
#367530000000
1!
1'
1/
#367540000000
0!
0'
0/
#367550000000
1!
1'
1/
#367560000000
0!
0'
0/
#367570000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#367580000000
0!
0'
0/
#367590000000
1!
1'
1/
#367600000000
0!
0'
0/
#367610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#367620000000
0!
0'
0/
#367630000000
1!
1'
1/
#367640000000
0!
0'
0/
#367650000000
#367660000000
1!
1'
1/
#367670000000
0!
0'
0/
#367680000000
1!
1'
1/
#367690000000
0!
1"
0'
1(
0/
10
#367700000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#367710000000
0!
0'
0/
#367720000000
1!
1'
1/
#367730000000
0!
0'
0/
#367740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#367750000000
0!
0'
0/
#367760000000
1!
1'
1/
#367770000000
0!
1"
0'
1(
0/
10
#367780000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#367790000000
0!
1$
0'
1+
0/
#367800000000
1!
1'
1/
#367810000000
0!
0'
0/
#367820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#367830000000
0!
0'
0/
#367840000000
1!
1'
1/
#367850000000
0!
0'
0/
#367860000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#367870000000
0!
0'
0/
#367880000000
1!
1'
1/
#367890000000
0!
0'
0/
#367900000000
1!
1'
1/
#367910000000
0!
0'
0/
#367920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#367930000000
0!
0'
0/
#367940000000
1!
1'
1/
#367950000000
0!
0'
0/
#367960000000
1!
1'
1/
#367970000000
0!
0'
0/
#367980000000
1!
1'
1/
#367990000000
0!
0'
0/
#368000000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#368010000000
0!
0'
0/
#368020000000
1!
1'
1/
#368030000000
0!
0'
0/
#368040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#368050000000
0!
0'
0/
#368060000000
1!
1'
1/
#368070000000
0!
0'
0/
#368080000000
#368090000000
1!
1'
1/
#368100000000
0!
0'
0/
#368110000000
1!
1'
1/
#368120000000
0!
1"
0'
1(
0/
10
#368130000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#368140000000
0!
0'
0/
#368150000000
1!
1'
1/
#368160000000
0!
0'
0/
#368170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#368180000000
0!
0'
0/
#368190000000
1!
1'
1/
#368200000000
0!
1"
0'
1(
0/
10
#368210000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#368220000000
0!
1$
0'
1+
0/
#368230000000
1!
1'
1/
#368240000000
0!
0'
0/
#368250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#368260000000
0!
0'
0/
#368270000000
1!
1'
1/
#368280000000
0!
0'
0/
#368290000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#368300000000
0!
0'
0/
#368310000000
1!
1'
1/
#368320000000
0!
0'
0/
#368330000000
1!
1'
1/
#368340000000
0!
0'
0/
#368350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#368360000000
0!
0'
0/
#368370000000
1!
1'
1/
#368380000000
0!
0'
0/
#368390000000
1!
1'
1/
#368400000000
0!
0'
0/
#368410000000
1!
1'
1/
#368420000000
0!
0'
0/
#368430000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#368440000000
0!
0'
0/
#368450000000
1!
1'
1/
#368460000000
0!
0'
0/
#368470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#368480000000
0!
0'
0/
#368490000000
1!
1'
1/
#368500000000
0!
0'
0/
#368510000000
#368520000000
1!
1'
1/
#368530000000
0!
0'
0/
#368540000000
1!
1'
1/
#368550000000
0!
1"
0'
1(
0/
10
#368560000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#368570000000
0!
0'
0/
#368580000000
1!
1'
1/
#368590000000
0!
0'
0/
#368600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#368610000000
0!
0'
0/
#368620000000
1!
1'
1/
#368630000000
0!
1"
0'
1(
0/
10
#368640000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#368650000000
0!
1$
0'
1+
0/
#368660000000
1!
1'
1/
#368670000000
0!
0'
0/
#368680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#368690000000
0!
0'
0/
#368700000000
1!
1'
1/
#368710000000
0!
0'
0/
#368720000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#368730000000
0!
0'
0/
#368740000000
1!
1'
1/
#368750000000
0!
0'
0/
#368760000000
1!
1'
1/
#368770000000
0!
0'
0/
#368780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#368790000000
0!
0'
0/
#368800000000
1!
1'
1/
#368810000000
0!
0'
0/
#368820000000
1!
1'
1/
#368830000000
0!
0'
0/
#368840000000
1!
1'
1/
#368850000000
0!
0'
0/
#368860000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#368870000000
0!
0'
0/
#368880000000
1!
1'
1/
#368890000000
0!
0'
0/
#368900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#368910000000
0!
0'
0/
#368920000000
1!
1'
1/
#368930000000
0!
0'
0/
#368940000000
#368950000000
1!
1'
1/
#368960000000
0!
0'
0/
#368970000000
1!
1'
1/
#368980000000
0!
1"
0'
1(
0/
10
#368990000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#369000000000
0!
0'
0/
#369010000000
1!
1'
1/
#369020000000
0!
0'
0/
#369030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#369040000000
0!
0'
0/
#369050000000
1!
1'
1/
#369060000000
0!
1"
0'
1(
0/
10
#369070000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#369080000000
0!
1$
0'
1+
0/
#369090000000
1!
1'
1/
#369100000000
0!
0'
0/
#369110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#369120000000
0!
0'
0/
#369130000000
1!
1'
1/
#369140000000
0!
0'
0/
#369150000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#369160000000
0!
0'
0/
#369170000000
1!
1'
1/
#369180000000
0!
0'
0/
#369190000000
1!
1'
1/
#369200000000
0!
0'
0/
#369210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#369220000000
0!
0'
0/
#369230000000
1!
1'
1/
#369240000000
0!
0'
0/
#369250000000
1!
1'
1/
#369260000000
0!
0'
0/
#369270000000
1!
1'
1/
#369280000000
0!
0'
0/
#369290000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#369300000000
0!
0'
0/
#369310000000
1!
1'
1/
#369320000000
0!
0'
0/
#369330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#369340000000
0!
0'
0/
#369350000000
1!
1'
1/
#369360000000
0!
0'
0/
#369370000000
#369380000000
1!
1'
1/
#369390000000
0!
0'
0/
#369400000000
1!
1'
1/
#369410000000
0!
1"
0'
1(
0/
10
#369420000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#369430000000
0!
0'
0/
#369440000000
1!
1'
1/
#369450000000
0!
0'
0/
#369460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#369470000000
0!
0'
0/
#369480000000
1!
1'
1/
#369490000000
0!
1"
0'
1(
0/
10
#369500000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#369510000000
0!
1$
0'
1+
0/
#369520000000
1!
1'
1/
#369530000000
0!
0'
0/
#369540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#369550000000
0!
0'
0/
#369560000000
1!
1'
1/
#369570000000
0!
0'
0/
#369580000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#369590000000
0!
0'
0/
#369600000000
1!
1'
1/
#369610000000
0!
0'
0/
#369620000000
1!
1'
1/
#369630000000
0!
0'
0/
#369640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#369650000000
0!
0'
0/
#369660000000
1!
1'
1/
#369670000000
0!
0'
0/
#369680000000
1!
1'
1/
#369690000000
0!
0'
0/
#369700000000
1!
1'
1/
#369710000000
0!
0'
0/
#369720000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#369730000000
0!
0'
0/
#369740000000
1!
1'
1/
#369750000000
0!
0'
0/
#369760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#369770000000
0!
0'
0/
#369780000000
1!
1'
1/
#369790000000
0!
0'
0/
#369800000000
#369810000000
1!
1'
1/
#369820000000
0!
0'
0/
#369830000000
1!
1'
1/
#369840000000
0!
1"
0'
1(
0/
10
#369850000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#369860000000
0!
0'
0/
#369870000000
1!
1'
1/
#369880000000
0!
0'
0/
#369890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#369900000000
0!
0'
0/
#369910000000
1!
1'
1/
#369920000000
0!
1"
0'
1(
0/
10
#369930000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#369940000000
0!
1$
0'
1+
0/
#369950000000
1!
1'
1/
#369960000000
0!
0'
0/
#369970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#369980000000
0!
0'
0/
#369990000000
1!
1'
1/
#370000000000
0!
0'
0/
#370010000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#370020000000
0!
0'
0/
#370030000000
1!
1'
1/
#370040000000
0!
0'
0/
#370050000000
1!
1'
1/
#370060000000
0!
0'
0/
#370070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#370080000000
0!
0'
0/
#370090000000
1!
1'
1/
#370100000000
0!
0'
0/
#370110000000
1!
1'
1/
#370120000000
0!
0'
0/
#370130000000
1!
1'
1/
#370140000000
0!
0'
0/
#370150000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#370160000000
0!
0'
0/
#370170000000
1!
1'
1/
#370180000000
0!
0'
0/
#370190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#370200000000
0!
0'
0/
#370210000000
1!
1'
1/
#370220000000
0!
0'
0/
#370230000000
#370240000000
1!
1'
1/
#370250000000
0!
0'
0/
#370260000000
1!
1'
1/
#370270000000
0!
1"
0'
1(
0/
10
#370280000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#370290000000
0!
0'
0/
#370300000000
1!
1'
1/
#370310000000
0!
0'
0/
#370320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#370330000000
0!
0'
0/
#370340000000
1!
1'
1/
#370350000000
0!
1"
0'
1(
0/
10
#370360000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#370370000000
0!
1$
0'
1+
0/
#370380000000
1!
1'
1/
#370390000000
0!
0'
0/
#370400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#370410000000
0!
0'
0/
#370420000000
1!
1'
1/
#370430000000
0!
0'
0/
#370440000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#370450000000
0!
0'
0/
#370460000000
1!
1'
1/
#370470000000
0!
0'
0/
#370480000000
1!
1'
1/
#370490000000
0!
0'
0/
#370500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#370510000000
0!
0'
0/
#370520000000
1!
1'
1/
#370530000000
0!
0'
0/
#370540000000
1!
1'
1/
#370550000000
0!
0'
0/
#370560000000
1!
1'
1/
#370570000000
0!
0'
0/
#370580000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#370590000000
0!
0'
0/
#370600000000
1!
1'
1/
#370610000000
0!
0'
0/
#370620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#370630000000
0!
0'
0/
#370640000000
1!
1'
1/
#370650000000
0!
0'
0/
#370660000000
#370670000000
1!
1'
1/
#370680000000
0!
0'
0/
#370690000000
1!
1'
1/
#370700000000
0!
1"
0'
1(
0/
10
#370710000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#370720000000
0!
0'
0/
#370730000000
1!
1'
1/
#370740000000
0!
0'
0/
#370750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#370760000000
0!
0'
0/
#370770000000
1!
1'
1/
#370780000000
0!
1"
0'
1(
0/
10
#370790000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#370800000000
0!
1$
0'
1+
0/
#370810000000
1!
1'
1/
#370820000000
0!
0'
0/
#370830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#370840000000
0!
0'
0/
#370850000000
1!
1'
1/
#370860000000
0!
0'
0/
#370870000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#370880000000
0!
0'
0/
#370890000000
1!
1'
1/
#370900000000
0!
0'
0/
#370910000000
1!
1'
1/
#370920000000
0!
0'
0/
#370930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#370940000000
0!
0'
0/
#370950000000
1!
1'
1/
#370960000000
0!
0'
0/
#370970000000
1!
1'
1/
#370980000000
0!
0'
0/
#370990000000
1!
1'
1/
#371000000000
0!
0'
0/
#371010000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#371020000000
0!
0'
0/
#371030000000
1!
1'
1/
#371040000000
0!
0'
0/
#371050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#371060000000
0!
0'
0/
#371070000000
1!
1'
1/
#371080000000
0!
0'
0/
#371090000000
#371100000000
1!
1'
1/
#371110000000
0!
0'
0/
#371120000000
1!
1'
1/
#371130000000
0!
1"
0'
1(
0/
10
#371140000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#371150000000
0!
0'
0/
#371160000000
1!
1'
1/
#371170000000
0!
0'
0/
#371180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#371190000000
0!
0'
0/
#371200000000
1!
1'
1/
#371210000000
0!
1"
0'
1(
0/
10
#371220000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#371230000000
0!
1$
0'
1+
0/
#371240000000
1!
1'
1/
#371250000000
0!
0'
0/
#371260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#371270000000
0!
0'
0/
#371280000000
1!
1'
1/
#371290000000
0!
0'
0/
#371300000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#371310000000
0!
0'
0/
#371320000000
1!
1'
1/
#371330000000
0!
0'
0/
#371340000000
1!
1'
1/
#371350000000
0!
0'
0/
#371360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#371370000000
0!
0'
0/
#371380000000
1!
1'
1/
#371390000000
0!
0'
0/
#371400000000
1!
1'
1/
#371410000000
0!
0'
0/
#371420000000
1!
1'
1/
#371430000000
0!
0'
0/
#371440000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#371450000000
0!
0'
0/
#371460000000
1!
1'
1/
#371470000000
0!
0'
0/
#371480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#371490000000
0!
0'
0/
#371500000000
1!
1'
1/
#371510000000
0!
0'
0/
#371520000000
#371530000000
1!
1'
1/
#371540000000
0!
0'
0/
#371550000000
1!
1'
1/
#371560000000
0!
1"
0'
1(
0/
10
#371570000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#371580000000
0!
0'
0/
#371590000000
1!
1'
1/
#371600000000
0!
0'
0/
#371610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#371620000000
0!
0'
0/
#371630000000
1!
1'
1/
#371640000000
0!
1"
0'
1(
0/
10
#371650000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#371660000000
0!
1$
0'
1+
0/
#371670000000
1!
1'
1/
#371680000000
0!
0'
0/
#371690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#371700000000
0!
0'
0/
#371710000000
1!
1'
1/
#371720000000
0!
0'
0/
#371730000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#371740000000
0!
0'
0/
#371750000000
1!
1'
1/
#371760000000
0!
0'
0/
#371770000000
1!
1'
1/
#371780000000
0!
0'
0/
#371790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#371800000000
0!
0'
0/
#371810000000
1!
1'
1/
#371820000000
0!
0'
0/
#371830000000
1!
1'
1/
#371840000000
0!
0'
0/
#371850000000
1!
1'
1/
#371860000000
0!
0'
0/
#371870000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#371880000000
0!
0'
0/
#371890000000
1!
1'
1/
#371900000000
0!
0'
0/
#371910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#371920000000
0!
0'
0/
#371930000000
1!
1'
1/
#371940000000
0!
0'
0/
#371950000000
#371960000000
1!
1'
1/
#371970000000
0!
0'
0/
#371980000000
1!
1'
1/
#371990000000
0!
1"
0'
1(
0/
10
#372000000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#372010000000
0!
0'
0/
#372020000000
1!
1'
1/
#372030000000
0!
0'
0/
#372040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#372050000000
0!
0'
0/
#372060000000
1!
1'
1/
#372070000000
0!
1"
0'
1(
0/
10
#372080000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#372090000000
0!
1$
0'
1+
0/
#372100000000
1!
1'
1/
#372110000000
0!
0'
0/
#372120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#372130000000
0!
0'
0/
#372140000000
1!
1'
1/
#372150000000
0!
0'
0/
#372160000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#372170000000
0!
0'
0/
#372180000000
1!
1'
1/
#372190000000
0!
0'
0/
#372200000000
1!
1'
1/
#372210000000
0!
0'
0/
#372220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#372230000000
0!
0'
0/
#372240000000
1!
1'
1/
#372250000000
0!
0'
0/
#372260000000
1!
1'
1/
#372270000000
0!
0'
0/
#372280000000
1!
1'
1/
#372290000000
0!
0'
0/
#372300000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#372310000000
0!
0'
0/
#372320000000
1!
1'
1/
#372330000000
0!
0'
0/
#372340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#372350000000
0!
0'
0/
#372360000000
1!
1'
1/
#372370000000
0!
0'
0/
#372380000000
#372390000000
1!
1'
1/
#372400000000
0!
0'
0/
#372410000000
1!
1'
1/
#372420000000
0!
1"
0'
1(
0/
10
#372430000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#372440000000
0!
0'
0/
#372450000000
1!
1'
1/
#372460000000
0!
0'
0/
#372470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#372480000000
0!
0'
0/
#372490000000
1!
1'
1/
#372500000000
0!
1"
0'
1(
0/
10
#372510000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#372520000000
0!
1$
0'
1+
0/
#372530000000
1!
1'
1/
#372540000000
0!
0'
0/
#372550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#372560000000
0!
0'
0/
#372570000000
1!
1'
1/
#372580000000
0!
0'
0/
#372590000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#372600000000
0!
0'
0/
#372610000000
1!
1'
1/
#372620000000
0!
0'
0/
#372630000000
1!
1'
1/
#372640000000
0!
0'
0/
#372650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#372660000000
0!
0'
0/
#372670000000
1!
1'
1/
#372680000000
0!
0'
0/
#372690000000
1!
1'
1/
#372700000000
0!
0'
0/
#372710000000
1!
1'
1/
#372720000000
0!
0'
0/
#372730000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#372740000000
0!
0'
0/
#372750000000
1!
1'
1/
#372760000000
0!
0'
0/
#372770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#372780000000
0!
0'
0/
#372790000000
1!
1'
1/
#372800000000
0!
0'
0/
#372810000000
#372820000000
1!
1'
1/
#372830000000
0!
0'
0/
#372840000000
1!
1'
1/
#372850000000
0!
1"
0'
1(
0/
10
#372860000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#372870000000
0!
0'
0/
#372880000000
1!
1'
1/
#372890000000
0!
0'
0/
#372900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#372910000000
0!
0'
0/
#372920000000
1!
1'
1/
#372930000000
0!
1"
0'
1(
0/
10
#372940000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#372950000000
0!
1$
0'
1+
0/
#372960000000
1!
1'
1/
#372970000000
0!
0'
0/
#372980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#372990000000
0!
0'
0/
#373000000000
1!
1'
1/
#373010000000
0!
0'
0/
#373020000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#373030000000
0!
0'
0/
#373040000000
1!
1'
1/
#373050000000
0!
0'
0/
#373060000000
1!
1'
1/
#373070000000
0!
0'
0/
#373080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#373090000000
0!
0'
0/
#373100000000
1!
1'
1/
#373110000000
0!
0'
0/
#373120000000
1!
1'
1/
#373130000000
0!
0'
0/
#373140000000
1!
1'
1/
#373150000000
0!
0'
0/
#373160000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#373170000000
0!
0'
0/
#373180000000
1!
1'
1/
#373190000000
0!
0'
0/
#373200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#373210000000
0!
0'
0/
#373220000000
1!
1'
1/
#373230000000
0!
0'
0/
#373240000000
#373250000000
1!
1'
1/
#373260000000
0!
0'
0/
#373270000000
1!
1'
1/
#373280000000
0!
1"
0'
1(
0/
10
#373290000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#373300000000
0!
0'
0/
#373310000000
1!
1'
1/
#373320000000
0!
0'
0/
#373330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#373340000000
0!
0'
0/
#373350000000
1!
1'
1/
#373360000000
0!
1"
0'
1(
0/
10
#373370000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#373380000000
0!
1$
0'
1+
0/
#373390000000
1!
1'
1/
#373400000000
0!
0'
0/
#373410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#373420000000
0!
0'
0/
#373430000000
1!
1'
1/
#373440000000
0!
0'
0/
#373450000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#373460000000
0!
0'
0/
#373470000000
1!
1'
1/
#373480000000
0!
0'
0/
#373490000000
1!
1'
1/
#373500000000
0!
0'
0/
#373510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#373520000000
0!
0'
0/
#373530000000
1!
1'
1/
#373540000000
0!
0'
0/
#373550000000
1!
1'
1/
#373560000000
0!
0'
0/
#373570000000
1!
1'
1/
#373580000000
0!
0'
0/
#373590000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#373600000000
0!
0'
0/
#373610000000
1!
1'
1/
#373620000000
0!
0'
0/
#373630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#373640000000
0!
0'
0/
#373650000000
1!
1'
1/
#373660000000
0!
0'
0/
#373670000000
#373680000000
1!
1'
1/
#373690000000
0!
0'
0/
#373700000000
1!
1'
1/
#373710000000
0!
1"
0'
1(
0/
10
#373720000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#373730000000
0!
0'
0/
#373740000000
1!
1'
1/
#373750000000
0!
0'
0/
#373760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#373770000000
0!
0'
0/
#373780000000
1!
1'
1/
#373790000000
0!
1"
0'
1(
0/
10
#373800000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#373810000000
0!
1$
0'
1+
0/
#373820000000
1!
1'
1/
#373830000000
0!
0'
0/
#373840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#373850000000
0!
0'
0/
#373860000000
1!
1'
1/
#373870000000
0!
0'
0/
#373880000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#373890000000
0!
0'
0/
#373900000000
1!
1'
1/
#373910000000
0!
0'
0/
#373920000000
1!
1'
1/
#373930000000
0!
0'
0/
#373940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#373950000000
0!
0'
0/
#373960000000
1!
1'
1/
#373970000000
0!
0'
0/
#373980000000
1!
1'
1/
#373990000000
0!
0'
0/
#374000000000
1!
1'
1/
#374010000000
0!
0'
0/
#374020000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#374030000000
0!
0'
0/
#374040000000
1!
1'
1/
#374050000000
0!
0'
0/
#374060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#374070000000
0!
0'
0/
#374080000000
1!
1'
1/
#374090000000
0!
0'
0/
#374100000000
#374110000000
1!
1'
1/
#374120000000
0!
0'
0/
#374130000000
1!
1'
1/
#374140000000
0!
1"
0'
1(
0/
10
#374150000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#374160000000
0!
0'
0/
#374170000000
1!
1'
1/
#374180000000
0!
0'
0/
#374190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#374200000000
0!
0'
0/
#374210000000
1!
1'
1/
#374220000000
0!
1"
0'
1(
0/
10
#374230000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#374240000000
0!
1$
0'
1+
0/
#374250000000
1!
1'
1/
#374260000000
0!
0'
0/
#374270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#374280000000
0!
0'
0/
#374290000000
1!
1'
1/
#374300000000
0!
0'
0/
#374310000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#374320000000
0!
0'
0/
#374330000000
1!
1'
1/
#374340000000
0!
0'
0/
#374350000000
1!
1'
1/
#374360000000
0!
0'
0/
#374370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#374380000000
0!
0'
0/
#374390000000
1!
1'
1/
#374400000000
0!
0'
0/
#374410000000
1!
1'
1/
#374420000000
0!
0'
0/
#374430000000
1!
1'
1/
#374440000000
0!
0'
0/
#374450000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#374460000000
0!
0'
0/
#374470000000
1!
1'
1/
#374480000000
0!
0'
0/
#374490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#374500000000
0!
0'
0/
#374510000000
1!
1'
1/
#374520000000
0!
0'
0/
#374530000000
#374540000000
1!
1'
1/
#374550000000
0!
0'
0/
#374560000000
1!
1'
1/
#374570000000
0!
1"
0'
1(
0/
10
#374580000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#374590000000
0!
0'
0/
#374600000000
1!
1'
1/
#374610000000
0!
0'
0/
#374620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#374630000000
0!
0'
0/
#374640000000
1!
1'
1/
#374650000000
0!
1"
0'
1(
0/
10
#374660000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#374670000000
0!
1$
0'
1+
0/
#374680000000
1!
1'
1/
#374690000000
0!
0'
0/
#374700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#374710000000
0!
0'
0/
#374720000000
1!
1'
1/
#374730000000
0!
0'
0/
#374740000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#374750000000
0!
0'
0/
#374760000000
1!
1'
1/
#374770000000
0!
0'
0/
#374780000000
1!
1'
1/
#374790000000
0!
0'
0/
#374800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#374810000000
0!
0'
0/
#374820000000
1!
1'
1/
#374830000000
0!
0'
0/
#374840000000
1!
1'
1/
#374850000000
0!
0'
0/
#374860000000
1!
1'
1/
#374870000000
0!
0'
0/
#374880000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#374890000000
0!
0'
0/
#374900000000
1!
1'
1/
#374910000000
0!
0'
0/
#374920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#374930000000
0!
0'
0/
#374940000000
1!
1'
1/
#374950000000
0!
0'
0/
#374960000000
#374970000000
1!
1'
1/
#374980000000
0!
0'
0/
#374990000000
1!
1'
1/
#375000000000
0!
1"
0'
1(
0/
10
#375010000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#375020000000
0!
0'
0/
#375030000000
1!
1'
1/
#375040000000
0!
0'
0/
#375050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#375060000000
0!
0'
0/
#375070000000
1!
1'
1/
#375080000000
0!
1"
0'
1(
0/
10
#375090000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#375100000000
0!
1$
0'
1+
0/
#375110000000
1!
1'
1/
#375120000000
0!
0'
0/
#375130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#375140000000
0!
0'
0/
#375150000000
1!
1'
1/
#375160000000
0!
0'
0/
#375170000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#375180000000
0!
0'
0/
#375190000000
1!
1'
1/
#375200000000
0!
0'
0/
#375210000000
1!
1'
1/
#375220000000
0!
0'
0/
#375230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#375240000000
0!
0'
0/
#375250000000
1!
1'
1/
#375260000000
0!
0'
0/
#375270000000
1!
1'
1/
#375280000000
0!
0'
0/
#375290000000
1!
1'
1/
#375300000000
0!
0'
0/
#375310000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#375320000000
0!
0'
0/
#375330000000
1!
1'
1/
#375340000000
0!
0'
0/
#375350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#375360000000
0!
0'
0/
#375370000000
1!
1'
1/
#375380000000
0!
0'
0/
#375390000000
#375400000000
1!
1'
1/
#375410000000
0!
0'
0/
#375420000000
1!
1'
1/
#375430000000
0!
1"
0'
1(
0/
10
#375440000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#375450000000
0!
0'
0/
#375460000000
1!
1'
1/
#375470000000
0!
0'
0/
#375480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#375490000000
0!
0'
0/
#375500000000
1!
1'
1/
#375510000000
0!
1"
0'
1(
0/
10
#375520000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#375530000000
0!
1$
0'
1+
0/
#375540000000
1!
1'
1/
#375550000000
0!
0'
0/
#375560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#375570000000
0!
0'
0/
#375580000000
1!
1'
1/
#375590000000
0!
0'
0/
#375600000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#375610000000
0!
0'
0/
#375620000000
1!
1'
1/
#375630000000
0!
0'
0/
#375640000000
1!
1'
1/
#375650000000
0!
0'
0/
#375660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#375670000000
0!
0'
0/
#375680000000
1!
1'
1/
#375690000000
0!
0'
0/
#375700000000
1!
1'
1/
#375710000000
0!
0'
0/
#375720000000
1!
1'
1/
#375730000000
0!
0'
0/
#375740000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#375750000000
0!
0'
0/
#375760000000
1!
1'
1/
#375770000000
0!
0'
0/
#375780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#375790000000
0!
0'
0/
#375800000000
1!
1'
1/
#375810000000
0!
0'
0/
#375820000000
#375830000000
1!
1'
1/
#375840000000
0!
0'
0/
#375850000000
1!
1'
1/
#375860000000
0!
1"
0'
1(
0/
10
#375870000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#375880000000
0!
0'
0/
#375890000000
1!
1'
1/
#375900000000
0!
0'
0/
#375910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#375920000000
0!
0'
0/
#375930000000
1!
1'
1/
#375940000000
0!
1"
0'
1(
0/
10
#375950000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#375960000000
0!
1$
0'
1+
0/
#375970000000
1!
1'
1/
#375980000000
0!
0'
0/
#375990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#376000000000
0!
0'
0/
#376010000000
1!
1'
1/
#376020000000
0!
0'
0/
#376030000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#376040000000
0!
0'
0/
#376050000000
1!
1'
1/
#376060000000
0!
0'
0/
#376070000000
1!
1'
1/
#376080000000
0!
0'
0/
#376090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#376100000000
0!
0'
0/
#376110000000
1!
1'
1/
#376120000000
0!
0'
0/
#376130000000
1!
1'
1/
#376140000000
0!
0'
0/
#376150000000
1!
1'
1/
#376160000000
0!
0'
0/
#376170000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#376180000000
0!
0'
0/
#376190000000
1!
1'
1/
#376200000000
0!
0'
0/
#376210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#376220000000
0!
0'
0/
#376230000000
1!
1'
1/
#376240000000
0!
0'
0/
#376250000000
#376260000000
1!
1'
1/
#376270000000
0!
0'
0/
#376280000000
1!
1'
1/
#376290000000
0!
1"
0'
1(
0/
10
#376300000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#376310000000
0!
0'
0/
#376320000000
1!
1'
1/
#376330000000
0!
0'
0/
#376340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#376350000000
0!
0'
0/
#376360000000
1!
1'
1/
#376370000000
0!
1"
0'
1(
0/
10
#376380000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#376390000000
0!
1$
0'
1+
0/
#376400000000
1!
1'
1/
#376410000000
0!
0'
0/
#376420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#376430000000
0!
0'
0/
#376440000000
1!
1'
1/
#376450000000
0!
0'
0/
#376460000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#376470000000
0!
0'
0/
#376480000000
1!
1'
1/
#376490000000
0!
0'
0/
#376500000000
1!
1'
1/
#376510000000
0!
0'
0/
#376520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#376530000000
0!
0'
0/
#376540000000
1!
1'
1/
#376550000000
0!
0'
0/
#376560000000
1!
1'
1/
#376570000000
0!
0'
0/
#376580000000
1!
1'
1/
#376590000000
0!
0'
0/
#376600000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#376610000000
0!
0'
0/
#376620000000
1!
1'
1/
#376630000000
0!
0'
0/
#376640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#376650000000
0!
0'
0/
#376660000000
1!
1'
1/
#376670000000
0!
0'
0/
#376680000000
#376690000000
1!
1'
1/
#376700000000
0!
0'
0/
#376710000000
1!
1'
1/
#376720000000
0!
1"
0'
1(
0/
10
#376730000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#376740000000
0!
0'
0/
#376750000000
1!
1'
1/
#376760000000
0!
0'
0/
#376770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#376780000000
0!
0'
0/
#376790000000
1!
1'
1/
#376800000000
0!
1"
0'
1(
0/
10
#376810000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#376820000000
0!
1$
0'
1+
0/
#376830000000
1!
1'
1/
#376840000000
0!
0'
0/
#376850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#376860000000
0!
0'
0/
#376870000000
1!
1'
1/
#376880000000
0!
0'
0/
#376890000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#376900000000
0!
0'
0/
#376910000000
1!
1'
1/
#376920000000
0!
0'
0/
#376930000000
1!
1'
1/
#376940000000
0!
0'
0/
#376950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#376960000000
0!
0'
0/
#376970000000
1!
1'
1/
#376980000000
0!
0'
0/
#376990000000
1!
1'
1/
#377000000000
0!
0'
0/
#377010000000
1!
1'
1/
#377020000000
0!
0'
0/
#377030000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#377040000000
0!
0'
0/
#377050000000
1!
1'
1/
#377060000000
0!
0'
0/
#377070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#377080000000
0!
0'
0/
#377090000000
1!
1'
1/
#377100000000
0!
0'
0/
#377110000000
#377120000000
1!
1'
1/
#377130000000
0!
0'
0/
#377140000000
1!
1'
1/
#377150000000
0!
1"
0'
1(
0/
10
#377160000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#377170000000
0!
0'
0/
#377180000000
1!
1'
1/
#377190000000
0!
0'
0/
#377200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#377210000000
0!
0'
0/
#377220000000
1!
1'
1/
#377230000000
0!
1"
0'
1(
0/
10
#377240000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#377250000000
0!
1$
0'
1+
0/
#377260000000
1!
1'
1/
#377270000000
0!
0'
0/
#377280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#377290000000
0!
0'
0/
#377300000000
1!
1'
1/
#377310000000
0!
0'
0/
#377320000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#377330000000
0!
0'
0/
#377340000000
1!
1'
1/
#377350000000
0!
0'
0/
#377360000000
1!
1'
1/
#377370000000
0!
0'
0/
#377380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#377390000000
0!
0'
0/
#377400000000
1!
1'
1/
#377410000000
0!
0'
0/
#377420000000
1!
1'
1/
#377430000000
0!
0'
0/
#377440000000
1!
1'
1/
#377450000000
0!
0'
0/
#377460000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#377470000000
0!
0'
0/
#377480000000
1!
1'
1/
#377490000000
0!
0'
0/
#377500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#377510000000
0!
0'
0/
#377520000000
1!
1'
1/
#377530000000
0!
0'
0/
#377540000000
#377550000000
1!
1'
1/
#377560000000
0!
0'
0/
#377570000000
1!
1'
1/
#377580000000
0!
1"
0'
1(
0/
10
#377590000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#377600000000
0!
0'
0/
#377610000000
1!
1'
1/
#377620000000
0!
0'
0/
#377630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#377640000000
0!
0'
0/
#377650000000
1!
1'
1/
#377660000000
0!
1"
0'
1(
0/
10
#377670000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#377680000000
0!
1$
0'
1+
0/
#377690000000
1!
1'
1/
#377700000000
0!
0'
0/
#377710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#377720000000
0!
0'
0/
#377730000000
1!
1'
1/
#377740000000
0!
0'
0/
#377750000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#377760000000
0!
0'
0/
#377770000000
1!
1'
1/
#377780000000
0!
0'
0/
#377790000000
1!
1'
1/
#377800000000
0!
0'
0/
#377810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#377820000000
0!
0'
0/
#377830000000
1!
1'
1/
#377840000000
0!
0'
0/
#377850000000
1!
1'
1/
#377860000000
0!
0'
0/
#377870000000
1!
1'
1/
#377880000000
0!
0'
0/
#377890000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#377900000000
0!
0'
0/
#377910000000
1!
1'
1/
#377920000000
0!
0'
0/
#377930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#377940000000
0!
0'
0/
#377950000000
1!
1'
1/
#377960000000
0!
0'
0/
#377970000000
#377980000000
1!
1'
1/
#377990000000
0!
0'
0/
#378000000000
1!
1'
1/
#378010000000
0!
1"
0'
1(
0/
10
#378020000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#378030000000
0!
0'
0/
#378040000000
1!
1'
1/
#378050000000
0!
0'
0/
#378060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#378070000000
0!
0'
0/
#378080000000
1!
1'
1/
#378090000000
0!
1"
0'
1(
0/
10
#378100000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#378110000000
0!
1$
0'
1+
0/
#378120000000
1!
1'
1/
#378130000000
0!
0'
0/
#378140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#378150000000
0!
0'
0/
#378160000000
1!
1'
1/
#378170000000
0!
0'
0/
#378180000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#378190000000
0!
0'
0/
#378200000000
1!
1'
1/
#378210000000
0!
0'
0/
#378220000000
1!
1'
1/
#378230000000
0!
0'
0/
#378240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#378250000000
0!
0'
0/
#378260000000
1!
1'
1/
#378270000000
0!
0'
0/
#378280000000
1!
1'
1/
#378290000000
0!
0'
0/
#378300000000
1!
1'
1/
#378310000000
0!
0'
0/
#378320000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#378330000000
0!
0'
0/
#378340000000
1!
1'
1/
#378350000000
0!
0'
0/
#378360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#378370000000
0!
0'
0/
#378380000000
1!
1'
1/
#378390000000
0!
0'
0/
#378400000000
#378410000000
1!
1'
1/
#378420000000
0!
0'
0/
#378430000000
1!
1'
1/
#378440000000
0!
1"
0'
1(
0/
10
#378450000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#378460000000
0!
0'
0/
#378470000000
1!
1'
1/
#378480000000
0!
0'
0/
#378490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#378500000000
0!
0'
0/
#378510000000
1!
1'
1/
#378520000000
0!
1"
0'
1(
0/
10
#378530000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#378540000000
0!
1$
0'
1+
0/
#378550000000
1!
1'
1/
#378560000000
0!
0'
0/
#378570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#378580000000
0!
0'
0/
#378590000000
1!
1'
1/
#378600000000
0!
0'
0/
#378610000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#378620000000
0!
0'
0/
#378630000000
1!
1'
1/
#378640000000
0!
0'
0/
#378650000000
1!
1'
1/
#378660000000
0!
0'
0/
#378670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#378680000000
0!
0'
0/
#378690000000
1!
1'
1/
#378700000000
0!
0'
0/
#378710000000
1!
1'
1/
#378720000000
0!
0'
0/
#378730000000
1!
1'
1/
#378740000000
0!
0'
0/
#378750000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#378760000000
0!
0'
0/
#378770000000
1!
1'
1/
#378780000000
0!
0'
0/
#378790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#378800000000
0!
0'
0/
#378810000000
1!
1'
1/
#378820000000
0!
0'
0/
#378830000000
#378840000000
1!
1'
1/
#378850000000
0!
0'
0/
#378860000000
1!
1'
1/
#378870000000
0!
1"
0'
1(
0/
10
#378880000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#378890000000
0!
0'
0/
#378900000000
1!
1'
1/
#378910000000
0!
0'
0/
#378920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#378930000000
0!
0'
0/
#378940000000
1!
1'
1/
#378950000000
0!
1"
0'
1(
0/
10
#378960000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#378970000000
0!
1$
0'
1+
0/
#378980000000
1!
1'
1/
#378990000000
0!
0'
0/
#379000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#379010000000
0!
0'
0/
#379020000000
1!
1'
1/
#379030000000
0!
0'
0/
#379040000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#379050000000
0!
0'
0/
#379060000000
1!
1'
1/
#379070000000
0!
0'
0/
#379080000000
1!
1'
1/
#379090000000
0!
0'
0/
#379100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#379110000000
0!
0'
0/
#379120000000
1!
1'
1/
#379130000000
0!
0'
0/
#379140000000
1!
1'
1/
#379150000000
0!
0'
0/
#379160000000
1!
1'
1/
#379170000000
0!
0'
0/
#379180000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#379190000000
0!
0'
0/
#379200000000
1!
1'
1/
#379210000000
0!
0'
0/
#379220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#379230000000
0!
0'
0/
#379240000000
1!
1'
1/
#379250000000
0!
0'
0/
#379260000000
#379270000000
1!
1'
1/
#379280000000
0!
0'
0/
#379290000000
1!
1'
1/
#379300000000
0!
1"
0'
1(
0/
10
#379310000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#379320000000
0!
0'
0/
#379330000000
1!
1'
1/
#379340000000
0!
0'
0/
#379350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#379360000000
0!
0'
0/
#379370000000
1!
1'
1/
#379380000000
0!
1"
0'
1(
0/
10
#379390000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#379400000000
0!
1$
0'
1+
0/
#379410000000
1!
1'
1/
#379420000000
0!
0'
0/
#379430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#379440000000
0!
0'
0/
#379450000000
1!
1'
1/
#379460000000
0!
0'
0/
#379470000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#379480000000
0!
0'
0/
#379490000000
1!
1'
1/
#379500000000
0!
0'
0/
#379510000000
1!
1'
1/
#379520000000
0!
0'
0/
#379530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#379540000000
0!
0'
0/
#379550000000
1!
1'
1/
#379560000000
0!
0'
0/
#379570000000
1!
1'
1/
#379580000000
0!
0'
0/
#379590000000
1!
1'
1/
#379600000000
0!
0'
0/
#379610000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#379620000000
0!
0'
0/
#379630000000
1!
1'
1/
#379640000000
0!
0'
0/
#379650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#379660000000
0!
0'
0/
#379670000000
1!
1'
1/
#379680000000
0!
0'
0/
#379690000000
#379700000000
1!
1'
1/
#379710000000
0!
0'
0/
#379720000000
1!
1'
1/
#379730000000
0!
1"
0'
1(
0/
10
#379740000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#379750000000
0!
0'
0/
#379760000000
1!
1'
1/
#379770000000
0!
0'
0/
#379780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#379790000000
0!
0'
0/
#379800000000
1!
1'
1/
#379810000000
0!
1"
0'
1(
0/
10
#379820000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#379830000000
0!
1$
0'
1+
0/
#379840000000
1!
1'
1/
#379850000000
0!
0'
0/
#379860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#379870000000
0!
0'
0/
#379880000000
1!
1'
1/
#379890000000
0!
0'
0/
#379900000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#379910000000
0!
0'
0/
#379920000000
1!
1'
1/
#379930000000
0!
0'
0/
#379940000000
1!
1'
1/
#379950000000
0!
0'
0/
#379960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#379970000000
0!
0'
0/
#379980000000
1!
1'
1/
#379990000000
0!
0'
0/
#380000000000
1!
1'
1/
#380010000000
0!
0'
0/
#380020000000
1!
1'
1/
#380030000000
0!
0'
0/
#380040000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#380050000000
0!
0'
0/
#380060000000
1!
1'
1/
#380070000000
0!
0'
0/
#380080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#380090000000
0!
0'
0/
#380100000000
1!
1'
1/
#380110000000
0!
0'
0/
#380120000000
#380130000000
1!
1'
1/
#380140000000
0!
0'
0/
#380150000000
1!
1'
1/
#380160000000
0!
1"
0'
1(
0/
10
#380170000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#380180000000
0!
0'
0/
#380190000000
1!
1'
1/
#380200000000
0!
0'
0/
#380210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#380220000000
0!
0'
0/
#380230000000
1!
1'
1/
#380240000000
0!
1"
0'
1(
0/
10
#380250000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#380260000000
0!
1$
0'
1+
0/
#380270000000
1!
1'
1/
#380280000000
0!
0'
0/
#380290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#380300000000
0!
0'
0/
#380310000000
1!
1'
1/
#380320000000
0!
0'
0/
#380330000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#380340000000
0!
0'
0/
#380350000000
1!
1'
1/
#380360000000
0!
0'
0/
#380370000000
1!
1'
1/
#380380000000
0!
0'
0/
#380390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#380400000000
0!
0'
0/
#380410000000
1!
1'
1/
#380420000000
0!
0'
0/
#380430000000
1!
1'
1/
#380440000000
0!
0'
0/
#380450000000
1!
1'
1/
#380460000000
0!
0'
0/
#380470000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#380480000000
0!
0'
0/
#380490000000
1!
1'
1/
#380500000000
0!
0'
0/
#380510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#380520000000
0!
0'
0/
#380530000000
1!
1'
1/
#380540000000
0!
0'
0/
#380550000000
#380560000000
1!
1'
1/
#380570000000
0!
0'
0/
#380580000000
1!
1'
1/
#380590000000
0!
1"
0'
1(
0/
10
#380600000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#380610000000
0!
0'
0/
#380620000000
1!
1'
1/
#380630000000
0!
0'
0/
#380640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#380650000000
0!
0'
0/
#380660000000
1!
1'
1/
#380670000000
0!
1"
0'
1(
0/
10
#380680000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#380690000000
0!
1$
0'
1+
0/
#380700000000
1!
1'
1/
#380710000000
0!
0'
0/
#380720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#380730000000
0!
0'
0/
#380740000000
1!
1'
1/
#380750000000
0!
0'
0/
#380760000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#380770000000
0!
0'
0/
#380780000000
1!
1'
1/
#380790000000
0!
0'
0/
#380800000000
1!
1'
1/
#380810000000
0!
0'
0/
#380820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#380830000000
0!
0'
0/
#380840000000
1!
1'
1/
#380850000000
0!
0'
0/
#380860000000
1!
1'
1/
#380870000000
0!
0'
0/
#380880000000
1!
1'
1/
#380890000000
0!
0'
0/
#380900000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#380910000000
0!
0'
0/
#380920000000
1!
1'
1/
#380930000000
0!
0'
0/
#380940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#380950000000
0!
0'
0/
#380960000000
1!
1'
1/
#380970000000
0!
0'
0/
#380980000000
#380990000000
1!
1'
1/
#381000000000
0!
0'
0/
#381010000000
1!
1'
1/
#381020000000
0!
1"
0'
1(
0/
10
#381030000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#381040000000
0!
0'
0/
#381050000000
1!
1'
1/
#381060000000
0!
0'
0/
#381070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#381080000000
0!
0'
0/
#381090000000
1!
1'
1/
#381100000000
0!
1"
0'
1(
0/
10
#381110000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#381120000000
0!
1$
0'
1+
0/
#381130000000
1!
1'
1/
#381140000000
0!
0'
0/
#381150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#381160000000
0!
0'
0/
#381170000000
1!
1'
1/
#381180000000
0!
0'
0/
#381190000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#381200000000
0!
0'
0/
#381210000000
1!
1'
1/
#381220000000
0!
0'
0/
#381230000000
1!
1'
1/
#381240000000
0!
0'
0/
#381250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#381260000000
0!
0'
0/
#381270000000
1!
1'
1/
#381280000000
0!
0'
0/
#381290000000
1!
1'
1/
#381300000000
0!
0'
0/
#381310000000
1!
1'
1/
#381320000000
0!
0'
0/
#381330000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#381340000000
0!
0'
0/
#381350000000
1!
1'
1/
#381360000000
0!
0'
0/
#381370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#381380000000
0!
0'
0/
#381390000000
1!
1'
1/
#381400000000
0!
0'
0/
#381410000000
#381420000000
1!
1'
1/
#381430000000
0!
0'
0/
#381440000000
1!
1'
1/
#381450000000
0!
1"
0'
1(
0/
10
#381460000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#381470000000
0!
0'
0/
#381480000000
1!
1'
1/
#381490000000
0!
0'
0/
#381500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#381510000000
0!
0'
0/
#381520000000
1!
1'
1/
#381530000000
0!
1"
0'
1(
0/
10
#381540000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#381550000000
0!
1$
0'
1+
0/
#381560000000
1!
1'
1/
#381570000000
0!
0'
0/
#381580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#381590000000
0!
0'
0/
#381600000000
1!
1'
1/
#381610000000
0!
0'
0/
#381620000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#381630000000
0!
0'
0/
#381640000000
1!
1'
1/
#381650000000
0!
0'
0/
#381660000000
1!
1'
1/
#381670000000
0!
0'
0/
#381680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#381690000000
0!
0'
0/
#381700000000
1!
1'
1/
#381710000000
0!
0'
0/
#381720000000
1!
1'
1/
#381730000000
0!
0'
0/
#381740000000
1!
1'
1/
#381750000000
0!
0'
0/
#381760000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#381770000000
0!
0'
0/
#381780000000
1!
1'
1/
#381790000000
0!
0'
0/
#381800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#381810000000
0!
0'
0/
#381820000000
1!
1'
1/
#381830000000
0!
0'
0/
#381840000000
#381850000000
1!
1'
1/
#381860000000
0!
0'
0/
#381870000000
1!
1'
1/
#381880000000
0!
1"
0'
1(
0/
10
#381890000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#381900000000
0!
0'
0/
#381910000000
1!
1'
1/
#381920000000
0!
0'
0/
#381930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#381940000000
0!
0'
0/
#381950000000
1!
1'
1/
#381960000000
0!
1"
0'
1(
0/
10
#381970000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#381980000000
0!
1$
0'
1+
0/
#381990000000
1!
1'
1/
#382000000000
0!
0'
0/
#382010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#382020000000
0!
0'
0/
#382030000000
1!
1'
1/
#382040000000
0!
0'
0/
#382050000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#382060000000
0!
0'
0/
#382070000000
1!
1'
1/
#382080000000
0!
0'
0/
#382090000000
1!
1'
1/
#382100000000
0!
0'
0/
#382110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#382120000000
0!
0'
0/
#382130000000
1!
1'
1/
#382140000000
0!
0'
0/
#382150000000
1!
1'
1/
#382160000000
0!
0'
0/
#382170000000
1!
1'
1/
#382180000000
0!
0'
0/
#382190000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#382200000000
0!
0'
0/
#382210000000
1!
1'
1/
#382220000000
0!
0'
0/
#382230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#382240000000
0!
0'
0/
#382250000000
1!
1'
1/
#382260000000
0!
0'
0/
#382270000000
#382280000000
1!
1'
1/
#382290000000
0!
0'
0/
#382300000000
1!
1'
1/
#382310000000
0!
1"
0'
1(
0/
10
#382320000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#382330000000
0!
0'
0/
#382340000000
1!
1'
1/
#382350000000
0!
0'
0/
#382360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#382370000000
0!
0'
0/
#382380000000
1!
1'
1/
#382390000000
0!
1"
0'
1(
0/
10
#382400000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#382410000000
0!
1$
0'
1+
0/
#382420000000
1!
1'
1/
#382430000000
0!
0'
0/
#382440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#382450000000
0!
0'
0/
#382460000000
1!
1'
1/
#382470000000
0!
0'
0/
#382480000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#382490000000
0!
0'
0/
#382500000000
1!
1'
1/
#382510000000
0!
0'
0/
#382520000000
1!
1'
1/
#382530000000
0!
0'
0/
#382540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#382550000000
0!
0'
0/
#382560000000
1!
1'
1/
#382570000000
0!
0'
0/
#382580000000
1!
1'
1/
#382590000000
0!
0'
0/
#382600000000
1!
1'
1/
#382610000000
0!
0'
0/
#382620000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#382630000000
0!
0'
0/
#382640000000
1!
1'
1/
#382650000000
0!
0'
0/
#382660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#382670000000
0!
0'
0/
#382680000000
1!
1'
1/
#382690000000
0!
0'
0/
#382700000000
#382710000000
1!
1'
1/
#382720000000
0!
0'
0/
#382730000000
1!
1'
1/
#382740000000
0!
1"
0'
1(
0/
10
#382750000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#382760000000
0!
0'
0/
#382770000000
1!
1'
1/
#382780000000
0!
0'
0/
#382790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#382800000000
0!
0'
0/
#382810000000
1!
1'
1/
#382820000000
0!
1"
0'
1(
0/
10
#382830000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#382840000000
0!
1$
0'
1+
0/
#382850000000
1!
1'
1/
#382860000000
0!
0'
0/
#382870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#382880000000
0!
0'
0/
#382890000000
1!
1'
1/
#382900000000
0!
0'
0/
#382910000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#382920000000
0!
0'
0/
#382930000000
1!
1'
1/
#382940000000
0!
0'
0/
#382950000000
1!
1'
1/
#382960000000
0!
0'
0/
#382970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#382980000000
0!
0'
0/
#382990000000
1!
1'
1/
#383000000000
0!
0'
0/
#383010000000
1!
1'
1/
#383020000000
0!
0'
0/
#383030000000
1!
1'
1/
#383040000000
0!
0'
0/
#383050000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#383060000000
0!
0'
0/
#383070000000
1!
1'
1/
#383080000000
0!
0'
0/
#383090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#383100000000
0!
0'
0/
#383110000000
1!
1'
1/
#383120000000
0!
0'
0/
#383130000000
#383140000000
1!
1'
1/
#383150000000
0!
0'
0/
#383160000000
1!
1'
1/
#383170000000
0!
1"
0'
1(
0/
10
#383180000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#383190000000
0!
0'
0/
#383200000000
1!
1'
1/
#383210000000
0!
0'
0/
#383220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#383230000000
0!
0'
0/
#383240000000
1!
1'
1/
#383250000000
0!
1"
0'
1(
0/
10
#383260000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#383270000000
0!
1$
0'
1+
0/
#383280000000
1!
1'
1/
#383290000000
0!
0'
0/
#383300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#383310000000
0!
0'
0/
#383320000000
1!
1'
1/
#383330000000
0!
0'
0/
#383340000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#383350000000
0!
0'
0/
#383360000000
1!
1'
1/
#383370000000
0!
0'
0/
#383380000000
1!
1'
1/
#383390000000
0!
0'
0/
#383400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#383410000000
0!
0'
0/
#383420000000
1!
1'
1/
#383430000000
0!
0'
0/
#383440000000
1!
1'
1/
#383450000000
0!
0'
0/
#383460000000
1!
1'
1/
#383470000000
0!
0'
0/
#383480000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#383490000000
0!
0'
0/
#383500000000
1!
1'
1/
#383510000000
0!
0'
0/
#383520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#383530000000
0!
0'
0/
#383540000000
1!
1'
1/
#383550000000
0!
0'
0/
#383560000000
#383570000000
1!
1'
1/
#383580000000
0!
0'
0/
#383590000000
1!
1'
1/
#383600000000
0!
1"
0'
1(
0/
10
#383610000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#383620000000
0!
0'
0/
#383630000000
1!
1'
1/
#383640000000
0!
0'
0/
#383650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#383660000000
0!
0'
0/
#383670000000
1!
1'
1/
#383680000000
0!
1"
0'
1(
0/
10
#383690000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#383700000000
0!
1$
0'
1+
0/
#383710000000
1!
1'
1/
#383720000000
0!
0'
0/
#383730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#383740000000
0!
0'
0/
#383750000000
1!
1'
1/
#383760000000
0!
0'
0/
#383770000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#383780000000
0!
0'
0/
#383790000000
1!
1'
1/
#383800000000
0!
0'
0/
#383810000000
1!
1'
1/
#383820000000
0!
0'
0/
#383830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#383840000000
0!
0'
0/
#383850000000
1!
1'
1/
#383860000000
0!
0'
0/
#383870000000
1!
1'
1/
#383880000000
0!
0'
0/
#383890000000
1!
1'
1/
#383900000000
0!
0'
0/
#383910000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#383920000000
0!
0'
0/
#383930000000
1!
1'
1/
#383940000000
0!
0'
0/
#383950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#383960000000
0!
0'
0/
#383970000000
1!
1'
1/
#383980000000
0!
0'
0/
#383990000000
#384000000000
1!
1'
1/
#384010000000
0!
0'
0/
#384020000000
1!
1'
1/
#384030000000
0!
1"
0'
1(
0/
10
#384040000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#384050000000
0!
0'
0/
#384060000000
1!
1'
1/
#384070000000
0!
0'
0/
#384080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#384090000000
0!
0'
0/
#384100000000
1!
1'
1/
#384110000000
0!
1"
0'
1(
0/
10
#384120000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#384130000000
0!
1$
0'
1+
0/
#384140000000
1!
1'
1/
#384150000000
0!
0'
0/
#384160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#384170000000
0!
0'
0/
#384180000000
1!
1'
1/
#384190000000
0!
0'
0/
#384200000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#384210000000
0!
0'
0/
#384220000000
1!
1'
1/
#384230000000
0!
0'
0/
#384240000000
1!
1'
1/
#384250000000
0!
0'
0/
#384260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#384270000000
0!
0'
0/
#384280000000
1!
1'
1/
#384290000000
0!
0'
0/
#384300000000
1!
1'
1/
#384310000000
0!
0'
0/
#384320000000
1!
1'
1/
#384330000000
0!
0'
0/
#384340000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#384350000000
0!
0'
0/
#384360000000
1!
1'
1/
#384370000000
0!
0'
0/
#384380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#384390000000
0!
0'
0/
#384400000000
1!
1'
1/
#384410000000
0!
0'
0/
#384420000000
#384430000000
1!
1'
1/
#384440000000
0!
0'
0/
#384450000000
1!
1'
1/
#384460000000
0!
1"
0'
1(
0/
10
#384470000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#384480000000
0!
0'
0/
#384490000000
1!
1'
1/
#384500000000
0!
0'
0/
#384510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#384520000000
0!
0'
0/
#384530000000
1!
1'
1/
#384540000000
0!
1"
0'
1(
0/
10
#384550000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#384560000000
0!
1$
0'
1+
0/
#384570000000
1!
1'
1/
#384580000000
0!
0'
0/
#384590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#384600000000
0!
0'
0/
#384610000000
1!
1'
1/
#384620000000
0!
0'
0/
#384630000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#384640000000
0!
0'
0/
#384650000000
1!
1'
1/
#384660000000
0!
0'
0/
#384670000000
1!
1'
1/
#384680000000
0!
0'
0/
#384690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#384700000000
0!
0'
0/
#384710000000
1!
1'
1/
#384720000000
0!
0'
0/
#384730000000
1!
1'
1/
#384740000000
0!
0'
0/
#384750000000
1!
1'
1/
#384760000000
0!
0'
0/
#384770000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#384780000000
0!
0'
0/
#384790000000
1!
1'
1/
#384800000000
0!
0'
0/
#384810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#384820000000
0!
0'
0/
#384830000000
1!
1'
1/
#384840000000
0!
0'
0/
#384850000000
#384860000000
1!
1'
1/
#384870000000
0!
0'
0/
#384880000000
1!
1'
1/
#384890000000
0!
1"
0'
1(
0/
10
#384900000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#384910000000
0!
0'
0/
#384920000000
1!
1'
1/
#384930000000
0!
0'
0/
#384940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#384950000000
0!
0'
0/
#384960000000
1!
1'
1/
#384970000000
0!
1"
0'
1(
0/
10
#384980000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#384990000000
0!
1$
0'
1+
0/
#385000000000
1!
1'
1/
#385010000000
0!
0'
0/
#385020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#385030000000
0!
0'
0/
#385040000000
1!
1'
1/
#385050000000
0!
0'
0/
#385060000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#385070000000
0!
0'
0/
#385080000000
1!
1'
1/
#385090000000
0!
0'
0/
#385100000000
1!
1'
1/
#385110000000
0!
0'
0/
#385120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#385130000000
0!
0'
0/
#385140000000
1!
1'
1/
#385150000000
0!
0'
0/
#385160000000
1!
1'
1/
#385170000000
0!
0'
0/
#385180000000
1!
1'
1/
#385190000000
0!
0'
0/
#385200000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#385210000000
0!
0'
0/
#385220000000
1!
1'
1/
#385230000000
0!
0'
0/
#385240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#385250000000
0!
0'
0/
#385260000000
1!
1'
1/
#385270000000
0!
0'
0/
#385280000000
#385290000000
1!
1'
1/
#385300000000
0!
0'
0/
#385310000000
1!
1'
1/
#385320000000
0!
1"
0'
1(
0/
10
#385330000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#385340000000
0!
0'
0/
#385350000000
1!
1'
1/
#385360000000
0!
0'
0/
#385370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#385380000000
0!
0'
0/
#385390000000
1!
1'
1/
#385400000000
0!
1"
0'
1(
0/
10
#385410000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#385420000000
0!
1$
0'
1+
0/
#385430000000
1!
1'
1/
#385440000000
0!
0'
0/
#385450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#385460000000
0!
0'
0/
#385470000000
1!
1'
1/
#385480000000
0!
0'
0/
#385490000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#385500000000
0!
0'
0/
#385510000000
1!
1'
1/
#385520000000
0!
0'
0/
#385530000000
1!
1'
1/
#385540000000
0!
0'
0/
#385550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#385560000000
0!
0'
0/
#385570000000
1!
1'
1/
#385580000000
0!
0'
0/
#385590000000
1!
1'
1/
#385600000000
0!
0'
0/
#385610000000
1!
1'
1/
#385620000000
0!
0'
0/
#385630000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#385640000000
0!
0'
0/
#385650000000
1!
1'
1/
#385660000000
0!
0'
0/
#385670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#385680000000
0!
0'
0/
#385690000000
1!
1'
1/
#385700000000
0!
0'
0/
#385710000000
#385720000000
1!
1'
1/
#385730000000
0!
0'
0/
#385740000000
1!
1'
1/
#385750000000
0!
1"
0'
1(
0/
10
#385760000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#385770000000
0!
0'
0/
#385780000000
1!
1'
1/
#385790000000
0!
0'
0/
#385800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#385810000000
0!
0'
0/
#385820000000
1!
1'
1/
#385830000000
0!
1"
0'
1(
0/
10
#385840000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#385850000000
0!
1$
0'
1+
0/
#385860000000
1!
1'
1/
#385870000000
0!
0'
0/
#385880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#385890000000
0!
0'
0/
#385900000000
1!
1'
1/
#385910000000
0!
0'
0/
#385920000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#385930000000
0!
0'
0/
#385940000000
1!
1'
1/
#385950000000
0!
0'
0/
#385960000000
1!
1'
1/
#385970000000
0!
0'
0/
#385980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#385990000000
0!
0'
0/
#386000000000
1!
1'
1/
#386010000000
0!
0'
0/
#386020000000
1!
1'
1/
#386030000000
0!
0'
0/
#386040000000
1!
1'
1/
#386050000000
0!
0'
0/
#386060000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#386070000000
0!
0'
0/
#386080000000
1!
1'
1/
#386090000000
0!
0'
0/
#386100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#386110000000
0!
0'
0/
#386120000000
1!
1'
1/
#386130000000
0!
0'
0/
#386140000000
#386150000000
1!
1'
1/
#386160000000
0!
0'
0/
#386170000000
1!
1'
1/
#386180000000
0!
1"
0'
1(
0/
10
#386190000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#386200000000
0!
0'
0/
#386210000000
1!
1'
1/
#386220000000
0!
0'
0/
#386230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#386240000000
0!
0'
0/
#386250000000
1!
1'
1/
#386260000000
0!
1"
0'
1(
0/
10
#386270000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#386280000000
0!
1$
0'
1+
0/
#386290000000
1!
1'
1/
#386300000000
0!
0'
0/
#386310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#386320000000
0!
0'
0/
#386330000000
1!
1'
1/
#386340000000
0!
0'
0/
#386350000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#386360000000
0!
0'
0/
#386370000000
1!
1'
1/
#386380000000
0!
0'
0/
#386390000000
1!
1'
1/
#386400000000
0!
0'
0/
#386410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#386420000000
0!
0'
0/
#386430000000
1!
1'
1/
#386440000000
0!
0'
0/
#386450000000
1!
1'
1/
#386460000000
0!
0'
0/
#386470000000
1!
1'
1/
#386480000000
0!
0'
0/
#386490000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#386500000000
0!
0'
0/
#386510000000
1!
1'
1/
#386520000000
0!
0'
0/
#386530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#386540000000
0!
0'
0/
#386550000000
1!
1'
1/
#386560000000
0!
0'
0/
#386570000000
#386580000000
1!
1'
1/
#386590000000
0!
0'
0/
#386600000000
1!
1'
1/
#386610000000
0!
1"
0'
1(
0/
10
#386620000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#386630000000
0!
0'
0/
#386640000000
1!
1'
1/
#386650000000
0!
0'
0/
#386660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#386670000000
0!
0'
0/
#386680000000
1!
1'
1/
#386690000000
0!
1"
0'
1(
0/
10
#386700000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#386710000000
0!
1$
0'
1+
0/
#386720000000
1!
1'
1/
#386730000000
0!
0'
0/
#386740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#386750000000
0!
0'
0/
#386760000000
1!
1'
1/
#386770000000
0!
0'
0/
#386780000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#386790000000
0!
0'
0/
#386800000000
1!
1'
1/
#386810000000
0!
0'
0/
#386820000000
1!
1'
1/
#386830000000
0!
0'
0/
#386840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#386850000000
0!
0'
0/
#386860000000
1!
1'
1/
#386870000000
0!
0'
0/
#386880000000
1!
1'
1/
#386890000000
0!
0'
0/
#386900000000
1!
1'
1/
#386910000000
0!
0'
0/
#386920000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#386930000000
0!
0'
0/
#386940000000
1!
1'
1/
#386950000000
0!
0'
0/
#386960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#386970000000
0!
0'
0/
#386980000000
1!
1'
1/
#386990000000
0!
0'
0/
#387000000000
#387010000000
1!
1'
1/
#387020000000
0!
0'
0/
#387030000000
1!
1'
1/
#387040000000
0!
1"
0'
1(
0/
10
#387050000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#387060000000
0!
0'
0/
#387070000000
1!
1'
1/
#387080000000
0!
0'
0/
#387090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#387100000000
0!
0'
0/
#387110000000
1!
1'
1/
#387120000000
0!
1"
0'
1(
0/
10
#387130000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#387140000000
0!
1$
0'
1+
0/
#387150000000
1!
1'
1/
#387160000000
0!
0'
0/
#387170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#387180000000
0!
0'
0/
#387190000000
1!
1'
1/
#387200000000
0!
0'
0/
#387210000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#387220000000
0!
0'
0/
#387230000000
1!
1'
1/
#387240000000
0!
0'
0/
#387250000000
1!
1'
1/
#387260000000
0!
0'
0/
#387270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#387280000000
0!
0'
0/
#387290000000
1!
1'
1/
#387300000000
0!
0'
0/
#387310000000
1!
1'
1/
#387320000000
0!
0'
0/
#387330000000
1!
1'
1/
#387340000000
0!
0'
0/
#387350000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#387360000000
0!
0'
0/
#387370000000
1!
1'
1/
#387380000000
0!
0'
0/
#387390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#387400000000
0!
0'
0/
#387410000000
1!
1'
1/
#387420000000
0!
0'
0/
#387430000000
#387440000000
1!
1'
1/
#387450000000
0!
0'
0/
#387460000000
1!
1'
1/
#387470000000
0!
1"
0'
1(
0/
10
#387480000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#387490000000
0!
0'
0/
#387500000000
1!
1'
1/
#387510000000
0!
0'
0/
#387520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#387530000000
0!
0'
0/
#387540000000
1!
1'
1/
#387550000000
0!
1"
0'
1(
0/
10
#387560000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#387570000000
0!
1$
0'
1+
0/
#387580000000
1!
1'
1/
#387590000000
0!
0'
0/
#387600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#387610000000
0!
0'
0/
#387620000000
1!
1'
1/
#387630000000
0!
0'
0/
#387640000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#387650000000
0!
0'
0/
#387660000000
1!
1'
1/
#387670000000
0!
0'
0/
#387680000000
1!
1'
1/
#387690000000
0!
0'
0/
#387700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#387710000000
0!
0'
0/
#387720000000
1!
1'
1/
#387730000000
0!
0'
0/
#387740000000
1!
1'
1/
#387750000000
0!
0'
0/
#387760000000
1!
1'
1/
#387770000000
0!
0'
0/
#387780000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#387790000000
0!
0'
0/
#387800000000
1!
1'
1/
#387810000000
0!
0'
0/
#387820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#387830000000
0!
0'
0/
#387840000000
1!
1'
1/
#387850000000
0!
0'
0/
#387860000000
#387870000000
1!
1'
1/
#387880000000
0!
0'
0/
#387890000000
1!
1'
1/
#387900000000
0!
1"
0'
1(
0/
10
#387910000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#387920000000
0!
0'
0/
#387930000000
1!
1'
1/
#387940000000
0!
0'
0/
#387950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#387960000000
0!
0'
0/
#387970000000
1!
1'
1/
#387980000000
0!
1"
0'
1(
0/
10
#387990000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#388000000000
0!
1$
0'
1+
0/
#388010000000
1!
1'
1/
#388020000000
0!
0'
0/
#388030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#388040000000
0!
0'
0/
#388050000000
1!
1'
1/
#388060000000
0!
0'
0/
#388070000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#388080000000
0!
0'
0/
#388090000000
1!
1'
1/
#388100000000
0!
0'
0/
#388110000000
1!
1'
1/
#388120000000
0!
0'
0/
#388130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#388140000000
0!
0'
0/
#388150000000
1!
1'
1/
#388160000000
0!
0'
0/
#388170000000
1!
1'
1/
#388180000000
0!
0'
0/
#388190000000
1!
1'
1/
#388200000000
0!
0'
0/
#388210000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#388220000000
0!
0'
0/
#388230000000
1!
1'
1/
#388240000000
0!
0'
0/
#388250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#388260000000
0!
0'
0/
#388270000000
1!
1'
1/
#388280000000
0!
0'
0/
#388290000000
#388300000000
1!
1'
1/
#388310000000
0!
0'
0/
#388320000000
1!
1'
1/
#388330000000
0!
1"
0'
1(
0/
10
#388340000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#388350000000
0!
0'
0/
#388360000000
1!
1'
1/
#388370000000
0!
0'
0/
#388380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#388390000000
0!
0'
0/
#388400000000
1!
1'
1/
#388410000000
0!
1"
0'
1(
0/
10
#388420000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#388430000000
0!
1$
0'
1+
0/
#388440000000
1!
1'
1/
#388450000000
0!
0'
0/
#388460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#388470000000
0!
0'
0/
#388480000000
1!
1'
1/
#388490000000
0!
0'
0/
#388500000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#388510000000
0!
0'
0/
#388520000000
1!
1'
1/
#388530000000
0!
0'
0/
#388540000000
1!
1'
1/
#388550000000
0!
0'
0/
#388560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#388570000000
0!
0'
0/
#388580000000
1!
1'
1/
#388590000000
0!
0'
0/
#388600000000
1!
1'
1/
#388610000000
0!
0'
0/
#388620000000
1!
1'
1/
#388630000000
0!
0'
0/
#388640000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#388650000000
0!
0'
0/
#388660000000
1!
1'
1/
#388670000000
0!
0'
0/
#388680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#388690000000
0!
0'
0/
#388700000000
1!
1'
1/
#388710000000
0!
0'
0/
#388720000000
#388730000000
1!
1'
1/
#388740000000
0!
0'
0/
#388750000000
1!
1'
1/
#388760000000
0!
1"
0'
1(
0/
10
#388770000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#388780000000
0!
0'
0/
#388790000000
1!
1'
1/
#388800000000
0!
0'
0/
#388810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#388820000000
0!
0'
0/
#388830000000
1!
1'
1/
#388840000000
0!
1"
0'
1(
0/
10
#388850000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#388860000000
0!
1$
0'
1+
0/
#388870000000
1!
1'
1/
#388880000000
0!
0'
0/
#388890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#388900000000
0!
0'
0/
#388910000000
1!
1'
1/
#388920000000
0!
0'
0/
#388930000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#388940000000
0!
0'
0/
#388950000000
1!
1'
1/
#388960000000
0!
0'
0/
#388970000000
1!
1'
1/
#388980000000
0!
0'
0/
#388990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#389000000000
0!
0'
0/
#389010000000
1!
1'
1/
#389020000000
0!
0'
0/
#389030000000
1!
1'
1/
#389040000000
0!
0'
0/
#389050000000
1!
1'
1/
#389060000000
0!
0'
0/
#389070000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#389080000000
0!
0'
0/
#389090000000
1!
1'
1/
#389100000000
0!
0'
0/
#389110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#389120000000
0!
0'
0/
#389130000000
1!
1'
1/
#389140000000
0!
0'
0/
#389150000000
#389160000000
1!
1'
1/
#389170000000
0!
0'
0/
#389180000000
1!
1'
1/
#389190000000
0!
1"
0'
1(
0/
10
#389200000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#389210000000
0!
0'
0/
#389220000000
1!
1'
1/
#389230000000
0!
0'
0/
#389240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#389250000000
0!
0'
0/
#389260000000
1!
1'
1/
#389270000000
0!
1"
0'
1(
0/
10
#389280000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#389290000000
0!
1$
0'
1+
0/
#389300000000
1!
1'
1/
#389310000000
0!
0'
0/
#389320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#389330000000
0!
0'
0/
#389340000000
1!
1'
1/
#389350000000
0!
0'
0/
#389360000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#389370000000
0!
0'
0/
#389380000000
1!
1'
1/
#389390000000
0!
0'
0/
#389400000000
1!
1'
1/
#389410000000
0!
0'
0/
#389420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#389430000000
0!
0'
0/
#389440000000
1!
1'
1/
#389450000000
0!
0'
0/
#389460000000
1!
1'
1/
#389470000000
0!
0'
0/
#389480000000
1!
1'
1/
#389490000000
0!
0'
0/
#389500000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#389510000000
0!
0'
0/
#389520000000
1!
1'
1/
#389530000000
0!
0'
0/
#389540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#389550000000
0!
0'
0/
#389560000000
1!
1'
1/
#389570000000
0!
0'
0/
#389580000000
#389590000000
1!
1'
1/
#389600000000
0!
0'
0/
#389610000000
1!
1'
1/
#389620000000
0!
1"
0'
1(
0/
10
#389630000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#389640000000
0!
0'
0/
#389650000000
1!
1'
1/
#389660000000
0!
0'
0/
#389670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#389680000000
0!
0'
0/
#389690000000
1!
1'
1/
#389700000000
0!
1"
0'
1(
0/
10
#389710000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#389720000000
0!
1$
0'
1+
0/
#389730000000
1!
1'
1/
#389740000000
0!
0'
0/
#389750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#389760000000
0!
0'
0/
#389770000000
1!
1'
1/
#389780000000
0!
0'
0/
#389790000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#389800000000
0!
0'
0/
#389810000000
1!
1'
1/
#389820000000
0!
0'
0/
#389830000000
1!
1'
1/
#389840000000
0!
0'
0/
#389850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#389860000000
0!
0'
0/
#389870000000
1!
1'
1/
#389880000000
0!
0'
0/
#389890000000
1!
1'
1/
#389900000000
0!
0'
0/
#389910000000
1!
1'
1/
#389920000000
0!
0'
0/
#389930000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#389940000000
0!
0'
0/
#389950000000
1!
1'
1/
#389960000000
0!
0'
0/
#389970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#389980000000
0!
0'
0/
#389990000000
1!
1'
1/
#390000000000
0!
0'
0/
#390010000000
#390020000000
1!
1'
1/
#390030000000
0!
0'
0/
#390040000000
1!
1'
1/
#390050000000
0!
1"
0'
1(
0/
10
#390060000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#390070000000
0!
0'
0/
#390080000000
1!
1'
1/
#390090000000
0!
0'
0/
#390100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#390110000000
0!
0'
0/
#390120000000
1!
1'
1/
#390130000000
0!
1"
0'
1(
0/
10
#390140000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#390150000000
0!
1$
0'
1+
0/
#390160000000
1!
1'
1/
#390170000000
0!
0'
0/
#390180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#390190000000
0!
0'
0/
#390200000000
1!
1'
1/
#390210000000
0!
0'
0/
#390220000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#390230000000
0!
0'
0/
#390240000000
1!
1'
1/
#390250000000
0!
0'
0/
#390260000000
1!
1'
1/
#390270000000
0!
0'
0/
#390280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#390290000000
0!
0'
0/
#390300000000
1!
1'
1/
#390310000000
0!
0'
0/
#390320000000
1!
1'
1/
#390330000000
0!
0'
0/
#390340000000
1!
1'
1/
#390350000000
0!
0'
0/
#390360000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#390370000000
0!
0'
0/
#390380000000
1!
1'
1/
#390390000000
0!
0'
0/
#390400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#390410000000
0!
0'
0/
#390420000000
1!
1'
1/
#390430000000
0!
0'
0/
#390440000000
#390450000000
1!
1'
1/
#390460000000
0!
0'
0/
#390470000000
1!
1'
1/
#390480000000
0!
1"
0'
1(
0/
10
#390490000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#390500000000
0!
0'
0/
#390510000000
1!
1'
1/
#390520000000
0!
0'
0/
#390530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#390540000000
0!
0'
0/
#390550000000
1!
1'
1/
#390560000000
0!
1"
0'
1(
0/
10
#390570000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#390580000000
0!
1$
0'
1+
0/
#390590000000
1!
1'
1/
#390600000000
0!
0'
0/
#390610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#390620000000
0!
0'
0/
#390630000000
1!
1'
1/
#390640000000
0!
0'
0/
#390650000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#390660000000
0!
0'
0/
#390670000000
1!
1'
1/
#390680000000
0!
0'
0/
#390690000000
1!
1'
1/
#390700000000
0!
0'
0/
#390710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#390720000000
0!
0'
0/
#390730000000
1!
1'
1/
#390740000000
0!
0'
0/
#390750000000
1!
1'
1/
#390760000000
0!
0'
0/
#390770000000
1!
1'
1/
#390780000000
0!
0'
0/
#390790000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#390800000000
0!
0'
0/
#390810000000
1!
1'
1/
#390820000000
0!
0'
0/
#390830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#390840000000
0!
0'
0/
#390850000000
1!
1'
1/
#390860000000
0!
0'
0/
#390870000000
#390880000000
1!
1'
1/
#390890000000
0!
0'
0/
#390900000000
1!
1'
1/
#390910000000
0!
1"
0'
1(
0/
10
#390920000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#390930000000
0!
0'
0/
#390940000000
1!
1'
1/
#390950000000
0!
0'
0/
#390960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#390970000000
0!
0'
0/
#390980000000
1!
1'
1/
#390990000000
0!
1"
0'
1(
0/
10
#391000000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#391010000000
0!
1$
0'
1+
0/
#391020000000
1!
1'
1/
#391030000000
0!
0'
0/
#391040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#391050000000
0!
0'
0/
#391060000000
1!
1'
1/
#391070000000
0!
0'
0/
#391080000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#391090000000
0!
0'
0/
#391100000000
1!
1'
1/
#391110000000
0!
0'
0/
#391120000000
1!
1'
1/
#391130000000
0!
0'
0/
#391140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#391150000000
0!
0'
0/
#391160000000
1!
1'
1/
#391170000000
0!
0'
0/
#391180000000
1!
1'
1/
#391190000000
0!
0'
0/
#391200000000
1!
1'
1/
#391210000000
0!
0'
0/
#391220000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#391230000000
0!
0'
0/
#391240000000
1!
1'
1/
#391250000000
0!
0'
0/
#391260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#391270000000
0!
0'
0/
#391280000000
1!
1'
1/
#391290000000
0!
0'
0/
#391300000000
#391310000000
1!
1'
1/
#391320000000
0!
0'
0/
#391330000000
1!
1'
1/
#391340000000
0!
1"
0'
1(
0/
10
#391350000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#391360000000
0!
0'
0/
#391370000000
1!
1'
1/
#391380000000
0!
0'
0/
#391390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#391400000000
0!
0'
0/
#391410000000
1!
1'
1/
#391420000000
0!
1"
0'
1(
0/
10
#391430000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#391440000000
0!
1$
0'
1+
0/
#391450000000
1!
1'
1/
#391460000000
0!
0'
0/
#391470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#391480000000
0!
0'
0/
#391490000000
1!
1'
1/
#391500000000
0!
0'
0/
#391510000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#391520000000
0!
0'
0/
#391530000000
1!
1'
1/
#391540000000
0!
0'
0/
#391550000000
1!
1'
1/
#391560000000
0!
0'
0/
#391570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#391580000000
0!
0'
0/
#391590000000
1!
1'
1/
#391600000000
0!
0'
0/
#391610000000
1!
1'
1/
#391620000000
0!
0'
0/
#391630000000
1!
1'
1/
#391640000000
0!
0'
0/
#391650000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#391660000000
0!
0'
0/
#391670000000
1!
1'
1/
#391680000000
0!
0'
0/
#391690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#391700000000
0!
0'
0/
#391710000000
1!
1'
1/
#391720000000
0!
0'
0/
#391730000000
#391740000000
1!
1'
1/
#391750000000
0!
0'
0/
#391760000000
1!
1'
1/
#391770000000
0!
1"
0'
1(
0/
10
#391780000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#391790000000
0!
0'
0/
#391800000000
1!
1'
1/
#391810000000
0!
0'
0/
#391820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#391830000000
0!
0'
0/
#391840000000
1!
1'
1/
#391850000000
0!
1"
0'
1(
0/
10
#391860000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#391870000000
0!
1$
0'
1+
0/
#391880000000
1!
1'
1/
#391890000000
0!
0'
0/
#391900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#391910000000
0!
0'
0/
#391920000000
1!
1'
1/
#391930000000
0!
0'
0/
#391940000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#391950000000
0!
0'
0/
#391960000000
1!
1'
1/
#391970000000
0!
0'
0/
#391980000000
1!
1'
1/
#391990000000
0!
0'
0/
#392000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#392010000000
0!
0'
0/
#392020000000
1!
1'
1/
#392030000000
0!
0'
0/
#392040000000
1!
1'
1/
#392050000000
0!
0'
0/
#392060000000
1!
1'
1/
#392070000000
0!
0'
0/
#392080000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#392090000000
0!
0'
0/
#392100000000
1!
1'
1/
#392110000000
0!
0'
0/
#392120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#392130000000
0!
0'
0/
#392140000000
1!
1'
1/
#392150000000
0!
0'
0/
#392160000000
#392170000000
1!
1'
1/
#392180000000
0!
0'
0/
#392190000000
1!
1'
1/
#392200000000
0!
1"
0'
1(
0/
10
#392210000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#392220000000
0!
0'
0/
#392230000000
1!
1'
1/
#392240000000
0!
0'
0/
#392250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#392260000000
0!
0'
0/
#392270000000
1!
1'
1/
#392280000000
0!
1"
0'
1(
0/
10
#392290000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#392300000000
0!
1$
0'
1+
0/
#392310000000
1!
1'
1/
#392320000000
0!
0'
0/
#392330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#392340000000
0!
0'
0/
#392350000000
1!
1'
1/
#392360000000
0!
0'
0/
#392370000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#392380000000
0!
0'
0/
#392390000000
1!
1'
1/
#392400000000
0!
0'
0/
#392410000000
1!
1'
1/
#392420000000
0!
0'
0/
#392430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#392440000000
0!
0'
0/
#392450000000
1!
1'
1/
#392460000000
0!
0'
0/
#392470000000
1!
1'
1/
#392480000000
0!
0'
0/
#392490000000
1!
1'
1/
#392500000000
0!
0'
0/
#392510000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#392520000000
0!
0'
0/
#392530000000
1!
1'
1/
#392540000000
0!
0'
0/
#392550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#392560000000
0!
0'
0/
#392570000000
1!
1'
1/
#392580000000
0!
0'
0/
#392590000000
#392600000000
1!
1'
1/
#392610000000
0!
0'
0/
#392620000000
1!
1'
1/
#392630000000
0!
1"
0'
1(
0/
10
#392640000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#392650000000
0!
0'
0/
#392660000000
1!
1'
1/
#392670000000
0!
0'
0/
#392680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#392690000000
0!
0'
0/
#392700000000
1!
1'
1/
#392710000000
0!
1"
0'
1(
0/
10
#392720000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#392730000000
0!
1$
0'
1+
0/
#392740000000
1!
1'
1/
#392750000000
0!
0'
0/
#392760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#392770000000
0!
0'
0/
#392780000000
1!
1'
1/
#392790000000
0!
0'
0/
#392800000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#392810000000
0!
0'
0/
#392820000000
1!
1'
1/
#392830000000
0!
0'
0/
#392840000000
1!
1'
1/
#392850000000
0!
0'
0/
#392860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#392870000000
0!
0'
0/
#392880000000
1!
1'
1/
#392890000000
0!
0'
0/
#392900000000
1!
1'
1/
#392910000000
0!
0'
0/
#392920000000
1!
1'
1/
#392930000000
0!
0'
0/
#392940000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#392950000000
0!
0'
0/
#392960000000
1!
1'
1/
#392970000000
0!
0'
0/
#392980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#392990000000
0!
0'
0/
#393000000000
1!
1'
1/
#393010000000
0!
0'
0/
#393020000000
#393030000000
1!
1'
1/
#393040000000
0!
0'
0/
#393050000000
1!
1'
1/
#393060000000
0!
1"
0'
1(
0/
10
#393070000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#393080000000
0!
0'
0/
#393090000000
1!
1'
1/
#393100000000
0!
0'
0/
#393110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#393120000000
0!
0'
0/
#393130000000
1!
1'
1/
#393140000000
0!
1"
0'
1(
0/
10
#393150000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#393160000000
0!
1$
0'
1+
0/
#393170000000
1!
1'
1/
#393180000000
0!
0'
0/
#393190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#393200000000
0!
0'
0/
#393210000000
1!
1'
1/
#393220000000
0!
0'
0/
#393230000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#393240000000
0!
0'
0/
#393250000000
1!
1'
1/
#393260000000
0!
0'
0/
#393270000000
1!
1'
1/
#393280000000
0!
0'
0/
#393290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#393300000000
0!
0'
0/
#393310000000
1!
1'
1/
#393320000000
0!
0'
0/
#393330000000
1!
1'
1/
#393340000000
0!
0'
0/
#393350000000
1!
1'
1/
#393360000000
0!
0'
0/
#393370000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#393380000000
0!
0'
0/
#393390000000
1!
1'
1/
#393400000000
0!
0'
0/
#393410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#393420000000
0!
0'
0/
#393430000000
1!
1'
1/
#393440000000
0!
0'
0/
#393450000000
#393460000000
1!
1'
1/
#393470000000
0!
0'
0/
#393480000000
1!
1'
1/
#393490000000
0!
1"
0'
1(
0/
10
#393500000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#393510000000
0!
0'
0/
#393520000000
1!
1'
1/
#393530000000
0!
0'
0/
#393540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#393550000000
0!
0'
0/
#393560000000
1!
1'
1/
#393570000000
0!
1"
0'
1(
0/
10
#393580000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#393590000000
0!
1$
0'
1+
0/
#393600000000
1!
1'
1/
#393610000000
0!
0'
0/
#393620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#393630000000
0!
0'
0/
#393640000000
1!
1'
1/
#393650000000
0!
0'
0/
#393660000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#393670000000
0!
0'
0/
#393680000000
1!
1'
1/
#393690000000
0!
0'
0/
#393700000000
1!
1'
1/
#393710000000
0!
0'
0/
#393720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#393730000000
0!
0'
0/
#393740000000
1!
1'
1/
#393750000000
0!
0'
0/
#393760000000
1!
1'
1/
#393770000000
0!
0'
0/
#393780000000
1!
1'
1/
#393790000000
0!
0'
0/
#393800000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#393810000000
0!
0'
0/
#393820000000
1!
1'
1/
#393830000000
0!
0'
0/
#393840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#393850000000
0!
0'
0/
#393860000000
1!
1'
1/
#393870000000
0!
0'
0/
#393880000000
#393890000000
1!
1'
1/
#393900000000
0!
0'
0/
#393910000000
1!
1'
1/
#393920000000
0!
1"
0'
1(
0/
10
#393930000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#393940000000
0!
0'
0/
#393950000000
1!
1'
1/
#393960000000
0!
0'
0/
#393970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#393980000000
0!
0'
0/
#393990000000
1!
1'
1/
#394000000000
0!
1"
0'
1(
0/
10
#394010000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#394020000000
0!
1$
0'
1+
0/
#394030000000
1!
1'
1/
#394040000000
0!
0'
0/
#394050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#394060000000
0!
0'
0/
#394070000000
1!
1'
1/
#394080000000
0!
0'
0/
#394090000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#394100000000
0!
0'
0/
#394110000000
1!
1'
1/
#394120000000
0!
0'
0/
#394130000000
1!
1'
1/
#394140000000
0!
0'
0/
#394150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#394160000000
0!
0'
0/
#394170000000
1!
1'
1/
#394180000000
0!
0'
0/
#394190000000
1!
1'
1/
#394200000000
0!
0'
0/
#394210000000
1!
1'
1/
#394220000000
0!
0'
0/
#394230000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#394240000000
0!
0'
0/
#394250000000
1!
1'
1/
#394260000000
0!
0'
0/
#394270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#394280000000
0!
0'
0/
#394290000000
1!
1'
1/
#394300000000
0!
0'
0/
#394310000000
#394320000000
1!
1'
1/
#394330000000
0!
0'
0/
#394340000000
1!
1'
1/
#394350000000
0!
1"
0'
1(
0/
10
#394360000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#394370000000
0!
0'
0/
#394380000000
1!
1'
1/
#394390000000
0!
0'
0/
#394400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#394410000000
0!
0'
0/
#394420000000
1!
1'
1/
#394430000000
0!
1"
0'
1(
0/
10
#394440000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#394450000000
0!
1$
0'
1+
0/
#394460000000
1!
1'
1/
#394470000000
0!
0'
0/
#394480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#394490000000
0!
0'
0/
#394500000000
1!
1'
1/
#394510000000
0!
0'
0/
#394520000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#394530000000
0!
0'
0/
#394540000000
1!
1'
1/
#394550000000
0!
0'
0/
#394560000000
1!
1'
1/
#394570000000
0!
0'
0/
#394580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#394590000000
0!
0'
0/
#394600000000
1!
1'
1/
#394610000000
0!
0'
0/
#394620000000
1!
1'
1/
#394630000000
0!
0'
0/
#394640000000
1!
1'
1/
#394650000000
0!
0'
0/
#394660000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#394670000000
0!
0'
0/
#394680000000
1!
1'
1/
#394690000000
0!
0'
0/
#394700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#394710000000
0!
0'
0/
#394720000000
1!
1'
1/
#394730000000
0!
0'
0/
#394740000000
#394750000000
1!
1'
1/
#394760000000
0!
0'
0/
#394770000000
1!
1'
1/
#394780000000
0!
1"
0'
1(
0/
10
#394790000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#394800000000
0!
0'
0/
#394810000000
1!
1'
1/
#394820000000
0!
0'
0/
#394830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#394840000000
0!
0'
0/
#394850000000
1!
1'
1/
#394860000000
0!
1"
0'
1(
0/
10
#394870000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#394880000000
0!
1$
0'
1+
0/
#394890000000
1!
1'
1/
#394900000000
0!
0'
0/
#394910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#394920000000
0!
0'
0/
#394930000000
1!
1'
1/
#394940000000
0!
0'
0/
#394950000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#394960000000
0!
0'
0/
#394970000000
1!
1'
1/
#394980000000
0!
0'
0/
#394990000000
1!
1'
1/
#395000000000
0!
0'
0/
#395010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#395020000000
0!
0'
0/
#395030000000
1!
1'
1/
#395040000000
0!
0'
0/
#395050000000
1!
1'
1/
#395060000000
0!
0'
0/
#395070000000
1!
1'
1/
#395080000000
0!
0'
0/
#395090000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#395100000000
0!
0'
0/
#395110000000
1!
1'
1/
#395120000000
0!
0'
0/
#395130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#395140000000
0!
0'
0/
#395150000000
1!
1'
1/
#395160000000
0!
0'
0/
#395170000000
#395180000000
1!
1'
1/
#395190000000
0!
0'
0/
#395200000000
1!
1'
1/
#395210000000
0!
1"
0'
1(
0/
10
#395220000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#395230000000
0!
0'
0/
#395240000000
1!
1'
1/
#395250000000
0!
0'
0/
#395260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#395270000000
0!
0'
0/
#395280000000
1!
1'
1/
#395290000000
0!
1"
0'
1(
0/
10
#395300000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#395310000000
0!
1$
0'
1+
0/
#395320000000
1!
1'
1/
#395330000000
0!
0'
0/
#395340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#395350000000
0!
0'
0/
#395360000000
1!
1'
1/
#395370000000
0!
0'
0/
#395380000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#395390000000
0!
0'
0/
#395400000000
1!
1'
1/
#395410000000
0!
0'
0/
#395420000000
1!
1'
1/
#395430000000
0!
0'
0/
#395440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#395450000000
0!
0'
0/
#395460000000
1!
1'
1/
#395470000000
0!
0'
0/
#395480000000
1!
1'
1/
#395490000000
0!
0'
0/
#395500000000
1!
1'
1/
#395510000000
0!
0'
0/
#395520000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#395530000000
0!
0'
0/
#395540000000
1!
1'
1/
#395550000000
0!
0'
0/
#395560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#395570000000
0!
0'
0/
#395580000000
1!
1'
1/
#395590000000
0!
0'
0/
#395600000000
#395610000000
1!
1'
1/
#395620000000
0!
0'
0/
#395630000000
1!
1'
1/
#395640000000
0!
1"
0'
1(
0/
10
#395650000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#395660000000
0!
0'
0/
#395670000000
1!
1'
1/
#395680000000
0!
0'
0/
#395690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#395700000000
0!
0'
0/
#395710000000
1!
1'
1/
#395720000000
0!
1"
0'
1(
0/
10
#395730000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#395740000000
0!
1$
0'
1+
0/
#395750000000
1!
1'
1/
#395760000000
0!
0'
0/
#395770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#395780000000
0!
0'
0/
#395790000000
1!
1'
1/
#395800000000
0!
0'
0/
#395810000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#395820000000
0!
0'
0/
#395830000000
1!
1'
1/
#395840000000
0!
0'
0/
#395850000000
1!
1'
1/
#395860000000
0!
0'
0/
#395870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#395880000000
0!
0'
0/
#395890000000
1!
1'
1/
#395900000000
0!
0'
0/
#395910000000
1!
1'
1/
#395920000000
0!
0'
0/
#395930000000
1!
1'
1/
#395940000000
0!
0'
0/
#395950000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#395960000000
0!
0'
0/
#395970000000
1!
1'
1/
#395980000000
0!
0'
0/
#395990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#396000000000
0!
0'
0/
#396010000000
1!
1'
1/
#396020000000
0!
0'
0/
#396030000000
#396040000000
1!
1'
1/
#396050000000
0!
0'
0/
#396060000000
1!
1'
1/
#396070000000
0!
1"
0'
1(
0/
10
#396080000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#396090000000
0!
0'
0/
#396100000000
1!
1'
1/
#396110000000
0!
0'
0/
#396120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#396130000000
0!
0'
0/
#396140000000
1!
1'
1/
#396150000000
0!
1"
0'
1(
0/
10
#396160000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#396170000000
0!
1$
0'
1+
0/
#396180000000
1!
1'
1/
#396190000000
0!
0'
0/
#396200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#396210000000
0!
0'
0/
#396220000000
1!
1'
1/
#396230000000
0!
0'
0/
#396240000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#396250000000
0!
0'
0/
#396260000000
1!
1'
1/
#396270000000
0!
0'
0/
#396280000000
1!
1'
1/
#396290000000
0!
0'
0/
#396300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#396310000000
0!
0'
0/
#396320000000
1!
1'
1/
#396330000000
0!
0'
0/
#396340000000
1!
1'
1/
#396350000000
0!
0'
0/
#396360000000
1!
1'
1/
#396370000000
0!
0'
0/
#396380000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#396390000000
0!
0'
0/
#396400000000
1!
1'
1/
#396410000000
0!
0'
0/
#396420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#396430000000
0!
0'
0/
#396440000000
1!
1'
1/
#396450000000
0!
0'
0/
#396460000000
#396470000000
1!
1'
1/
#396480000000
0!
0'
0/
#396490000000
1!
1'
1/
#396500000000
0!
1"
0'
1(
0/
10
#396510000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#396520000000
0!
0'
0/
#396530000000
1!
1'
1/
#396540000000
0!
0'
0/
#396550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#396560000000
0!
0'
0/
#396570000000
1!
1'
1/
#396580000000
0!
1"
0'
1(
0/
10
#396590000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#396600000000
0!
1$
0'
1+
0/
#396610000000
1!
1'
1/
#396620000000
0!
0'
0/
#396630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#396640000000
0!
0'
0/
#396650000000
1!
1'
1/
#396660000000
0!
0'
0/
#396670000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#396680000000
0!
0'
0/
#396690000000
1!
1'
1/
#396700000000
0!
0'
0/
#396710000000
1!
1'
1/
#396720000000
0!
0'
0/
#396730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#396740000000
0!
0'
0/
#396750000000
1!
1'
1/
#396760000000
0!
0'
0/
#396770000000
1!
1'
1/
#396780000000
0!
0'
0/
#396790000000
1!
1'
1/
#396800000000
0!
0'
0/
#396810000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#396820000000
0!
0'
0/
#396830000000
1!
1'
1/
#396840000000
0!
0'
0/
#396850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#396860000000
0!
0'
0/
#396870000000
1!
1'
1/
#396880000000
0!
0'
0/
#396890000000
#396900000000
1!
1'
1/
#396910000000
0!
0'
0/
#396920000000
1!
1'
1/
#396930000000
0!
1"
0'
1(
0/
10
#396940000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#396950000000
0!
0'
0/
#396960000000
1!
1'
1/
#396970000000
0!
0'
0/
#396980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#396990000000
0!
0'
0/
#397000000000
1!
1'
1/
#397010000000
0!
1"
0'
1(
0/
10
#397020000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#397030000000
0!
1$
0'
1+
0/
#397040000000
1!
1'
1/
#397050000000
0!
0'
0/
#397060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#397070000000
0!
0'
0/
#397080000000
1!
1'
1/
#397090000000
0!
0'
0/
#397100000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#397110000000
0!
0'
0/
#397120000000
1!
1'
1/
#397130000000
0!
0'
0/
#397140000000
1!
1'
1/
#397150000000
0!
0'
0/
#397160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#397170000000
0!
0'
0/
#397180000000
1!
1'
1/
#397190000000
0!
0'
0/
#397200000000
1!
1'
1/
#397210000000
0!
0'
0/
#397220000000
1!
1'
1/
#397230000000
0!
0'
0/
#397240000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#397250000000
0!
0'
0/
#397260000000
1!
1'
1/
#397270000000
0!
0'
0/
#397280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#397290000000
0!
0'
0/
#397300000000
1!
1'
1/
#397310000000
0!
0'
0/
#397320000000
#397330000000
1!
1'
1/
#397340000000
0!
0'
0/
#397350000000
1!
1'
1/
#397360000000
0!
1"
0'
1(
0/
10
#397370000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#397380000000
0!
0'
0/
#397390000000
1!
1'
1/
#397400000000
0!
0'
0/
#397410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#397420000000
0!
0'
0/
#397430000000
1!
1'
1/
#397440000000
0!
1"
0'
1(
0/
10
#397450000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#397460000000
0!
1$
0'
1+
0/
#397470000000
1!
1'
1/
#397480000000
0!
0'
0/
#397490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#397500000000
0!
0'
0/
#397510000000
1!
1'
1/
#397520000000
0!
0'
0/
#397530000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#397540000000
0!
0'
0/
#397550000000
1!
1'
1/
#397560000000
0!
0'
0/
#397570000000
1!
1'
1/
#397580000000
0!
0'
0/
#397590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#397600000000
0!
0'
0/
#397610000000
1!
1'
1/
#397620000000
0!
0'
0/
#397630000000
1!
1'
1/
#397640000000
0!
0'
0/
#397650000000
1!
1'
1/
#397660000000
0!
0'
0/
#397670000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#397680000000
0!
0'
0/
#397690000000
1!
1'
1/
#397700000000
0!
0'
0/
#397710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#397720000000
0!
0'
0/
#397730000000
1!
1'
1/
#397740000000
0!
0'
0/
#397750000000
#397760000000
1!
1'
1/
#397770000000
0!
0'
0/
#397780000000
1!
1'
1/
#397790000000
0!
1"
0'
1(
0/
10
#397800000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#397810000000
0!
0'
0/
#397820000000
1!
1'
1/
#397830000000
0!
0'
0/
#397840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#397850000000
0!
0'
0/
#397860000000
1!
1'
1/
#397870000000
0!
1"
0'
1(
0/
10
#397880000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#397890000000
0!
1$
0'
1+
0/
#397900000000
1!
1'
1/
#397910000000
0!
0'
0/
#397920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#397930000000
0!
0'
0/
#397940000000
1!
1'
1/
#397950000000
0!
0'
0/
#397960000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#397970000000
0!
0'
0/
#397980000000
1!
1'
1/
#397990000000
0!
0'
0/
#398000000000
1!
1'
1/
#398010000000
0!
0'
0/
#398020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#398030000000
0!
0'
0/
#398040000000
1!
1'
1/
#398050000000
0!
0'
0/
#398060000000
1!
1'
1/
#398070000000
0!
0'
0/
#398080000000
1!
1'
1/
#398090000000
0!
0'
0/
#398100000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#398110000000
0!
0'
0/
#398120000000
1!
1'
1/
#398130000000
0!
0'
0/
#398140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#398150000000
0!
0'
0/
#398160000000
1!
1'
1/
#398170000000
0!
0'
0/
#398180000000
#398190000000
1!
1'
1/
#398200000000
0!
0'
0/
#398210000000
1!
1'
1/
#398220000000
0!
1"
0'
1(
0/
10
#398230000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#398240000000
0!
0'
0/
#398250000000
1!
1'
1/
#398260000000
0!
0'
0/
#398270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#398280000000
0!
0'
0/
#398290000000
1!
1'
1/
#398300000000
0!
1"
0'
1(
0/
10
#398310000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#398320000000
0!
1$
0'
1+
0/
#398330000000
1!
1'
1/
#398340000000
0!
0'
0/
#398350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#398360000000
0!
0'
0/
#398370000000
1!
1'
1/
#398380000000
0!
0'
0/
#398390000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#398400000000
0!
0'
0/
#398410000000
1!
1'
1/
#398420000000
0!
0'
0/
#398430000000
1!
1'
1/
#398440000000
0!
0'
0/
#398450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#398460000000
0!
0'
0/
#398470000000
1!
1'
1/
#398480000000
0!
0'
0/
#398490000000
1!
1'
1/
#398500000000
0!
0'
0/
#398510000000
1!
1'
1/
#398520000000
0!
0'
0/
#398530000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#398540000000
0!
0'
0/
#398550000000
1!
1'
1/
#398560000000
0!
0'
0/
#398570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#398580000000
0!
0'
0/
#398590000000
1!
1'
1/
#398600000000
0!
0'
0/
#398610000000
#398620000000
1!
1'
1/
#398630000000
0!
0'
0/
#398640000000
1!
1'
1/
#398650000000
0!
1"
0'
1(
0/
10
#398660000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#398670000000
0!
0'
0/
#398680000000
1!
1'
1/
#398690000000
0!
0'
0/
#398700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#398710000000
0!
0'
0/
#398720000000
1!
1'
1/
#398730000000
0!
1"
0'
1(
0/
10
#398740000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#398750000000
0!
1$
0'
1+
0/
#398760000000
1!
1'
1/
#398770000000
0!
0'
0/
#398780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#398790000000
0!
0'
0/
#398800000000
1!
1'
1/
#398810000000
0!
0'
0/
#398820000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#398830000000
0!
0'
0/
#398840000000
1!
1'
1/
#398850000000
0!
0'
0/
#398860000000
1!
1'
1/
#398870000000
0!
0'
0/
#398880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#398890000000
0!
0'
0/
#398900000000
1!
1'
1/
#398910000000
0!
0'
0/
#398920000000
1!
1'
1/
#398930000000
0!
0'
0/
#398940000000
1!
1'
1/
#398950000000
0!
0'
0/
#398960000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#398970000000
0!
0'
0/
#398980000000
1!
1'
1/
#398990000000
0!
0'
0/
#399000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#399010000000
0!
0'
0/
#399020000000
1!
1'
1/
#399030000000
0!
0'
0/
#399040000000
#399050000000
1!
1'
1/
#399060000000
0!
0'
0/
#399070000000
1!
1'
1/
#399080000000
0!
1"
0'
1(
0/
10
#399090000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#399100000000
0!
0'
0/
#399110000000
1!
1'
1/
#399120000000
0!
0'
0/
#399130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#399140000000
0!
0'
0/
#399150000000
1!
1'
1/
#399160000000
0!
1"
0'
1(
0/
10
#399170000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#399180000000
0!
1$
0'
1+
0/
#399190000000
1!
1'
1/
#399200000000
0!
0'
0/
#399210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#399220000000
0!
0'
0/
#399230000000
1!
1'
1/
#399240000000
0!
0'
0/
#399250000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#399260000000
0!
0'
0/
#399270000000
1!
1'
1/
#399280000000
0!
0'
0/
#399290000000
1!
1'
1/
#399300000000
0!
0'
0/
#399310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#399320000000
0!
0'
0/
#399330000000
1!
1'
1/
#399340000000
0!
0'
0/
#399350000000
1!
1'
1/
#399360000000
0!
0'
0/
#399370000000
1!
1'
1/
#399380000000
0!
0'
0/
#399390000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#399400000000
0!
0'
0/
#399410000000
1!
1'
1/
#399420000000
0!
0'
0/
#399430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#399440000000
0!
0'
0/
#399450000000
1!
1'
1/
#399460000000
0!
0'
0/
#399470000000
#399480000000
1!
1'
1/
#399490000000
0!
0'
0/
#399500000000
1!
1'
1/
#399510000000
0!
1"
0'
1(
0/
10
#399520000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#399530000000
0!
0'
0/
#399540000000
1!
1'
1/
#399550000000
0!
0'
0/
#399560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#399570000000
0!
0'
0/
#399580000000
1!
1'
1/
#399590000000
0!
1"
0'
1(
0/
10
#399600000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#399610000000
0!
1$
0'
1+
0/
#399620000000
1!
1'
1/
#399630000000
0!
0'
0/
#399640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#399650000000
0!
0'
0/
#399660000000
1!
1'
1/
#399670000000
0!
0'
0/
#399680000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#399690000000
0!
0'
0/
#399700000000
1!
1'
1/
#399710000000
0!
0'
0/
#399720000000
1!
1'
1/
#399730000000
0!
0'
0/
#399740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#399750000000
0!
0'
0/
#399760000000
1!
1'
1/
#399770000000
0!
0'
0/
#399780000000
1!
1'
1/
#399790000000
0!
0'
0/
#399800000000
1!
1'
1/
#399810000000
0!
0'
0/
#399820000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#399830000000
0!
0'
0/
#399840000000
1!
1'
1/
#399850000000
0!
0'
0/
#399860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#399870000000
0!
0'
0/
#399880000000
1!
1'
1/
#399890000000
0!
0'
0/
#399900000000
#399910000000
1!
1'
1/
#399920000000
0!
0'
0/
#399930000000
1!
1'
1/
#399940000000
0!
1"
0'
1(
0/
10
#399950000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#399960000000
0!
0'
0/
#399970000000
1!
1'
1/
#399980000000
0!
0'
0/
#399990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#400000000000
0!
0'
0/
#400010000000
1!
1'
1/
#400020000000
0!
1"
0'
1(
0/
10
#400030000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#400040000000
0!
1$
0'
1+
0/
#400050000000
1!
1'
1/
#400060000000
0!
0'
0/
#400070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#400080000000
0!
0'
0/
#400090000000
1!
1'
1/
#400100000000
0!
0'
0/
#400110000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#400120000000
0!
0'
0/
#400130000000
1!
1'
1/
#400140000000
0!
0'
0/
#400150000000
1!
1'
1/
#400160000000
0!
0'
0/
#400170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#400180000000
0!
0'
0/
#400190000000
1!
1'
1/
#400200000000
0!
0'
0/
#400210000000
1!
1'
1/
#400220000000
0!
0'
0/
#400230000000
1!
1'
1/
#400240000000
0!
0'
0/
#400250000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#400260000000
0!
0'
0/
#400270000000
1!
1'
1/
#400280000000
0!
0'
0/
#400290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#400300000000
0!
0'
0/
#400310000000
1!
1'
1/
#400320000000
0!
0'
0/
#400330000000
#400340000000
1!
1'
1/
#400350000000
0!
0'
0/
#400360000000
1!
1'
1/
#400370000000
0!
1"
0'
1(
0/
10
#400380000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#400390000000
0!
0'
0/
#400400000000
1!
1'
1/
#400410000000
0!
0'
0/
#400420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#400430000000
0!
0'
0/
#400440000000
1!
1'
1/
#400450000000
0!
1"
0'
1(
0/
10
#400460000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#400470000000
0!
1$
0'
1+
0/
#400480000000
1!
1'
1/
#400490000000
0!
0'
0/
#400500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#400510000000
0!
0'
0/
#400520000000
1!
1'
1/
#400530000000
0!
0'
0/
#400540000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#400550000000
0!
0'
0/
#400560000000
1!
1'
1/
#400570000000
0!
0'
0/
#400580000000
1!
1'
1/
#400590000000
0!
0'
0/
#400600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#400610000000
0!
0'
0/
#400620000000
1!
1'
1/
#400630000000
0!
0'
0/
#400640000000
1!
1'
1/
#400650000000
0!
0'
0/
#400660000000
1!
1'
1/
#400670000000
0!
0'
0/
#400680000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#400690000000
0!
0'
0/
#400700000000
1!
1'
1/
#400710000000
0!
0'
0/
#400720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#400730000000
0!
0'
0/
#400740000000
1!
1'
1/
#400750000000
0!
0'
0/
#400760000000
#400770000000
1!
1'
1/
#400780000000
0!
0'
0/
#400790000000
1!
1'
1/
#400800000000
0!
1"
0'
1(
0/
10
#400810000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#400820000000
0!
0'
0/
#400830000000
1!
1'
1/
#400840000000
0!
0'
0/
#400850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#400860000000
0!
0'
0/
#400870000000
1!
1'
1/
#400880000000
0!
1"
0'
1(
0/
10
#400890000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#400900000000
0!
1$
0'
1+
0/
#400910000000
1!
1'
1/
#400920000000
0!
0'
0/
#400930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#400940000000
0!
0'
0/
#400950000000
1!
1'
1/
#400960000000
0!
0'
0/
#400970000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#400980000000
0!
0'
0/
#400990000000
1!
1'
1/
#401000000000
0!
0'
0/
#401010000000
1!
1'
1/
#401020000000
0!
0'
0/
#401030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#401040000000
0!
0'
0/
#401050000000
1!
1'
1/
#401060000000
0!
0'
0/
#401070000000
1!
1'
1/
#401080000000
0!
0'
0/
#401090000000
1!
1'
1/
#401100000000
0!
0'
0/
#401110000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#401120000000
0!
0'
0/
#401130000000
1!
1'
1/
#401140000000
0!
0'
0/
#401150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#401160000000
0!
0'
0/
#401170000000
1!
1'
1/
#401180000000
0!
0'
0/
#401190000000
#401200000000
1!
1'
1/
#401210000000
0!
0'
0/
#401220000000
1!
1'
1/
#401230000000
0!
1"
0'
1(
0/
10
#401240000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#401250000000
0!
0'
0/
#401260000000
1!
1'
1/
#401270000000
0!
0'
0/
#401280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#401290000000
0!
0'
0/
#401300000000
1!
1'
1/
#401310000000
0!
1"
0'
1(
0/
10
#401320000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#401330000000
0!
1$
0'
1+
0/
#401340000000
1!
1'
1/
#401350000000
0!
0'
0/
#401360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#401370000000
0!
0'
0/
#401380000000
1!
1'
1/
#401390000000
0!
0'
0/
#401400000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#401410000000
0!
0'
0/
#401420000000
1!
1'
1/
#401430000000
0!
0'
0/
#401440000000
1!
1'
1/
#401450000000
0!
0'
0/
#401460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#401470000000
0!
0'
0/
#401480000000
1!
1'
1/
#401490000000
0!
0'
0/
#401500000000
1!
1'
1/
#401510000000
0!
0'
0/
#401520000000
1!
1'
1/
#401530000000
0!
0'
0/
#401540000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#401550000000
0!
0'
0/
#401560000000
1!
1'
1/
#401570000000
0!
0'
0/
#401580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#401590000000
0!
0'
0/
#401600000000
1!
1'
1/
#401610000000
0!
0'
0/
#401620000000
#401630000000
1!
1'
1/
#401640000000
0!
0'
0/
#401650000000
1!
1'
1/
#401660000000
0!
1"
0'
1(
0/
10
#401670000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#401680000000
0!
0'
0/
#401690000000
1!
1'
1/
#401700000000
0!
0'
0/
#401710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#401720000000
0!
0'
0/
#401730000000
1!
1'
1/
#401740000000
0!
1"
0'
1(
0/
10
#401750000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#401760000000
0!
1$
0'
1+
0/
#401770000000
1!
1'
1/
#401780000000
0!
0'
0/
#401790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#401800000000
0!
0'
0/
#401810000000
1!
1'
1/
#401820000000
0!
0'
0/
#401830000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#401840000000
0!
0'
0/
#401850000000
1!
1'
1/
#401860000000
0!
0'
0/
#401870000000
1!
1'
1/
#401880000000
0!
0'
0/
#401890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#401900000000
0!
0'
0/
#401910000000
1!
1'
1/
#401920000000
0!
0'
0/
#401930000000
1!
1'
1/
#401940000000
0!
0'
0/
#401950000000
1!
1'
1/
#401960000000
0!
0'
0/
#401970000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#401980000000
0!
0'
0/
#401990000000
1!
1'
1/
#402000000000
0!
0'
0/
#402010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#402020000000
0!
0'
0/
#402030000000
1!
1'
1/
#402040000000
0!
0'
0/
#402050000000
#402060000000
1!
1'
1/
#402070000000
0!
0'
0/
#402080000000
1!
1'
1/
#402090000000
0!
1"
0'
1(
0/
10
#402100000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#402110000000
0!
0'
0/
#402120000000
1!
1'
1/
#402130000000
0!
0'
0/
#402140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#402150000000
0!
0'
0/
#402160000000
1!
1'
1/
#402170000000
0!
1"
0'
1(
0/
10
#402180000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#402190000000
0!
1$
0'
1+
0/
#402200000000
1!
1'
1/
#402210000000
0!
0'
0/
#402220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#402230000000
0!
0'
0/
#402240000000
1!
1'
1/
#402250000000
0!
0'
0/
#402260000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#402270000000
0!
0'
0/
#402280000000
1!
1'
1/
#402290000000
0!
0'
0/
#402300000000
1!
1'
1/
#402310000000
0!
0'
0/
#402320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#402330000000
0!
0'
0/
#402340000000
1!
1'
1/
#402350000000
0!
0'
0/
#402360000000
1!
1'
1/
#402370000000
0!
0'
0/
#402380000000
1!
1'
1/
#402390000000
0!
0'
0/
#402400000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#402410000000
0!
0'
0/
#402420000000
1!
1'
1/
#402430000000
0!
0'
0/
#402440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#402450000000
0!
0'
0/
#402460000000
1!
1'
1/
#402470000000
0!
0'
0/
#402480000000
#402490000000
1!
1'
1/
#402500000000
0!
0'
0/
#402510000000
1!
1'
1/
#402520000000
0!
1"
0'
1(
0/
10
#402530000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#402540000000
0!
0'
0/
#402550000000
1!
1'
1/
#402560000000
0!
0'
0/
#402570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#402580000000
0!
0'
0/
#402590000000
1!
1'
1/
#402600000000
0!
1"
0'
1(
0/
10
#402610000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#402620000000
0!
1$
0'
1+
0/
#402630000000
1!
1'
1/
#402640000000
0!
0'
0/
#402650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#402660000000
0!
0'
0/
#402670000000
1!
1'
1/
#402680000000
0!
0'
0/
#402690000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#402700000000
0!
0'
0/
#402710000000
1!
1'
1/
#402720000000
0!
0'
0/
#402730000000
1!
1'
1/
#402740000000
0!
0'
0/
#402750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#402760000000
0!
0'
0/
#402770000000
1!
1'
1/
#402780000000
0!
0'
0/
#402790000000
1!
1'
1/
#402800000000
0!
0'
0/
#402810000000
1!
1'
1/
#402820000000
0!
0'
0/
#402830000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#402840000000
0!
0'
0/
#402850000000
1!
1'
1/
#402860000000
0!
0'
0/
#402870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#402880000000
0!
0'
0/
#402890000000
1!
1'
1/
#402900000000
0!
0'
0/
#402910000000
#402920000000
1!
1'
1/
#402930000000
0!
0'
0/
#402940000000
1!
1'
1/
#402950000000
0!
1"
0'
1(
0/
10
#402960000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#402970000000
0!
0'
0/
#402980000000
1!
1'
1/
#402990000000
0!
0'
0/
#403000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#403010000000
0!
0'
0/
#403020000000
1!
1'
1/
#403030000000
0!
1"
0'
1(
0/
10
#403040000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#403050000000
0!
1$
0'
1+
0/
#403060000000
1!
1'
1/
#403070000000
0!
0'
0/
#403080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#403090000000
0!
0'
0/
#403100000000
1!
1'
1/
#403110000000
0!
0'
0/
#403120000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#403130000000
0!
0'
0/
#403140000000
1!
1'
1/
#403150000000
0!
0'
0/
#403160000000
1!
1'
1/
#403170000000
0!
0'
0/
#403180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#403190000000
0!
0'
0/
#403200000000
1!
1'
1/
#403210000000
0!
0'
0/
#403220000000
1!
1'
1/
#403230000000
0!
0'
0/
#403240000000
1!
1'
1/
#403250000000
0!
0'
0/
#403260000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#403270000000
0!
0'
0/
#403280000000
1!
1'
1/
#403290000000
0!
0'
0/
#403300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#403310000000
0!
0'
0/
#403320000000
1!
1'
1/
#403330000000
0!
0'
0/
#403340000000
#403350000000
1!
1'
1/
#403360000000
0!
0'
0/
#403370000000
1!
1'
1/
#403380000000
0!
1"
0'
1(
0/
10
#403390000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#403400000000
0!
0'
0/
#403410000000
1!
1'
1/
#403420000000
0!
0'
0/
#403430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#403440000000
0!
0'
0/
#403450000000
1!
1'
1/
#403460000000
0!
1"
0'
1(
0/
10
#403470000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#403480000000
0!
1$
0'
1+
0/
#403490000000
1!
1'
1/
#403500000000
0!
0'
0/
#403510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#403520000000
0!
0'
0/
#403530000000
1!
1'
1/
#403540000000
0!
0'
0/
#403550000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#403560000000
0!
0'
0/
#403570000000
1!
1'
1/
#403580000000
0!
0'
0/
#403590000000
1!
1'
1/
#403600000000
0!
0'
0/
#403610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#403620000000
0!
0'
0/
#403630000000
1!
1'
1/
#403640000000
0!
0'
0/
#403650000000
1!
1'
1/
#403660000000
0!
0'
0/
#403670000000
1!
1'
1/
#403680000000
0!
0'
0/
#403690000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#403700000000
0!
0'
0/
#403710000000
1!
1'
1/
#403720000000
0!
0'
0/
#403730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#403740000000
0!
0'
0/
#403750000000
1!
1'
1/
#403760000000
0!
0'
0/
#403770000000
#403780000000
1!
1'
1/
#403790000000
0!
0'
0/
#403800000000
1!
1'
1/
#403810000000
0!
1"
0'
1(
0/
10
#403820000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#403830000000
0!
0'
0/
#403840000000
1!
1'
1/
#403850000000
0!
0'
0/
#403860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#403870000000
0!
0'
0/
#403880000000
1!
1'
1/
#403890000000
0!
1"
0'
1(
0/
10
#403900000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#403910000000
0!
1$
0'
1+
0/
#403920000000
1!
1'
1/
#403930000000
0!
0'
0/
#403940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#403950000000
0!
0'
0/
#403960000000
1!
1'
1/
#403970000000
0!
0'
0/
#403980000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#403990000000
0!
0'
0/
#404000000000
1!
1'
1/
#404010000000
0!
0'
0/
#404020000000
1!
1'
1/
#404030000000
0!
0'
0/
#404040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#404050000000
0!
0'
0/
#404060000000
1!
1'
1/
#404070000000
0!
0'
0/
#404080000000
1!
1'
1/
#404090000000
0!
0'
0/
#404100000000
1!
1'
1/
#404110000000
0!
0'
0/
#404120000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#404130000000
0!
0'
0/
#404140000000
1!
1'
1/
#404150000000
0!
0'
0/
#404160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#404170000000
0!
0'
0/
#404180000000
1!
1'
1/
#404190000000
0!
0'
0/
#404200000000
#404210000000
1!
1'
1/
#404220000000
0!
0'
0/
#404230000000
1!
1'
1/
#404240000000
0!
1"
0'
1(
0/
10
#404250000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#404260000000
0!
0'
0/
#404270000000
1!
1'
1/
#404280000000
0!
0'
0/
#404290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#404300000000
0!
0'
0/
#404310000000
1!
1'
1/
#404320000000
0!
1"
0'
1(
0/
10
#404330000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#404340000000
0!
1$
0'
1+
0/
#404350000000
1!
1'
1/
#404360000000
0!
0'
0/
#404370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#404380000000
0!
0'
0/
#404390000000
1!
1'
1/
#404400000000
0!
0'
0/
#404410000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#404420000000
0!
0'
0/
#404430000000
1!
1'
1/
#404440000000
0!
0'
0/
#404450000000
1!
1'
1/
#404460000000
0!
0'
0/
#404470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#404480000000
0!
0'
0/
#404490000000
1!
1'
1/
#404500000000
0!
0'
0/
#404510000000
1!
1'
1/
#404520000000
0!
0'
0/
#404530000000
1!
1'
1/
#404540000000
0!
0'
0/
#404550000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#404560000000
0!
0'
0/
#404570000000
1!
1'
1/
#404580000000
0!
0'
0/
#404590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#404600000000
0!
0'
0/
#404610000000
1!
1'
1/
#404620000000
0!
0'
0/
#404630000000
#404640000000
1!
1'
1/
#404650000000
0!
0'
0/
#404660000000
1!
1'
1/
#404670000000
0!
1"
0'
1(
0/
10
#404680000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#404690000000
0!
0'
0/
#404700000000
1!
1'
1/
#404710000000
0!
0'
0/
#404720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#404730000000
0!
0'
0/
#404740000000
1!
1'
1/
#404750000000
0!
1"
0'
1(
0/
10
#404760000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#404770000000
0!
1$
0'
1+
0/
#404780000000
1!
1'
1/
#404790000000
0!
0'
0/
#404800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#404810000000
0!
0'
0/
#404820000000
1!
1'
1/
#404830000000
0!
0'
0/
#404840000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#404850000000
0!
0'
0/
#404860000000
1!
1'
1/
#404870000000
0!
0'
0/
#404880000000
1!
1'
1/
#404890000000
0!
0'
0/
#404900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#404910000000
0!
0'
0/
#404920000000
1!
1'
1/
#404930000000
0!
0'
0/
#404940000000
1!
1'
1/
#404950000000
0!
0'
0/
#404960000000
1!
1'
1/
#404970000000
0!
0'
0/
#404980000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#404990000000
0!
0'
0/
#405000000000
1!
1'
1/
#405010000000
0!
0'
0/
#405020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#405030000000
0!
0'
0/
#405040000000
1!
1'
1/
#405050000000
0!
0'
0/
#405060000000
#405070000000
1!
1'
1/
#405080000000
0!
0'
0/
#405090000000
1!
1'
1/
#405100000000
0!
1"
0'
1(
0/
10
#405110000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#405120000000
0!
0'
0/
#405130000000
1!
1'
1/
#405140000000
0!
0'
0/
#405150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#405160000000
0!
0'
0/
#405170000000
1!
1'
1/
#405180000000
0!
1"
0'
1(
0/
10
#405190000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#405200000000
0!
1$
0'
1+
0/
#405210000000
1!
1'
1/
#405220000000
0!
0'
0/
#405230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#405240000000
0!
0'
0/
#405250000000
1!
1'
1/
#405260000000
0!
0'
0/
#405270000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#405280000000
0!
0'
0/
#405290000000
1!
1'
1/
#405300000000
0!
0'
0/
#405310000000
1!
1'
1/
#405320000000
0!
0'
0/
#405330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#405340000000
0!
0'
0/
#405350000000
1!
1'
1/
#405360000000
0!
0'
0/
#405370000000
1!
1'
1/
#405380000000
0!
0'
0/
#405390000000
1!
1'
1/
#405400000000
0!
0'
0/
#405410000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#405420000000
0!
0'
0/
#405430000000
1!
1'
1/
#405440000000
0!
0'
0/
#405450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#405460000000
0!
0'
0/
#405470000000
1!
1'
1/
#405480000000
0!
0'
0/
#405490000000
#405500000000
1!
1'
1/
#405510000000
0!
0'
0/
#405520000000
1!
1'
1/
#405530000000
0!
1"
0'
1(
0/
10
#405540000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#405550000000
0!
0'
0/
#405560000000
1!
1'
1/
#405570000000
0!
0'
0/
#405580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#405590000000
0!
0'
0/
#405600000000
1!
1'
1/
#405610000000
0!
1"
0'
1(
0/
10
#405620000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#405630000000
0!
1$
0'
1+
0/
#405640000000
1!
1'
1/
#405650000000
0!
0'
0/
#405660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#405670000000
0!
0'
0/
#405680000000
1!
1'
1/
#405690000000
0!
0'
0/
#405700000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#405710000000
0!
0'
0/
#405720000000
1!
1'
1/
#405730000000
0!
0'
0/
#405740000000
1!
1'
1/
#405750000000
0!
0'
0/
#405760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#405770000000
0!
0'
0/
#405780000000
1!
1'
1/
#405790000000
0!
0'
0/
#405800000000
1!
1'
1/
#405810000000
0!
0'
0/
#405820000000
1!
1'
1/
#405830000000
0!
0'
0/
#405840000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#405850000000
0!
0'
0/
#405860000000
1!
1'
1/
#405870000000
0!
0'
0/
#405880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#405890000000
0!
0'
0/
#405900000000
1!
1'
1/
#405910000000
0!
0'
0/
#405920000000
#405930000000
1!
1'
1/
#405940000000
0!
0'
0/
#405950000000
1!
1'
1/
#405960000000
0!
1"
0'
1(
0/
10
#405970000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#405980000000
0!
0'
0/
#405990000000
1!
1'
1/
#406000000000
0!
0'
0/
#406010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#406020000000
0!
0'
0/
#406030000000
1!
1'
1/
#406040000000
0!
1"
0'
1(
0/
10
#406050000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#406060000000
0!
1$
0'
1+
0/
#406070000000
1!
1'
1/
#406080000000
0!
0'
0/
#406090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#406100000000
0!
0'
0/
#406110000000
1!
1'
1/
#406120000000
0!
0'
0/
#406130000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#406140000000
0!
0'
0/
#406150000000
1!
1'
1/
#406160000000
0!
0'
0/
#406170000000
1!
1'
1/
#406180000000
0!
0'
0/
#406190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#406200000000
0!
0'
0/
#406210000000
1!
1'
1/
#406220000000
0!
0'
0/
#406230000000
1!
1'
1/
#406240000000
0!
0'
0/
#406250000000
1!
1'
1/
#406260000000
0!
0'
0/
#406270000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#406280000000
0!
0'
0/
#406290000000
1!
1'
1/
#406300000000
0!
0'
0/
#406310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#406320000000
0!
0'
0/
#406330000000
1!
1'
1/
#406340000000
0!
0'
0/
#406350000000
#406360000000
1!
1'
1/
#406370000000
0!
0'
0/
#406380000000
1!
1'
1/
#406390000000
0!
1"
0'
1(
0/
10
#406400000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#406410000000
0!
0'
0/
#406420000000
1!
1'
1/
#406430000000
0!
0'
0/
#406440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#406450000000
0!
0'
0/
#406460000000
1!
1'
1/
#406470000000
0!
1"
0'
1(
0/
10
#406480000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#406490000000
0!
1$
0'
1+
0/
#406500000000
1!
1'
1/
#406510000000
0!
0'
0/
#406520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#406530000000
0!
0'
0/
#406540000000
1!
1'
1/
#406550000000
0!
0'
0/
#406560000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#406570000000
0!
0'
0/
#406580000000
1!
1'
1/
#406590000000
0!
0'
0/
#406600000000
1!
1'
1/
#406610000000
0!
0'
0/
#406620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#406630000000
0!
0'
0/
#406640000000
1!
1'
1/
#406650000000
0!
0'
0/
#406660000000
1!
1'
1/
#406670000000
0!
0'
0/
#406680000000
1!
1'
1/
#406690000000
0!
0'
0/
#406700000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#406710000000
0!
0'
0/
#406720000000
1!
1'
1/
#406730000000
0!
0'
0/
#406740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#406750000000
0!
0'
0/
#406760000000
1!
1'
1/
#406770000000
0!
0'
0/
#406780000000
#406790000000
1!
1'
1/
#406800000000
0!
0'
0/
#406810000000
1!
1'
1/
#406820000000
0!
1"
0'
1(
0/
10
#406830000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#406840000000
0!
0'
0/
#406850000000
1!
1'
1/
#406860000000
0!
0'
0/
#406870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#406880000000
0!
0'
0/
#406890000000
1!
1'
1/
#406900000000
0!
1"
0'
1(
0/
10
#406910000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#406920000000
0!
1$
0'
1+
0/
#406930000000
1!
1'
1/
#406940000000
0!
0'
0/
#406950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#406960000000
0!
0'
0/
#406970000000
1!
1'
1/
#406980000000
0!
0'
0/
#406990000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#407000000000
0!
0'
0/
#407010000000
1!
1'
1/
#407020000000
0!
0'
0/
#407030000000
1!
1'
1/
#407040000000
0!
0'
0/
#407050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#407060000000
0!
0'
0/
#407070000000
1!
1'
1/
#407080000000
0!
0'
0/
#407090000000
1!
1'
1/
#407100000000
0!
0'
0/
#407110000000
1!
1'
1/
#407120000000
0!
0'
0/
#407130000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#407140000000
0!
0'
0/
#407150000000
1!
1'
1/
#407160000000
0!
0'
0/
#407170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#407180000000
0!
0'
0/
#407190000000
1!
1'
1/
#407200000000
0!
0'
0/
#407210000000
#407220000000
1!
1'
1/
#407230000000
0!
0'
0/
#407240000000
1!
1'
1/
#407250000000
0!
1"
0'
1(
0/
10
#407260000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#407270000000
0!
0'
0/
#407280000000
1!
1'
1/
#407290000000
0!
0'
0/
#407300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#407310000000
0!
0'
0/
#407320000000
1!
1'
1/
#407330000000
0!
1"
0'
1(
0/
10
#407340000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#407350000000
0!
1$
0'
1+
0/
#407360000000
1!
1'
1/
#407370000000
0!
0'
0/
#407380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#407390000000
0!
0'
0/
#407400000000
1!
1'
1/
#407410000000
0!
0'
0/
#407420000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#407430000000
0!
0'
0/
#407440000000
1!
1'
1/
#407450000000
0!
0'
0/
#407460000000
1!
1'
1/
#407470000000
0!
0'
0/
#407480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#407490000000
0!
0'
0/
#407500000000
1!
1'
1/
#407510000000
0!
0'
0/
#407520000000
1!
1'
1/
#407530000000
0!
0'
0/
#407540000000
1!
1'
1/
#407550000000
0!
0'
0/
#407560000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#407570000000
0!
0'
0/
#407580000000
1!
1'
1/
#407590000000
0!
0'
0/
#407600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#407610000000
0!
0'
0/
#407620000000
1!
1'
1/
#407630000000
0!
0'
0/
#407640000000
#407650000000
1!
1'
1/
#407660000000
0!
0'
0/
#407670000000
1!
1'
1/
#407680000000
0!
1"
0'
1(
0/
10
#407690000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#407700000000
0!
0'
0/
#407710000000
1!
1'
1/
#407720000000
0!
0'
0/
#407730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#407740000000
0!
0'
0/
#407750000000
1!
1'
1/
#407760000000
0!
1"
0'
1(
0/
10
#407770000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#407780000000
0!
1$
0'
1+
0/
#407790000000
1!
1'
1/
#407800000000
0!
0'
0/
#407810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#407820000000
0!
0'
0/
#407830000000
1!
1'
1/
#407840000000
0!
0'
0/
#407850000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#407860000000
0!
0'
0/
#407870000000
1!
1'
1/
#407880000000
0!
0'
0/
#407890000000
1!
1'
1/
#407900000000
0!
0'
0/
#407910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#407920000000
0!
0'
0/
#407930000000
1!
1'
1/
#407940000000
0!
0'
0/
#407950000000
1!
1'
1/
#407960000000
0!
0'
0/
#407970000000
1!
1'
1/
#407980000000
0!
0'
0/
#407990000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#408000000000
0!
0'
0/
#408010000000
1!
1'
1/
#408020000000
0!
0'
0/
#408030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#408040000000
0!
0'
0/
#408050000000
1!
1'
1/
#408060000000
0!
0'
0/
#408070000000
#408080000000
1!
1'
1/
#408090000000
0!
0'
0/
#408100000000
1!
1'
1/
#408110000000
0!
1"
0'
1(
0/
10
#408120000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#408130000000
0!
0'
0/
#408140000000
1!
1'
1/
#408150000000
0!
0'
0/
#408160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#408170000000
0!
0'
0/
#408180000000
1!
1'
1/
#408190000000
0!
1"
0'
1(
0/
10
#408200000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#408210000000
0!
1$
0'
1+
0/
#408220000000
1!
1'
1/
#408230000000
0!
0'
0/
#408240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#408250000000
0!
0'
0/
#408260000000
1!
1'
1/
#408270000000
0!
0'
0/
#408280000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#408290000000
0!
0'
0/
#408300000000
1!
1'
1/
#408310000000
0!
0'
0/
#408320000000
1!
1'
1/
#408330000000
0!
0'
0/
#408340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#408350000000
0!
0'
0/
#408360000000
1!
1'
1/
#408370000000
0!
0'
0/
#408380000000
1!
1'
1/
#408390000000
0!
0'
0/
#408400000000
1!
1'
1/
#408410000000
0!
0'
0/
#408420000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#408430000000
0!
0'
0/
#408440000000
1!
1'
1/
#408450000000
0!
0'
0/
#408460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#408470000000
0!
0'
0/
#408480000000
1!
1'
1/
#408490000000
0!
0'
0/
#408500000000
#408510000000
1!
1'
1/
#408520000000
0!
0'
0/
#408530000000
1!
1'
1/
#408540000000
0!
1"
0'
1(
0/
10
#408550000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#408560000000
0!
0'
0/
#408570000000
1!
1'
1/
#408580000000
0!
0'
0/
#408590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#408600000000
0!
0'
0/
#408610000000
1!
1'
1/
#408620000000
0!
1"
0'
1(
0/
10
#408630000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#408640000000
0!
1$
0'
1+
0/
#408650000000
1!
1'
1/
#408660000000
0!
0'
0/
#408670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#408680000000
0!
0'
0/
#408690000000
1!
1'
1/
#408700000000
0!
0'
0/
#408710000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#408720000000
0!
0'
0/
#408730000000
1!
1'
1/
#408740000000
0!
0'
0/
#408750000000
1!
1'
1/
#408760000000
0!
0'
0/
#408770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#408780000000
0!
0'
0/
#408790000000
1!
1'
1/
#408800000000
0!
0'
0/
#408810000000
1!
1'
1/
#408820000000
0!
0'
0/
#408830000000
1!
1'
1/
#408840000000
0!
0'
0/
#408850000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#408860000000
0!
0'
0/
#408870000000
1!
1'
1/
#408880000000
0!
0'
0/
#408890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#408900000000
0!
0'
0/
#408910000000
1!
1'
1/
#408920000000
0!
0'
0/
#408930000000
#408940000000
1!
1'
1/
#408950000000
0!
0'
0/
#408960000000
1!
1'
1/
#408970000000
0!
1"
0'
1(
0/
10
#408980000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#408990000000
0!
0'
0/
#409000000000
1!
1'
1/
#409010000000
0!
0'
0/
#409020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#409030000000
0!
0'
0/
#409040000000
1!
1'
1/
#409050000000
0!
1"
0'
1(
0/
10
#409060000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#409070000000
0!
1$
0'
1+
0/
#409080000000
1!
1'
1/
#409090000000
0!
0'
0/
#409100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#409110000000
0!
0'
0/
#409120000000
1!
1'
1/
#409130000000
0!
0'
0/
#409140000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#409150000000
0!
0'
0/
#409160000000
1!
1'
1/
#409170000000
0!
0'
0/
#409180000000
1!
1'
1/
#409190000000
0!
0'
0/
#409200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#409210000000
0!
0'
0/
#409220000000
1!
1'
1/
#409230000000
0!
0'
0/
#409240000000
1!
1'
1/
#409250000000
0!
0'
0/
#409260000000
1!
1'
1/
#409270000000
0!
0'
0/
#409280000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#409290000000
0!
0'
0/
#409300000000
1!
1'
1/
#409310000000
0!
0'
0/
#409320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#409330000000
0!
0'
0/
#409340000000
1!
1'
1/
#409350000000
0!
0'
0/
#409360000000
#409370000000
1!
1'
1/
#409380000000
0!
0'
0/
#409390000000
1!
1'
1/
#409400000000
0!
1"
0'
1(
0/
10
#409410000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#409420000000
0!
0'
0/
#409430000000
1!
1'
1/
#409440000000
0!
0'
0/
#409450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#409460000000
0!
0'
0/
#409470000000
1!
1'
1/
#409480000000
0!
1"
0'
1(
0/
10
#409490000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#409500000000
0!
1$
0'
1+
0/
#409510000000
1!
1'
1/
#409520000000
0!
0'
0/
#409530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#409540000000
0!
0'
0/
#409550000000
1!
1'
1/
#409560000000
0!
0'
0/
#409570000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#409580000000
0!
0'
0/
#409590000000
1!
1'
1/
#409600000000
0!
0'
0/
#409610000000
1!
1'
1/
#409620000000
0!
0'
0/
#409630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#409640000000
0!
0'
0/
#409650000000
1!
1'
1/
#409660000000
0!
0'
0/
#409670000000
1!
1'
1/
#409680000000
0!
0'
0/
#409690000000
1!
1'
1/
#409700000000
0!
0'
0/
#409710000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#409720000000
0!
0'
0/
#409730000000
1!
1'
1/
#409740000000
0!
0'
0/
#409750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#409760000000
0!
0'
0/
#409770000000
1!
1'
1/
#409780000000
0!
0'
0/
#409790000000
#409800000000
1!
1'
1/
#409810000000
0!
0'
0/
#409820000000
1!
1'
1/
#409830000000
0!
1"
0'
1(
0/
10
#409840000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#409850000000
0!
0'
0/
#409860000000
1!
1'
1/
#409870000000
0!
0'
0/
#409880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#409890000000
0!
0'
0/
#409900000000
1!
1'
1/
#409910000000
0!
1"
0'
1(
0/
10
#409920000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#409930000000
0!
1$
0'
1+
0/
#409940000000
1!
1'
1/
#409950000000
0!
0'
0/
#409960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#409970000000
0!
0'
0/
#409980000000
1!
1'
1/
#409990000000
0!
0'
0/
#410000000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#410010000000
0!
0'
0/
#410020000000
1!
1'
1/
#410030000000
0!
0'
0/
#410040000000
1!
1'
1/
#410050000000
0!
0'
0/
#410060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#410070000000
0!
0'
0/
#410080000000
1!
1'
1/
#410090000000
0!
0'
0/
#410100000000
1!
1'
1/
#410110000000
0!
0'
0/
#410120000000
1!
1'
1/
#410130000000
0!
0'
0/
#410140000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#410150000000
0!
0'
0/
#410160000000
1!
1'
1/
#410170000000
0!
0'
0/
#410180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#410190000000
0!
0'
0/
#410200000000
1!
1'
1/
#410210000000
0!
0'
0/
#410220000000
#410230000000
1!
1'
1/
#410240000000
0!
0'
0/
#410250000000
1!
1'
1/
#410260000000
0!
1"
0'
1(
0/
10
#410270000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#410280000000
0!
0'
0/
#410290000000
1!
1'
1/
#410300000000
0!
0'
0/
#410310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#410320000000
0!
0'
0/
#410330000000
1!
1'
1/
#410340000000
0!
1"
0'
1(
0/
10
#410350000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#410360000000
0!
1$
0'
1+
0/
#410370000000
1!
1'
1/
#410380000000
0!
0'
0/
#410390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#410400000000
0!
0'
0/
#410410000000
1!
1'
1/
#410420000000
0!
0'
0/
#410430000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#410440000000
0!
0'
0/
#410450000000
1!
1'
1/
#410460000000
0!
0'
0/
#410470000000
1!
1'
1/
#410480000000
0!
0'
0/
#410490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#410500000000
0!
0'
0/
#410510000000
1!
1'
1/
#410520000000
0!
0'
0/
#410530000000
1!
1'
1/
#410540000000
0!
0'
0/
#410550000000
1!
1'
1/
#410560000000
0!
0'
0/
#410570000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#410580000000
0!
0'
0/
#410590000000
1!
1'
1/
#410600000000
0!
0'
0/
#410610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#410620000000
0!
0'
0/
#410630000000
1!
1'
1/
#410640000000
0!
0'
0/
#410650000000
#410660000000
1!
1'
1/
#410670000000
0!
0'
0/
#410680000000
1!
1'
1/
#410690000000
0!
1"
0'
1(
0/
10
#410700000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#410710000000
0!
0'
0/
#410720000000
1!
1'
1/
#410730000000
0!
0'
0/
#410740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#410750000000
0!
0'
0/
#410760000000
1!
1'
1/
#410770000000
0!
1"
0'
1(
0/
10
#410780000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#410790000000
0!
1$
0'
1+
0/
#410800000000
1!
1'
1/
#410810000000
0!
0'
0/
#410820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#410830000000
0!
0'
0/
#410840000000
1!
1'
1/
#410850000000
0!
0'
0/
#410860000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#410870000000
0!
0'
0/
#410880000000
1!
1'
1/
#410890000000
0!
0'
0/
#410900000000
1!
1'
1/
#410910000000
0!
0'
0/
#410920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#410930000000
0!
0'
0/
#410940000000
1!
1'
1/
#410950000000
0!
0'
0/
#410960000000
1!
1'
1/
#410970000000
0!
0'
0/
#410980000000
1!
1'
1/
#410990000000
0!
0'
0/
#411000000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#411010000000
0!
0'
0/
#411020000000
1!
1'
1/
#411030000000
0!
0'
0/
#411040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#411050000000
0!
0'
0/
#411060000000
1!
1'
1/
#411070000000
0!
0'
0/
#411080000000
#411090000000
1!
1'
1/
#411100000000
0!
0'
0/
#411110000000
1!
1'
1/
#411120000000
0!
1"
0'
1(
0/
10
#411130000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#411140000000
0!
0'
0/
#411150000000
1!
1'
1/
#411160000000
0!
0'
0/
#411170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#411180000000
0!
0'
0/
#411190000000
1!
1'
1/
#411200000000
0!
1"
0'
1(
0/
10
#411210000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#411220000000
0!
1$
0'
1+
0/
#411230000000
1!
1'
1/
#411240000000
0!
0'
0/
#411250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#411260000000
0!
0'
0/
#411270000000
1!
1'
1/
#411280000000
0!
0'
0/
#411290000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#411300000000
0!
0'
0/
#411310000000
1!
1'
1/
#411320000000
0!
0'
0/
#411330000000
1!
1'
1/
#411340000000
0!
0'
0/
#411350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#411360000000
0!
0'
0/
#411370000000
1!
1'
1/
#411380000000
0!
0'
0/
#411390000000
1!
1'
1/
#411400000000
0!
0'
0/
#411410000000
1!
1'
1/
#411420000000
0!
0'
0/
#411430000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#411440000000
0!
0'
0/
#411450000000
1!
1'
1/
#411460000000
0!
0'
0/
#411470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#411480000000
0!
0'
0/
#411490000000
1!
1'
1/
#411500000000
0!
0'
0/
#411510000000
#411520000000
1!
1'
1/
#411530000000
0!
0'
0/
#411540000000
1!
1'
1/
#411550000000
0!
1"
0'
1(
0/
10
#411560000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#411570000000
0!
0'
0/
#411580000000
1!
1'
1/
#411590000000
0!
0'
0/
#411600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#411610000000
0!
0'
0/
#411620000000
1!
1'
1/
#411630000000
0!
1"
0'
1(
0/
10
#411640000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#411650000000
0!
1$
0'
1+
0/
#411660000000
1!
1'
1/
#411670000000
0!
0'
0/
#411680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#411690000000
0!
0'
0/
#411700000000
1!
1'
1/
#411710000000
0!
0'
0/
#411720000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#411730000000
0!
0'
0/
#411740000000
1!
1'
1/
#411750000000
0!
0'
0/
#411760000000
1!
1'
1/
#411770000000
0!
0'
0/
#411780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#411790000000
0!
0'
0/
#411800000000
1!
1'
1/
#411810000000
0!
0'
0/
#411820000000
1!
1'
1/
#411830000000
0!
0'
0/
#411840000000
1!
1'
1/
#411850000000
0!
0'
0/
#411860000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#411870000000
0!
0'
0/
#411880000000
1!
1'
1/
#411890000000
0!
0'
0/
#411900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#411910000000
0!
0'
0/
#411920000000
1!
1'
1/
#411930000000
0!
0'
0/
#411940000000
#411950000000
1!
1'
1/
#411960000000
0!
0'
0/
#411970000000
1!
1'
1/
#411980000000
0!
1"
0'
1(
0/
10
#411990000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#412000000000
0!
0'
0/
#412010000000
1!
1'
1/
#412020000000
0!
0'
0/
#412030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#412040000000
0!
0'
0/
#412050000000
1!
1'
1/
#412060000000
0!
1"
0'
1(
0/
10
#412070000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#412080000000
0!
1$
0'
1+
0/
#412090000000
1!
1'
1/
#412100000000
0!
0'
0/
#412110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#412120000000
0!
0'
0/
#412130000000
1!
1'
1/
#412140000000
0!
0'
0/
#412150000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#412160000000
0!
0'
0/
#412170000000
1!
1'
1/
#412180000000
0!
0'
0/
#412190000000
1!
1'
1/
#412200000000
0!
0'
0/
#412210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#412220000000
0!
0'
0/
#412230000000
1!
1'
1/
#412240000000
0!
0'
0/
#412250000000
1!
1'
1/
#412260000000
0!
0'
0/
#412270000000
1!
1'
1/
#412280000000
0!
0'
0/
#412290000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#412300000000
0!
0'
0/
#412310000000
1!
1'
1/
#412320000000
0!
0'
0/
#412330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#412340000000
0!
0'
0/
#412350000000
1!
1'
1/
#412360000000
0!
0'
0/
#412370000000
#412380000000
1!
1'
1/
#412390000000
0!
0'
0/
#412400000000
1!
1'
1/
#412410000000
0!
1"
0'
1(
0/
10
#412420000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#412430000000
0!
0'
0/
#412440000000
1!
1'
1/
#412450000000
0!
0'
0/
#412460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#412470000000
0!
0'
0/
#412480000000
1!
1'
1/
#412490000000
0!
1"
0'
1(
0/
10
#412500000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#412510000000
0!
1$
0'
1+
0/
#412520000000
1!
1'
1/
#412530000000
0!
0'
0/
#412540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#412550000000
0!
0'
0/
#412560000000
1!
1'
1/
#412570000000
0!
0'
0/
#412580000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#412590000000
0!
0'
0/
#412600000000
1!
1'
1/
#412610000000
0!
0'
0/
#412620000000
1!
1'
1/
#412630000000
0!
0'
0/
#412640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#412650000000
0!
0'
0/
#412660000000
1!
1'
1/
#412670000000
0!
0'
0/
#412680000000
1!
1'
1/
#412690000000
0!
0'
0/
#412700000000
1!
1'
1/
#412710000000
0!
0'
0/
#412720000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#412730000000
0!
0'
0/
#412740000000
1!
1'
1/
#412750000000
0!
0'
0/
#412760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#412770000000
0!
0'
0/
#412780000000
1!
1'
1/
#412790000000
0!
0'
0/
#412800000000
#412810000000
1!
1'
1/
#412820000000
0!
0'
0/
#412830000000
1!
1'
1/
#412840000000
0!
1"
0'
1(
0/
10
#412850000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#412860000000
0!
0'
0/
#412870000000
1!
1'
1/
#412880000000
0!
0'
0/
#412890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#412900000000
0!
0'
0/
#412910000000
1!
1'
1/
#412920000000
0!
1"
0'
1(
0/
10
#412930000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#412940000000
0!
1$
0'
1+
0/
#412950000000
1!
1'
1/
#412960000000
0!
0'
0/
#412970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#412980000000
0!
0'
0/
#412990000000
1!
1'
1/
#413000000000
0!
0'
0/
#413010000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#413020000000
0!
0'
0/
#413030000000
1!
1'
1/
#413040000000
0!
0'
0/
#413050000000
1!
1'
1/
#413060000000
0!
0'
0/
#413070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#413080000000
0!
0'
0/
#413090000000
1!
1'
1/
#413100000000
0!
0'
0/
#413110000000
1!
1'
1/
#413120000000
0!
0'
0/
#413130000000
1!
1'
1/
#413140000000
0!
0'
0/
#413150000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#413160000000
0!
0'
0/
#413170000000
1!
1'
1/
#413180000000
0!
0'
0/
#413190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#413200000000
0!
0'
0/
#413210000000
1!
1'
1/
#413220000000
0!
0'
0/
#413230000000
#413240000000
1!
1'
1/
#413250000000
0!
0'
0/
#413260000000
1!
1'
1/
#413270000000
0!
1"
0'
1(
0/
10
#413280000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#413290000000
0!
0'
0/
#413300000000
1!
1'
1/
#413310000000
0!
0'
0/
#413320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#413330000000
0!
0'
0/
#413340000000
1!
1'
1/
#413350000000
0!
1"
0'
1(
0/
10
#413360000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#413370000000
0!
1$
0'
1+
0/
#413380000000
1!
1'
1/
#413390000000
0!
0'
0/
#413400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#413410000000
0!
0'
0/
#413420000000
1!
1'
1/
#413430000000
0!
0'
0/
#413440000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#413450000000
0!
0'
0/
#413460000000
1!
1'
1/
#413470000000
0!
0'
0/
#413480000000
1!
1'
1/
#413490000000
0!
0'
0/
#413500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#413510000000
0!
0'
0/
#413520000000
1!
1'
1/
#413530000000
0!
0'
0/
#413540000000
1!
1'
1/
#413550000000
0!
0'
0/
#413560000000
1!
1'
1/
#413570000000
0!
0'
0/
#413580000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#413590000000
0!
0'
0/
#413600000000
1!
1'
1/
#413610000000
0!
0'
0/
#413620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#413630000000
0!
0'
0/
#413640000000
1!
1'
1/
#413650000000
0!
0'
0/
#413660000000
#413670000000
1!
1'
1/
#413680000000
0!
0'
0/
#413690000000
1!
1'
1/
#413700000000
0!
1"
0'
1(
0/
10
#413710000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#413720000000
0!
0'
0/
#413730000000
1!
1'
1/
#413740000000
0!
0'
0/
#413750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#413760000000
0!
0'
0/
#413770000000
1!
1'
1/
#413780000000
0!
1"
0'
1(
0/
10
#413790000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#413800000000
0!
1$
0'
1+
0/
#413810000000
1!
1'
1/
#413820000000
0!
0'
0/
#413830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#413840000000
0!
0'
0/
#413850000000
1!
1'
1/
#413860000000
0!
0'
0/
#413870000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#413880000000
0!
0'
0/
#413890000000
1!
1'
1/
#413900000000
0!
0'
0/
#413910000000
1!
1'
1/
#413920000000
0!
0'
0/
#413930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#413940000000
0!
0'
0/
#413950000000
1!
1'
1/
#413960000000
0!
0'
0/
#413970000000
1!
1'
1/
#413980000000
0!
0'
0/
#413990000000
1!
1'
1/
#414000000000
0!
0'
0/
#414010000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#414020000000
0!
0'
0/
#414030000000
1!
1'
1/
#414040000000
0!
0'
0/
#414050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#414060000000
0!
0'
0/
#414070000000
1!
1'
1/
#414080000000
0!
0'
0/
#414090000000
#414100000000
1!
1'
1/
#414110000000
0!
0'
0/
#414120000000
1!
1'
1/
#414130000000
0!
1"
0'
1(
0/
10
#414140000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#414150000000
0!
0'
0/
#414160000000
1!
1'
1/
#414170000000
0!
0'
0/
#414180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#414190000000
0!
0'
0/
#414200000000
1!
1'
1/
#414210000000
0!
1"
0'
1(
0/
10
#414220000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#414230000000
0!
1$
0'
1+
0/
#414240000000
1!
1'
1/
#414250000000
0!
0'
0/
#414260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#414270000000
0!
0'
0/
#414280000000
1!
1'
1/
#414290000000
0!
0'
0/
#414300000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#414310000000
0!
0'
0/
#414320000000
1!
1'
1/
#414330000000
0!
0'
0/
#414340000000
1!
1'
1/
#414350000000
0!
0'
0/
#414360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#414370000000
0!
0'
0/
#414380000000
1!
1'
1/
#414390000000
0!
0'
0/
#414400000000
1!
1'
1/
#414410000000
0!
0'
0/
#414420000000
1!
1'
1/
#414430000000
0!
0'
0/
#414440000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#414450000000
0!
0'
0/
#414460000000
1!
1'
1/
#414470000000
0!
0'
0/
#414480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#414490000000
0!
0'
0/
#414500000000
1!
1'
1/
#414510000000
0!
0'
0/
#414520000000
#414530000000
1!
1'
1/
#414540000000
0!
0'
0/
#414550000000
1!
1'
1/
#414560000000
0!
1"
0'
1(
0/
10
#414570000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#414580000000
0!
0'
0/
#414590000000
1!
1'
1/
#414600000000
0!
0'
0/
#414610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#414620000000
0!
0'
0/
#414630000000
1!
1'
1/
#414640000000
0!
1"
0'
1(
0/
10
#414650000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#414660000000
0!
1$
0'
1+
0/
#414670000000
1!
1'
1/
#414680000000
0!
0'
0/
#414690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#414700000000
0!
0'
0/
#414710000000
1!
1'
1/
#414720000000
0!
0'
0/
#414730000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#414740000000
0!
0'
0/
#414750000000
1!
1'
1/
#414760000000
0!
0'
0/
#414770000000
1!
1'
1/
#414780000000
0!
0'
0/
#414790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#414800000000
0!
0'
0/
#414810000000
1!
1'
1/
#414820000000
0!
0'
0/
#414830000000
1!
1'
1/
#414840000000
0!
0'
0/
#414850000000
1!
1'
1/
#414860000000
0!
0'
0/
#414870000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#414880000000
0!
0'
0/
#414890000000
1!
1'
1/
#414900000000
0!
0'
0/
#414910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#414920000000
0!
0'
0/
#414930000000
1!
1'
1/
#414940000000
0!
0'
0/
#414950000000
#414960000000
1!
1'
1/
#414970000000
0!
0'
0/
#414980000000
1!
1'
1/
#414990000000
0!
1"
0'
1(
0/
10
#415000000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#415010000000
0!
0'
0/
#415020000000
1!
1'
1/
#415030000000
0!
0'
0/
#415040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#415050000000
0!
0'
0/
#415060000000
1!
1'
1/
#415070000000
0!
1"
0'
1(
0/
10
#415080000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#415090000000
0!
1$
0'
1+
0/
#415100000000
1!
1'
1/
#415110000000
0!
0'
0/
#415120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#415130000000
0!
0'
0/
#415140000000
1!
1'
1/
#415150000000
0!
0'
0/
#415160000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#415170000000
0!
0'
0/
#415180000000
1!
1'
1/
#415190000000
0!
0'
0/
#415200000000
1!
1'
1/
#415210000000
0!
0'
0/
#415220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#415230000000
0!
0'
0/
#415240000000
1!
1'
1/
#415250000000
0!
0'
0/
#415260000000
1!
1'
1/
#415270000000
0!
0'
0/
#415280000000
1!
1'
1/
#415290000000
0!
0'
0/
#415300000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#415310000000
0!
0'
0/
#415320000000
1!
1'
1/
#415330000000
0!
0'
0/
#415340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#415350000000
0!
0'
0/
#415360000000
1!
1'
1/
#415370000000
0!
0'
0/
#415380000000
#415390000000
1!
1'
1/
#415400000000
0!
0'
0/
#415410000000
1!
1'
1/
#415420000000
0!
1"
0'
1(
0/
10
#415430000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#415440000000
0!
0'
0/
#415450000000
1!
1'
1/
#415460000000
0!
0'
0/
#415470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#415480000000
0!
0'
0/
#415490000000
1!
1'
1/
#415500000000
0!
1"
0'
1(
0/
10
#415510000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#415520000000
0!
1$
0'
1+
0/
#415530000000
1!
1'
1/
#415540000000
0!
0'
0/
#415550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#415560000000
0!
0'
0/
#415570000000
1!
1'
1/
#415580000000
0!
0'
0/
#415590000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#415600000000
0!
0'
0/
#415610000000
1!
1'
1/
#415620000000
0!
0'
0/
#415630000000
1!
1'
1/
#415640000000
0!
0'
0/
#415650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#415660000000
0!
0'
0/
#415670000000
1!
1'
1/
#415680000000
0!
0'
0/
#415690000000
1!
1'
1/
#415700000000
0!
0'
0/
#415710000000
1!
1'
1/
#415720000000
0!
0'
0/
#415730000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#415740000000
0!
0'
0/
#415750000000
1!
1'
1/
#415760000000
0!
0'
0/
#415770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#415780000000
0!
0'
0/
#415790000000
1!
1'
1/
#415800000000
0!
0'
0/
#415810000000
#415820000000
1!
1'
1/
#415830000000
0!
0'
0/
#415840000000
1!
1'
1/
#415850000000
0!
1"
0'
1(
0/
10
#415860000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#415870000000
0!
0'
0/
#415880000000
1!
1'
1/
#415890000000
0!
0'
0/
#415900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#415910000000
0!
0'
0/
#415920000000
1!
1'
1/
#415930000000
0!
1"
0'
1(
0/
10
#415940000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#415950000000
0!
1$
0'
1+
0/
#415960000000
1!
1'
1/
#415970000000
0!
0'
0/
#415980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#415990000000
0!
0'
0/
#416000000000
1!
1'
1/
#416010000000
0!
0'
0/
#416020000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#416030000000
0!
0'
0/
#416040000000
1!
1'
1/
#416050000000
0!
0'
0/
#416060000000
1!
1'
1/
#416070000000
0!
0'
0/
#416080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#416090000000
0!
0'
0/
#416100000000
1!
1'
1/
#416110000000
0!
0'
0/
#416120000000
1!
1'
1/
#416130000000
0!
0'
0/
#416140000000
1!
1'
1/
#416150000000
0!
0'
0/
#416160000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#416170000000
0!
0'
0/
#416180000000
1!
1'
1/
#416190000000
0!
0'
0/
#416200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#416210000000
0!
0'
0/
#416220000000
1!
1'
1/
#416230000000
0!
0'
0/
#416240000000
#416250000000
1!
1'
1/
#416260000000
0!
0'
0/
#416270000000
1!
1'
1/
#416280000000
0!
1"
0'
1(
0/
10
#416290000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#416300000000
0!
0'
0/
#416310000000
1!
1'
1/
#416320000000
0!
0'
0/
#416330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#416340000000
0!
0'
0/
#416350000000
1!
1'
1/
#416360000000
0!
1"
0'
1(
0/
10
#416370000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#416380000000
0!
1$
0'
1+
0/
#416390000000
1!
1'
1/
#416400000000
0!
0'
0/
#416410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#416420000000
0!
0'
0/
#416430000000
1!
1'
1/
#416440000000
0!
0'
0/
#416450000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#416460000000
0!
0'
0/
#416470000000
1!
1'
1/
#416480000000
0!
0'
0/
#416490000000
1!
1'
1/
#416500000000
0!
0'
0/
#416510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#416520000000
0!
0'
0/
#416530000000
1!
1'
1/
#416540000000
0!
0'
0/
#416550000000
1!
1'
1/
#416560000000
0!
0'
0/
#416570000000
1!
1'
1/
#416580000000
0!
0'
0/
#416590000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#416600000000
0!
0'
0/
#416610000000
1!
1'
1/
#416620000000
0!
0'
0/
#416630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#416640000000
0!
0'
0/
#416650000000
1!
1'
1/
#416660000000
0!
0'
0/
#416670000000
#416680000000
1!
1'
1/
#416690000000
0!
0'
0/
#416700000000
1!
1'
1/
#416710000000
0!
1"
0'
1(
0/
10
#416720000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#416730000000
0!
0'
0/
#416740000000
1!
1'
1/
#416750000000
0!
0'
0/
#416760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#416770000000
0!
0'
0/
#416780000000
1!
1'
1/
#416790000000
0!
1"
0'
1(
0/
10
#416800000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#416810000000
0!
1$
0'
1+
0/
#416820000000
1!
1'
1/
#416830000000
0!
0'
0/
#416840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#416850000000
0!
0'
0/
#416860000000
1!
1'
1/
#416870000000
0!
0'
0/
#416880000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#416890000000
0!
0'
0/
#416900000000
1!
1'
1/
#416910000000
0!
0'
0/
#416920000000
1!
1'
1/
#416930000000
0!
0'
0/
#416940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#416950000000
0!
0'
0/
#416960000000
1!
1'
1/
#416970000000
0!
0'
0/
#416980000000
1!
1'
1/
#416990000000
0!
0'
0/
#417000000000
1!
1'
1/
#417010000000
0!
0'
0/
#417020000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#417030000000
0!
0'
0/
#417040000000
1!
1'
1/
#417050000000
0!
0'
0/
#417060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#417070000000
0!
0'
0/
#417080000000
1!
1'
1/
#417090000000
0!
0'
0/
#417100000000
#417110000000
1!
1'
1/
#417120000000
0!
0'
0/
#417130000000
1!
1'
1/
#417140000000
0!
1"
0'
1(
0/
10
#417150000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#417160000000
0!
0'
0/
#417170000000
1!
1'
1/
#417180000000
0!
0'
0/
#417190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#417200000000
0!
0'
0/
#417210000000
1!
1'
1/
#417220000000
0!
1"
0'
1(
0/
10
#417230000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#417240000000
0!
1$
0'
1+
0/
#417250000000
1!
1'
1/
#417260000000
0!
0'
0/
#417270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#417280000000
0!
0'
0/
#417290000000
1!
1'
1/
#417300000000
0!
0'
0/
#417310000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#417320000000
0!
0'
0/
#417330000000
1!
1'
1/
#417340000000
0!
0'
0/
#417350000000
1!
1'
1/
#417360000000
0!
0'
0/
#417370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#417380000000
0!
0'
0/
#417390000000
1!
1'
1/
#417400000000
0!
0'
0/
#417410000000
1!
1'
1/
#417420000000
0!
0'
0/
#417430000000
1!
1'
1/
#417440000000
0!
0'
0/
#417450000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#417460000000
0!
0'
0/
#417470000000
1!
1'
1/
#417480000000
0!
0'
0/
#417490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#417500000000
0!
0'
0/
#417510000000
1!
1'
1/
#417520000000
0!
0'
0/
#417530000000
#417540000000
1!
1'
1/
#417550000000
0!
0'
0/
#417560000000
1!
1'
1/
#417570000000
0!
1"
0'
1(
0/
10
#417580000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#417590000000
0!
0'
0/
#417600000000
1!
1'
1/
#417610000000
0!
0'
0/
#417620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#417630000000
0!
0'
0/
#417640000000
1!
1'
1/
#417650000000
0!
1"
0'
1(
0/
10
#417660000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#417670000000
0!
1$
0'
1+
0/
#417680000000
1!
1'
1/
#417690000000
0!
0'
0/
#417700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#417710000000
0!
0'
0/
#417720000000
1!
1'
1/
#417730000000
0!
0'
0/
#417740000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#417750000000
0!
0'
0/
#417760000000
1!
1'
1/
#417770000000
0!
0'
0/
#417780000000
1!
1'
1/
#417790000000
0!
0'
0/
#417800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#417810000000
0!
0'
0/
#417820000000
1!
1'
1/
#417830000000
0!
0'
0/
#417840000000
1!
1'
1/
#417850000000
0!
0'
0/
#417860000000
1!
1'
1/
#417870000000
0!
0'
0/
#417880000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#417890000000
0!
0'
0/
#417900000000
1!
1'
1/
#417910000000
0!
0'
0/
#417920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#417930000000
0!
0'
0/
#417940000000
1!
1'
1/
#417950000000
0!
0'
0/
#417960000000
#417970000000
1!
1'
1/
#417980000000
0!
0'
0/
#417990000000
1!
1'
1/
#418000000000
0!
1"
0'
1(
0/
10
#418010000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#418020000000
0!
0'
0/
#418030000000
1!
1'
1/
#418040000000
0!
0'
0/
#418050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#418060000000
0!
0'
0/
#418070000000
1!
1'
1/
#418080000000
0!
1"
0'
1(
0/
10
#418090000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#418100000000
0!
1$
0'
1+
0/
#418110000000
1!
1'
1/
#418120000000
0!
0'
0/
#418130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#418140000000
0!
0'
0/
#418150000000
1!
1'
1/
#418160000000
0!
0'
0/
#418170000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#418180000000
0!
0'
0/
#418190000000
1!
1'
1/
#418200000000
0!
0'
0/
#418210000000
1!
1'
1/
#418220000000
0!
0'
0/
#418230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#418240000000
0!
0'
0/
#418250000000
1!
1'
1/
#418260000000
0!
0'
0/
#418270000000
1!
1'
1/
#418280000000
0!
0'
0/
#418290000000
1!
1'
1/
#418300000000
0!
0'
0/
#418310000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#418320000000
0!
0'
0/
#418330000000
1!
1'
1/
#418340000000
0!
0'
0/
#418350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#418360000000
0!
0'
0/
#418370000000
1!
1'
1/
#418380000000
0!
0'
0/
#418390000000
#418400000000
1!
1'
1/
#418410000000
0!
0'
0/
#418420000000
1!
1'
1/
#418430000000
0!
1"
0'
1(
0/
10
#418440000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#418450000000
0!
0'
0/
#418460000000
1!
1'
1/
#418470000000
0!
0'
0/
#418480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#418490000000
0!
0'
0/
#418500000000
1!
1'
1/
#418510000000
0!
1"
0'
1(
0/
10
#418520000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#418530000000
0!
1$
0'
1+
0/
#418540000000
1!
1'
1/
#418550000000
0!
0'
0/
#418560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#418570000000
0!
0'
0/
#418580000000
1!
1'
1/
#418590000000
0!
0'
0/
#418600000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#418610000000
0!
0'
0/
#418620000000
1!
1'
1/
#418630000000
0!
0'
0/
#418640000000
1!
1'
1/
#418650000000
0!
0'
0/
#418660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#418670000000
0!
0'
0/
#418680000000
1!
1'
1/
#418690000000
0!
0'
0/
#418700000000
1!
1'
1/
#418710000000
0!
0'
0/
#418720000000
1!
1'
1/
#418730000000
0!
0'
0/
#418740000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#418750000000
0!
0'
0/
#418760000000
1!
1'
1/
#418770000000
0!
0'
0/
#418780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#418790000000
0!
0'
0/
#418800000000
1!
1'
1/
#418810000000
0!
0'
0/
#418820000000
#418830000000
1!
1'
1/
#418840000000
0!
0'
0/
#418850000000
1!
1'
1/
#418860000000
0!
1"
0'
1(
0/
10
#418870000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#418880000000
0!
0'
0/
#418890000000
1!
1'
1/
#418900000000
0!
0'
0/
#418910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#418920000000
0!
0'
0/
#418930000000
1!
1'
1/
#418940000000
0!
1"
0'
1(
0/
10
#418950000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#418960000000
0!
1$
0'
1+
0/
#418970000000
1!
1'
1/
#418980000000
0!
0'
0/
#418990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#419000000000
0!
0'
0/
#419010000000
1!
1'
1/
#419020000000
0!
0'
0/
#419030000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#419040000000
0!
0'
0/
#419050000000
1!
1'
1/
#419060000000
0!
0'
0/
#419070000000
1!
1'
1/
#419080000000
0!
0'
0/
#419090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#419100000000
0!
0'
0/
#419110000000
1!
1'
1/
#419120000000
0!
0'
0/
#419130000000
1!
1'
1/
#419140000000
0!
0'
0/
#419150000000
1!
1'
1/
#419160000000
0!
0'
0/
#419170000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#419180000000
0!
0'
0/
#419190000000
1!
1'
1/
#419200000000
0!
0'
0/
#419210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#419220000000
0!
0'
0/
#419230000000
1!
1'
1/
#419240000000
0!
0'
0/
#419250000000
#419260000000
1!
1'
1/
#419270000000
0!
0'
0/
#419280000000
1!
1'
1/
#419290000000
0!
1"
0'
1(
0/
10
#419300000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#419310000000
0!
0'
0/
#419320000000
1!
1'
1/
#419330000000
0!
0'
0/
#419340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#419350000000
0!
0'
0/
#419360000000
1!
1'
1/
#419370000000
0!
1"
0'
1(
0/
10
#419380000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#419390000000
0!
1$
0'
1+
0/
#419400000000
1!
1'
1/
#419410000000
0!
0'
0/
#419420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#419430000000
0!
0'
0/
#419440000000
1!
1'
1/
#419450000000
0!
0'
0/
#419460000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#419470000000
0!
0'
0/
#419480000000
1!
1'
1/
#419490000000
0!
0'
0/
#419500000000
1!
1'
1/
#419510000000
0!
0'
0/
#419520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#419530000000
0!
0'
0/
#419540000000
1!
1'
1/
#419550000000
0!
0'
0/
#419560000000
1!
1'
1/
#419570000000
0!
0'
0/
#419580000000
1!
1'
1/
#419590000000
0!
0'
0/
#419600000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#419610000000
0!
0'
0/
#419620000000
1!
1'
1/
#419630000000
0!
0'
0/
#419640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#419650000000
0!
0'
0/
#419660000000
1!
1'
1/
#419670000000
0!
0'
0/
#419680000000
#419690000000
1!
1'
1/
#419700000000
0!
0'
0/
#419710000000
1!
1'
1/
#419720000000
0!
1"
0'
1(
0/
10
#419730000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#419740000000
0!
0'
0/
#419750000000
1!
1'
1/
#419760000000
0!
0'
0/
#419770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#419780000000
0!
0'
0/
#419790000000
1!
1'
1/
#419800000000
0!
1"
0'
1(
0/
10
#419810000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#419820000000
0!
1$
0'
1+
0/
#419830000000
1!
1'
1/
#419840000000
0!
0'
0/
#419850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#419860000000
0!
0'
0/
#419870000000
1!
1'
1/
#419880000000
0!
0'
0/
#419890000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#419900000000
0!
0'
0/
#419910000000
1!
1'
1/
#419920000000
0!
0'
0/
#419930000000
1!
1'
1/
#419940000000
0!
0'
0/
#419950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#419960000000
0!
0'
0/
#419970000000
1!
1'
1/
#419980000000
0!
0'
0/
#419990000000
1!
1'
1/
#420000000000
0!
0'
0/
#420010000000
1!
1'
1/
#420020000000
0!
0'
0/
#420030000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#420040000000
0!
0'
0/
#420050000000
1!
1'
1/
#420060000000
0!
0'
0/
#420070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#420080000000
0!
0'
0/
#420090000000
1!
1'
1/
#420100000000
0!
0'
0/
#420110000000
#420120000000
1!
1'
1/
#420130000000
0!
0'
0/
#420140000000
1!
1'
1/
#420150000000
0!
1"
0'
1(
0/
10
#420160000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#420170000000
0!
0'
0/
#420180000000
1!
1'
1/
#420190000000
0!
0'
0/
#420200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#420210000000
0!
0'
0/
#420220000000
1!
1'
1/
#420230000000
0!
1"
0'
1(
0/
10
#420240000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#420250000000
0!
1$
0'
1+
0/
#420260000000
1!
1'
1/
#420270000000
0!
0'
0/
#420280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#420290000000
0!
0'
0/
#420300000000
1!
1'
1/
#420310000000
0!
0'
0/
#420320000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#420330000000
0!
0'
0/
#420340000000
1!
1'
1/
#420350000000
0!
0'
0/
#420360000000
1!
1'
1/
#420370000000
0!
0'
0/
#420380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#420390000000
0!
0'
0/
#420400000000
1!
1'
1/
#420410000000
0!
0'
0/
#420420000000
1!
1'
1/
#420430000000
0!
0'
0/
#420440000000
1!
1'
1/
#420450000000
0!
0'
0/
#420460000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#420470000000
0!
0'
0/
#420480000000
1!
1'
1/
#420490000000
0!
0'
0/
#420500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#420510000000
0!
0'
0/
#420520000000
1!
1'
1/
#420530000000
0!
0'
0/
#420540000000
#420550000000
1!
1'
1/
#420560000000
0!
0'
0/
#420570000000
1!
1'
1/
#420580000000
0!
1"
0'
1(
0/
10
#420590000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#420600000000
0!
0'
0/
#420610000000
1!
1'
1/
#420620000000
0!
0'
0/
#420630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#420640000000
0!
0'
0/
#420650000000
1!
1'
1/
#420660000000
0!
1"
0'
1(
0/
10
#420670000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#420680000000
0!
1$
0'
1+
0/
#420690000000
1!
1'
1/
#420700000000
0!
0'
0/
#420710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#420720000000
0!
0'
0/
#420730000000
1!
1'
1/
#420740000000
0!
0'
0/
#420750000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#420760000000
0!
0'
0/
#420770000000
1!
1'
1/
#420780000000
0!
0'
0/
#420790000000
1!
1'
1/
#420800000000
0!
0'
0/
#420810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#420820000000
0!
0'
0/
#420830000000
1!
1'
1/
#420840000000
0!
0'
0/
#420850000000
1!
1'
1/
#420860000000
0!
0'
0/
#420870000000
1!
1'
1/
#420880000000
0!
0'
0/
#420890000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#420900000000
0!
0'
0/
#420910000000
1!
1'
1/
#420920000000
0!
0'
0/
#420930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#420940000000
0!
0'
0/
#420950000000
1!
1'
1/
#420960000000
0!
0'
0/
#420970000000
#420980000000
1!
1'
1/
#420990000000
0!
0'
0/
#421000000000
1!
1'
1/
#421010000000
0!
1"
0'
1(
0/
10
#421020000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#421030000000
0!
0'
0/
#421040000000
1!
1'
1/
#421050000000
0!
0'
0/
#421060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#421070000000
0!
0'
0/
#421080000000
1!
1'
1/
#421090000000
0!
1"
0'
1(
0/
10
#421100000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#421110000000
0!
1$
0'
1+
0/
#421120000000
1!
1'
1/
#421130000000
0!
0'
0/
#421140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#421150000000
0!
0'
0/
#421160000000
1!
1'
1/
#421170000000
0!
0'
0/
#421180000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#421190000000
0!
0'
0/
#421200000000
1!
1'
1/
#421210000000
0!
0'
0/
#421220000000
1!
1'
1/
#421230000000
0!
0'
0/
#421240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#421250000000
0!
0'
0/
#421260000000
1!
1'
1/
#421270000000
0!
0'
0/
#421280000000
1!
1'
1/
#421290000000
0!
0'
0/
#421300000000
1!
1'
1/
#421310000000
0!
0'
0/
#421320000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#421330000000
0!
0'
0/
#421340000000
1!
1'
1/
#421350000000
0!
0'
0/
#421360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#421370000000
0!
0'
0/
#421380000000
1!
1'
1/
#421390000000
0!
0'
0/
#421400000000
#421410000000
1!
1'
1/
#421420000000
0!
0'
0/
#421430000000
1!
1'
1/
#421440000000
0!
1"
0'
1(
0/
10
#421450000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#421460000000
0!
0'
0/
#421470000000
1!
1'
1/
#421480000000
0!
0'
0/
#421490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#421500000000
0!
0'
0/
#421510000000
1!
1'
1/
#421520000000
0!
1"
0'
1(
0/
10
#421530000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#421540000000
0!
1$
0'
1+
0/
#421550000000
1!
1'
1/
#421560000000
0!
0'
0/
#421570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#421580000000
0!
0'
0/
#421590000000
1!
1'
1/
#421600000000
0!
0'
0/
#421610000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#421620000000
0!
0'
0/
#421630000000
1!
1'
1/
#421640000000
0!
0'
0/
#421650000000
1!
1'
1/
#421660000000
0!
0'
0/
#421670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#421680000000
0!
0'
0/
#421690000000
1!
1'
1/
#421700000000
0!
0'
0/
#421710000000
1!
1'
1/
#421720000000
0!
0'
0/
#421730000000
1!
1'
1/
#421740000000
0!
0'
0/
#421750000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#421760000000
0!
0'
0/
#421770000000
1!
1'
1/
#421780000000
0!
0'
0/
#421790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#421800000000
0!
0'
0/
#421810000000
1!
1'
1/
#421820000000
0!
0'
0/
#421830000000
#421840000000
1!
1'
1/
#421850000000
0!
0'
0/
#421860000000
1!
1'
1/
#421870000000
0!
1"
0'
1(
0/
10
#421880000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#421890000000
0!
0'
0/
#421900000000
1!
1'
1/
#421910000000
0!
0'
0/
#421920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#421930000000
0!
0'
0/
#421940000000
1!
1'
1/
#421950000000
0!
1"
0'
1(
0/
10
#421960000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#421970000000
0!
1$
0'
1+
0/
#421980000000
1!
1'
1/
#421990000000
0!
0'
0/
#422000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#422010000000
0!
0'
0/
#422020000000
1!
1'
1/
#422030000000
0!
0'
0/
#422040000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#422050000000
0!
0'
0/
#422060000000
1!
1'
1/
#422070000000
0!
0'
0/
#422080000000
1!
1'
1/
#422090000000
0!
0'
0/
#422100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#422110000000
0!
0'
0/
#422120000000
1!
1'
1/
#422130000000
0!
0'
0/
#422140000000
1!
1'
1/
#422150000000
0!
0'
0/
#422160000000
1!
1'
1/
#422170000000
0!
0'
0/
#422180000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#422190000000
0!
0'
0/
#422200000000
1!
1'
1/
#422210000000
0!
0'
0/
#422220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#422230000000
0!
0'
0/
#422240000000
1!
1'
1/
#422250000000
0!
0'
0/
#422260000000
#422270000000
1!
1'
1/
#422280000000
0!
0'
0/
#422290000000
1!
1'
1/
#422300000000
0!
1"
0'
1(
0/
10
#422310000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#422320000000
0!
0'
0/
#422330000000
1!
1'
1/
#422340000000
0!
0'
0/
#422350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#422360000000
0!
0'
0/
#422370000000
1!
1'
1/
#422380000000
0!
1"
0'
1(
0/
10
#422390000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#422400000000
0!
1$
0'
1+
0/
#422410000000
1!
1'
1/
#422420000000
0!
0'
0/
#422430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#422440000000
0!
0'
0/
#422450000000
1!
1'
1/
#422460000000
0!
0'
0/
#422470000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#422480000000
0!
0'
0/
#422490000000
1!
1'
1/
#422500000000
0!
0'
0/
#422510000000
1!
1'
1/
#422520000000
0!
0'
0/
#422530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#422540000000
0!
0'
0/
#422550000000
1!
1'
1/
#422560000000
0!
0'
0/
#422570000000
1!
1'
1/
#422580000000
0!
0'
0/
#422590000000
1!
1'
1/
#422600000000
0!
0'
0/
#422610000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#422620000000
0!
0'
0/
#422630000000
1!
1'
1/
#422640000000
0!
0'
0/
#422650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#422660000000
0!
0'
0/
#422670000000
1!
1'
1/
#422680000000
0!
0'
0/
#422690000000
#422700000000
1!
1'
1/
#422710000000
0!
0'
0/
#422720000000
1!
1'
1/
#422730000000
0!
1"
0'
1(
0/
10
#422740000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#422750000000
0!
0'
0/
#422760000000
1!
1'
1/
#422770000000
0!
0'
0/
#422780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#422790000000
0!
0'
0/
#422800000000
1!
1'
1/
#422810000000
0!
1"
0'
1(
0/
10
#422820000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#422830000000
0!
1$
0'
1+
0/
#422840000000
1!
1'
1/
#422850000000
0!
0'
0/
#422860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#422870000000
0!
0'
0/
#422880000000
1!
1'
1/
#422890000000
0!
0'
0/
#422900000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#422910000000
0!
0'
0/
#422920000000
1!
1'
1/
#422930000000
0!
0'
0/
#422940000000
1!
1'
1/
#422950000000
0!
0'
0/
#422960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#422970000000
0!
0'
0/
#422980000000
1!
1'
1/
#422990000000
0!
0'
0/
#423000000000
1!
1'
1/
#423010000000
0!
0'
0/
#423020000000
1!
1'
1/
#423030000000
0!
0'
0/
#423040000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#423050000000
0!
0'
0/
#423060000000
1!
1'
1/
#423070000000
0!
0'
0/
#423080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#423090000000
0!
0'
0/
#423100000000
1!
1'
1/
#423110000000
0!
0'
0/
#423120000000
#423130000000
1!
1'
1/
#423140000000
0!
0'
0/
#423150000000
1!
1'
1/
#423160000000
0!
1"
0'
1(
0/
10
#423170000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#423180000000
0!
0'
0/
#423190000000
1!
1'
1/
#423200000000
0!
0'
0/
#423210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#423220000000
0!
0'
0/
#423230000000
1!
1'
1/
#423240000000
0!
1"
0'
1(
0/
10
#423250000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#423260000000
0!
1$
0'
1+
0/
#423270000000
1!
1'
1/
#423280000000
0!
0'
0/
#423290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#423300000000
0!
0'
0/
#423310000000
1!
1'
1/
#423320000000
0!
0'
0/
#423330000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#423340000000
0!
0'
0/
#423350000000
1!
1'
1/
#423360000000
0!
0'
0/
#423370000000
1!
1'
1/
#423380000000
0!
0'
0/
#423390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#423400000000
0!
0'
0/
#423410000000
1!
1'
1/
#423420000000
0!
0'
0/
#423430000000
1!
1'
1/
#423440000000
0!
0'
0/
#423450000000
1!
1'
1/
#423460000000
0!
0'
0/
#423470000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#423480000000
0!
0'
0/
#423490000000
1!
1'
1/
#423500000000
0!
0'
0/
#423510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#423520000000
0!
0'
0/
#423530000000
1!
1'
1/
#423540000000
0!
0'
0/
#423550000000
#423560000000
1!
1'
1/
#423570000000
0!
0'
0/
#423580000000
1!
1'
1/
#423590000000
0!
1"
0'
1(
0/
10
#423600000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#423610000000
0!
0'
0/
#423620000000
1!
1'
1/
#423630000000
0!
0'
0/
#423640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#423650000000
0!
0'
0/
#423660000000
1!
1'
1/
#423670000000
0!
1"
0'
1(
0/
10
#423680000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#423690000000
0!
1$
0'
1+
0/
#423700000000
1!
1'
1/
#423710000000
0!
0'
0/
#423720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#423730000000
0!
0'
0/
#423740000000
1!
1'
1/
#423750000000
0!
0'
0/
#423760000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#423770000000
0!
0'
0/
#423780000000
1!
1'
1/
#423790000000
0!
0'
0/
#423800000000
1!
1'
1/
#423810000000
0!
0'
0/
#423820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#423830000000
0!
0'
0/
#423840000000
1!
1'
1/
#423850000000
0!
0'
0/
#423860000000
1!
1'
1/
#423870000000
0!
0'
0/
#423880000000
1!
1'
1/
#423890000000
0!
0'
0/
#423900000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#423910000000
0!
0'
0/
#423920000000
1!
1'
1/
#423930000000
0!
0'
0/
#423940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#423950000000
0!
0'
0/
#423960000000
1!
1'
1/
#423970000000
0!
0'
0/
#423980000000
#423990000000
1!
1'
1/
#424000000000
0!
0'
0/
#424010000000
1!
1'
1/
#424020000000
0!
1"
0'
1(
0/
10
#424030000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#424040000000
0!
0'
0/
#424050000000
1!
1'
1/
#424060000000
0!
0'
0/
#424070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#424080000000
0!
0'
0/
#424090000000
1!
1'
1/
#424100000000
0!
1"
0'
1(
0/
10
#424110000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#424120000000
0!
1$
0'
1+
0/
#424130000000
1!
1'
1/
#424140000000
0!
0'
0/
#424150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#424160000000
0!
0'
0/
#424170000000
1!
1'
1/
#424180000000
0!
0'
0/
#424190000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#424200000000
0!
0'
0/
#424210000000
1!
1'
1/
#424220000000
0!
0'
0/
#424230000000
1!
1'
1/
#424240000000
0!
0'
0/
#424250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#424260000000
0!
0'
0/
#424270000000
1!
1'
1/
#424280000000
0!
0'
0/
#424290000000
1!
1'
1/
#424300000000
0!
0'
0/
#424310000000
1!
1'
1/
#424320000000
0!
0'
0/
#424330000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#424340000000
0!
0'
0/
#424350000000
1!
1'
1/
#424360000000
0!
0'
0/
#424370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#424380000000
0!
0'
0/
#424390000000
1!
1'
1/
#424400000000
0!
0'
0/
#424410000000
#424420000000
1!
1'
1/
#424430000000
0!
0'
0/
#424440000000
1!
1'
1/
#424450000000
0!
1"
0'
1(
0/
10
#424460000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#424470000000
0!
0'
0/
#424480000000
1!
1'
1/
#424490000000
0!
0'
0/
#424500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#424510000000
0!
0'
0/
#424520000000
1!
1'
1/
#424530000000
0!
1"
0'
1(
0/
10
#424540000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#424550000000
0!
1$
0'
1+
0/
#424560000000
1!
1'
1/
#424570000000
0!
0'
0/
#424580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#424590000000
0!
0'
0/
#424600000000
1!
1'
1/
#424610000000
0!
0'
0/
#424620000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#424630000000
0!
0'
0/
#424640000000
1!
1'
1/
#424650000000
0!
0'
0/
#424660000000
1!
1'
1/
#424670000000
0!
0'
0/
#424680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#424690000000
0!
0'
0/
#424700000000
1!
1'
1/
#424710000000
0!
0'
0/
#424720000000
1!
1'
1/
#424730000000
0!
0'
0/
#424740000000
1!
1'
1/
#424750000000
0!
0'
0/
#424760000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#424770000000
0!
0'
0/
#424780000000
1!
1'
1/
#424790000000
0!
0'
0/
#424800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#424810000000
0!
0'
0/
#424820000000
1!
1'
1/
#424830000000
0!
0'
0/
#424840000000
#424850000000
1!
1'
1/
#424860000000
0!
0'
0/
#424870000000
1!
1'
1/
#424880000000
0!
1"
0'
1(
0/
10
#424890000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#424900000000
0!
0'
0/
#424910000000
1!
1'
1/
#424920000000
0!
0'
0/
#424930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#424940000000
0!
0'
0/
#424950000000
1!
1'
1/
#424960000000
0!
1"
0'
1(
0/
10
#424970000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#424980000000
0!
1$
0'
1+
0/
#424990000000
1!
1'
1/
#425000000000
0!
0'
0/
#425010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#425020000000
0!
0'
0/
#425030000000
1!
1'
1/
#425040000000
0!
0'
0/
#425050000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#425060000000
0!
0'
0/
#425070000000
1!
1'
1/
#425080000000
0!
0'
0/
#425090000000
1!
1'
1/
#425100000000
0!
0'
0/
#425110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#425120000000
0!
0'
0/
#425130000000
1!
1'
1/
#425140000000
0!
0'
0/
#425150000000
1!
1'
1/
#425160000000
0!
0'
0/
#425170000000
1!
1'
1/
#425180000000
0!
0'
0/
#425190000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#425200000000
0!
0'
0/
#425210000000
1!
1'
1/
#425220000000
0!
0'
0/
#425230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#425240000000
0!
0'
0/
#425250000000
1!
1'
1/
#425260000000
0!
0'
0/
#425270000000
#425280000000
1!
1'
1/
#425290000000
0!
0'
0/
#425300000000
1!
1'
1/
#425310000000
0!
1"
0'
1(
0/
10
#425320000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#425330000000
0!
0'
0/
#425340000000
1!
1'
1/
#425350000000
0!
0'
0/
#425360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#425370000000
0!
0'
0/
#425380000000
1!
1'
1/
#425390000000
0!
1"
0'
1(
0/
10
#425400000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#425410000000
0!
1$
0'
1+
0/
#425420000000
1!
1'
1/
#425430000000
0!
0'
0/
#425440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#425450000000
0!
0'
0/
#425460000000
1!
1'
1/
#425470000000
0!
0'
0/
#425480000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#425490000000
0!
0'
0/
#425500000000
1!
1'
1/
#425510000000
0!
0'
0/
#425520000000
1!
1'
1/
#425530000000
0!
0'
0/
#425540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#425550000000
0!
0'
0/
#425560000000
1!
1'
1/
#425570000000
0!
0'
0/
#425580000000
1!
1'
1/
#425590000000
0!
0'
0/
#425600000000
1!
1'
1/
#425610000000
0!
0'
0/
#425620000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#425630000000
0!
0'
0/
#425640000000
1!
1'
1/
#425650000000
0!
0'
0/
#425660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#425670000000
0!
0'
0/
#425680000000
1!
1'
1/
#425690000000
0!
0'
0/
#425700000000
#425710000000
1!
1'
1/
#425720000000
0!
0'
0/
#425730000000
1!
1'
1/
#425740000000
0!
1"
0'
1(
0/
10
#425750000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#425760000000
0!
0'
0/
#425770000000
1!
1'
1/
#425780000000
0!
0'
0/
#425790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#425800000000
0!
0'
0/
#425810000000
1!
1'
1/
#425820000000
0!
1"
0'
1(
0/
10
#425830000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#425840000000
0!
1$
0'
1+
0/
#425850000000
1!
1'
1/
#425860000000
0!
0'
0/
#425870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#425880000000
0!
0'
0/
#425890000000
1!
1'
1/
#425900000000
0!
0'
0/
#425910000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#425920000000
0!
0'
0/
#425930000000
1!
1'
1/
#425940000000
0!
0'
0/
#425950000000
1!
1'
1/
#425960000000
0!
0'
0/
#425970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#425980000000
0!
0'
0/
#425990000000
1!
1'
1/
#426000000000
0!
0'
0/
#426010000000
1!
1'
1/
#426020000000
0!
0'
0/
#426030000000
1!
1'
1/
#426040000000
0!
0'
0/
#426050000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#426060000000
0!
0'
0/
#426070000000
1!
1'
1/
#426080000000
0!
0'
0/
#426090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#426100000000
0!
0'
0/
#426110000000
1!
1'
1/
#426120000000
0!
0'
0/
#426130000000
#426140000000
1!
1'
1/
#426150000000
0!
0'
0/
#426160000000
1!
1'
1/
#426170000000
0!
1"
0'
1(
0/
10
#426180000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#426190000000
0!
0'
0/
#426200000000
1!
1'
1/
#426210000000
0!
0'
0/
#426220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#426230000000
0!
0'
0/
#426240000000
1!
1'
1/
#426250000000
0!
1"
0'
1(
0/
10
#426260000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#426270000000
0!
1$
0'
1+
0/
#426280000000
1!
1'
1/
#426290000000
0!
0'
0/
#426300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#426310000000
0!
0'
0/
#426320000000
1!
1'
1/
#426330000000
0!
0'
0/
#426340000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#426350000000
0!
0'
0/
#426360000000
1!
1'
1/
#426370000000
0!
0'
0/
#426380000000
1!
1'
1/
#426390000000
0!
0'
0/
#426400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#426410000000
0!
0'
0/
#426420000000
1!
1'
1/
#426430000000
0!
0'
0/
#426440000000
1!
1'
1/
#426450000000
0!
0'
0/
#426460000000
1!
1'
1/
#426470000000
0!
0'
0/
#426480000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#426490000000
0!
0'
0/
#426500000000
1!
1'
1/
#426510000000
0!
0'
0/
#426520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#426530000000
0!
0'
0/
#426540000000
1!
1'
1/
#426550000000
0!
0'
0/
#426560000000
#426570000000
1!
1'
1/
#426580000000
0!
0'
0/
#426590000000
1!
1'
1/
#426600000000
0!
1"
0'
1(
0/
10
#426610000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#426620000000
0!
0'
0/
#426630000000
1!
1'
1/
#426640000000
0!
0'
0/
#426650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#426660000000
0!
0'
0/
#426670000000
1!
1'
1/
#426680000000
0!
1"
0'
1(
0/
10
#426690000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#426700000000
0!
1$
0'
1+
0/
#426710000000
1!
1'
1/
#426720000000
0!
0'
0/
#426730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#426740000000
0!
0'
0/
#426750000000
1!
1'
1/
#426760000000
0!
0'
0/
#426770000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#426780000000
0!
0'
0/
#426790000000
1!
1'
1/
#426800000000
0!
0'
0/
#426810000000
1!
1'
1/
#426820000000
0!
0'
0/
#426830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#426840000000
0!
0'
0/
#426850000000
1!
1'
1/
#426860000000
0!
0'
0/
#426870000000
1!
1'
1/
#426880000000
0!
0'
0/
#426890000000
1!
1'
1/
#426900000000
0!
0'
0/
#426910000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#426920000000
0!
0'
0/
#426930000000
1!
1'
1/
#426940000000
0!
0'
0/
#426950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#426960000000
0!
0'
0/
#426970000000
1!
1'
1/
#426980000000
0!
0'
0/
#426990000000
#427000000000
1!
1'
1/
#427010000000
0!
0'
0/
#427020000000
1!
1'
1/
#427030000000
0!
1"
0'
1(
0/
10
#427040000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#427050000000
0!
0'
0/
#427060000000
1!
1'
1/
#427070000000
0!
0'
0/
#427080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#427090000000
0!
0'
0/
#427100000000
1!
1'
1/
#427110000000
0!
1"
0'
1(
0/
10
#427120000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#427130000000
0!
1$
0'
1+
0/
#427140000000
1!
1'
1/
#427150000000
0!
0'
0/
#427160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#427170000000
0!
0'
0/
#427180000000
1!
1'
1/
#427190000000
0!
0'
0/
#427200000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#427210000000
0!
0'
0/
#427220000000
1!
1'
1/
#427230000000
0!
0'
0/
#427240000000
1!
1'
1/
#427250000000
0!
0'
0/
#427260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#427270000000
0!
0'
0/
#427280000000
1!
1'
1/
#427290000000
0!
0'
0/
#427300000000
1!
1'
1/
#427310000000
0!
0'
0/
#427320000000
1!
1'
1/
#427330000000
0!
0'
0/
#427340000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#427350000000
0!
0'
0/
#427360000000
1!
1'
1/
#427370000000
0!
0'
0/
#427380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#427390000000
0!
0'
0/
#427400000000
1!
1'
1/
#427410000000
0!
0'
0/
#427420000000
#427430000000
1!
1'
1/
#427440000000
0!
0'
0/
#427450000000
1!
1'
1/
#427460000000
0!
1"
0'
1(
0/
10
#427470000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#427480000000
0!
0'
0/
#427490000000
1!
1'
1/
#427500000000
0!
0'
0/
#427510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#427520000000
0!
0'
0/
#427530000000
1!
1'
1/
#427540000000
0!
1"
0'
1(
0/
10
#427550000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#427560000000
0!
1$
0'
1+
0/
#427570000000
1!
1'
1/
#427580000000
0!
0'
0/
#427590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#427600000000
0!
0'
0/
#427610000000
1!
1'
1/
#427620000000
0!
0'
0/
#427630000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#427640000000
0!
0'
0/
#427650000000
1!
1'
1/
#427660000000
0!
0'
0/
#427670000000
1!
1'
1/
#427680000000
0!
0'
0/
#427690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#427700000000
0!
0'
0/
#427710000000
1!
1'
1/
#427720000000
0!
0'
0/
#427730000000
1!
1'
1/
#427740000000
0!
0'
0/
#427750000000
1!
1'
1/
#427760000000
0!
0'
0/
#427770000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#427780000000
0!
0'
0/
#427790000000
1!
1'
1/
#427800000000
0!
0'
0/
#427810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#427820000000
0!
0'
0/
#427830000000
1!
1'
1/
#427840000000
0!
0'
0/
#427850000000
#427860000000
1!
1'
1/
#427870000000
0!
0'
0/
#427880000000
1!
1'
1/
#427890000000
0!
1"
0'
1(
0/
10
#427900000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#427910000000
0!
0'
0/
#427920000000
1!
1'
1/
#427930000000
0!
0'
0/
#427940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#427950000000
0!
0'
0/
#427960000000
1!
1'
1/
#427970000000
0!
1"
0'
1(
0/
10
#427980000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#427990000000
0!
1$
0'
1+
0/
#428000000000
1!
1'
1/
#428010000000
0!
0'
0/
#428020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#428030000000
0!
0'
0/
#428040000000
1!
1'
1/
#428050000000
0!
0'
0/
#428060000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#428070000000
0!
0'
0/
#428080000000
1!
1'
1/
#428090000000
0!
0'
0/
#428100000000
1!
1'
1/
#428110000000
0!
0'
0/
#428120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#428130000000
0!
0'
0/
#428140000000
1!
1'
1/
#428150000000
0!
0'
0/
#428160000000
1!
1'
1/
#428170000000
0!
0'
0/
#428180000000
1!
1'
1/
#428190000000
0!
0'
0/
#428200000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#428210000000
0!
0'
0/
#428220000000
1!
1'
1/
#428230000000
0!
0'
0/
#428240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#428250000000
0!
0'
0/
#428260000000
1!
1'
1/
#428270000000
0!
0'
0/
#428280000000
#428290000000
1!
1'
1/
#428300000000
0!
0'
0/
#428310000000
1!
1'
1/
#428320000000
0!
1"
0'
1(
0/
10
#428330000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#428340000000
0!
0'
0/
#428350000000
1!
1'
1/
#428360000000
0!
0'
0/
#428370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#428380000000
0!
0'
0/
#428390000000
1!
1'
1/
#428400000000
0!
1"
0'
1(
0/
10
#428410000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#428420000000
0!
1$
0'
1+
0/
#428430000000
1!
1'
1/
#428440000000
0!
0'
0/
#428450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#428460000000
0!
0'
0/
#428470000000
1!
1'
1/
#428480000000
0!
0'
0/
#428490000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#428500000000
0!
0'
0/
#428510000000
1!
1'
1/
#428520000000
0!
0'
0/
#428530000000
1!
1'
1/
#428540000000
0!
0'
0/
#428550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#428560000000
0!
0'
0/
#428570000000
1!
1'
1/
#428580000000
0!
0'
0/
#428590000000
1!
1'
1/
#428600000000
0!
0'
0/
#428610000000
1!
1'
1/
#428620000000
0!
0'
0/
#428630000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#428640000000
0!
0'
0/
#428650000000
1!
1'
1/
#428660000000
0!
0'
0/
#428670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#428680000000
0!
0'
0/
#428690000000
1!
1'
1/
#428700000000
0!
0'
0/
#428710000000
#428720000000
1!
1'
1/
#428730000000
0!
0'
0/
#428740000000
1!
1'
1/
#428750000000
0!
1"
0'
1(
0/
10
#428760000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#428770000000
0!
0'
0/
#428780000000
1!
1'
1/
#428790000000
0!
0'
0/
#428800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#428810000000
0!
0'
0/
#428820000000
1!
1'
1/
#428830000000
0!
1"
0'
1(
0/
10
#428840000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#428850000000
0!
1$
0'
1+
0/
#428860000000
1!
1'
1/
#428870000000
0!
0'
0/
#428880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#428890000000
0!
0'
0/
#428900000000
1!
1'
1/
#428910000000
0!
0'
0/
#428920000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#428930000000
0!
0'
0/
#428940000000
1!
1'
1/
#428950000000
0!
0'
0/
#428960000000
1!
1'
1/
#428970000000
0!
0'
0/
#428980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#428990000000
0!
0'
0/
#429000000000
1!
1'
1/
#429010000000
0!
0'
0/
#429020000000
1!
1'
1/
#429030000000
0!
0'
0/
#429040000000
1!
1'
1/
#429050000000
0!
0'
0/
#429060000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#429070000000
0!
0'
0/
#429080000000
1!
1'
1/
#429090000000
0!
0'
0/
#429100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#429110000000
0!
0'
0/
#429120000000
1!
1'
1/
#429130000000
0!
0'
0/
#429140000000
#429150000000
1!
1'
1/
#429160000000
0!
0'
0/
#429170000000
1!
1'
1/
#429180000000
0!
1"
0'
1(
0/
10
#429190000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#429200000000
0!
0'
0/
#429210000000
1!
1'
1/
#429220000000
0!
0'
0/
#429230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#429240000000
0!
0'
0/
#429250000000
1!
1'
1/
#429260000000
0!
1"
0'
1(
0/
10
#429270000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#429280000000
0!
1$
0'
1+
0/
#429290000000
1!
1'
1/
#429300000000
0!
0'
0/
#429310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#429320000000
0!
0'
0/
#429330000000
1!
1'
1/
#429340000000
0!
0'
0/
#429350000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#429360000000
0!
0'
0/
#429370000000
1!
1'
1/
#429380000000
0!
0'
0/
#429390000000
1!
1'
1/
#429400000000
0!
0'
0/
#429410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#429420000000
0!
0'
0/
#429430000000
1!
1'
1/
#429440000000
0!
0'
0/
#429450000000
1!
1'
1/
#429460000000
0!
0'
0/
#429470000000
1!
1'
1/
#429480000000
0!
0'
0/
#429490000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#429500000000
0!
0'
0/
#429510000000
1!
1'
1/
#429520000000
0!
0'
0/
#429530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#429540000000
0!
0'
0/
#429550000000
1!
1'
1/
#429560000000
0!
0'
0/
#429570000000
#429580000000
1!
1'
1/
#429590000000
0!
0'
0/
#429600000000
1!
1'
1/
#429610000000
0!
1"
0'
1(
0/
10
#429620000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#429630000000
0!
0'
0/
#429640000000
1!
1'
1/
#429650000000
0!
0'
0/
#429660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#429670000000
0!
0'
0/
#429680000000
1!
1'
1/
#429690000000
0!
1"
0'
1(
0/
10
#429700000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#429710000000
0!
1$
0'
1+
0/
#429720000000
1!
1'
1/
#429730000000
0!
0'
0/
#429740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#429750000000
0!
0'
0/
#429760000000
1!
1'
1/
#429770000000
0!
0'
0/
#429780000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#429790000000
0!
0'
0/
#429800000000
1!
1'
1/
#429810000000
0!
0'
0/
#429820000000
1!
1'
1/
#429830000000
0!
0'
0/
#429840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#429850000000
0!
0'
0/
#429860000000
1!
1'
1/
#429870000000
0!
0'
0/
#429880000000
1!
1'
1/
#429890000000
0!
0'
0/
#429900000000
1!
1'
1/
#429910000000
0!
0'
0/
#429920000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#429930000000
0!
0'
0/
#429940000000
1!
1'
1/
#429950000000
0!
0'
0/
#429960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#429970000000
0!
0'
0/
#429980000000
1!
1'
1/
#429990000000
0!
0'
0/
#430000000000
#430010000000
1!
1'
1/
#430020000000
0!
0'
0/
#430030000000
1!
1'
1/
#430040000000
0!
1"
0'
1(
0/
10
#430050000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#430060000000
0!
0'
0/
#430070000000
1!
1'
1/
#430080000000
0!
0'
0/
#430090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#430100000000
0!
0'
0/
#430110000000
1!
1'
1/
#430120000000
0!
1"
0'
1(
0/
10
#430130000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#430140000000
0!
1$
0'
1+
0/
#430150000000
1!
1'
1/
#430160000000
0!
0'
0/
#430170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#430180000000
0!
0'
0/
#430190000000
1!
1'
1/
#430200000000
0!
0'
0/
#430210000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#430220000000
0!
0'
0/
#430230000000
1!
1'
1/
#430240000000
0!
0'
0/
#430250000000
1!
1'
1/
#430260000000
0!
0'
0/
#430270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#430280000000
0!
0'
0/
#430290000000
1!
1'
1/
#430300000000
0!
0'
0/
#430310000000
1!
1'
1/
#430320000000
0!
0'
0/
#430330000000
1!
1'
1/
#430340000000
0!
0'
0/
#430350000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#430360000000
0!
0'
0/
#430370000000
1!
1'
1/
#430380000000
0!
0'
0/
#430390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#430400000000
0!
0'
0/
#430410000000
1!
1'
1/
#430420000000
0!
0'
0/
#430430000000
#430440000000
1!
1'
1/
#430450000000
0!
0'
0/
#430460000000
1!
1'
1/
#430470000000
0!
1"
0'
1(
0/
10
#430480000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#430490000000
0!
0'
0/
#430500000000
1!
1'
1/
#430510000000
0!
0'
0/
#430520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#430530000000
0!
0'
0/
#430540000000
1!
1'
1/
#430550000000
0!
1"
0'
1(
0/
10
#430560000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#430570000000
0!
1$
0'
1+
0/
#430580000000
1!
1'
1/
#430590000000
0!
0'
0/
#430600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#430610000000
0!
0'
0/
#430620000000
1!
1'
1/
#430630000000
0!
0'
0/
#430640000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#430650000000
0!
0'
0/
#430660000000
1!
1'
1/
#430670000000
0!
0'
0/
#430680000000
1!
1'
1/
#430690000000
0!
0'
0/
#430700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#430710000000
0!
0'
0/
#430720000000
1!
1'
1/
#430730000000
0!
0'
0/
#430740000000
1!
1'
1/
#430750000000
0!
0'
0/
#430760000000
1!
1'
1/
#430770000000
0!
0'
0/
#430780000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#430790000000
0!
0'
0/
#430800000000
1!
1'
1/
#430810000000
0!
0'
0/
#430820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#430830000000
0!
0'
0/
#430840000000
1!
1'
1/
#430850000000
0!
0'
0/
#430860000000
#430870000000
1!
1'
1/
#430880000000
0!
0'
0/
#430890000000
1!
1'
1/
#430900000000
0!
1"
0'
1(
0/
10
#430910000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#430920000000
0!
0'
0/
#430930000000
1!
1'
1/
#430940000000
0!
0'
0/
#430950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#430960000000
0!
0'
0/
#430970000000
1!
1'
1/
#430980000000
0!
1"
0'
1(
0/
10
#430990000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#431000000000
0!
1$
0'
1+
0/
#431010000000
1!
1'
1/
#431020000000
0!
0'
0/
#431030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#431040000000
0!
0'
0/
#431050000000
1!
1'
1/
#431060000000
0!
0'
0/
#431070000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#431080000000
0!
0'
0/
#431090000000
1!
1'
1/
#431100000000
0!
0'
0/
#431110000000
1!
1'
1/
#431120000000
0!
0'
0/
#431130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#431140000000
0!
0'
0/
#431150000000
1!
1'
1/
#431160000000
0!
0'
0/
#431170000000
1!
1'
1/
#431180000000
0!
0'
0/
#431190000000
1!
1'
1/
#431200000000
0!
0'
0/
#431210000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#431220000000
0!
0'
0/
#431230000000
1!
1'
1/
#431240000000
0!
0'
0/
#431250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#431260000000
0!
0'
0/
#431270000000
1!
1'
1/
#431280000000
0!
0'
0/
#431290000000
#431300000000
1!
1'
1/
#431310000000
0!
0'
0/
#431320000000
1!
1'
1/
#431330000000
0!
1"
0'
1(
0/
10
#431340000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#431350000000
0!
0'
0/
#431360000000
1!
1'
1/
#431370000000
0!
0'
0/
#431380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#431390000000
0!
0'
0/
#431400000000
1!
1'
1/
#431410000000
0!
1"
0'
1(
0/
10
#431420000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#431430000000
0!
1$
0'
1+
0/
#431440000000
1!
1'
1/
#431450000000
0!
0'
0/
#431460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#431470000000
0!
0'
0/
#431480000000
1!
1'
1/
#431490000000
0!
0'
0/
#431500000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#431510000000
0!
0'
0/
#431520000000
1!
1'
1/
#431530000000
0!
0'
0/
#431540000000
1!
1'
1/
#431550000000
0!
0'
0/
#431560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#431570000000
0!
0'
0/
#431580000000
1!
1'
1/
#431590000000
0!
0'
0/
#431600000000
1!
1'
1/
#431610000000
0!
0'
0/
#431620000000
1!
1'
1/
#431630000000
0!
0'
0/
#431640000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#431650000000
0!
0'
0/
#431660000000
1!
1'
1/
#431670000000
0!
0'
0/
#431680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#431690000000
0!
0'
0/
#431700000000
1!
1'
1/
#431710000000
0!
0'
0/
#431720000000
#431730000000
1!
1'
1/
#431740000000
0!
0'
0/
#431750000000
1!
1'
1/
#431760000000
0!
1"
0'
1(
0/
10
#431770000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#431780000000
0!
0'
0/
#431790000000
1!
1'
1/
#431800000000
0!
0'
0/
#431810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#431820000000
0!
0'
0/
#431830000000
1!
1'
1/
#431840000000
0!
1"
0'
1(
0/
10
#431850000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#431860000000
0!
1$
0'
1+
0/
#431870000000
1!
1'
1/
#431880000000
0!
0'
0/
#431890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#431900000000
0!
0'
0/
#431910000000
1!
1'
1/
#431920000000
0!
0'
0/
#431930000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#431940000000
0!
0'
0/
#431950000000
1!
1'
1/
#431960000000
0!
0'
0/
#431970000000
1!
1'
1/
#431980000000
0!
0'
0/
#431990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#432000000000
0!
0'
0/
#432010000000
1!
1'
1/
#432020000000
0!
0'
0/
#432030000000
1!
1'
1/
#432040000000
0!
0'
0/
#432050000000
1!
1'
1/
#432060000000
0!
0'
0/
#432070000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#432080000000
0!
0'
0/
#432090000000
1!
1'
1/
#432100000000
0!
0'
0/
#432110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#432120000000
0!
0'
0/
#432130000000
1!
1'
1/
#432140000000
0!
0'
0/
#432150000000
#432160000000
1!
1'
1/
#432170000000
0!
0'
0/
#432180000000
1!
1'
1/
#432190000000
0!
1"
0'
1(
0/
10
#432200000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#432210000000
0!
0'
0/
#432220000000
1!
1'
1/
#432230000000
0!
0'
0/
#432240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#432250000000
0!
0'
0/
#432260000000
1!
1'
1/
#432270000000
0!
1"
0'
1(
0/
10
#432280000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#432290000000
0!
1$
0'
1+
0/
#432300000000
1!
1'
1/
#432310000000
0!
0'
0/
#432320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#432330000000
0!
0'
0/
#432340000000
1!
1'
1/
#432350000000
0!
0'
0/
#432360000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#432370000000
0!
0'
0/
#432380000000
1!
1'
1/
#432390000000
0!
0'
0/
#432400000000
1!
1'
1/
#432410000000
0!
0'
0/
#432420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#432430000000
0!
0'
0/
#432440000000
1!
1'
1/
#432450000000
0!
0'
0/
#432460000000
1!
1'
1/
#432470000000
0!
0'
0/
#432480000000
1!
1'
1/
#432490000000
0!
0'
0/
#432500000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#432510000000
0!
0'
0/
#432520000000
1!
1'
1/
#432530000000
0!
0'
0/
#432540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#432550000000
0!
0'
0/
#432560000000
1!
1'
1/
#432570000000
0!
0'
0/
#432580000000
#432590000000
1!
1'
1/
#432600000000
0!
0'
0/
#432610000000
1!
1'
1/
#432620000000
0!
1"
0'
1(
0/
10
#432630000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#432640000000
0!
0'
0/
#432650000000
1!
1'
1/
#432660000000
0!
0'
0/
#432670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#432680000000
0!
0'
0/
#432690000000
1!
1'
1/
#432700000000
0!
1"
0'
1(
0/
10
#432710000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#432720000000
0!
1$
0'
1+
0/
#432730000000
1!
1'
1/
#432740000000
0!
0'
0/
#432750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#432760000000
0!
0'
0/
#432770000000
1!
1'
1/
#432780000000
0!
0'
0/
#432790000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#432800000000
0!
0'
0/
#432810000000
1!
1'
1/
#432820000000
0!
0'
0/
#432830000000
1!
1'
1/
#432840000000
0!
0'
0/
#432850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#432860000000
0!
0'
0/
#432870000000
1!
1'
1/
#432880000000
0!
0'
0/
#432890000000
1!
1'
1/
#432900000000
0!
0'
0/
#432910000000
1!
1'
1/
#432920000000
0!
0'
0/
#432930000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#432940000000
0!
0'
0/
#432950000000
1!
1'
1/
#432960000000
0!
0'
0/
#432970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#432980000000
0!
0'
0/
#432990000000
1!
1'
1/
#433000000000
0!
0'
0/
#433010000000
#433020000000
1!
1'
1/
#433030000000
0!
0'
0/
#433040000000
1!
1'
1/
#433050000000
0!
1"
0'
1(
0/
10
#433060000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#433070000000
0!
0'
0/
#433080000000
1!
1'
1/
#433090000000
0!
0'
0/
#433100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#433110000000
0!
0'
0/
#433120000000
1!
1'
1/
#433130000000
0!
1"
0'
1(
0/
10
#433140000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#433150000000
0!
1$
0'
1+
0/
#433160000000
1!
1'
1/
#433170000000
0!
0'
0/
#433180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#433190000000
0!
0'
0/
#433200000000
1!
1'
1/
#433210000000
0!
0'
0/
#433220000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#433230000000
0!
0'
0/
#433240000000
1!
1'
1/
#433250000000
0!
0'
0/
#433260000000
1!
1'
1/
#433270000000
0!
0'
0/
#433280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#433290000000
0!
0'
0/
#433300000000
1!
1'
1/
#433310000000
0!
0'
0/
#433320000000
1!
1'
1/
#433330000000
0!
0'
0/
#433340000000
1!
1'
1/
#433350000000
0!
0'
0/
#433360000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#433370000000
0!
0'
0/
#433380000000
1!
1'
1/
#433390000000
0!
0'
0/
#433400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#433410000000
0!
0'
0/
#433420000000
1!
1'
1/
#433430000000
0!
0'
0/
#433440000000
#433450000000
1!
1'
1/
#433460000000
0!
0'
0/
#433470000000
1!
1'
1/
#433480000000
0!
1"
0'
1(
0/
10
#433490000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#433500000000
0!
0'
0/
#433510000000
1!
1'
1/
#433520000000
0!
0'
0/
#433530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#433540000000
0!
0'
0/
#433550000000
1!
1'
1/
#433560000000
0!
1"
0'
1(
0/
10
#433570000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#433580000000
0!
1$
0'
1+
0/
#433590000000
1!
1'
1/
#433600000000
0!
0'
0/
#433610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#433620000000
0!
0'
0/
#433630000000
1!
1'
1/
#433640000000
0!
0'
0/
#433650000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#433660000000
0!
0'
0/
#433670000000
1!
1'
1/
#433680000000
0!
0'
0/
#433690000000
1!
1'
1/
#433700000000
0!
0'
0/
#433710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#433720000000
0!
0'
0/
#433730000000
1!
1'
1/
#433740000000
0!
0'
0/
#433750000000
1!
1'
1/
#433760000000
0!
0'
0/
#433770000000
1!
1'
1/
#433780000000
0!
0'
0/
#433790000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#433800000000
0!
0'
0/
#433810000000
1!
1'
1/
#433820000000
0!
0'
0/
#433830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#433840000000
0!
0'
0/
#433850000000
1!
1'
1/
#433860000000
0!
0'
0/
#433870000000
#433880000000
1!
1'
1/
#433890000000
0!
0'
0/
#433900000000
1!
1'
1/
#433910000000
0!
1"
0'
1(
0/
10
#433920000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#433930000000
0!
0'
0/
#433940000000
1!
1'
1/
#433950000000
0!
0'
0/
#433960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#433970000000
0!
0'
0/
#433980000000
1!
1'
1/
#433990000000
0!
1"
0'
1(
0/
10
#434000000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#434010000000
0!
1$
0'
1+
0/
#434020000000
1!
1'
1/
#434030000000
0!
0'
0/
#434040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#434050000000
0!
0'
0/
#434060000000
1!
1'
1/
#434070000000
0!
0'
0/
#434080000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#434090000000
0!
0'
0/
#434100000000
1!
1'
1/
#434110000000
0!
0'
0/
#434120000000
1!
1'
1/
#434130000000
0!
0'
0/
#434140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#434150000000
0!
0'
0/
#434160000000
1!
1'
1/
#434170000000
0!
0'
0/
#434180000000
1!
1'
1/
#434190000000
0!
0'
0/
#434200000000
1!
1'
1/
#434210000000
0!
0'
0/
#434220000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#434230000000
0!
0'
0/
#434240000000
1!
1'
1/
#434250000000
0!
0'
0/
#434260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#434270000000
0!
0'
0/
#434280000000
1!
1'
1/
#434290000000
0!
0'
0/
#434300000000
#434310000000
1!
1'
1/
#434320000000
0!
0'
0/
#434330000000
1!
1'
1/
#434340000000
0!
1"
0'
1(
0/
10
#434350000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#434360000000
0!
0'
0/
#434370000000
1!
1'
1/
#434380000000
0!
0'
0/
#434390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#434400000000
0!
0'
0/
#434410000000
1!
1'
1/
#434420000000
0!
1"
0'
1(
0/
10
#434430000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#434440000000
0!
1$
0'
1+
0/
#434450000000
1!
1'
1/
#434460000000
0!
0'
0/
#434470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#434480000000
0!
0'
0/
#434490000000
1!
1'
1/
#434500000000
0!
0'
0/
#434510000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#434520000000
0!
0'
0/
#434530000000
1!
1'
1/
#434540000000
0!
0'
0/
#434550000000
1!
1'
1/
#434560000000
0!
0'
0/
#434570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#434580000000
0!
0'
0/
#434590000000
1!
1'
1/
#434600000000
0!
0'
0/
#434610000000
1!
1'
1/
#434620000000
0!
0'
0/
#434630000000
1!
1'
1/
#434640000000
0!
0'
0/
#434650000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#434660000000
0!
0'
0/
#434670000000
1!
1'
1/
#434680000000
0!
0'
0/
#434690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#434700000000
0!
0'
0/
#434710000000
1!
1'
1/
#434720000000
0!
0'
0/
#434730000000
#434740000000
1!
1'
1/
#434750000000
0!
0'
0/
#434760000000
1!
1'
1/
#434770000000
0!
1"
0'
1(
0/
10
#434780000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#434790000000
0!
0'
0/
#434800000000
1!
1'
1/
#434810000000
0!
0'
0/
#434820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#434830000000
0!
0'
0/
#434840000000
1!
1'
1/
#434850000000
0!
1"
0'
1(
0/
10
#434860000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#434870000000
0!
1$
0'
1+
0/
#434880000000
1!
1'
1/
#434890000000
0!
0'
0/
#434900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#434910000000
0!
0'
0/
#434920000000
1!
1'
1/
#434930000000
0!
0'
0/
#434940000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#434950000000
0!
0'
0/
#434960000000
1!
1'
1/
#434970000000
0!
0'
0/
#434980000000
1!
1'
1/
#434990000000
0!
0'
0/
#435000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#435010000000
0!
0'
0/
#435020000000
1!
1'
1/
#435030000000
0!
0'
0/
#435040000000
1!
1'
1/
#435050000000
0!
0'
0/
#435060000000
1!
1'
1/
#435070000000
0!
0'
0/
#435080000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#435090000000
0!
0'
0/
#435100000000
1!
1'
1/
#435110000000
0!
0'
0/
#435120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#435130000000
0!
0'
0/
#435140000000
1!
1'
1/
#435150000000
0!
0'
0/
#435160000000
#435170000000
1!
1'
1/
#435180000000
0!
0'
0/
#435190000000
1!
1'
1/
#435200000000
0!
1"
0'
1(
0/
10
#435210000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#435220000000
0!
0'
0/
#435230000000
1!
1'
1/
#435240000000
0!
0'
0/
#435250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#435260000000
0!
0'
0/
#435270000000
1!
1'
1/
#435280000000
0!
1"
0'
1(
0/
10
#435290000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#435300000000
0!
1$
0'
1+
0/
#435310000000
1!
1'
1/
#435320000000
0!
0'
0/
#435330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#435340000000
0!
0'
0/
#435350000000
1!
1'
1/
#435360000000
0!
0'
0/
#435370000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#435380000000
0!
0'
0/
#435390000000
1!
1'
1/
#435400000000
0!
0'
0/
#435410000000
1!
1'
1/
#435420000000
0!
0'
0/
#435430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#435440000000
0!
0'
0/
#435450000000
1!
1'
1/
#435460000000
0!
0'
0/
#435470000000
1!
1'
1/
#435480000000
0!
0'
0/
#435490000000
1!
1'
1/
#435500000000
0!
0'
0/
#435510000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#435520000000
0!
0'
0/
#435530000000
1!
1'
1/
#435540000000
0!
0'
0/
#435550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#435560000000
0!
0'
0/
#435570000000
1!
1'
1/
#435580000000
0!
0'
0/
#435590000000
#435600000000
1!
1'
1/
#435610000000
0!
0'
0/
#435620000000
1!
1'
1/
#435630000000
0!
1"
0'
1(
0/
10
#435640000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#435650000000
0!
0'
0/
#435660000000
1!
1'
1/
#435670000000
0!
0'
0/
#435680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#435690000000
0!
0'
0/
#435700000000
1!
1'
1/
#435710000000
0!
1"
0'
1(
0/
10
#435720000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#435730000000
0!
1$
0'
1+
0/
#435740000000
1!
1'
1/
#435750000000
0!
0'
0/
#435760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#435770000000
0!
0'
0/
#435780000000
1!
1'
1/
#435790000000
0!
0'
0/
#435800000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#435810000000
0!
0'
0/
#435820000000
1!
1'
1/
#435830000000
0!
0'
0/
#435840000000
1!
1'
1/
#435850000000
0!
0'
0/
#435860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#435870000000
0!
0'
0/
#435880000000
1!
1'
1/
#435890000000
0!
0'
0/
#435900000000
1!
1'
1/
#435910000000
0!
0'
0/
#435920000000
1!
1'
1/
#435930000000
0!
0'
0/
#435940000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#435950000000
0!
0'
0/
#435960000000
1!
1'
1/
#435970000000
0!
0'
0/
#435980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#435990000000
0!
0'
0/
#436000000000
1!
1'
1/
#436010000000
0!
0'
0/
#436020000000
#436030000000
1!
1'
1/
#436040000000
0!
0'
0/
#436050000000
1!
1'
1/
#436060000000
0!
1"
0'
1(
0/
10
#436070000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#436080000000
0!
0'
0/
#436090000000
1!
1'
1/
#436100000000
0!
0'
0/
#436110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#436120000000
0!
0'
0/
#436130000000
1!
1'
1/
#436140000000
0!
1"
0'
1(
0/
10
#436150000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#436160000000
0!
1$
0'
1+
0/
#436170000000
1!
1'
1/
#436180000000
0!
0'
0/
#436190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#436200000000
0!
0'
0/
#436210000000
1!
1'
1/
#436220000000
0!
0'
0/
#436230000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#436240000000
0!
0'
0/
#436250000000
1!
1'
1/
#436260000000
0!
0'
0/
#436270000000
1!
1'
1/
#436280000000
0!
0'
0/
#436290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#436300000000
0!
0'
0/
#436310000000
1!
1'
1/
#436320000000
0!
0'
0/
#436330000000
1!
1'
1/
#436340000000
0!
0'
0/
#436350000000
1!
1'
1/
#436360000000
0!
0'
0/
#436370000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#436380000000
0!
0'
0/
#436390000000
1!
1'
1/
#436400000000
0!
0'
0/
#436410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#436420000000
0!
0'
0/
#436430000000
1!
1'
1/
#436440000000
0!
0'
0/
#436450000000
#436460000000
1!
1'
1/
#436470000000
0!
0'
0/
#436480000000
1!
1'
1/
#436490000000
0!
1"
0'
1(
0/
10
#436500000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#436510000000
0!
0'
0/
#436520000000
1!
1'
1/
#436530000000
0!
0'
0/
#436540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#436550000000
0!
0'
0/
#436560000000
1!
1'
1/
#436570000000
0!
1"
0'
1(
0/
10
#436580000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#436590000000
0!
1$
0'
1+
0/
#436600000000
1!
1'
1/
#436610000000
0!
0'
0/
#436620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#436630000000
0!
0'
0/
#436640000000
1!
1'
1/
#436650000000
0!
0'
0/
#436660000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#436670000000
0!
0'
0/
#436680000000
1!
1'
1/
#436690000000
0!
0'
0/
#436700000000
1!
1'
1/
#436710000000
0!
0'
0/
#436720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#436730000000
0!
0'
0/
#436740000000
1!
1'
1/
#436750000000
0!
0'
0/
#436760000000
1!
1'
1/
#436770000000
0!
0'
0/
#436780000000
1!
1'
1/
#436790000000
0!
0'
0/
#436800000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#436810000000
0!
0'
0/
#436820000000
1!
1'
1/
#436830000000
0!
0'
0/
#436840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#436850000000
0!
0'
0/
#436860000000
1!
1'
1/
#436870000000
0!
0'
0/
#436880000000
#436890000000
1!
1'
1/
#436900000000
0!
0'
0/
#436910000000
1!
1'
1/
#436920000000
0!
1"
0'
1(
0/
10
#436930000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#436940000000
0!
0'
0/
#436950000000
1!
1'
1/
#436960000000
0!
0'
0/
#436970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#436980000000
0!
0'
0/
#436990000000
1!
1'
1/
#437000000000
0!
1"
0'
1(
0/
10
#437010000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#437020000000
0!
1$
0'
1+
0/
#437030000000
1!
1'
1/
#437040000000
0!
0'
0/
#437050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#437060000000
0!
0'
0/
#437070000000
1!
1'
1/
#437080000000
0!
0'
0/
#437090000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#437100000000
0!
0'
0/
#437110000000
1!
1'
1/
#437120000000
0!
0'
0/
#437130000000
1!
1'
1/
#437140000000
0!
0'
0/
#437150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#437160000000
0!
0'
0/
#437170000000
1!
1'
1/
#437180000000
0!
0'
0/
#437190000000
1!
1'
1/
#437200000000
0!
0'
0/
#437210000000
1!
1'
1/
#437220000000
0!
0'
0/
#437230000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#437240000000
0!
0'
0/
#437250000000
1!
1'
1/
#437260000000
0!
0'
0/
#437270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#437280000000
0!
0'
0/
#437290000000
1!
1'
1/
#437300000000
0!
0'
0/
#437310000000
#437320000000
1!
1'
1/
#437330000000
0!
0'
0/
#437340000000
1!
1'
1/
#437350000000
0!
1"
0'
1(
0/
10
#437360000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#437370000000
0!
0'
0/
#437380000000
1!
1'
1/
#437390000000
0!
0'
0/
#437400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#437410000000
0!
0'
0/
#437420000000
1!
1'
1/
#437430000000
0!
1"
0'
1(
0/
10
#437440000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#437450000000
0!
1$
0'
1+
0/
#437460000000
1!
1'
1/
#437470000000
0!
0'
0/
#437480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#437490000000
0!
0'
0/
#437500000000
1!
1'
1/
#437510000000
0!
0'
0/
#437520000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#437530000000
0!
0'
0/
#437540000000
1!
1'
1/
#437550000000
0!
0'
0/
#437560000000
1!
1'
1/
#437570000000
0!
0'
0/
#437580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#437590000000
0!
0'
0/
#437600000000
1!
1'
1/
#437610000000
0!
0'
0/
#437620000000
1!
1'
1/
#437630000000
0!
0'
0/
#437640000000
1!
1'
1/
#437650000000
0!
0'
0/
#437660000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#437670000000
0!
0'
0/
#437680000000
1!
1'
1/
#437690000000
0!
0'
0/
#437700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#437710000000
0!
0'
0/
#437720000000
1!
1'
1/
#437730000000
0!
0'
0/
#437740000000
#437750000000
1!
1'
1/
#437760000000
0!
0'
0/
#437770000000
1!
1'
1/
#437780000000
0!
1"
0'
1(
0/
10
#437790000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#437800000000
0!
0'
0/
#437810000000
1!
1'
1/
#437820000000
0!
0'
0/
#437830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#437840000000
0!
0'
0/
#437850000000
1!
1'
1/
#437860000000
0!
1"
0'
1(
0/
10
#437870000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#437880000000
0!
1$
0'
1+
0/
#437890000000
1!
1'
1/
#437900000000
0!
0'
0/
#437910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#437920000000
0!
0'
0/
#437930000000
1!
1'
1/
#437940000000
0!
0'
0/
#437950000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#437960000000
0!
0'
0/
#437970000000
1!
1'
1/
#437980000000
0!
0'
0/
#437990000000
1!
1'
1/
#438000000000
0!
0'
0/
#438010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#438020000000
0!
0'
0/
#438030000000
1!
1'
1/
#438040000000
0!
0'
0/
#438050000000
1!
1'
1/
#438060000000
0!
0'
0/
#438070000000
1!
1'
1/
#438080000000
0!
0'
0/
#438090000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#438100000000
0!
0'
0/
#438110000000
1!
1'
1/
#438120000000
0!
0'
0/
#438130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#438140000000
0!
0'
0/
#438150000000
1!
1'
1/
#438160000000
0!
0'
0/
#438170000000
#438180000000
1!
1'
1/
#438190000000
0!
0'
0/
#438200000000
1!
1'
1/
#438210000000
0!
1"
0'
1(
0/
10
#438220000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#438230000000
0!
0'
0/
#438240000000
1!
1'
1/
#438250000000
0!
0'
0/
#438260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#438270000000
0!
0'
0/
#438280000000
1!
1'
1/
#438290000000
0!
1"
0'
1(
0/
10
#438300000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#438310000000
0!
1$
0'
1+
0/
#438320000000
1!
1'
1/
#438330000000
0!
0'
0/
#438340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#438350000000
0!
0'
0/
#438360000000
1!
1'
1/
#438370000000
0!
0'
0/
#438380000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#438390000000
0!
0'
0/
#438400000000
1!
1'
1/
#438410000000
0!
0'
0/
#438420000000
1!
1'
1/
#438430000000
0!
0'
0/
#438440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#438450000000
0!
0'
0/
#438460000000
1!
1'
1/
#438470000000
0!
0'
0/
#438480000000
1!
1'
1/
#438490000000
0!
0'
0/
#438500000000
1!
1'
1/
#438510000000
0!
0'
0/
#438520000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#438530000000
0!
0'
0/
#438540000000
1!
1'
1/
#438550000000
0!
0'
0/
#438560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#438570000000
0!
0'
0/
#438580000000
1!
1'
1/
#438590000000
0!
0'
0/
#438600000000
#438610000000
1!
1'
1/
#438620000000
0!
0'
0/
#438630000000
1!
1'
1/
#438640000000
0!
1"
0'
1(
0/
10
#438650000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#438660000000
0!
0'
0/
#438670000000
1!
1'
1/
#438680000000
0!
0'
0/
#438690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#438700000000
0!
0'
0/
#438710000000
1!
1'
1/
#438720000000
0!
1"
0'
1(
0/
10
#438730000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#438740000000
0!
1$
0'
1+
0/
#438750000000
1!
1'
1/
#438760000000
0!
0'
0/
#438770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#438780000000
0!
0'
0/
#438790000000
1!
1'
1/
#438800000000
0!
0'
0/
#438810000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#438820000000
0!
0'
0/
#438830000000
1!
1'
1/
#438840000000
0!
0'
0/
#438850000000
1!
1'
1/
#438860000000
0!
0'
0/
#438870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#438880000000
0!
0'
0/
#438890000000
1!
1'
1/
#438900000000
0!
0'
0/
#438910000000
1!
1'
1/
#438920000000
0!
0'
0/
#438930000000
1!
1'
1/
#438940000000
0!
0'
0/
#438950000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#438960000000
0!
0'
0/
#438970000000
1!
1'
1/
#438980000000
0!
0'
0/
#438990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#439000000000
0!
0'
0/
#439010000000
1!
1'
1/
#439020000000
0!
0'
0/
#439030000000
#439040000000
1!
1'
1/
#439050000000
0!
0'
0/
#439060000000
1!
1'
1/
#439070000000
0!
1"
0'
1(
0/
10
#439080000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#439090000000
0!
0'
0/
#439100000000
1!
1'
1/
#439110000000
0!
0'
0/
#439120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#439130000000
0!
0'
0/
#439140000000
1!
1'
1/
#439150000000
0!
1"
0'
1(
0/
10
#439160000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#439170000000
0!
1$
0'
1+
0/
#439180000000
1!
1'
1/
#439190000000
0!
0'
0/
#439200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#439210000000
0!
0'
0/
#439220000000
1!
1'
1/
#439230000000
0!
0'
0/
#439240000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#439250000000
0!
0'
0/
#439260000000
1!
1'
1/
#439270000000
0!
0'
0/
#439280000000
1!
1'
1/
#439290000000
0!
0'
0/
#439300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#439310000000
0!
0'
0/
#439320000000
1!
1'
1/
#439330000000
0!
0'
0/
#439340000000
1!
1'
1/
#439350000000
0!
0'
0/
#439360000000
1!
1'
1/
#439370000000
0!
0'
0/
#439380000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#439390000000
0!
0'
0/
#439400000000
1!
1'
1/
#439410000000
0!
0'
0/
#439420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#439430000000
0!
0'
0/
#439440000000
1!
1'
1/
#439450000000
0!
0'
0/
#439460000000
#439470000000
1!
1'
1/
#439480000000
0!
0'
0/
#439490000000
1!
1'
1/
#439500000000
0!
1"
0'
1(
0/
10
#439510000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#439520000000
0!
0'
0/
#439530000000
1!
1'
1/
#439540000000
0!
0'
0/
#439550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#439560000000
0!
0'
0/
#439570000000
1!
1'
1/
#439580000000
0!
1"
0'
1(
0/
10
#439590000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#439600000000
0!
1$
0'
1+
0/
#439610000000
1!
1'
1/
#439620000000
0!
0'
0/
#439630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#439640000000
0!
0'
0/
#439650000000
1!
1'
1/
#439660000000
0!
0'
0/
#439670000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#439680000000
0!
0'
0/
#439690000000
1!
1'
1/
#439700000000
0!
0'
0/
#439710000000
1!
1'
1/
#439720000000
0!
0'
0/
#439730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#439740000000
0!
0'
0/
#439750000000
1!
1'
1/
#439760000000
0!
0'
0/
#439770000000
1!
1'
1/
#439780000000
0!
0'
0/
#439790000000
1!
1'
1/
#439800000000
0!
0'
0/
#439810000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#439820000000
0!
0'
0/
#439830000000
1!
1'
1/
#439840000000
0!
0'
0/
#439850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#439860000000
0!
0'
0/
#439870000000
1!
1'
1/
#439880000000
0!
0'
0/
#439890000000
#439900000000
1!
1'
1/
#439910000000
0!
0'
0/
#439920000000
1!
1'
1/
#439930000000
0!
1"
0'
1(
0/
10
#439940000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#439950000000
0!
0'
0/
#439960000000
1!
1'
1/
#439970000000
0!
0'
0/
#439980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#439990000000
0!
0'
0/
#440000000000
1!
1'
1/
#440010000000
0!
1"
0'
1(
0/
10
#440020000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#440030000000
0!
1$
0'
1+
0/
#440040000000
1!
1'
1/
#440050000000
0!
0'
0/
#440060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#440070000000
0!
0'
0/
#440080000000
1!
1'
1/
#440090000000
0!
0'
0/
#440100000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#440110000000
0!
0'
0/
#440120000000
1!
1'
1/
#440130000000
0!
0'
0/
#440140000000
1!
1'
1/
#440150000000
0!
0'
0/
#440160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#440170000000
0!
0'
0/
#440180000000
1!
1'
1/
#440190000000
0!
0'
0/
#440200000000
1!
1'
1/
#440210000000
0!
0'
0/
#440220000000
1!
1'
1/
#440230000000
0!
0'
0/
#440240000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#440250000000
0!
0'
0/
#440260000000
1!
1'
1/
#440270000000
0!
0'
0/
#440280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#440290000000
0!
0'
0/
#440300000000
1!
1'
1/
#440310000000
0!
0'
0/
#440320000000
#440330000000
1!
1'
1/
#440340000000
0!
0'
0/
#440350000000
1!
1'
1/
#440360000000
0!
1"
0'
1(
0/
10
#440370000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#440380000000
0!
0'
0/
#440390000000
1!
1'
1/
#440400000000
0!
0'
0/
#440410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#440420000000
0!
0'
0/
#440430000000
1!
1'
1/
#440440000000
0!
1"
0'
1(
0/
10
#440450000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#440460000000
0!
1$
0'
1+
0/
#440470000000
1!
1'
1/
#440480000000
0!
0'
0/
#440490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#440500000000
0!
0'
0/
#440510000000
1!
1'
1/
#440520000000
0!
0'
0/
#440530000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#440540000000
0!
0'
0/
#440550000000
1!
1'
1/
#440560000000
0!
0'
0/
#440570000000
1!
1'
1/
#440580000000
0!
0'
0/
#440590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#440600000000
0!
0'
0/
#440610000000
1!
1'
1/
#440620000000
0!
0'
0/
#440630000000
1!
1'
1/
#440640000000
0!
0'
0/
#440650000000
1!
1'
1/
#440660000000
0!
0'
0/
#440670000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#440680000000
0!
0'
0/
#440690000000
1!
1'
1/
#440700000000
0!
0'
0/
#440710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#440720000000
0!
0'
0/
#440730000000
1!
1'
1/
#440740000000
0!
0'
0/
#440750000000
#440760000000
1!
1'
1/
#440770000000
0!
0'
0/
#440780000000
1!
1'
1/
#440790000000
0!
1"
0'
1(
0/
10
#440800000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#440810000000
0!
0'
0/
#440820000000
1!
1'
1/
#440830000000
0!
0'
0/
#440840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#440850000000
0!
0'
0/
#440860000000
1!
1'
1/
#440870000000
0!
1"
0'
1(
0/
10
#440880000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#440890000000
0!
1$
0'
1+
0/
#440900000000
1!
1'
1/
#440910000000
0!
0'
0/
#440920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#440930000000
0!
0'
0/
#440940000000
1!
1'
1/
#440950000000
0!
0'
0/
#440960000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#440970000000
0!
0'
0/
#440980000000
1!
1'
1/
#440990000000
0!
0'
0/
#441000000000
1!
1'
1/
#441010000000
0!
0'
0/
#441020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#441030000000
0!
0'
0/
#441040000000
1!
1'
1/
#441050000000
0!
0'
0/
#441060000000
1!
1'
1/
#441070000000
0!
0'
0/
#441080000000
1!
1'
1/
#441090000000
0!
0'
0/
#441100000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#441110000000
0!
0'
0/
#441120000000
1!
1'
1/
#441130000000
0!
0'
0/
#441140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#441150000000
0!
0'
0/
#441160000000
1!
1'
1/
#441170000000
0!
0'
0/
#441180000000
#441190000000
1!
1'
1/
#441200000000
0!
0'
0/
#441210000000
1!
1'
1/
#441220000000
0!
1"
0'
1(
0/
10
#441230000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#441240000000
0!
0'
0/
#441250000000
1!
1'
1/
#441260000000
0!
0'
0/
#441270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#441280000000
0!
0'
0/
#441290000000
1!
1'
1/
#441300000000
0!
1"
0'
1(
0/
10
#441310000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#441320000000
0!
1$
0'
1+
0/
#441330000000
1!
1'
1/
#441340000000
0!
0'
0/
#441350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#441360000000
0!
0'
0/
#441370000000
1!
1'
1/
#441380000000
0!
0'
0/
#441390000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#441400000000
0!
0'
0/
#441410000000
1!
1'
1/
#441420000000
0!
0'
0/
#441430000000
1!
1'
1/
#441440000000
0!
0'
0/
#441450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#441460000000
0!
0'
0/
#441470000000
1!
1'
1/
#441480000000
0!
0'
0/
#441490000000
1!
1'
1/
#441500000000
0!
0'
0/
#441510000000
1!
1'
1/
#441520000000
0!
0'
0/
#441530000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#441540000000
0!
0'
0/
#441550000000
1!
1'
1/
#441560000000
0!
0'
0/
#441570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#441580000000
0!
0'
0/
#441590000000
1!
1'
1/
#441600000000
0!
0'
0/
#441610000000
#441620000000
1!
1'
1/
#441630000000
0!
0'
0/
#441640000000
1!
1'
1/
#441650000000
0!
1"
0'
1(
0/
10
#441660000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#441670000000
0!
0'
0/
#441680000000
1!
1'
1/
#441690000000
0!
0'
0/
#441700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#441710000000
0!
0'
0/
#441720000000
1!
1'
1/
#441730000000
0!
1"
0'
1(
0/
10
#441740000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#441750000000
0!
1$
0'
1+
0/
#441760000000
1!
1'
1/
#441770000000
0!
0'
0/
#441780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#441790000000
0!
0'
0/
#441800000000
1!
1'
1/
#441810000000
0!
0'
0/
#441820000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#441830000000
0!
0'
0/
#441840000000
1!
1'
1/
#441850000000
0!
0'
0/
#441860000000
1!
1'
1/
#441870000000
0!
0'
0/
#441880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#441890000000
0!
0'
0/
#441900000000
1!
1'
1/
#441910000000
0!
0'
0/
#441920000000
1!
1'
1/
#441930000000
0!
0'
0/
#441940000000
1!
1'
1/
#441950000000
0!
0'
0/
#441960000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#441970000000
0!
0'
0/
#441980000000
1!
1'
1/
#441990000000
0!
0'
0/
#442000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#442010000000
0!
0'
0/
#442020000000
1!
1'
1/
#442030000000
0!
0'
0/
#442040000000
#442050000000
1!
1'
1/
#442060000000
0!
0'
0/
#442070000000
1!
1'
1/
#442080000000
0!
1"
0'
1(
0/
10
#442090000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#442100000000
0!
0'
0/
#442110000000
1!
1'
1/
#442120000000
0!
0'
0/
#442130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#442140000000
0!
0'
0/
#442150000000
1!
1'
1/
#442160000000
0!
1"
0'
1(
0/
10
#442170000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#442180000000
0!
1$
0'
1+
0/
#442190000000
1!
1'
1/
#442200000000
0!
0'
0/
#442210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#442220000000
0!
0'
0/
#442230000000
1!
1'
1/
#442240000000
0!
0'
0/
#442250000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#442260000000
0!
0'
0/
#442270000000
1!
1'
1/
#442280000000
0!
0'
0/
#442290000000
1!
1'
1/
#442300000000
0!
0'
0/
#442310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#442320000000
0!
0'
0/
#442330000000
1!
1'
1/
#442340000000
0!
0'
0/
#442350000000
1!
1'
1/
#442360000000
0!
0'
0/
#442370000000
1!
1'
1/
#442380000000
0!
0'
0/
#442390000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#442400000000
0!
0'
0/
#442410000000
1!
1'
1/
#442420000000
0!
0'
0/
#442430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#442440000000
0!
0'
0/
#442450000000
1!
1'
1/
#442460000000
0!
0'
0/
#442470000000
#442480000000
1!
1'
1/
#442490000000
0!
0'
0/
#442500000000
1!
1'
1/
#442510000000
0!
1"
0'
1(
0/
10
#442520000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#442530000000
0!
0'
0/
#442540000000
1!
1'
1/
#442550000000
0!
0'
0/
#442560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#442570000000
0!
0'
0/
#442580000000
1!
1'
1/
#442590000000
0!
1"
0'
1(
0/
10
#442600000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#442610000000
0!
1$
0'
1+
0/
#442620000000
1!
1'
1/
#442630000000
0!
0'
0/
#442640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#442650000000
0!
0'
0/
#442660000000
1!
1'
1/
#442670000000
0!
0'
0/
#442680000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#442690000000
0!
0'
0/
#442700000000
1!
1'
1/
#442710000000
0!
0'
0/
#442720000000
1!
1'
1/
#442730000000
0!
0'
0/
#442740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#442750000000
0!
0'
0/
#442760000000
1!
1'
1/
#442770000000
0!
0'
0/
#442780000000
1!
1'
1/
#442790000000
0!
0'
0/
#442800000000
1!
1'
1/
#442810000000
0!
0'
0/
#442820000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#442830000000
0!
0'
0/
#442840000000
1!
1'
1/
#442850000000
0!
0'
0/
#442860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#442870000000
0!
0'
0/
#442880000000
1!
1'
1/
#442890000000
0!
0'
0/
#442900000000
#442910000000
1!
1'
1/
#442920000000
0!
0'
0/
#442930000000
1!
1'
1/
#442940000000
0!
1"
0'
1(
0/
10
#442950000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#442960000000
0!
0'
0/
#442970000000
1!
1'
1/
#442980000000
0!
0'
0/
#442990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#443000000000
0!
0'
0/
#443010000000
1!
1'
1/
#443020000000
0!
1"
0'
1(
0/
10
#443030000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#443040000000
0!
1$
0'
1+
0/
#443050000000
1!
1'
1/
#443060000000
0!
0'
0/
#443070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#443080000000
0!
0'
0/
#443090000000
1!
1'
1/
#443100000000
0!
0'
0/
#443110000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#443120000000
0!
0'
0/
#443130000000
1!
1'
1/
#443140000000
0!
0'
0/
#443150000000
1!
1'
1/
#443160000000
0!
0'
0/
#443170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#443180000000
0!
0'
0/
#443190000000
1!
1'
1/
#443200000000
0!
0'
0/
#443210000000
1!
1'
1/
#443220000000
0!
0'
0/
#443230000000
1!
1'
1/
#443240000000
0!
0'
0/
#443250000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#443260000000
0!
0'
0/
#443270000000
1!
1'
1/
#443280000000
0!
0'
0/
#443290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#443300000000
0!
0'
0/
#443310000000
1!
1'
1/
#443320000000
0!
0'
0/
#443330000000
#443340000000
1!
1'
1/
#443350000000
0!
0'
0/
#443360000000
1!
1'
1/
#443370000000
0!
1"
0'
1(
0/
10
#443380000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#443390000000
0!
0'
0/
#443400000000
1!
1'
1/
#443410000000
0!
0'
0/
#443420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#443430000000
0!
0'
0/
#443440000000
1!
1'
1/
#443450000000
0!
1"
0'
1(
0/
10
#443460000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#443470000000
0!
1$
0'
1+
0/
#443480000000
1!
1'
1/
#443490000000
0!
0'
0/
#443500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#443510000000
0!
0'
0/
#443520000000
1!
1'
1/
#443530000000
0!
0'
0/
#443540000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#443550000000
0!
0'
0/
#443560000000
1!
1'
1/
#443570000000
0!
0'
0/
#443580000000
1!
1'
1/
#443590000000
0!
0'
0/
#443600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#443610000000
0!
0'
0/
#443620000000
1!
1'
1/
#443630000000
0!
0'
0/
#443640000000
1!
1'
1/
#443650000000
0!
0'
0/
#443660000000
1!
1'
1/
#443670000000
0!
0'
0/
#443680000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#443690000000
0!
0'
0/
#443700000000
1!
1'
1/
#443710000000
0!
0'
0/
#443720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#443730000000
0!
0'
0/
#443740000000
1!
1'
1/
#443750000000
0!
0'
0/
#443760000000
#443770000000
1!
1'
1/
#443780000000
0!
0'
0/
#443790000000
1!
1'
1/
#443800000000
0!
1"
0'
1(
0/
10
#443810000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#443820000000
0!
0'
0/
#443830000000
1!
1'
1/
#443840000000
0!
0'
0/
#443850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#443860000000
0!
0'
0/
#443870000000
1!
1'
1/
#443880000000
0!
1"
0'
1(
0/
10
#443890000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#443900000000
0!
1$
0'
1+
0/
#443910000000
1!
1'
1/
#443920000000
0!
0'
0/
#443930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#443940000000
0!
0'
0/
#443950000000
1!
1'
1/
#443960000000
0!
0'
0/
#443970000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#443980000000
0!
0'
0/
#443990000000
1!
1'
1/
#444000000000
0!
0'
0/
#444010000000
1!
1'
1/
#444020000000
0!
0'
0/
#444030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#444040000000
0!
0'
0/
#444050000000
1!
1'
1/
#444060000000
0!
0'
0/
#444070000000
1!
1'
1/
#444080000000
0!
0'
0/
#444090000000
1!
1'
1/
#444100000000
0!
0'
0/
#444110000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#444120000000
0!
0'
0/
#444130000000
1!
1'
1/
#444140000000
0!
0'
0/
#444150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#444160000000
0!
0'
0/
#444170000000
1!
1'
1/
#444180000000
0!
0'
0/
#444190000000
#444200000000
1!
1'
1/
#444210000000
0!
0'
0/
#444220000000
1!
1'
1/
#444230000000
0!
1"
0'
1(
0/
10
#444240000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#444250000000
0!
0'
0/
#444260000000
1!
1'
1/
#444270000000
0!
0'
0/
#444280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#444290000000
0!
0'
0/
#444300000000
1!
1'
1/
#444310000000
0!
1"
0'
1(
0/
10
#444320000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#444330000000
0!
1$
0'
1+
0/
#444340000000
1!
1'
1/
#444350000000
0!
0'
0/
#444360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#444370000000
0!
0'
0/
#444380000000
1!
1'
1/
#444390000000
0!
0'
0/
#444400000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#444410000000
0!
0'
0/
#444420000000
1!
1'
1/
#444430000000
0!
0'
0/
#444440000000
1!
1'
1/
#444450000000
0!
0'
0/
#444460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#444470000000
0!
0'
0/
#444480000000
1!
1'
1/
#444490000000
0!
0'
0/
#444500000000
1!
1'
1/
#444510000000
0!
0'
0/
#444520000000
1!
1'
1/
#444530000000
0!
0'
0/
#444540000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#444550000000
0!
0'
0/
#444560000000
1!
1'
1/
#444570000000
0!
0'
0/
#444580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#444590000000
0!
0'
0/
#444600000000
1!
1'
1/
#444610000000
0!
0'
0/
#444620000000
#444630000000
1!
1'
1/
#444640000000
0!
0'
0/
#444650000000
1!
1'
1/
#444660000000
0!
1"
0'
1(
0/
10
#444670000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#444680000000
0!
0'
0/
#444690000000
1!
1'
1/
#444700000000
0!
0'
0/
#444710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#444720000000
0!
0'
0/
#444730000000
1!
1'
1/
#444740000000
0!
1"
0'
1(
0/
10
#444750000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#444760000000
0!
1$
0'
1+
0/
#444770000000
1!
1'
1/
#444780000000
0!
0'
0/
#444790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#444800000000
0!
0'
0/
#444810000000
1!
1'
1/
#444820000000
0!
0'
0/
#444830000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#444840000000
0!
0'
0/
#444850000000
1!
1'
1/
#444860000000
0!
0'
0/
#444870000000
1!
1'
1/
#444880000000
0!
0'
0/
#444890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#444900000000
0!
0'
0/
#444910000000
1!
1'
1/
#444920000000
0!
0'
0/
#444930000000
1!
1'
1/
#444940000000
0!
0'
0/
#444950000000
1!
1'
1/
#444960000000
0!
0'
0/
#444970000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#444980000000
0!
0'
0/
#444990000000
1!
1'
1/
#445000000000
0!
0'
0/
#445010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#445020000000
0!
0'
0/
#445030000000
1!
1'
1/
#445040000000
0!
0'
0/
#445050000000
#445060000000
1!
1'
1/
#445070000000
0!
0'
0/
#445080000000
1!
1'
1/
#445090000000
0!
1"
0'
1(
0/
10
#445100000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#445110000000
0!
0'
0/
#445120000000
1!
1'
1/
#445130000000
0!
0'
0/
#445140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#445150000000
0!
0'
0/
#445160000000
1!
1'
1/
#445170000000
0!
1"
0'
1(
0/
10
#445180000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#445190000000
0!
1$
0'
1+
0/
#445200000000
1!
1'
1/
#445210000000
0!
0'
0/
#445220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#445230000000
0!
0'
0/
#445240000000
1!
1'
1/
#445250000000
0!
0'
0/
#445260000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#445270000000
0!
0'
0/
#445280000000
1!
1'
1/
#445290000000
0!
0'
0/
#445300000000
1!
1'
1/
#445310000000
0!
0'
0/
#445320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#445330000000
0!
0'
0/
#445340000000
1!
1'
1/
#445350000000
0!
0'
0/
#445360000000
1!
1'
1/
#445370000000
0!
0'
0/
#445380000000
1!
1'
1/
#445390000000
0!
0'
0/
#445400000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#445410000000
0!
0'
0/
#445420000000
1!
1'
1/
#445430000000
0!
0'
0/
#445440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#445450000000
0!
0'
0/
#445460000000
1!
1'
1/
#445470000000
0!
0'
0/
#445480000000
#445490000000
1!
1'
1/
#445500000000
0!
0'
0/
#445510000000
1!
1'
1/
#445520000000
0!
1"
0'
1(
0/
10
#445530000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#445540000000
0!
0'
0/
#445550000000
1!
1'
1/
#445560000000
0!
0'
0/
#445570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#445580000000
0!
0'
0/
#445590000000
1!
1'
1/
#445600000000
0!
1"
0'
1(
0/
10
#445610000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#445620000000
0!
1$
0'
1+
0/
#445630000000
1!
1'
1/
#445640000000
0!
0'
0/
#445650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#445660000000
0!
0'
0/
#445670000000
1!
1'
1/
#445680000000
0!
0'
0/
#445690000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#445700000000
0!
0'
0/
#445710000000
1!
1'
1/
#445720000000
0!
0'
0/
#445730000000
1!
1'
1/
#445740000000
0!
0'
0/
#445750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#445760000000
0!
0'
0/
#445770000000
1!
1'
1/
#445780000000
0!
0'
0/
#445790000000
1!
1'
1/
#445800000000
0!
0'
0/
#445810000000
1!
1'
1/
#445820000000
0!
0'
0/
#445830000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#445840000000
0!
0'
0/
#445850000000
1!
1'
1/
#445860000000
0!
0'
0/
#445870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#445880000000
0!
0'
0/
#445890000000
1!
1'
1/
#445900000000
0!
0'
0/
#445910000000
#445920000000
1!
1'
1/
#445930000000
0!
0'
0/
#445940000000
1!
1'
1/
#445950000000
0!
1"
0'
1(
0/
10
#445960000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#445970000000
0!
0'
0/
#445980000000
1!
1'
1/
#445990000000
0!
0'
0/
#446000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#446010000000
0!
0'
0/
#446020000000
1!
1'
1/
#446030000000
0!
1"
0'
1(
0/
10
#446040000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#446050000000
0!
1$
0'
1+
0/
#446060000000
1!
1'
1/
#446070000000
0!
0'
0/
#446080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#446090000000
0!
0'
0/
#446100000000
1!
1'
1/
#446110000000
0!
0'
0/
#446120000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#446130000000
0!
0'
0/
#446140000000
1!
1'
1/
#446150000000
0!
0'
0/
#446160000000
1!
1'
1/
#446170000000
0!
0'
0/
#446180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#446190000000
0!
0'
0/
#446200000000
1!
1'
1/
#446210000000
0!
0'
0/
#446220000000
1!
1'
1/
#446230000000
0!
0'
0/
#446240000000
1!
1'
1/
#446250000000
0!
0'
0/
#446260000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#446270000000
0!
0'
0/
#446280000000
1!
1'
1/
#446290000000
0!
0'
0/
#446300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#446310000000
0!
0'
0/
#446320000000
1!
1'
1/
#446330000000
0!
0'
0/
#446340000000
#446350000000
1!
1'
1/
#446360000000
0!
0'
0/
#446370000000
1!
1'
1/
#446380000000
0!
1"
0'
1(
0/
10
#446390000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#446400000000
0!
0'
0/
#446410000000
1!
1'
1/
#446420000000
0!
0'
0/
#446430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#446440000000
0!
0'
0/
#446450000000
1!
1'
1/
#446460000000
0!
1"
0'
1(
0/
10
#446470000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#446480000000
0!
1$
0'
1+
0/
#446490000000
1!
1'
1/
#446500000000
0!
0'
0/
#446510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#446520000000
0!
0'
0/
#446530000000
1!
1'
1/
#446540000000
0!
0'
0/
#446550000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#446560000000
0!
0'
0/
#446570000000
1!
1'
1/
#446580000000
0!
0'
0/
#446590000000
1!
1'
1/
#446600000000
0!
0'
0/
#446610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#446620000000
0!
0'
0/
#446630000000
1!
1'
1/
#446640000000
0!
0'
0/
#446650000000
1!
1'
1/
#446660000000
0!
0'
0/
#446670000000
1!
1'
1/
#446680000000
0!
0'
0/
#446690000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#446700000000
0!
0'
0/
#446710000000
1!
1'
1/
#446720000000
0!
0'
0/
#446730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#446740000000
0!
0'
0/
#446750000000
1!
1'
1/
#446760000000
0!
0'
0/
#446770000000
#446780000000
1!
1'
1/
#446790000000
0!
0'
0/
#446800000000
1!
1'
1/
#446810000000
0!
1"
0'
1(
0/
10
#446820000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#446830000000
0!
0'
0/
#446840000000
1!
1'
1/
#446850000000
0!
0'
0/
#446860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#446870000000
0!
0'
0/
#446880000000
1!
1'
1/
#446890000000
0!
1"
0'
1(
0/
10
#446900000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#446910000000
0!
1$
0'
1+
0/
#446920000000
1!
1'
1/
#446930000000
0!
0'
0/
#446940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#446950000000
0!
0'
0/
#446960000000
1!
1'
1/
#446970000000
0!
0'
0/
#446980000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#446990000000
0!
0'
0/
#447000000000
1!
1'
1/
#447010000000
0!
0'
0/
#447020000000
1!
1'
1/
#447030000000
0!
0'
0/
#447040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#447050000000
0!
0'
0/
#447060000000
1!
1'
1/
#447070000000
0!
0'
0/
#447080000000
1!
1'
1/
#447090000000
0!
0'
0/
#447100000000
1!
1'
1/
#447110000000
0!
0'
0/
#447120000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#447130000000
0!
0'
0/
#447140000000
1!
1'
1/
#447150000000
0!
0'
0/
#447160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#447170000000
0!
0'
0/
#447180000000
1!
1'
1/
#447190000000
0!
0'
0/
#447200000000
#447210000000
1!
1'
1/
#447220000000
0!
0'
0/
#447230000000
1!
1'
1/
#447240000000
0!
1"
0'
1(
0/
10
#447250000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#447260000000
0!
0'
0/
#447270000000
1!
1'
1/
#447280000000
0!
0'
0/
#447290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#447300000000
0!
0'
0/
#447310000000
1!
1'
1/
#447320000000
0!
1"
0'
1(
0/
10
#447330000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#447340000000
0!
1$
0'
1+
0/
#447350000000
1!
1'
1/
#447360000000
0!
0'
0/
#447370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#447380000000
0!
0'
0/
#447390000000
1!
1'
1/
#447400000000
0!
0'
0/
#447410000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#447420000000
0!
0'
0/
#447430000000
1!
1'
1/
#447440000000
0!
0'
0/
#447450000000
1!
1'
1/
#447460000000
0!
0'
0/
#447470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#447480000000
0!
0'
0/
#447490000000
1!
1'
1/
#447500000000
0!
0'
0/
#447510000000
1!
1'
1/
#447520000000
0!
0'
0/
#447530000000
1!
1'
1/
#447540000000
0!
0'
0/
#447550000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#447560000000
0!
0'
0/
#447570000000
1!
1'
1/
#447580000000
0!
0'
0/
#447590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#447600000000
0!
0'
0/
#447610000000
1!
1'
1/
#447620000000
0!
0'
0/
#447630000000
#447640000000
1!
1'
1/
#447650000000
0!
0'
0/
#447660000000
1!
1'
1/
#447670000000
0!
1"
0'
1(
0/
10
#447680000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#447690000000
0!
0'
0/
#447700000000
1!
1'
1/
#447710000000
0!
0'
0/
#447720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#447730000000
0!
0'
0/
#447740000000
1!
1'
1/
#447750000000
0!
1"
0'
1(
0/
10
#447760000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#447770000000
0!
1$
0'
1+
0/
#447780000000
1!
1'
1/
#447790000000
0!
0'
0/
#447800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#447810000000
0!
0'
0/
#447820000000
1!
1'
1/
#447830000000
0!
0'
0/
#447840000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#447850000000
0!
0'
0/
#447860000000
1!
1'
1/
#447870000000
0!
0'
0/
#447880000000
1!
1'
1/
#447890000000
0!
0'
0/
#447900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#447910000000
0!
0'
0/
#447920000000
1!
1'
1/
#447930000000
0!
0'
0/
#447940000000
1!
1'
1/
#447950000000
0!
0'
0/
#447960000000
1!
1'
1/
#447970000000
0!
0'
0/
#447980000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#447990000000
0!
0'
0/
#448000000000
1!
1'
1/
#448010000000
0!
0'
0/
#448020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#448030000000
0!
0'
0/
#448040000000
1!
1'
1/
#448050000000
0!
0'
0/
#448060000000
#448070000000
1!
1'
1/
#448080000000
0!
0'
0/
#448090000000
1!
1'
1/
#448100000000
0!
1"
0'
1(
0/
10
#448110000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#448120000000
0!
0'
0/
#448130000000
1!
1'
1/
#448140000000
0!
0'
0/
#448150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#448160000000
0!
0'
0/
#448170000000
1!
1'
1/
#448180000000
0!
1"
0'
1(
0/
10
#448190000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#448200000000
0!
1$
0'
1+
0/
#448210000000
1!
1'
1/
#448220000000
0!
0'
0/
#448230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#448240000000
0!
0'
0/
#448250000000
1!
1'
1/
#448260000000
0!
0'
0/
#448270000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#448280000000
0!
0'
0/
#448290000000
1!
1'
1/
#448300000000
0!
0'
0/
#448310000000
1!
1'
1/
#448320000000
0!
0'
0/
#448330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#448340000000
0!
0'
0/
#448350000000
1!
1'
1/
#448360000000
0!
0'
0/
#448370000000
1!
1'
1/
#448380000000
0!
0'
0/
#448390000000
1!
1'
1/
#448400000000
0!
0'
0/
#448410000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#448420000000
0!
0'
0/
#448430000000
1!
1'
1/
#448440000000
0!
0'
0/
#448450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#448460000000
0!
0'
0/
#448470000000
1!
1'
1/
#448480000000
0!
0'
0/
#448490000000
#448500000000
1!
1'
1/
#448510000000
0!
0'
0/
#448520000000
1!
1'
1/
#448530000000
0!
1"
0'
1(
0/
10
#448540000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#448550000000
0!
0'
0/
#448560000000
1!
1'
1/
#448570000000
0!
0'
0/
#448580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#448590000000
0!
0'
0/
#448600000000
1!
1'
1/
#448610000000
0!
1"
0'
1(
0/
10
#448620000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#448630000000
0!
1$
0'
1+
0/
#448640000000
1!
1'
1/
#448650000000
0!
0'
0/
#448660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#448670000000
0!
0'
0/
#448680000000
1!
1'
1/
#448690000000
0!
0'
0/
#448700000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#448710000000
0!
0'
0/
#448720000000
1!
1'
1/
#448730000000
0!
0'
0/
#448740000000
1!
1'
1/
#448750000000
0!
0'
0/
#448760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#448770000000
0!
0'
0/
#448780000000
1!
1'
1/
#448790000000
0!
0'
0/
#448800000000
1!
1'
1/
#448810000000
0!
0'
0/
#448820000000
1!
1'
1/
#448830000000
0!
0'
0/
#448840000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#448850000000
0!
0'
0/
#448860000000
1!
1'
1/
#448870000000
0!
0'
0/
#448880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#448890000000
0!
0'
0/
#448900000000
1!
1'
1/
#448910000000
0!
0'
0/
#448920000000
#448930000000
1!
1'
1/
#448940000000
0!
0'
0/
#448950000000
1!
1'
1/
#448960000000
0!
1"
0'
1(
0/
10
#448970000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#448980000000
0!
0'
0/
#448990000000
1!
1'
1/
#449000000000
0!
0'
0/
#449010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#449020000000
0!
0'
0/
#449030000000
1!
1'
1/
#449040000000
0!
1"
0'
1(
0/
10
#449050000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#449060000000
0!
1$
0'
1+
0/
#449070000000
1!
1'
1/
#449080000000
0!
0'
0/
#449090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#449100000000
0!
0'
0/
#449110000000
1!
1'
1/
#449120000000
0!
0'
0/
#449130000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#449140000000
0!
0'
0/
#449150000000
1!
1'
1/
#449160000000
0!
0'
0/
#449170000000
1!
1'
1/
#449180000000
0!
0'
0/
#449190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#449200000000
0!
0'
0/
#449210000000
1!
1'
1/
#449220000000
0!
0'
0/
#449230000000
1!
1'
1/
#449240000000
0!
0'
0/
#449250000000
1!
1'
1/
#449260000000
0!
0'
0/
#449270000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#449280000000
0!
0'
0/
#449290000000
1!
1'
1/
#449300000000
0!
0'
0/
#449310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#449320000000
0!
0'
0/
#449330000000
1!
1'
1/
#449340000000
0!
0'
0/
#449350000000
#449360000000
1!
1'
1/
#449370000000
0!
0'
0/
#449380000000
1!
1'
1/
#449390000000
0!
1"
0'
1(
0/
10
#449400000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#449410000000
0!
0'
0/
#449420000000
1!
1'
1/
#449430000000
0!
0'
0/
#449440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#449450000000
0!
0'
0/
#449460000000
1!
1'
1/
#449470000000
0!
1"
0'
1(
0/
10
#449480000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#449490000000
0!
1$
0'
1+
0/
#449500000000
1!
1'
1/
#449510000000
0!
0'
0/
#449520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#449530000000
0!
0'
0/
#449540000000
1!
1'
1/
#449550000000
0!
0'
0/
#449560000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#449570000000
0!
0'
0/
#449580000000
1!
1'
1/
#449590000000
0!
0'
0/
#449600000000
1!
1'
1/
#449610000000
0!
0'
0/
#449620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#449630000000
0!
0'
0/
#449640000000
1!
1'
1/
#449650000000
0!
0'
0/
#449660000000
1!
1'
1/
#449670000000
0!
0'
0/
#449680000000
1!
1'
1/
#449690000000
0!
0'
0/
#449700000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#449710000000
0!
0'
0/
#449720000000
1!
1'
1/
#449730000000
0!
0'
0/
#449740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#449750000000
0!
0'
0/
#449760000000
1!
1'
1/
#449770000000
0!
0'
0/
#449780000000
#449790000000
1!
1'
1/
#449800000000
0!
0'
0/
#449810000000
1!
1'
1/
#449820000000
0!
1"
0'
1(
0/
10
#449830000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#449840000000
0!
0'
0/
#449850000000
1!
1'
1/
#449860000000
0!
0'
0/
#449870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#449880000000
0!
0'
0/
#449890000000
1!
1'
1/
#449900000000
0!
1"
0'
1(
0/
10
#449910000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#449920000000
0!
1$
0'
1+
0/
#449930000000
1!
1'
1/
#449940000000
0!
0'
0/
#449950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#449960000000
0!
0'
0/
#449970000000
1!
1'
1/
#449980000000
0!
0'
0/
#449990000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#450000000000
0!
0'
0/
#450010000000
1!
1'
1/
#450020000000
0!
0'
0/
#450030000000
1!
1'
1/
#450040000000
0!
0'
0/
#450050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#450060000000
0!
0'
0/
#450070000000
1!
1'
1/
#450080000000
0!
0'
0/
#450090000000
1!
1'
1/
#450100000000
0!
0'
0/
#450110000000
1!
1'
1/
#450120000000
0!
0'
0/
#450130000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#450140000000
0!
0'
0/
#450150000000
1!
1'
1/
#450160000000
0!
0'
0/
#450170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#450180000000
0!
0'
0/
#450190000000
1!
1'
1/
#450200000000
0!
0'
0/
#450210000000
#450220000000
1!
1'
1/
#450230000000
0!
0'
0/
#450240000000
1!
1'
1/
#450250000000
0!
1"
0'
1(
0/
10
#450260000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#450270000000
0!
0'
0/
#450280000000
1!
1'
1/
#450290000000
0!
0'
0/
#450300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#450310000000
0!
0'
0/
#450320000000
1!
1'
1/
#450330000000
0!
1"
0'
1(
0/
10
#450340000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#450350000000
0!
1$
0'
1+
0/
#450360000000
1!
1'
1/
#450370000000
0!
0'
0/
#450380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#450390000000
0!
0'
0/
#450400000000
1!
1'
1/
#450410000000
0!
0'
0/
#450420000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#450430000000
0!
0'
0/
#450440000000
1!
1'
1/
#450450000000
0!
0'
0/
#450460000000
1!
1'
1/
#450470000000
0!
0'
0/
#450480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#450490000000
0!
0'
0/
#450500000000
1!
1'
1/
#450510000000
0!
0'
0/
#450520000000
1!
1'
1/
#450530000000
0!
0'
0/
#450540000000
1!
1'
1/
#450550000000
0!
0'
0/
#450560000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#450570000000
0!
0'
0/
#450580000000
1!
1'
1/
#450590000000
0!
0'
0/
#450600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#450610000000
0!
0'
0/
#450620000000
1!
1'
1/
#450630000000
0!
0'
0/
#450640000000
#450650000000
1!
1'
1/
#450660000000
0!
0'
0/
#450670000000
1!
1'
1/
#450680000000
0!
1"
0'
1(
0/
10
#450690000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#450700000000
0!
0'
0/
#450710000000
1!
1'
1/
#450720000000
0!
0'
0/
#450730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#450740000000
0!
0'
0/
#450750000000
1!
1'
1/
#450760000000
0!
1"
0'
1(
0/
10
#450770000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#450780000000
0!
1$
0'
1+
0/
#450790000000
1!
1'
1/
#450800000000
0!
0'
0/
#450810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#450820000000
0!
0'
0/
#450830000000
1!
1'
1/
#450840000000
0!
0'
0/
#450850000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#450860000000
0!
0'
0/
#450870000000
1!
1'
1/
#450880000000
0!
0'
0/
#450890000000
1!
1'
1/
#450900000000
0!
0'
0/
#450910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#450920000000
0!
0'
0/
#450930000000
1!
1'
1/
#450940000000
0!
0'
0/
#450950000000
1!
1'
1/
#450960000000
0!
0'
0/
#450970000000
1!
1'
1/
#450980000000
0!
0'
0/
#450990000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#451000000000
0!
0'
0/
#451010000000
1!
1'
1/
#451020000000
0!
0'
0/
#451030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#451040000000
0!
0'
0/
#451050000000
1!
1'
1/
#451060000000
0!
0'
0/
#451070000000
#451080000000
1!
1'
1/
#451090000000
0!
0'
0/
#451100000000
1!
1'
1/
#451110000000
0!
1"
0'
1(
0/
10
#451120000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#451130000000
0!
0'
0/
#451140000000
1!
1'
1/
#451150000000
0!
0'
0/
#451160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#451170000000
0!
0'
0/
#451180000000
1!
1'
1/
#451190000000
0!
1"
0'
1(
0/
10
#451200000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#451210000000
0!
1$
0'
1+
0/
#451220000000
1!
1'
1/
#451230000000
0!
0'
0/
#451240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#451250000000
0!
0'
0/
#451260000000
1!
1'
1/
#451270000000
0!
0'
0/
#451280000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#451290000000
0!
0'
0/
#451300000000
1!
1'
1/
#451310000000
0!
0'
0/
#451320000000
1!
1'
1/
#451330000000
0!
0'
0/
#451340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#451350000000
0!
0'
0/
#451360000000
1!
1'
1/
#451370000000
0!
0'
0/
#451380000000
1!
1'
1/
#451390000000
0!
0'
0/
#451400000000
1!
1'
1/
#451410000000
0!
0'
0/
#451420000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#451430000000
0!
0'
0/
#451440000000
1!
1'
1/
#451450000000
0!
0'
0/
#451460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#451470000000
0!
0'
0/
#451480000000
1!
1'
1/
#451490000000
0!
0'
0/
#451500000000
#451510000000
1!
1'
1/
#451520000000
0!
0'
0/
#451530000000
1!
1'
1/
#451540000000
0!
1"
0'
1(
0/
10
#451550000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#451560000000
0!
0'
0/
#451570000000
1!
1'
1/
#451580000000
0!
0'
0/
#451590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#451600000000
0!
0'
0/
#451610000000
1!
1'
1/
#451620000000
0!
1"
0'
1(
0/
10
#451630000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#451640000000
0!
1$
0'
1+
0/
#451650000000
1!
1'
1/
#451660000000
0!
0'
0/
#451670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#451680000000
0!
0'
0/
#451690000000
1!
1'
1/
#451700000000
0!
0'
0/
#451710000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#451720000000
0!
0'
0/
#451730000000
1!
1'
1/
#451740000000
0!
0'
0/
#451750000000
1!
1'
1/
#451760000000
0!
0'
0/
#451770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#451780000000
0!
0'
0/
#451790000000
1!
1'
1/
#451800000000
0!
0'
0/
#451810000000
1!
1'
1/
#451820000000
0!
0'
0/
#451830000000
1!
1'
1/
#451840000000
0!
0'
0/
#451850000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#451860000000
0!
0'
0/
#451870000000
1!
1'
1/
#451880000000
0!
0'
0/
#451890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#451900000000
0!
0'
0/
#451910000000
1!
1'
1/
#451920000000
0!
0'
0/
#451930000000
#451940000000
1!
1'
1/
#451950000000
0!
0'
0/
#451960000000
1!
1'
1/
#451970000000
0!
1"
0'
1(
0/
10
#451980000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#451990000000
0!
0'
0/
#452000000000
1!
1'
1/
#452010000000
0!
0'
0/
#452020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#452030000000
0!
0'
0/
#452040000000
1!
1'
1/
#452050000000
0!
1"
0'
1(
0/
10
#452060000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#452070000000
0!
1$
0'
1+
0/
#452080000000
1!
1'
1/
#452090000000
0!
0'
0/
#452100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#452110000000
0!
0'
0/
#452120000000
1!
1'
1/
#452130000000
0!
0'
0/
#452140000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#452150000000
0!
0'
0/
#452160000000
1!
1'
1/
#452170000000
0!
0'
0/
#452180000000
1!
1'
1/
#452190000000
0!
0'
0/
#452200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#452210000000
0!
0'
0/
#452220000000
1!
1'
1/
#452230000000
0!
0'
0/
#452240000000
1!
1'
1/
#452250000000
0!
0'
0/
#452260000000
1!
1'
1/
#452270000000
0!
0'
0/
#452280000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#452290000000
0!
0'
0/
#452300000000
1!
1'
1/
#452310000000
0!
0'
0/
#452320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#452330000000
0!
0'
0/
#452340000000
1!
1'
1/
#452350000000
0!
0'
0/
#452360000000
#452370000000
1!
1'
1/
#452380000000
0!
0'
0/
#452390000000
1!
1'
1/
#452400000000
0!
1"
0'
1(
0/
10
#452410000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#452420000000
0!
0'
0/
#452430000000
1!
1'
1/
#452440000000
0!
0'
0/
#452450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#452460000000
0!
0'
0/
#452470000000
1!
1'
1/
#452480000000
0!
1"
0'
1(
0/
10
#452490000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#452500000000
0!
1$
0'
1+
0/
#452510000000
1!
1'
1/
#452520000000
0!
0'
0/
#452530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#452540000000
0!
0'
0/
#452550000000
1!
1'
1/
#452560000000
0!
0'
0/
#452570000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#452580000000
0!
0'
0/
#452590000000
1!
1'
1/
#452600000000
0!
0'
0/
#452610000000
1!
1'
1/
#452620000000
0!
0'
0/
#452630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#452640000000
0!
0'
0/
#452650000000
1!
1'
1/
#452660000000
0!
0'
0/
#452670000000
1!
1'
1/
#452680000000
0!
0'
0/
#452690000000
1!
1'
1/
#452700000000
0!
0'
0/
#452710000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#452720000000
0!
0'
0/
#452730000000
1!
1'
1/
#452740000000
0!
0'
0/
#452750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#452760000000
0!
0'
0/
#452770000000
1!
1'
1/
#452780000000
0!
0'
0/
#452790000000
#452800000000
1!
1'
1/
#452810000000
0!
0'
0/
#452820000000
1!
1'
1/
#452830000000
0!
1"
0'
1(
0/
10
#452840000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#452850000000
0!
0'
0/
#452860000000
1!
1'
1/
#452870000000
0!
0'
0/
#452880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#452890000000
0!
0'
0/
#452900000000
1!
1'
1/
#452910000000
0!
1"
0'
1(
0/
10
#452920000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#452930000000
0!
1$
0'
1+
0/
#452940000000
1!
1'
1/
#452950000000
0!
0'
0/
#452960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#452970000000
0!
0'
0/
#452980000000
1!
1'
1/
#452990000000
0!
0'
0/
#453000000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#453010000000
0!
0'
0/
#453020000000
1!
1'
1/
#453030000000
0!
0'
0/
#453040000000
1!
1'
1/
#453050000000
0!
0'
0/
#453060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#453070000000
0!
0'
0/
#453080000000
1!
1'
1/
#453090000000
0!
0'
0/
#453100000000
1!
1'
1/
#453110000000
0!
0'
0/
#453120000000
1!
1'
1/
#453130000000
0!
0'
0/
#453140000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#453150000000
0!
0'
0/
#453160000000
1!
1'
1/
#453170000000
0!
0'
0/
#453180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#453190000000
0!
0'
0/
#453200000000
1!
1'
1/
#453210000000
0!
0'
0/
#453220000000
#453230000000
1!
1'
1/
#453240000000
0!
0'
0/
#453250000000
1!
1'
1/
#453260000000
0!
1"
0'
1(
0/
10
#453270000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#453280000000
0!
0'
0/
#453290000000
1!
1'
1/
#453300000000
0!
0'
0/
#453310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#453320000000
0!
0'
0/
#453330000000
1!
1'
1/
#453340000000
0!
1"
0'
1(
0/
10
#453350000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#453360000000
0!
1$
0'
1+
0/
#453370000000
1!
1'
1/
#453380000000
0!
0'
0/
#453390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#453400000000
0!
0'
0/
#453410000000
1!
1'
1/
#453420000000
0!
0'
0/
#453430000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#453440000000
0!
0'
0/
#453450000000
1!
1'
1/
#453460000000
0!
0'
0/
#453470000000
1!
1'
1/
#453480000000
0!
0'
0/
#453490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#453500000000
0!
0'
0/
#453510000000
1!
1'
1/
#453520000000
0!
0'
0/
#453530000000
1!
1'
1/
#453540000000
0!
0'
0/
#453550000000
1!
1'
1/
#453560000000
0!
0'
0/
#453570000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#453580000000
0!
0'
0/
#453590000000
1!
1'
1/
#453600000000
0!
0'
0/
#453610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#453620000000
0!
0'
0/
#453630000000
1!
1'
1/
#453640000000
0!
0'
0/
#453650000000
#453660000000
1!
1'
1/
#453670000000
0!
0'
0/
#453680000000
1!
1'
1/
#453690000000
0!
1"
0'
1(
0/
10
#453700000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#453710000000
0!
0'
0/
#453720000000
1!
1'
1/
#453730000000
0!
0'
0/
#453740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#453750000000
0!
0'
0/
#453760000000
1!
1'
1/
#453770000000
0!
1"
0'
1(
0/
10
#453780000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#453790000000
0!
1$
0'
1+
0/
#453800000000
1!
1'
1/
#453810000000
0!
0'
0/
#453820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#453830000000
0!
0'
0/
#453840000000
1!
1'
1/
#453850000000
0!
0'
0/
#453860000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#453870000000
0!
0'
0/
#453880000000
1!
1'
1/
#453890000000
0!
0'
0/
#453900000000
1!
1'
1/
#453910000000
0!
0'
0/
#453920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#453930000000
0!
0'
0/
#453940000000
1!
1'
1/
#453950000000
0!
0'
0/
#453960000000
1!
1'
1/
#453970000000
0!
0'
0/
#453980000000
1!
1'
1/
#453990000000
0!
0'
0/
#454000000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#454010000000
0!
0'
0/
#454020000000
1!
1'
1/
#454030000000
0!
0'
0/
#454040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#454050000000
0!
0'
0/
#454060000000
1!
1'
1/
#454070000000
0!
0'
0/
#454080000000
#454090000000
1!
1'
1/
#454100000000
0!
0'
0/
#454110000000
1!
1'
1/
#454120000000
0!
1"
0'
1(
0/
10
#454130000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#454140000000
0!
0'
0/
#454150000000
1!
1'
1/
#454160000000
0!
0'
0/
#454170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#454180000000
0!
0'
0/
#454190000000
1!
1'
1/
#454200000000
0!
1"
0'
1(
0/
10
#454210000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#454220000000
0!
1$
0'
1+
0/
#454230000000
1!
1'
1/
#454240000000
0!
0'
0/
#454250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#454260000000
0!
0'
0/
#454270000000
1!
1'
1/
#454280000000
0!
0'
0/
#454290000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#454300000000
0!
0'
0/
#454310000000
1!
1'
1/
#454320000000
0!
0'
0/
#454330000000
1!
1'
1/
#454340000000
0!
0'
0/
#454350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#454360000000
0!
0'
0/
#454370000000
1!
1'
1/
#454380000000
0!
0'
0/
#454390000000
1!
1'
1/
#454400000000
0!
0'
0/
#454410000000
1!
1'
1/
#454420000000
0!
0'
0/
#454430000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#454440000000
0!
0'
0/
#454450000000
1!
1'
1/
#454460000000
0!
0'
0/
#454470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#454480000000
0!
0'
0/
#454490000000
1!
1'
1/
#454500000000
0!
0'
0/
#454510000000
#454520000000
1!
1'
1/
#454530000000
0!
0'
0/
#454540000000
1!
1'
1/
#454550000000
0!
1"
0'
1(
0/
10
#454560000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#454570000000
0!
0'
0/
#454580000000
1!
1'
1/
#454590000000
0!
0'
0/
#454600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#454610000000
0!
0'
0/
#454620000000
1!
1'
1/
#454630000000
0!
1"
0'
1(
0/
10
#454640000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#454650000000
0!
1$
0'
1+
0/
#454660000000
1!
1'
1/
#454670000000
0!
0'
0/
#454680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#454690000000
0!
0'
0/
#454700000000
1!
1'
1/
#454710000000
0!
0'
0/
#454720000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#454730000000
0!
0'
0/
#454740000000
1!
1'
1/
#454750000000
0!
0'
0/
#454760000000
1!
1'
1/
#454770000000
0!
0'
0/
#454780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#454790000000
0!
0'
0/
#454800000000
1!
1'
1/
#454810000000
0!
0'
0/
#454820000000
1!
1'
1/
#454830000000
0!
0'
0/
#454840000000
1!
1'
1/
#454850000000
0!
0'
0/
#454860000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#454870000000
0!
0'
0/
#454880000000
1!
1'
1/
#454890000000
0!
0'
0/
#454900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#454910000000
0!
0'
0/
#454920000000
1!
1'
1/
#454930000000
0!
0'
0/
#454940000000
#454950000000
1!
1'
1/
#454960000000
0!
0'
0/
#454970000000
1!
1'
1/
#454980000000
0!
1"
0'
1(
0/
10
#454990000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#455000000000
0!
0'
0/
#455010000000
1!
1'
1/
#455020000000
0!
0'
0/
#455030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#455040000000
0!
0'
0/
#455050000000
1!
1'
1/
#455060000000
0!
1"
0'
1(
0/
10
#455070000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#455080000000
0!
1$
0'
1+
0/
#455090000000
1!
1'
1/
#455100000000
0!
0'
0/
#455110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#455120000000
0!
0'
0/
#455130000000
1!
1'
1/
#455140000000
0!
0'
0/
#455150000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#455160000000
0!
0'
0/
#455170000000
1!
1'
1/
#455180000000
0!
0'
0/
#455190000000
1!
1'
1/
#455200000000
0!
0'
0/
#455210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#455220000000
0!
0'
0/
#455230000000
1!
1'
1/
#455240000000
0!
0'
0/
#455250000000
1!
1'
1/
#455260000000
0!
0'
0/
#455270000000
1!
1'
1/
#455280000000
0!
0'
0/
#455290000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#455300000000
0!
0'
0/
#455310000000
1!
1'
1/
#455320000000
0!
0'
0/
#455330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#455340000000
0!
0'
0/
#455350000000
1!
1'
1/
#455360000000
0!
0'
0/
#455370000000
#455380000000
1!
1'
1/
#455390000000
0!
0'
0/
#455400000000
1!
1'
1/
#455410000000
0!
1"
0'
1(
0/
10
#455420000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#455430000000
0!
0'
0/
#455440000000
1!
1'
1/
#455450000000
0!
0'
0/
#455460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#455470000000
0!
0'
0/
#455480000000
1!
1'
1/
#455490000000
0!
1"
0'
1(
0/
10
#455500000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#455510000000
0!
1$
0'
1+
0/
#455520000000
1!
1'
1/
#455530000000
0!
0'
0/
#455540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#455550000000
0!
0'
0/
#455560000000
1!
1'
1/
#455570000000
0!
0'
0/
#455580000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#455590000000
0!
0'
0/
#455600000000
1!
1'
1/
#455610000000
0!
0'
0/
#455620000000
1!
1'
1/
#455630000000
0!
0'
0/
#455640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#455650000000
0!
0'
0/
#455660000000
1!
1'
1/
#455670000000
0!
0'
0/
#455680000000
1!
1'
1/
#455690000000
0!
0'
0/
#455700000000
1!
1'
1/
#455710000000
0!
0'
0/
#455720000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#455730000000
0!
0'
0/
#455740000000
1!
1'
1/
#455750000000
0!
0'
0/
#455760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#455770000000
0!
0'
0/
#455780000000
1!
1'
1/
#455790000000
0!
0'
0/
#455800000000
#455810000000
1!
1'
1/
#455820000000
0!
0'
0/
#455830000000
1!
1'
1/
#455840000000
0!
1"
0'
1(
0/
10
#455850000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#455860000000
0!
0'
0/
#455870000000
1!
1'
1/
#455880000000
0!
0'
0/
#455890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#455900000000
0!
0'
0/
#455910000000
1!
1'
1/
#455920000000
0!
1"
0'
1(
0/
10
#455930000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#455940000000
0!
1$
0'
1+
0/
#455950000000
1!
1'
1/
#455960000000
0!
0'
0/
#455970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#455980000000
0!
0'
0/
#455990000000
1!
1'
1/
#456000000000
0!
0'
0/
#456010000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#456020000000
0!
0'
0/
#456030000000
1!
1'
1/
#456040000000
0!
0'
0/
#456050000000
1!
1'
1/
#456060000000
0!
0'
0/
#456070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#456080000000
0!
0'
0/
#456090000000
1!
1'
1/
#456100000000
0!
0'
0/
#456110000000
1!
1'
1/
#456120000000
0!
0'
0/
#456130000000
1!
1'
1/
#456140000000
0!
0'
0/
#456150000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#456160000000
0!
0'
0/
#456170000000
1!
1'
1/
#456180000000
0!
0'
0/
#456190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#456200000000
0!
0'
0/
#456210000000
1!
1'
1/
#456220000000
0!
0'
0/
#456230000000
#456240000000
1!
1'
1/
#456250000000
0!
0'
0/
#456260000000
1!
1'
1/
#456270000000
0!
1"
0'
1(
0/
10
#456280000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#456290000000
0!
0'
0/
#456300000000
1!
1'
1/
#456310000000
0!
0'
0/
#456320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#456330000000
0!
0'
0/
#456340000000
1!
1'
1/
#456350000000
0!
1"
0'
1(
0/
10
#456360000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#456370000000
0!
1$
0'
1+
0/
#456380000000
1!
1'
1/
#456390000000
0!
0'
0/
#456400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#456410000000
0!
0'
0/
#456420000000
1!
1'
1/
#456430000000
0!
0'
0/
#456440000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#456450000000
0!
0'
0/
#456460000000
1!
1'
1/
#456470000000
0!
0'
0/
#456480000000
1!
1'
1/
#456490000000
0!
0'
0/
#456500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#456510000000
0!
0'
0/
#456520000000
1!
1'
1/
#456530000000
0!
0'
0/
#456540000000
1!
1'
1/
#456550000000
0!
0'
0/
#456560000000
1!
1'
1/
#456570000000
0!
0'
0/
#456580000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#456590000000
0!
0'
0/
#456600000000
1!
1'
1/
#456610000000
0!
0'
0/
#456620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#456630000000
0!
0'
0/
#456640000000
1!
1'
1/
#456650000000
0!
0'
0/
#456660000000
#456670000000
1!
1'
1/
#456680000000
0!
0'
0/
#456690000000
1!
1'
1/
#456700000000
0!
1"
0'
1(
0/
10
#456710000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#456720000000
0!
0'
0/
#456730000000
1!
1'
1/
#456740000000
0!
0'
0/
#456750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#456760000000
0!
0'
0/
#456770000000
1!
1'
1/
#456780000000
0!
1"
0'
1(
0/
10
#456790000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#456800000000
0!
1$
0'
1+
0/
#456810000000
1!
1'
1/
#456820000000
0!
0'
0/
#456830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#456840000000
0!
0'
0/
#456850000000
1!
1'
1/
#456860000000
0!
0'
0/
#456870000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#456880000000
0!
0'
0/
#456890000000
1!
1'
1/
#456900000000
0!
0'
0/
#456910000000
1!
1'
1/
#456920000000
0!
0'
0/
#456930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#456940000000
0!
0'
0/
#456950000000
1!
1'
1/
#456960000000
0!
0'
0/
#456970000000
1!
1'
1/
#456980000000
0!
0'
0/
#456990000000
1!
1'
1/
#457000000000
0!
0'
0/
#457010000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#457020000000
0!
0'
0/
#457030000000
1!
1'
1/
#457040000000
0!
0'
0/
#457050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#457060000000
0!
0'
0/
#457070000000
1!
1'
1/
#457080000000
0!
0'
0/
#457090000000
#457100000000
1!
1'
1/
#457110000000
0!
0'
0/
#457120000000
1!
1'
1/
#457130000000
0!
1"
0'
1(
0/
10
#457140000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#457150000000
0!
0'
0/
#457160000000
1!
1'
1/
#457170000000
0!
0'
0/
#457180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#457190000000
0!
0'
0/
#457200000000
1!
1'
1/
#457210000000
0!
1"
0'
1(
0/
10
#457220000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#457230000000
0!
1$
0'
1+
0/
#457240000000
1!
1'
1/
#457250000000
0!
0'
0/
#457260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#457270000000
0!
0'
0/
#457280000000
1!
1'
1/
#457290000000
0!
0'
0/
#457300000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#457310000000
0!
0'
0/
#457320000000
1!
1'
1/
#457330000000
0!
0'
0/
#457340000000
1!
1'
1/
#457350000000
0!
0'
0/
#457360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#457370000000
0!
0'
0/
#457380000000
1!
1'
1/
#457390000000
0!
0'
0/
#457400000000
1!
1'
1/
#457410000000
0!
0'
0/
#457420000000
1!
1'
1/
#457430000000
0!
0'
0/
#457440000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#457450000000
0!
0'
0/
#457460000000
1!
1'
1/
#457470000000
0!
0'
0/
#457480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#457490000000
0!
0'
0/
#457500000000
1!
1'
1/
#457510000000
0!
0'
0/
#457520000000
#457530000000
1!
1'
1/
#457540000000
0!
0'
0/
#457550000000
1!
1'
1/
#457560000000
0!
1"
0'
1(
0/
10
#457570000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#457580000000
0!
0'
0/
#457590000000
1!
1'
1/
#457600000000
0!
0'
0/
#457610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#457620000000
0!
0'
0/
#457630000000
1!
1'
1/
#457640000000
0!
1"
0'
1(
0/
10
#457650000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#457660000000
0!
1$
0'
1+
0/
#457670000000
1!
1'
1/
#457680000000
0!
0'
0/
#457690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#457700000000
0!
0'
0/
#457710000000
1!
1'
1/
#457720000000
0!
0'
0/
#457730000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#457740000000
0!
0'
0/
#457750000000
1!
1'
1/
#457760000000
0!
0'
0/
#457770000000
1!
1'
1/
#457780000000
0!
0'
0/
#457790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#457800000000
0!
0'
0/
#457810000000
1!
1'
1/
#457820000000
0!
0'
0/
#457830000000
1!
1'
1/
#457840000000
0!
0'
0/
#457850000000
1!
1'
1/
#457860000000
0!
0'
0/
#457870000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#457880000000
0!
0'
0/
#457890000000
1!
1'
1/
#457900000000
0!
0'
0/
#457910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#457920000000
0!
0'
0/
#457930000000
1!
1'
1/
#457940000000
0!
0'
0/
#457950000000
#457960000000
1!
1'
1/
#457970000000
0!
0'
0/
#457980000000
1!
1'
1/
#457990000000
0!
1"
0'
1(
0/
10
#458000000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#458010000000
0!
0'
0/
#458020000000
1!
1'
1/
#458030000000
0!
0'
0/
#458040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#458050000000
0!
0'
0/
#458060000000
1!
1'
1/
#458070000000
0!
1"
0'
1(
0/
10
#458080000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#458090000000
0!
1$
0'
1+
0/
#458100000000
1!
1'
1/
#458110000000
0!
0'
0/
#458120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#458130000000
0!
0'
0/
#458140000000
1!
1'
1/
#458150000000
0!
0'
0/
#458160000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#458170000000
0!
0'
0/
#458180000000
1!
1'
1/
#458190000000
0!
0'
0/
#458200000000
1!
1'
1/
#458210000000
0!
0'
0/
#458220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#458230000000
0!
0'
0/
#458240000000
1!
1'
1/
#458250000000
0!
0'
0/
#458260000000
1!
1'
1/
#458270000000
0!
0'
0/
#458280000000
1!
1'
1/
#458290000000
0!
0'
0/
#458300000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#458310000000
0!
0'
0/
#458320000000
1!
1'
1/
#458330000000
0!
0'
0/
#458340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#458350000000
0!
0'
0/
#458360000000
1!
1'
1/
#458370000000
0!
0'
0/
#458380000000
#458390000000
1!
1'
1/
#458400000000
0!
0'
0/
#458410000000
1!
1'
1/
#458420000000
0!
1"
0'
1(
0/
10
#458430000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#458440000000
0!
0'
0/
#458450000000
1!
1'
1/
#458460000000
0!
0'
0/
#458470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#458480000000
0!
0'
0/
#458490000000
1!
1'
1/
#458500000000
0!
1"
0'
1(
0/
10
#458510000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#458520000000
0!
1$
0'
1+
0/
#458530000000
1!
1'
1/
#458540000000
0!
0'
0/
#458550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#458560000000
0!
0'
0/
#458570000000
1!
1'
1/
#458580000000
0!
0'
0/
#458590000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#458600000000
0!
0'
0/
#458610000000
1!
1'
1/
#458620000000
0!
0'
0/
#458630000000
1!
1'
1/
#458640000000
0!
0'
0/
#458650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#458660000000
0!
0'
0/
#458670000000
1!
1'
1/
#458680000000
0!
0'
0/
#458690000000
1!
1'
1/
#458700000000
0!
0'
0/
#458710000000
1!
1'
1/
#458720000000
0!
0'
0/
#458730000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#458740000000
0!
0'
0/
#458750000000
1!
1'
1/
#458760000000
0!
0'
0/
#458770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#458780000000
0!
0'
0/
#458790000000
1!
1'
1/
#458800000000
0!
0'
0/
#458810000000
#458820000000
1!
1'
1/
#458830000000
0!
0'
0/
#458840000000
1!
1'
1/
#458850000000
0!
1"
0'
1(
0/
10
#458860000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#458870000000
0!
0'
0/
#458880000000
1!
1'
1/
#458890000000
0!
0'
0/
#458900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#458910000000
0!
0'
0/
#458920000000
1!
1'
1/
#458930000000
0!
1"
0'
1(
0/
10
#458940000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#458950000000
0!
1$
0'
1+
0/
#458960000000
1!
1'
1/
#458970000000
0!
0'
0/
#458980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#458990000000
0!
0'
0/
#459000000000
1!
1'
1/
#459010000000
0!
0'
0/
#459020000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#459030000000
0!
0'
0/
#459040000000
1!
1'
1/
#459050000000
0!
0'
0/
#459060000000
1!
1'
1/
#459070000000
0!
0'
0/
#459080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#459090000000
0!
0'
0/
#459100000000
1!
1'
1/
#459110000000
0!
0'
0/
#459120000000
1!
1'
1/
#459130000000
0!
0'
0/
#459140000000
1!
1'
1/
#459150000000
0!
0'
0/
#459160000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#459170000000
0!
0'
0/
#459180000000
1!
1'
1/
#459190000000
0!
0'
0/
#459200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#459210000000
0!
0'
0/
#459220000000
1!
1'
1/
#459230000000
0!
0'
0/
#459240000000
#459250000000
1!
1'
1/
#459260000000
0!
0'
0/
#459270000000
1!
1'
1/
#459280000000
0!
1"
0'
1(
0/
10
#459290000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#459300000000
0!
0'
0/
#459310000000
1!
1'
1/
#459320000000
0!
0'
0/
#459330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#459340000000
0!
0'
0/
#459350000000
1!
1'
1/
#459360000000
0!
1"
0'
1(
0/
10
#459370000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#459380000000
0!
1$
0'
1+
0/
#459390000000
1!
1'
1/
#459400000000
0!
0'
0/
#459410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#459420000000
0!
0'
0/
#459430000000
1!
1'
1/
#459440000000
0!
0'
0/
#459450000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#459460000000
0!
0'
0/
#459470000000
1!
1'
1/
#459480000000
0!
0'
0/
#459490000000
1!
1'
1/
#459500000000
0!
0'
0/
#459510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#459520000000
0!
0'
0/
#459530000000
1!
1'
1/
#459540000000
0!
0'
0/
#459550000000
1!
1'
1/
#459560000000
0!
0'
0/
#459570000000
1!
1'
1/
#459580000000
0!
0'
0/
#459590000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#459600000000
0!
0'
0/
#459610000000
1!
1'
1/
#459620000000
0!
0'
0/
#459630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#459640000000
0!
0'
0/
#459650000000
1!
1'
1/
#459660000000
0!
0'
0/
#459670000000
#459680000000
1!
1'
1/
#459690000000
0!
0'
0/
#459700000000
1!
1'
1/
#459710000000
0!
1"
0'
1(
0/
10
#459720000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#459730000000
0!
0'
0/
#459740000000
1!
1'
1/
#459750000000
0!
0'
0/
#459760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#459770000000
0!
0'
0/
#459780000000
1!
1'
1/
#459790000000
0!
1"
0'
1(
0/
10
#459800000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#459810000000
0!
1$
0'
1+
0/
#459820000000
1!
1'
1/
#459830000000
0!
0'
0/
#459840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#459850000000
0!
0'
0/
#459860000000
1!
1'
1/
#459870000000
0!
0'
0/
#459880000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#459890000000
0!
0'
0/
#459900000000
1!
1'
1/
#459910000000
0!
0'
0/
#459920000000
1!
1'
1/
#459930000000
0!
0'
0/
#459940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#459950000000
0!
0'
0/
#459960000000
1!
1'
1/
#459970000000
0!
0'
0/
#459980000000
1!
1'
1/
#459990000000
0!
0'
0/
#460000000000
1!
1'
1/
#460010000000
0!
0'
0/
#460020000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#460030000000
0!
0'
0/
#460040000000
1!
1'
1/
#460050000000
0!
0'
0/
#460060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#460070000000
0!
0'
0/
#460080000000
1!
1'
1/
#460090000000
0!
0'
0/
#460100000000
#460110000000
1!
1'
1/
#460120000000
0!
0'
0/
#460130000000
1!
1'
1/
#460140000000
0!
1"
0'
1(
0/
10
#460150000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#460160000000
0!
0'
0/
#460170000000
1!
1'
1/
#460180000000
0!
0'
0/
#460190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#460200000000
0!
0'
0/
#460210000000
1!
1'
1/
#460220000000
0!
1"
0'
1(
0/
10
#460230000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#460240000000
0!
1$
0'
1+
0/
#460250000000
1!
1'
1/
#460260000000
0!
0'
0/
#460270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#460280000000
0!
0'
0/
#460290000000
1!
1'
1/
#460300000000
0!
0'
0/
#460310000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#460320000000
0!
0'
0/
#460330000000
1!
1'
1/
#460340000000
0!
0'
0/
#460350000000
1!
1'
1/
#460360000000
0!
0'
0/
#460370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#460380000000
0!
0'
0/
#460390000000
1!
1'
1/
#460400000000
0!
0'
0/
#460410000000
1!
1'
1/
#460420000000
0!
0'
0/
#460430000000
1!
1'
1/
#460440000000
0!
0'
0/
#460450000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#460460000000
0!
0'
0/
#460470000000
1!
1'
1/
#460480000000
0!
0'
0/
#460490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#460500000000
0!
0'
0/
#460510000000
1!
1'
1/
#460520000000
0!
0'
0/
#460530000000
#460540000000
1!
1'
1/
#460550000000
0!
0'
0/
#460560000000
1!
1'
1/
#460570000000
0!
1"
0'
1(
0/
10
#460580000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#460590000000
0!
0'
0/
#460600000000
1!
1'
1/
#460610000000
0!
0'
0/
#460620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#460630000000
0!
0'
0/
#460640000000
1!
1'
1/
#460650000000
0!
1"
0'
1(
0/
10
#460660000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#460670000000
0!
1$
0'
1+
0/
#460680000000
1!
1'
1/
#460690000000
0!
0'
0/
#460700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#460710000000
0!
0'
0/
#460720000000
1!
1'
1/
#460730000000
0!
0'
0/
#460740000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#460750000000
0!
0'
0/
#460760000000
1!
1'
1/
#460770000000
0!
0'
0/
#460780000000
1!
1'
1/
#460790000000
0!
0'
0/
#460800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#460810000000
0!
0'
0/
#460820000000
1!
1'
1/
#460830000000
0!
0'
0/
#460840000000
1!
1'
1/
#460850000000
0!
0'
0/
#460860000000
1!
1'
1/
#460870000000
0!
0'
0/
#460880000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#460890000000
0!
0'
0/
#460900000000
1!
1'
1/
#460910000000
0!
0'
0/
#460920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#460930000000
0!
0'
0/
#460940000000
1!
1'
1/
#460950000000
0!
0'
0/
#460960000000
#460970000000
1!
1'
1/
#460980000000
0!
0'
0/
#460990000000
1!
1'
1/
#461000000000
0!
1"
0'
1(
0/
10
#461010000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#461020000000
0!
0'
0/
#461030000000
1!
1'
1/
#461040000000
0!
0'
0/
#461050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#461060000000
0!
0'
0/
#461070000000
1!
1'
1/
#461080000000
0!
1"
0'
1(
0/
10
#461090000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#461100000000
0!
1$
0'
1+
0/
#461110000000
1!
1'
1/
#461120000000
0!
0'
0/
#461130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#461140000000
0!
0'
0/
#461150000000
1!
1'
1/
#461160000000
0!
0'
0/
#461170000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#461180000000
0!
0'
0/
#461190000000
1!
1'
1/
#461200000000
0!
0'
0/
#461210000000
1!
1'
1/
#461220000000
0!
0'
0/
#461230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#461240000000
0!
0'
0/
#461250000000
1!
1'
1/
#461260000000
0!
0'
0/
#461270000000
1!
1'
1/
#461280000000
0!
0'
0/
#461290000000
1!
1'
1/
#461300000000
0!
0'
0/
#461310000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#461320000000
0!
0'
0/
#461330000000
1!
1'
1/
#461340000000
0!
0'
0/
#461350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#461360000000
0!
0'
0/
#461370000000
1!
1'
1/
#461380000000
0!
0'
0/
#461390000000
#461400000000
1!
1'
1/
#461410000000
0!
0'
0/
#461420000000
1!
1'
1/
#461430000000
0!
1"
0'
1(
0/
10
#461440000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#461450000000
0!
0'
0/
#461460000000
1!
1'
1/
#461470000000
0!
0'
0/
#461480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#461490000000
0!
0'
0/
#461500000000
1!
1'
1/
#461510000000
0!
1"
0'
1(
0/
10
#461520000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#461530000000
0!
1$
0'
1+
0/
#461540000000
1!
1'
1/
#461550000000
0!
0'
0/
#461560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#461570000000
0!
0'
0/
#461580000000
1!
1'
1/
#461590000000
0!
0'
0/
#461600000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#461610000000
0!
0'
0/
#461620000000
1!
1'
1/
#461630000000
0!
0'
0/
#461640000000
1!
1'
1/
#461650000000
0!
0'
0/
#461660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#461670000000
0!
0'
0/
#461680000000
1!
1'
1/
#461690000000
0!
0'
0/
#461700000000
1!
1'
1/
#461710000000
0!
0'
0/
#461720000000
1!
1'
1/
#461730000000
0!
0'
0/
#461740000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#461750000000
0!
0'
0/
#461760000000
1!
1'
1/
#461770000000
0!
0'
0/
#461780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#461790000000
0!
0'
0/
#461800000000
1!
1'
1/
#461810000000
0!
0'
0/
#461820000000
#461830000000
1!
1'
1/
#461840000000
0!
0'
0/
#461850000000
1!
1'
1/
#461860000000
0!
1"
0'
1(
0/
10
#461870000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#461880000000
0!
0'
0/
#461890000000
1!
1'
1/
#461900000000
0!
0'
0/
#461910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#461920000000
0!
0'
0/
#461930000000
1!
1'
1/
#461940000000
0!
1"
0'
1(
0/
10
#461950000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#461960000000
0!
1$
0'
1+
0/
#461970000000
1!
1'
1/
#461980000000
0!
0'
0/
#461990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#462000000000
0!
0'
0/
#462010000000
1!
1'
1/
#462020000000
0!
0'
0/
#462030000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#462040000000
0!
0'
0/
#462050000000
1!
1'
1/
#462060000000
0!
0'
0/
#462070000000
1!
1'
1/
#462080000000
0!
0'
0/
#462090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#462100000000
0!
0'
0/
#462110000000
1!
1'
1/
#462120000000
0!
0'
0/
#462130000000
1!
1'
1/
#462140000000
0!
0'
0/
#462150000000
1!
1'
1/
#462160000000
0!
0'
0/
#462170000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#462180000000
0!
0'
0/
#462190000000
1!
1'
1/
#462200000000
0!
0'
0/
#462210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#462220000000
0!
0'
0/
#462230000000
1!
1'
1/
#462240000000
0!
0'
0/
#462250000000
#462260000000
1!
1'
1/
#462270000000
0!
0'
0/
#462280000000
1!
1'
1/
#462290000000
0!
1"
0'
1(
0/
10
#462300000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#462310000000
0!
0'
0/
#462320000000
1!
1'
1/
#462330000000
0!
0'
0/
#462340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#462350000000
0!
0'
0/
#462360000000
1!
1'
1/
#462370000000
0!
1"
0'
1(
0/
10
#462380000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#462390000000
0!
1$
0'
1+
0/
#462400000000
1!
1'
1/
#462410000000
0!
0'
0/
#462420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#462430000000
0!
0'
0/
#462440000000
1!
1'
1/
#462450000000
0!
0'
0/
#462460000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#462470000000
0!
0'
0/
#462480000000
1!
1'
1/
#462490000000
0!
0'
0/
#462500000000
1!
1'
1/
#462510000000
0!
0'
0/
#462520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#462530000000
0!
0'
0/
#462540000000
1!
1'
1/
#462550000000
0!
0'
0/
#462560000000
1!
1'
1/
#462570000000
0!
0'
0/
#462580000000
1!
1'
1/
#462590000000
0!
0'
0/
#462600000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#462610000000
0!
0'
0/
#462620000000
1!
1'
1/
#462630000000
0!
0'
0/
#462640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#462650000000
0!
0'
0/
#462660000000
1!
1'
1/
#462670000000
0!
0'
0/
#462680000000
#462690000000
1!
1'
1/
#462700000000
0!
0'
0/
#462710000000
1!
1'
1/
#462720000000
0!
1"
0'
1(
0/
10
#462730000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#462740000000
0!
0'
0/
#462750000000
1!
1'
1/
#462760000000
0!
0'
0/
#462770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#462780000000
0!
0'
0/
#462790000000
1!
1'
1/
#462800000000
0!
1"
0'
1(
0/
10
#462810000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#462820000000
0!
1$
0'
1+
0/
#462830000000
1!
1'
1/
#462840000000
0!
0'
0/
#462850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#462860000000
0!
0'
0/
#462870000000
1!
1'
1/
#462880000000
0!
0'
0/
#462890000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#462900000000
0!
0'
0/
#462910000000
1!
1'
1/
#462920000000
0!
0'
0/
#462930000000
1!
1'
1/
#462940000000
0!
0'
0/
#462950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#462960000000
0!
0'
0/
#462970000000
1!
1'
1/
#462980000000
0!
0'
0/
#462990000000
1!
1'
1/
#463000000000
0!
0'
0/
#463010000000
1!
1'
1/
#463020000000
0!
0'
0/
#463030000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#463040000000
0!
0'
0/
#463050000000
1!
1'
1/
#463060000000
0!
0'
0/
#463070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#463080000000
0!
0'
0/
#463090000000
1!
1'
1/
#463100000000
0!
0'
0/
#463110000000
#463120000000
1!
1'
1/
#463130000000
0!
0'
0/
#463140000000
1!
1'
1/
#463150000000
0!
1"
0'
1(
0/
10
#463160000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#463170000000
0!
0'
0/
#463180000000
1!
1'
1/
#463190000000
0!
0'
0/
#463200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#463210000000
0!
0'
0/
#463220000000
1!
1'
1/
#463230000000
0!
1"
0'
1(
0/
10
#463240000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#463250000000
0!
1$
0'
1+
0/
#463260000000
1!
1'
1/
#463270000000
0!
0'
0/
#463280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#463290000000
0!
0'
0/
#463300000000
1!
1'
1/
#463310000000
0!
0'
0/
#463320000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#463330000000
0!
0'
0/
#463340000000
1!
1'
1/
#463350000000
0!
0'
0/
#463360000000
1!
1'
1/
#463370000000
0!
0'
0/
#463380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#463390000000
0!
0'
0/
#463400000000
1!
1'
1/
#463410000000
0!
0'
0/
#463420000000
1!
1'
1/
#463430000000
0!
0'
0/
#463440000000
1!
1'
1/
#463450000000
0!
0'
0/
#463460000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#463470000000
0!
0'
0/
#463480000000
1!
1'
1/
#463490000000
0!
0'
0/
#463500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#463510000000
0!
0'
0/
#463520000000
1!
1'
1/
#463530000000
0!
0'
0/
#463540000000
#463550000000
1!
1'
1/
#463560000000
0!
0'
0/
#463570000000
1!
1'
1/
#463580000000
0!
1"
0'
1(
0/
10
#463590000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#463600000000
0!
0'
0/
#463610000000
1!
1'
1/
#463620000000
0!
0'
0/
#463630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#463640000000
0!
0'
0/
#463650000000
1!
1'
1/
#463660000000
0!
1"
0'
1(
0/
10
#463670000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#463680000000
0!
1$
0'
1+
0/
#463690000000
1!
1'
1/
#463700000000
0!
0'
0/
#463710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#463720000000
0!
0'
0/
#463730000000
1!
1'
1/
#463740000000
0!
0'
0/
#463750000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#463760000000
0!
0'
0/
#463770000000
1!
1'
1/
#463780000000
0!
0'
0/
#463790000000
1!
1'
1/
#463800000000
0!
0'
0/
#463810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#463820000000
0!
0'
0/
#463830000000
1!
1'
1/
#463840000000
0!
0'
0/
#463850000000
1!
1'
1/
#463860000000
0!
0'
0/
#463870000000
1!
1'
1/
#463880000000
0!
0'
0/
#463890000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#463900000000
0!
0'
0/
#463910000000
1!
1'
1/
#463920000000
0!
0'
0/
#463930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#463940000000
0!
0'
0/
#463950000000
1!
1'
1/
#463960000000
0!
0'
0/
#463970000000
#463980000000
1!
1'
1/
#463990000000
0!
0'
0/
#464000000000
1!
1'
1/
#464010000000
0!
1"
0'
1(
0/
10
#464020000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#464030000000
0!
0'
0/
#464040000000
1!
1'
1/
#464050000000
0!
0'
0/
#464060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#464070000000
0!
0'
0/
#464080000000
1!
1'
1/
#464090000000
0!
1"
0'
1(
0/
10
#464100000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#464110000000
0!
1$
0'
1+
0/
#464120000000
1!
1'
1/
#464130000000
0!
0'
0/
#464140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#464150000000
0!
0'
0/
#464160000000
1!
1'
1/
#464170000000
0!
0'
0/
#464180000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#464190000000
0!
0'
0/
#464200000000
1!
1'
1/
#464210000000
0!
0'
0/
#464220000000
1!
1'
1/
#464230000000
0!
0'
0/
#464240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#464250000000
0!
0'
0/
#464260000000
1!
1'
1/
#464270000000
0!
0'
0/
#464280000000
1!
1'
1/
#464290000000
0!
0'
0/
#464300000000
1!
1'
1/
#464310000000
0!
0'
0/
#464320000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#464330000000
0!
0'
0/
#464340000000
1!
1'
1/
#464350000000
0!
0'
0/
#464360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#464370000000
0!
0'
0/
#464380000000
1!
1'
1/
#464390000000
0!
0'
0/
#464400000000
#464410000000
1!
1'
1/
#464420000000
0!
0'
0/
#464430000000
1!
1'
1/
#464440000000
0!
1"
0'
1(
0/
10
#464450000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#464460000000
0!
0'
0/
#464470000000
1!
1'
1/
#464480000000
0!
0'
0/
#464490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#464500000000
0!
0'
0/
#464510000000
1!
1'
1/
#464520000000
0!
1"
0'
1(
0/
10
#464530000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#464540000000
0!
1$
0'
1+
0/
#464550000000
1!
1'
1/
#464560000000
0!
0'
0/
#464570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#464580000000
0!
0'
0/
#464590000000
1!
1'
1/
#464600000000
0!
0'
0/
#464610000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#464620000000
0!
0'
0/
#464630000000
1!
1'
1/
#464640000000
0!
0'
0/
#464650000000
1!
1'
1/
#464660000000
0!
0'
0/
#464670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#464680000000
0!
0'
0/
#464690000000
1!
1'
1/
#464700000000
0!
0'
0/
#464710000000
1!
1'
1/
#464720000000
0!
0'
0/
#464730000000
1!
1'
1/
#464740000000
0!
0'
0/
#464750000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#464760000000
0!
0'
0/
#464770000000
1!
1'
1/
#464780000000
0!
0'
0/
#464790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#464800000000
0!
0'
0/
#464810000000
1!
1'
1/
#464820000000
0!
0'
0/
#464830000000
#464840000000
1!
1'
1/
#464850000000
0!
0'
0/
#464860000000
1!
1'
1/
#464870000000
0!
1"
0'
1(
0/
10
#464880000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#464890000000
0!
0'
0/
#464900000000
1!
1'
1/
#464910000000
0!
0'
0/
#464920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#464930000000
0!
0'
0/
#464940000000
1!
1'
1/
#464950000000
0!
1"
0'
1(
0/
10
#464960000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#464970000000
0!
1$
0'
1+
0/
#464980000000
1!
1'
1/
#464990000000
0!
0'
0/
#465000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#465010000000
0!
0'
0/
#465020000000
1!
1'
1/
#465030000000
0!
0'
0/
#465040000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#465050000000
0!
0'
0/
#465060000000
1!
1'
1/
#465070000000
0!
0'
0/
#465080000000
1!
1'
1/
#465090000000
0!
0'
0/
#465100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#465110000000
0!
0'
0/
#465120000000
1!
1'
1/
#465130000000
0!
0'
0/
#465140000000
1!
1'
1/
#465150000000
0!
0'
0/
#465160000000
1!
1'
1/
#465170000000
0!
0'
0/
#465180000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#465190000000
0!
0'
0/
#465200000000
1!
1'
1/
#465210000000
0!
0'
0/
#465220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#465230000000
0!
0'
0/
#465240000000
1!
1'
1/
#465250000000
0!
0'
0/
#465260000000
#465270000000
1!
1'
1/
#465280000000
0!
0'
0/
#465290000000
1!
1'
1/
#465300000000
0!
1"
0'
1(
0/
10
#465310000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#465320000000
0!
0'
0/
#465330000000
1!
1'
1/
#465340000000
0!
0'
0/
#465350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#465360000000
0!
0'
0/
#465370000000
1!
1'
1/
#465380000000
0!
1"
0'
1(
0/
10
#465390000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#465400000000
0!
1$
0'
1+
0/
#465410000000
1!
1'
1/
#465420000000
0!
0'
0/
#465430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#465440000000
0!
0'
0/
#465450000000
1!
1'
1/
#465460000000
0!
0'
0/
#465470000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#465480000000
0!
0'
0/
#465490000000
1!
1'
1/
#465500000000
0!
0'
0/
#465510000000
1!
1'
1/
#465520000000
0!
0'
0/
#465530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#465540000000
0!
0'
0/
#465550000000
1!
1'
1/
#465560000000
0!
0'
0/
#465570000000
1!
1'
1/
#465580000000
0!
0'
0/
#465590000000
1!
1'
1/
#465600000000
0!
0'
0/
#465610000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#465620000000
0!
0'
0/
#465630000000
1!
1'
1/
#465640000000
0!
0'
0/
#465650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#465660000000
0!
0'
0/
#465670000000
1!
1'
1/
#465680000000
0!
0'
0/
#465690000000
#465700000000
1!
1'
1/
#465710000000
0!
0'
0/
#465720000000
1!
1'
1/
#465730000000
0!
1"
0'
1(
0/
10
#465740000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#465750000000
0!
0'
0/
#465760000000
1!
1'
1/
#465770000000
0!
0'
0/
#465780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#465790000000
0!
0'
0/
#465800000000
1!
1'
1/
#465810000000
0!
1"
0'
1(
0/
10
#465820000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#465830000000
0!
1$
0'
1+
0/
#465840000000
1!
1'
1/
#465850000000
0!
0'
0/
#465860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#465870000000
0!
0'
0/
#465880000000
1!
1'
1/
#465890000000
0!
0'
0/
#465900000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#465910000000
0!
0'
0/
#465920000000
1!
1'
1/
#465930000000
0!
0'
0/
#465940000000
1!
1'
1/
#465950000000
0!
0'
0/
#465960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#465970000000
0!
0'
0/
#465980000000
1!
1'
1/
#465990000000
0!
0'
0/
#466000000000
1!
1'
1/
#466010000000
0!
0'
0/
#466020000000
1!
1'
1/
#466030000000
0!
0'
0/
#466040000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#466050000000
0!
0'
0/
#466060000000
1!
1'
1/
#466070000000
0!
0'
0/
#466080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#466090000000
0!
0'
0/
#466100000000
1!
1'
1/
#466110000000
0!
0'
0/
#466120000000
#466130000000
1!
1'
1/
#466140000000
0!
0'
0/
#466150000000
1!
1'
1/
#466160000000
0!
1"
0'
1(
0/
10
#466170000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#466180000000
0!
0'
0/
#466190000000
1!
1'
1/
#466200000000
0!
0'
0/
#466210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#466220000000
0!
0'
0/
#466230000000
1!
1'
1/
#466240000000
0!
1"
0'
1(
0/
10
#466250000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#466260000000
0!
1$
0'
1+
0/
#466270000000
1!
1'
1/
#466280000000
0!
0'
0/
#466290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#466300000000
0!
0'
0/
#466310000000
1!
1'
1/
#466320000000
0!
0'
0/
#466330000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#466340000000
0!
0'
0/
#466350000000
1!
1'
1/
#466360000000
0!
0'
0/
#466370000000
1!
1'
1/
#466380000000
0!
0'
0/
#466390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#466400000000
0!
0'
0/
#466410000000
1!
1'
1/
#466420000000
0!
0'
0/
#466430000000
1!
1'
1/
#466440000000
0!
0'
0/
#466450000000
1!
1'
1/
#466460000000
0!
0'
0/
#466470000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#466480000000
0!
0'
0/
#466490000000
1!
1'
1/
#466500000000
0!
0'
0/
#466510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#466520000000
0!
0'
0/
#466530000000
1!
1'
1/
#466540000000
0!
0'
0/
#466550000000
#466560000000
1!
1'
1/
#466570000000
0!
0'
0/
#466580000000
1!
1'
1/
#466590000000
0!
1"
0'
1(
0/
10
#466600000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#466610000000
0!
0'
0/
#466620000000
1!
1'
1/
#466630000000
0!
0'
0/
#466640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#466650000000
0!
0'
0/
#466660000000
1!
1'
1/
#466670000000
0!
1"
0'
1(
0/
10
#466680000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#466690000000
0!
1$
0'
1+
0/
#466700000000
1!
1'
1/
#466710000000
0!
0'
0/
#466720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#466730000000
0!
0'
0/
#466740000000
1!
1'
1/
#466750000000
0!
0'
0/
#466760000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#466770000000
0!
0'
0/
#466780000000
1!
1'
1/
#466790000000
0!
0'
0/
#466800000000
1!
1'
1/
#466810000000
0!
0'
0/
#466820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#466830000000
0!
0'
0/
#466840000000
1!
1'
1/
#466850000000
0!
0'
0/
#466860000000
1!
1'
1/
#466870000000
0!
0'
0/
#466880000000
1!
1'
1/
#466890000000
0!
0'
0/
#466900000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#466910000000
0!
0'
0/
#466920000000
1!
1'
1/
#466930000000
0!
0'
0/
#466940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#466950000000
0!
0'
0/
#466960000000
1!
1'
1/
#466970000000
0!
0'
0/
#466980000000
#466990000000
1!
1'
1/
#467000000000
0!
0'
0/
#467010000000
1!
1'
1/
#467020000000
0!
1"
0'
1(
0/
10
#467030000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#467040000000
0!
0'
0/
#467050000000
1!
1'
1/
#467060000000
0!
0'
0/
#467070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#467080000000
0!
0'
0/
#467090000000
1!
1'
1/
#467100000000
0!
1"
0'
1(
0/
10
#467110000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#467120000000
0!
1$
0'
1+
0/
#467130000000
1!
1'
1/
#467140000000
0!
0'
0/
#467150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#467160000000
0!
0'
0/
#467170000000
1!
1'
1/
#467180000000
0!
0'
0/
#467190000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#467200000000
0!
0'
0/
#467210000000
1!
1'
1/
#467220000000
0!
0'
0/
#467230000000
1!
1'
1/
#467240000000
0!
0'
0/
#467250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#467260000000
0!
0'
0/
#467270000000
1!
1'
1/
#467280000000
0!
0'
0/
#467290000000
1!
1'
1/
#467300000000
0!
0'
0/
#467310000000
1!
1'
1/
#467320000000
0!
0'
0/
#467330000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#467340000000
0!
0'
0/
#467350000000
1!
1'
1/
#467360000000
0!
0'
0/
#467370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#467380000000
0!
0'
0/
#467390000000
1!
1'
1/
#467400000000
0!
0'
0/
#467410000000
#467420000000
1!
1'
1/
#467430000000
0!
0'
0/
#467440000000
1!
1'
1/
#467450000000
0!
1"
0'
1(
0/
10
#467460000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#467470000000
0!
0'
0/
#467480000000
1!
1'
1/
#467490000000
0!
0'
0/
#467500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#467510000000
0!
0'
0/
#467520000000
1!
1'
1/
#467530000000
0!
1"
0'
1(
0/
10
#467540000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#467550000000
0!
1$
0'
1+
0/
#467560000000
1!
1'
1/
#467570000000
0!
0'
0/
#467580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#467590000000
0!
0'
0/
#467600000000
1!
1'
1/
#467610000000
0!
0'
0/
#467620000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#467630000000
0!
0'
0/
#467640000000
1!
1'
1/
#467650000000
0!
0'
0/
#467660000000
1!
1'
1/
#467670000000
0!
0'
0/
#467680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#467690000000
0!
0'
0/
#467700000000
1!
1'
1/
#467710000000
0!
0'
0/
#467720000000
1!
1'
1/
#467730000000
0!
0'
0/
#467740000000
1!
1'
1/
#467750000000
0!
0'
0/
#467760000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#467770000000
0!
0'
0/
#467780000000
1!
1'
1/
#467790000000
0!
0'
0/
#467800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#467810000000
0!
0'
0/
#467820000000
1!
1'
1/
#467830000000
0!
0'
0/
#467840000000
#467850000000
1!
1'
1/
#467860000000
0!
0'
0/
#467870000000
1!
1'
1/
#467880000000
0!
1"
0'
1(
0/
10
#467890000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#467900000000
0!
0'
0/
#467910000000
1!
1'
1/
#467920000000
0!
0'
0/
#467930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#467940000000
0!
0'
0/
#467950000000
1!
1'
1/
#467960000000
0!
1"
0'
1(
0/
10
#467970000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#467980000000
0!
1$
0'
1+
0/
#467990000000
1!
1'
1/
#468000000000
0!
0'
0/
#468010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#468020000000
0!
0'
0/
#468030000000
1!
1'
1/
#468040000000
0!
0'
0/
#468050000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#468060000000
0!
0'
0/
#468070000000
1!
1'
1/
#468080000000
0!
0'
0/
#468090000000
1!
1'
1/
#468100000000
0!
0'
0/
#468110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#468120000000
0!
0'
0/
#468130000000
1!
1'
1/
#468140000000
0!
0'
0/
#468150000000
1!
1'
1/
#468160000000
0!
0'
0/
#468170000000
1!
1'
1/
#468180000000
0!
0'
0/
#468190000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#468200000000
0!
0'
0/
#468210000000
1!
1'
1/
#468220000000
0!
0'
0/
#468230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#468240000000
0!
0'
0/
#468250000000
1!
1'
1/
#468260000000
0!
0'
0/
#468270000000
#468280000000
1!
1'
1/
#468290000000
0!
0'
0/
#468300000000
1!
1'
1/
#468310000000
0!
1"
0'
1(
0/
10
#468320000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#468330000000
0!
0'
0/
#468340000000
1!
1'
1/
#468350000000
0!
0'
0/
#468360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#468370000000
0!
0'
0/
#468380000000
1!
1'
1/
#468390000000
0!
1"
0'
1(
0/
10
#468400000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#468410000000
0!
1$
0'
1+
0/
#468420000000
1!
1'
1/
#468430000000
0!
0'
0/
#468440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#468450000000
0!
0'
0/
#468460000000
1!
1'
1/
#468470000000
0!
0'
0/
#468480000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#468490000000
0!
0'
0/
#468500000000
1!
1'
1/
#468510000000
0!
0'
0/
#468520000000
1!
1'
1/
#468530000000
0!
0'
0/
#468540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#468550000000
0!
0'
0/
#468560000000
1!
1'
1/
#468570000000
0!
0'
0/
#468580000000
1!
1'
1/
#468590000000
0!
0'
0/
#468600000000
1!
1'
1/
#468610000000
0!
0'
0/
#468620000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#468630000000
0!
0'
0/
#468640000000
1!
1'
1/
#468650000000
0!
0'
0/
#468660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#468670000000
0!
0'
0/
#468680000000
1!
1'
1/
#468690000000
0!
0'
0/
#468700000000
#468710000000
1!
1'
1/
#468720000000
0!
0'
0/
#468730000000
1!
1'
1/
#468740000000
0!
1"
0'
1(
0/
10
#468750000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#468760000000
0!
0'
0/
#468770000000
1!
1'
1/
#468780000000
0!
0'
0/
#468790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#468800000000
0!
0'
0/
#468810000000
1!
1'
1/
#468820000000
0!
1"
0'
1(
0/
10
#468830000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#468840000000
0!
1$
0'
1+
0/
#468850000000
1!
1'
1/
#468860000000
0!
0'
0/
#468870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#468880000000
0!
0'
0/
#468890000000
1!
1'
1/
#468900000000
0!
0'
0/
#468910000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#468920000000
0!
0'
0/
#468930000000
1!
1'
1/
#468940000000
0!
0'
0/
#468950000000
1!
1'
1/
#468960000000
0!
0'
0/
#468970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#468980000000
0!
0'
0/
#468990000000
1!
1'
1/
#469000000000
0!
0'
0/
#469010000000
1!
1'
1/
#469020000000
0!
0'
0/
#469030000000
1!
1'
1/
#469040000000
0!
0'
0/
#469050000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#469060000000
0!
0'
0/
#469070000000
1!
1'
1/
#469080000000
0!
0'
0/
#469090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#469100000000
0!
0'
0/
#469110000000
1!
1'
1/
#469120000000
0!
0'
0/
#469130000000
#469140000000
1!
1'
1/
#469150000000
0!
0'
0/
#469160000000
1!
1'
1/
#469170000000
0!
1"
0'
1(
0/
10
#469180000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#469190000000
0!
0'
0/
#469200000000
1!
1'
1/
#469210000000
0!
0'
0/
#469220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#469230000000
0!
0'
0/
#469240000000
1!
1'
1/
#469250000000
0!
1"
0'
1(
0/
10
#469260000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#469270000000
0!
1$
0'
1+
0/
#469280000000
1!
1'
1/
#469290000000
0!
0'
0/
#469300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#469310000000
0!
0'
0/
#469320000000
1!
1'
1/
#469330000000
0!
0'
0/
#469340000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#469350000000
0!
0'
0/
#469360000000
1!
1'
1/
#469370000000
0!
0'
0/
#469380000000
1!
1'
1/
#469390000000
0!
0'
0/
#469400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#469410000000
0!
0'
0/
#469420000000
1!
1'
1/
#469430000000
0!
0'
0/
#469440000000
1!
1'
1/
#469450000000
0!
0'
0/
#469460000000
1!
1'
1/
#469470000000
0!
0'
0/
#469480000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#469490000000
0!
0'
0/
#469500000000
1!
1'
1/
#469510000000
0!
0'
0/
#469520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#469530000000
0!
0'
0/
#469540000000
1!
1'
1/
#469550000000
0!
0'
0/
#469560000000
#469570000000
1!
1'
1/
#469580000000
0!
0'
0/
#469590000000
1!
1'
1/
#469600000000
0!
1"
0'
1(
0/
10
#469610000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#469620000000
0!
0'
0/
#469630000000
1!
1'
1/
#469640000000
0!
0'
0/
#469650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#469660000000
0!
0'
0/
#469670000000
1!
1'
1/
#469680000000
0!
1"
0'
1(
0/
10
#469690000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#469700000000
0!
1$
0'
1+
0/
#469710000000
1!
1'
1/
#469720000000
0!
0'
0/
#469730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#469740000000
0!
0'
0/
#469750000000
1!
1'
1/
#469760000000
0!
0'
0/
#469770000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#469780000000
0!
0'
0/
#469790000000
1!
1'
1/
#469800000000
0!
0'
0/
#469810000000
1!
1'
1/
#469820000000
0!
0'
0/
#469830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#469840000000
0!
0'
0/
#469850000000
1!
1'
1/
#469860000000
0!
0'
0/
#469870000000
1!
1'
1/
#469880000000
0!
0'
0/
#469890000000
1!
1'
1/
#469900000000
0!
0'
0/
#469910000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#469920000000
0!
0'
0/
#469930000000
1!
1'
1/
#469940000000
0!
0'
0/
#469950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#469960000000
0!
0'
0/
#469970000000
1!
1'
1/
#469980000000
0!
0'
0/
#469990000000
#470000000000
1!
1'
1/
#470010000000
0!
0'
0/
#470020000000
1!
1'
1/
#470030000000
0!
1"
0'
1(
0/
10
#470040000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#470050000000
0!
0'
0/
#470060000000
1!
1'
1/
#470070000000
0!
0'
0/
#470080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#470090000000
0!
0'
0/
#470100000000
1!
1'
1/
#470110000000
0!
1"
0'
1(
0/
10
#470120000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#470130000000
0!
1$
0'
1+
0/
#470140000000
1!
1'
1/
#470150000000
0!
0'
0/
#470160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#470170000000
0!
0'
0/
#470180000000
1!
1'
1/
#470190000000
0!
0'
0/
#470200000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#470210000000
0!
0'
0/
#470220000000
1!
1'
1/
#470230000000
0!
0'
0/
#470240000000
1!
1'
1/
#470250000000
0!
0'
0/
#470260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#470270000000
0!
0'
0/
#470280000000
1!
1'
1/
#470290000000
0!
0'
0/
#470300000000
1!
1'
1/
#470310000000
0!
0'
0/
#470320000000
1!
1'
1/
#470330000000
0!
0'
0/
#470340000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#470350000000
0!
0'
0/
#470360000000
1!
1'
1/
#470370000000
0!
0'
0/
#470380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#470390000000
0!
0'
0/
#470400000000
1!
1'
1/
#470410000000
0!
0'
0/
#470420000000
#470430000000
1!
1'
1/
#470440000000
0!
0'
0/
#470450000000
1!
1'
1/
#470460000000
0!
1"
0'
1(
0/
10
#470470000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#470480000000
0!
0'
0/
#470490000000
1!
1'
1/
#470500000000
0!
0'
0/
#470510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#470520000000
0!
0'
0/
#470530000000
1!
1'
1/
#470540000000
0!
1"
0'
1(
0/
10
#470550000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#470560000000
0!
1$
0'
1+
0/
#470570000000
1!
1'
1/
#470580000000
0!
0'
0/
#470590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#470600000000
0!
0'
0/
#470610000000
1!
1'
1/
#470620000000
0!
0'
0/
#470630000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#470640000000
0!
0'
0/
#470650000000
1!
1'
1/
#470660000000
0!
0'
0/
#470670000000
1!
1'
1/
#470680000000
0!
0'
0/
#470690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#470700000000
0!
0'
0/
#470710000000
1!
1'
1/
#470720000000
0!
0'
0/
#470730000000
1!
1'
1/
#470740000000
0!
0'
0/
#470750000000
1!
1'
1/
#470760000000
0!
0'
0/
#470770000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#470780000000
0!
0'
0/
#470790000000
1!
1'
1/
#470800000000
0!
0'
0/
#470810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#470820000000
0!
0'
0/
#470830000000
1!
1'
1/
#470840000000
0!
0'
0/
#470850000000
#470860000000
1!
1'
1/
#470870000000
0!
0'
0/
#470880000000
1!
1'
1/
#470890000000
0!
1"
0'
1(
0/
10
#470900000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#470910000000
0!
0'
0/
#470920000000
1!
1'
1/
#470930000000
0!
0'
0/
#470940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#470950000000
0!
0'
0/
#470960000000
1!
1'
1/
#470970000000
0!
1"
0'
1(
0/
10
#470980000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#470990000000
0!
1$
0'
1+
0/
#471000000000
1!
1'
1/
#471010000000
0!
0'
0/
#471020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#471030000000
0!
0'
0/
#471040000000
1!
1'
1/
#471050000000
0!
0'
0/
#471060000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#471070000000
0!
0'
0/
#471080000000
1!
1'
1/
#471090000000
0!
0'
0/
#471100000000
1!
1'
1/
#471110000000
0!
0'
0/
#471120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#471130000000
0!
0'
0/
#471140000000
1!
1'
1/
#471150000000
0!
0'
0/
#471160000000
1!
1'
1/
#471170000000
0!
0'
0/
#471180000000
1!
1'
1/
#471190000000
0!
0'
0/
#471200000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#471210000000
0!
0'
0/
#471220000000
1!
1'
1/
#471230000000
0!
0'
0/
#471240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#471250000000
0!
0'
0/
#471260000000
1!
1'
1/
#471270000000
0!
0'
0/
#471280000000
#471290000000
1!
1'
1/
#471300000000
0!
0'
0/
#471310000000
1!
1'
1/
#471320000000
0!
1"
0'
1(
0/
10
#471330000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#471340000000
0!
0'
0/
#471350000000
1!
1'
1/
#471360000000
0!
0'
0/
#471370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#471380000000
0!
0'
0/
#471390000000
1!
1'
1/
#471400000000
0!
1"
0'
1(
0/
10
#471410000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#471420000000
0!
1$
0'
1+
0/
#471430000000
1!
1'
1/
#471440000000
0!
0'
0/
#471450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#471460000000
0!
0'
0/
#471470000000
1!
1'
1/
#471480000000
0!
0'
0/
#471490000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#471500000000
0!
0'
0/
#471510000000
1!
1'
1/
#471520000000
0!
0'
0/
#471530000000
1!
1'
1/
#471540000000
0!
0'
0/
#471550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#471560000000
0!
0'
0/
#471570000000
1!
1'
1/
#471580000000
0!
0'
0/
#471590000000
1!
1'
1/
#471600000000
0!
0'
0/
#471610000000
1!
1'
1/
#471620000000
0!
0'
0/
#471630000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#471640000000
0!
0'
0/
#471650000000
1!
1'
1/
#471660000000
0!
0'
0/
#471670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#471680000000
0!
0'
0/
#471690000000
1!
1'
1/
#471700000000
0!
0'
0/
#471710000000
#471720000000
1!
1'
1/
#471730000000
0!
0'
0/
#471740000000
1!
1'
1/
#471750000000
0!
1"
0'
1(
0/
10
#471760000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#471770000000
0!
0'
0/
#471780000000
1!
1'
1/
#471790000000
0!
0'
0/
#471800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#471810000000
0!
0'
0/
#471820000000
1!
1'
1/
#471830000000
0!
1"
0'
1(
0/
10
#471840000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#471850000000
0!
1$
0'
1+
0/
#471860000000
1!
1'
1/
#471870000000
0!
0'
0/
#471880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#471890000000
0!
0'
0/
#471900000000
1!
1'
1/
#471910000000
0!
0'
0/
#471920000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#471930000000
0!
0'
0/
#471940000000
1!
1'
1/
#471950000000
0!
0'
0/
#471960000000
1!
1'
1/
#471970000000
0!
0'
0/
#471980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#471990000000
0!
0'
0/
#472000000000
1!
1'
1/
#472010000000
0!
0'
0/
#472020000000
1!
1'
1/
#472030000000
0!
0'
0/
#472040000000
1!
1'
1/
#472050000000
0!
0'
0/
#472060000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#472070000000
0!
0'
0/
#472080000000
1!
1'
1/
#472090000000
0!
0'
0/
#472100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#472110000000
0!
0'
0/
#472120000000
1!
1'
1/
#472130000000
0!
0'
0/
#472140000000
#472150000000
1!
1'
1/
#472160000000
0!
0'
0/
#472170000000
1!
1'
1/
#472180000000
0!
1"
0'
1(
0/
10
#472190000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#472200000000
0!
0'
0/
#472210000000
1!
1'
1/
#472220000000
0!
0'
0/
#472230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#472240000000
0!
0'
0/
#472250000000
1!
1'
1/
#472260000000
0!
1"
0'
1(
0/
10
#472270000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#472280000000
0!
1$
0'
1+
0/
#472290000000
1!
1'
1/
#472300000000
0!
0'
0/
#472310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#472320000000
0!
0'
0/
#472330000000
1!
1'
1/
#472340000000
0!
0'
0/
#472350000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#472360000000
0!
0'
0/
#472370000000
1!
1'
1/
#472380000000
0!
0'
0/
#472390000000
1!
1'
1/
#472400000000
0!
0'
0/
#472410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#472420000000
0!
0'
0/
#472430000000
1!
1'
1/
#472440000000
0!
0'
0/
#472450000000
1!
1'
1/
#472460000000
0!
0'
0/
#472470000000
1!
1'
1/
#472480000000
0!
0'
0/
#472490000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#472500000000
0!
0'
0/
#472510000000
1!
1'
1/
#472520000000
0!
0'
0/
#472530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#472540000000
0!
0'
0/
#472550000000
1!
1'
1/
#472560000000
0!
0'
0/
#472570000000
#472580000000
1!
1'
1/
#472590000000
0!
0'
0/
#472600000000
1!
1'
1/
#472610000000
0!
1"
0'
1(
0/
10
#472620000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#472630000000
0!
0'
0/
#472640000000
1!
1'
1/
#472650000000
0!
0'
0/
#472660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#472670000000
0!
0'
0/
#472680000000
1!
1'
1/
#472690000000
0!
1"
0'
1(
0/
10
#472700000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#472710000000
0!
1$
0'
1+
0/
#472720000000
1!
1'
1/
#472730000000
0!
0'
0/
#472740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#472750000000
0!
0'
0/
#472760000000
1!
1'
1/
#472770000000
0!
0'
0/
#472780000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#472790000000
0!
0'
0/
#472800000000
1!
1'
1/
#472810000000
0!
0'
0/
#472820000000
1!
1'
1/
#472830000000
0!
0'
0/
#472840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#472850000000
0!
0'
0/
#472860000000
1!
1'
1/
#472870000000
0!
0'
0/
#472880000000
1!
1'
1/
#472890000000
0!
0'
0/
#472900000000
1!
1'
1/
#472910000000
0!
0'
0/
#472920000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#472930000000
0!
0'
0/
#472940000000
1!
1'
1/
#472950000000
0!
0'
0/
#472960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#472970000000
0!
0'
0/
#472980000000
1!
1'
1/
#472990000000
0!
0'
0/
#473000000000
#473010000000
1!
1'
1/
#473020000000
0!
0'
0/
#473030000000
1!
1'
1/
#473040000000
0!
1"
0'
1(
0/
10
#473050000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#473060000000
0!
0'
0/
#473070000000
1!
1'
1/
#473080000000
0!
0'
0/
#473090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#473100000000
0!
0'
0/
#473110000000
1!
1'
1/
#473120000000
0!
1"
0'
1(
0/
10
#473130000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#473140000000
0!
1$
0'
1+
0/
#473150000000
1!
1'
1/
#473160000000
0!
0'
0/
#473170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#473180000000
0!
0'
0/
#473190000000
1!
1'
1/
#473200000000
0!
0'
0/
#473210000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#473220000000
0!
0'
0/
#473230000000
1!
1'
1/
#473240000000
0!
0'
0/
#473250000000
1!
1'
1/
#473260000000
0!
0'
0/
#473270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#473280000000
0!
0'
0/
#473290000000
1!
1'
1/
#473300000000
0!
0'
0/
#473310000000
1!
1'
1/
#473320000000
0!
0'
0/
#473330000000
1!
1'
1/
#473340000000
0!
0'
0/
#473350000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#473360000000
0!
0'
0/
#473370000000
1!
1'
1/
#473380000000
0!
0'
0/
#473390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#473400000000
0!
0'
0/
#473410000000
1!
1'
1/
#473420000000
0!
0'
0/
#473430000000
#473440000000
1!
1'
1/
#473450000000
0!
0'
0/
#473460000000
1!
1'
1/
#473470000000
0!
1"
0'
1(
0/
10
#473480000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#473490000000
0!
0'
0/
#473500000000
1!
1'
1/
#473510000000
0!
0'
0/
#473520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#473530000000
0!
0'
0/
#473540000000
1!
1'
1/
#473550000000
0!
1"
0'
1(
0/
10
#473560000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#473570000000
0!
1$
0'
1+
0/
#473580000000
1!
1'
1/
#473590000000
0!
0'
0/
#473600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#473610000000
0!
0'
0/
#473620000000
1!
1'
1/
#473630000000
0!
0'
0/
#473640000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#473650000000
0!
0'
0/
#473660000000
1!
1'
1/
#473670000000
0!
0'
0/
#473680000000
1!
1'
1/
#473690000000
0!
0'
0/
#473700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#473710000000
0!
0'
0/
#473720000000
1!
1'
1/
#473730000000
0!
0'
0/
#473740000000
1!
1'
1/
#473750000000
0!
0'
0/
#473760000000
1!
1'
1/
#473770000000
0!
0'
0/
#473780000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#473790000000
0!
0'
0/
#473800000000
1!
1'
1/
#473810000000
0!
0'
0/
#473820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#473830000000
0!
0'
0/
#473840000000
1!
1'
1/
#473850000000
0!
0'
0/
#473860000000
#473870000000
1!
1'
1/
#473880000000
0!
0'
0/
#473890000000
1!
1'
1/
#473900000000
0!
1"
0'
1(
0/
10
#473910000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#473920000000
0!
0'
0/
#473930000000
1!
1'
1/
#473940000000
0!
0'
0/
#473950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#473960000000
0!
0'
0/
#473970000000
1!
1'
1/
#473980000000
0!
1"
0'
1(
0/
10
#473990000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#474000000000
0!
1$
0'
1+
0/
#474010000000
1!
1'
1/
#474020000000
0!
0'
0/
#474030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#474040000000
0!
0'
0/
#474050000000
1!
1'
1/
#474060000000
0!
0'
0/
#474070000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#474080000000
0!
0'
0/
#474090000000
1!
1'
1/
#474100000000
0!
0'
0/
#474110000000
1!
1'
1/
#474120000000
0!
0'
0/
#474130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#474140000000
0!
0'
0/
#474150000000
1!
1'
1/
#474160000000
0!
0'
0/
#474170000000
1!
1'
1/
#474180000000
0!
0'
0/
#474190000000
1!
1'
1/
#474200000000
0!
0'
0/
#474210000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#474220000000
0!
0'
0/
#474230000000
1!
1'
1/
#474240000000
0!
0'
0/
#474250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#474260000000
0!
0'
0/
#474270000000
1!
1'
1/
#474280000000
0!
0'
0/
#474290000000
#474300000000
1!
1'
1/
#474310000000
0!
0'
0/
#474320000000
1!
1'
1/
#474330000000
0!
1"
0'
1(
0/
10
#474340000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#474350000000
0!
0'
0/
#474360000000
1!
1'
1/
#474370000000
0!
0'
0/
#474380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#474390000000
0!
0'
0/
#474400000000
1!
1'
1/
#474410000000
0!
1"
0'
1(
0/
10
#474420000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#474430000000
0!
1$
0'
1+
0/
#474440000000
1!
1'
1/
#474450000000
0!
0'
0/
#474460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#474470000000
0!
0'
0/
#474480000000
1!
1'
1/
#474490000000
0!
0'
0/
#474500000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#474510000000
0!
0'
0/
#474520000000
1!
1'
1/
#474530000000
0!
0'
0/
#474540000000
1!
1'
1/
#474550000000
0!
0'
0/
#474560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#474570000000
0!
0'
0/
#474580000000
1!
1'
1/
#474590000000
0!
0'
0/
#474600000000
1!
1'
1/
#474610000000
0!
0'
0/
#474620000000
1!
1'
1/
#474630000000
0!
0'
0/
#474640000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#474650000000
0!
0'
0/
#474660000000
1!
1'
1/
#474670000000
0!
0'
0/
#474680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#474690000000
0!
0'
0/
#474700000000
1!
1'
1/
#474710000000
0!
0'
0/
#474720000000
#474730000000
1!
1'
1/
#474740000000
0!
0'
0/
#474750000000
1!
1'
1/
#474760000000
0!
1"
0'
1(
0/
10
#474770000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#474780000000
0!
0'
0/
#474790000000
1!
1'
1/
#474800000000
0!
0'
0/
#474810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#474820000000
0!
0'
0/
#474830000000
1!
1'
1/
#474840000000
0!
1"
0'
1(
0/
10
#474850000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#474860000000
0!
1$
0'
1+
0/
#474870000000
1!
1'
1/
#474880000000
0!
0'
0/
#474890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#474900000000
0!
0'
0/
#474910000000
1!
1'
1/
#474920000000
0!
0'
0/
#474930000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#474940000000
0!
0'
0/
#474950000000
1!
1'
1/
#474960000000
0!
0'
0/
#474970000000
1!
1'
1/
#474980000000
0!
0'
0/
#474990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#475000000000
0!
0'
0/
#475010000000
1!
1'
1/
#475020000000
0!
0'
0/
#475030000000
1!
1'
1/
#475040000000
0!
0'
0/
#475050000000
1!
1'
1/
#475060000000
0!
0'
0/
#475070000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#475080000000
0!
0'
0/
#475090000000
1!
1'
1/
#475100000000
0!
0'
0/
#475110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#475120000000
0!
0'
0/
#475130000000
1!
1'
1/
#475140000000
0!
0'
0/
#475150000000
#475160000000
1!
1'
1/
#475170000000
0!
0'
0/
#475180000000
1!
1'
1/
#475190000000
0!
1"
0'
1(
0/
10
#475200000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#475210000000
0!
0'
0/
#475220000000
1!
1'
1/
#475230000000
0!
0'
0/
#475240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#475250000000
0!
0'
0/
#475260000000
1!
1'
1/
#475270000000
0!
1"
0'
1(
0/
10
#475280000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#475290000000
0!
1$
0'
1+
0/
#475300000000
1!
1'
1/
#475310000000
0!
0'
0/
#475320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#475330000000
0!
0'
0/
#475340000000
1!
1'
1/
#475350000000
0!
0'
0/
#475360000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#475370000000
0!
0'
0/
#475380000000
1!
1'
1/
#475390000000
0!
0'
0/
#475400000000
1!
1'
1/
#475410000000
0!
0'
0/
#475420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#475430000000
0!
0'
0/
#475440000000
1!
1'
1/
#475450000000
0!
0'
0/
#475460000000
1!
1'
1/
#475470000000
0!
0'
0/
#475480000000
1!
1'
1/
#475490000000
0!
0'
0/
#475500000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#475510000000
0!
0'
0/
#475520000000
1!
1'
1/
#475530000000
0!
0'
0/
#475540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#475550000000
0!
0'
0/
#475560000000
1!
1'
1/
#475570000000
0!
0'
0/
#475580000000
#475590000000
1!
1'
1/
#475600000000
0!
0'
0/
#475610000000
1!
1'
1/
#475620000000
0!
1"
0'
1(
0/
10
#475630000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#475640000000
0!
0'
0/
#475650000000
1!
1'
1/
#475660000000
0!
0'
0/
#475670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#475680000000
0!
0'
0/
#475690000000
1!
1'
1/
#475700000000
0!
1"
0'
1(
0/
10
#475710000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#475720000000
0!
1$
0'
1+
0/
#475730000000
1!
1'
1/
#475740000000
0!
0'
0/
#475750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#475760000000
0!
0'
0/
#475770000000
1!
1'
1/
#475780000000
0!
0'
0/
#475790000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#475800000000
0!
0'
0/
#475810000000
1!
1'
1/
#475820000000
0!
0'
0/
#475830000000
1!
1'
1/
#475840000000
0!
0'
0/
#475850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#475860000000
0!
0'
0/
#475870000000
1!
1'
1/
#475880000000
0!
0'
0/
#475890000000
1!
1'
1/
#475900000000
0!
0'
0/
#475910000000
1!
1'
1/
#475920000000
0!
0'
0/
#475930000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#475940000000
0!
0'
0/
#475950000000
1!
1'
1/
#475960000000
0!
0'
0/
#475970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#475980000000
0!
0'
0/
#475990000000
1!
1'
1/
#476000000000
0!
0'
0/
#476010000000
#476020000000
1!
1'
1/
#476030000000
0!
0'
0/
#476040000000
1!
1'
1/
#476050000000
0!
1"
0'
1(
0/
10
#476060000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#476070000000
0!
0'
0/
#476080000000
1!
1'
1/
#476090000000
0!
0'
0/
#476100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#476110000000
0!
0'
0/
#476120000000
1!
1'
1/
#476130000000
0!
1"
0'
1(
0/
10
#476140000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#476150000000
0!
1$
0'
1+
0/
#476160000000
1!
1'
1/
#476170000000
0!
0'
0/
#476180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#476190000000
0!
0'
0/
#476200000000
1!
1'
1/
#476210000000
0!
0'
0/
#476220000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#476230000000
0!
0'
0/
#476240000000
1!
1'
1/
#476250000000
0!
0'
0/
#476260000000
1!
1'
1/
#476270000000
0!
0'
0/
#476280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#476290000000
0!
0'
0/
#476300000000
1!
1'
1/
#476310000000
0!
0'
0/
#476320000000
1!
1'
1/
#476330000000
0!
0'
0/
#476340000000
1!
1'
1/
#476350000000
0!
0'
0/
#476360000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#476370000000
0!
0'
0/
#476380000000
1!
1'
1/
#476390000000
0!
0'
0/
#476400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#476410000000
0!
0'
0/
#476420000000
1!
1'
1/
#476430000000
0!
0'
0/
#476440000000
#476450000000
1!
1'
1/
#476460000000
0!
0'
0/
#476470000000
1!
1'
1/
#476480000000
0!
1"
0'
1(
0/
10
#476490000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#476500000000
0!
0'
0/
#476510000000
1!
1'
1/
#476520000000
0!
0'
0/
#476530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#476540000000
0!
0'
0/
#476550000000
1!
1'
1/
#476560000000
0!
1"
0'
1(
0/
10
#476570000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#476580000000
0!
1$
0'
1+
0/
#476590000000
1!
1'
1/
#476600000000
0!
0'
0/
#476610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#476620000000
0!
0'
0/
#476630000000
1!
1'
1/
#476640000000
0!
0'
0/
#476650000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#476660000000
0!
0'
0/
#476670000000
1!
1'
1/
#476680000000
0!
0'
0/
#476690000000
1!
1'
1/
#476700000000
0!
0'
0/
#476710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#476720000000
0!
0'
0/
#476730000000
1!
1'
1/
#476740000000
0!
0'
0/
#476750000000
1!
1'
1/
#476760000000
0!
0'
0/
#476770000000
1!
1'
1/
#476780000000
0!
0'
0/
#476790000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#476800000000
0!
0'
0/
#476810000000
1!
1'
1/
#476820000000
0!
0'
0/
#476830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#476840000000
0!
0'
0/
#476850000000
1!
1'
1/
#476860000000
0!
0'
0/
#476870000000
#476880000000
1!
1'
1/
#476890000000
0!
0'
0/
#476900000000
1!
1'
1/
#476910000000
0!
1"
0'
1(
0/
10
#476920000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#476930000000
0!
0'
0/
#476940000000
1!
1'
1/
#476950000000
0!
0'
0/
#476960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#476970000000
0!
0'
0/
#476980000000
1!
1'
1/
#476990000000
0!
1"
0'
1(
0/
10
#477000000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#477010000000
0!
1$
0'
1+
0/
#477020000000
1!
1'
1/
#477030000000
0!
0'
0/
#477040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#477050000000
0!
0'
0/
#477060000000
1!
1'
1/
#477070000000
0!
0'
0/
#477080000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#477090000000
0!
0'
0/
#477100000000
1!
1'
1/
#477110000000
0!
0'
0/
#477120000000
1!
1'
1/
#477130000000
0!
0'
0/
#477140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#477150000000
0!
0'
0/
#477160000000
1!
1'
1/
#477170000000
0!
0'
0/
#477180000000
1!
1'
1/
#477190000000
0!
0'
0/
#477200000000
1!
1'
1/
#477210000000
0!
0'
0/
#477220000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#477230000000
0!
0'
0/
#477240000000
1!
1'
1/
#477250000000
0!
0'
0/
#477260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#477270000000
0!
0'
0/
#477280000000
1!
1'
1/
#477290000000
0!
0'
0/
#477300000000
#477310000000
1!
1'
1/
#477320000000
0!
0'
0/
#477330000000
1!
1'
1/
#477340000000
0!
1"
0'
1(
0/
10
#477350000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#477360000000
0!
0'
0/
#477370000000
1!
1'
1/
#477380000000
0!
0'
0/
#477390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#477400000000
0!
0'
0/
#477410000000
1!
1'
1/
#477420000000
0!
1"
0'
1(
0/
10
#477430000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#477440000000
0!
1$
0'
1+
0/
#477450000000
1!
1'
1/
#477460000000
0!
0'
0/
#477470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#477480000000
0!
0'
0/
#477490000000
1!
1'
1/
#477500000000
0!
0'
0/
#477510000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#477520000000
0!
0'
0/
#477530000000
1!
1'
1/
#477540000000
0!
0'
0/
#477550000000
1!
1'
1/
#477560000000
0!
0'
0/
#477570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#477580000000
0!
0'
0/
#477590000000
1!
1'
1/
#477600000000
0!
0'
0/
#477610000000
1!
1'
1/
#477620000000
0!
0'
0/
#477630000000
1!
1'
1/
#477640000000
0!
0'
0/
#477650000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#477660000000
0!
0'
0/
#477670000000
1!
1'
1/
#477680000000
0!
0'
0/
#477690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#477700000000
0!
0'
0/
#477710000000
1!
1'
1/
#477720000000
0!
0'
0/
#477730000000
#477740000000
1!
1'
1/
#477750000000
0!
0'
0/
#477760000000
1!
1'
1/
#477770000000
0!
1"
0'
1(
0/
10
#477780000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#477790000000
0!
0'
0/
#477800000000
1!
1'
1/
#477810000000
0!
0'
0/
#477820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#477830000000
0!
0'
0/
#477840000000
1!
1'
1/
#477850000000
0!
1"
0'
1(
0/
10
#477860000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#477870000000
0!
1$
0'
1+
0/
#477880000000
1!
1'
1/
#477890000000
0!
0'
0/
#477900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#477910000000
0!
0'
0/
#477920000000
1!
1'
1/
#477930000000
0!
0'
0/
#477940000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#477950000000
0!
0'
0/
#477960000000
1!
1'
1/
#477970000000
0!
0'
0/
#477980000000
1!
1'
1/
#477990000000
0!
0'
0/
#478000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#478010000000
0!
0'
0/
#478020000000
1!
1'
1/
#478030000000
0!
0'
0/
#478040000000
1!
1'
1/
#478050000000
0!
0'
0/
#478060000000
1!
1'
1/
#478070000000
0!
0'
0/
#478080000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#478090000000
0!
0'
0/
#478100000000
1!
1'
1/
#478110000000
0!
0'
0/
#478120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#478130000000
0!
0'
0/
#478140000000
1!
1'
1/
#478150000000
0!
0'
0/
#478160000000
#478170000000
1!
1'
1/
#478180000000
0!
0'
0/
#478190000000
1!
1'
1/
#478200000000
0!
1"
0'
1(
0/
10
#478210000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#478220000000
0!
0'
0/
#478230000000
1!
1'
1/
#478240000000
0!
0'
0/
#478250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#478260000000
0!
0'
0/
#478270000000
1!
1'
1/
#478280000000
0!
1"
0'
1(
0/
10
#478290000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#478300000000
0!
1$
0'
1+
0/
#478310000000
1!
1'
1/
#478320000000
0!
0'
0/
#478330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#478340000000
0!
0'
0/
#478350000000
1!
1'
1/
#478360000000
0!
0'
0/
#478370000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#478380000000
0!
0'
0/
#478390000000
1!
1'
1/
#478400000000
0!
0'
0/
#478410000000
1!
1'
1/
#478420000000
0!
0'
0/
#478430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#478440000000
0!
0'
0/
#478450000000
1!
1'
1/
#478460000000
0!
0'
0/
#478470000000
1!
1'
1/
#478480000000
0!
0'
0/
#478490000000
1!
1'
1/
#478500000000
0!
0'
0/
#478510000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#478520000000
0!
0'
0/
#478530000000
1!
1'
1/
#478540000000
0!
0'
0/
#478550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#478560000000
0!
0'
0/
#478570000000
1!
1'
1/
#478580000000
0!
0'
0/
#478590000000
#478600000000
1!
1'
1/
#478610000000
0!
0'
0/
#478620000000
1!
1'
1/
#478630000000
0!
1"
0'
1(
0/
10
#478640000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#478650000000
0!
0'
0/
#478660000000
1!
1'
1/
#478670000000
0!
0'
0/
#478680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#478690000000
0!
0'
0/
#478700000000
1!
1'
1/
#478710000000
0!
1"
0'
1(
0/
10
#478720000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#478730000000
0!
1$
0'
1+
0/
#478740000000
1!
1'
1/
#478750000000
0!
0'
0/
#478760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#478770000000
0!
0'
0/
#478780000000
1!
1'
1/
#478790000000
0!
0'
0/
#478800000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#478810000000
0!
0'
0/
#478820000000
1!
1'
1/
#478830000000
0!
0'
0/
#478840000000
1!
1'
1/
#478850000000
0!
0'
0/
#478860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#478870000000
0!
0'
0/
#478880000000
1!
1'
1/
#478890000000
0!
0'
0/
#478900000000
1!
1'
1/
#478910000000
0!
0'
0/
#478920000000
1!
1'
1/
#478930000000
0!
0'
0/
#478940000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#478950000000
0!
0'
0/
#478960000000
1!
1'
1/
#478970000000
0!
0'
0/
#478980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#478990000000
0!
0'
0/
#479000000000
1!
1'
1/
#479010000000
0!
0'
0/
#479020000000
#479030000000
1!
1'
1/
#479040000000
0!
0'
0/
#479050000000
1!
1'
1/
#479060000000
0!
1"
0'
1(
0/
10
#479070000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#479080000000
0!
0'
0/
#479090000000
1!
1'
1/
#479100000000
0!
0'
0/
#479110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#479120000000
0!
0'
0/
#479130000000
1!
1'
1/
#479140000000
0!
1"
0'
1(
0/
10
#479150000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#479160000000
0!
1$
0'
1+
0/
#479170000000
1!
1'
1/
#479180000000
0!
0'
0/
#479190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#479200000000
0!
0'
0/
#479210000000
1!
1'
1/
#479220000000
0!
0'
0/
#479230000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#479240000000
0!
0'
0/
#479250000000
1!
1'
1/
#479260000000
0!
0'
0/
#479270000000
1!
1'
1/
#479280000000
0!
0'
0/
#479290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#479300000000
0!
0'
0/
#479310000000
1!
1'
1/
#479320000000
0!
0'
0/
#479330000000
1!
1'
1/
#479340000000
0!
0'
0/
#479350000000
1!
1'
1/
#479360000000
0!
0'
0/
#479370000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#479380000000
0!
0'
0/
#479390000000
1!
1'
1/
#479400000000
0!
0'
0/
#479410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#479420000000
0!
0'
0/
#479430000000
1!
1'
1/
#479440000000
0!
0'
0/
#479450000000
#479460000000
1!
1'
1/
#479470000000
0!
0'
0/
#479480000000
1!
1'
1/
#479490000000
0!
1"
0'
1(
0/
10
#479500000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#479510000000
0!
0'
0/
#479520000000
1!
1'
1/
#479530000000
0!
0'
0/
#479540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#479550000000
0!
0'
0/
#479560000000
1!
1'
1/
#479570000000
0!
1"
0'
1(
0/
10
#479580000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#479590000000
0!
1$
0'
1+
0/
#479600000000
1!
1'
1/
#479610000000
0!
0'
0/
#479620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#479630000000
0!
0'
0/
#479640000000
1!
1'
1/
#479650000000
0!
0'
0/
#479660000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#479670000000
0!
0'
0/
#479680000000
1!
1'
1/
#479690000000
0!
0'
0/
#479700000000
1!
1'
1/
#479710000000
0!
0'
0/
#479720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#479730000000
0!
0'
0/
#479740000000
1!
1'
1/
#479750000000
0!
0'
0/
#479760000000
1!
1'
1/
#479770000000
0!
0'
0/
#479780000000
1!
1'
1/
#479790000000
0!
0'
0/
#479800000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#479810000000
0!
0'
0/
#479820000000
1!
1'
1/
#479830000000
0!
0'
0/
#479840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#479850000000
0!
0'
0/
#479860000000
1!
1'
1/
#479870000000
0!
0'
0/
#479880000000
#479890000000
1!
1'
1/
#479900000000
0!
0'
0/
#479910000000
1!
1'
1/
#479920000000
0!
1"
0'
1(
0/
10
#479930000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#479940000000
0!
0'
0/
#479950000000
1!
1'
1/
#479960000000
0!
0'
0/
#479970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#479980000000
0!
0'
0/
#479990000000
1!
1'
1/
#480000000000
0!
1"
0'
1(
0/
10
#480010000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#480020000000
0!
1$
0'
1+
0/
#480030000000
1!
1'
1/
#480040000000
0!
0'
0/
#480050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#480060000000
0!
0'
0/
#480070000000
1!
1'
1/
#480080000000
0!
0'
0/
#480090000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#480100000000
0!
0'
0/
#480110000000
1!
1'
1/
#480120000000
0!
0'
0/
#480130000000
1!
1'
1/
#480140000000
0!
0'
0/
#480150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#480160000000
0!
0'
0/
#480170000000
1!
1'
1/
#480180000000
0!
0'
0/
#480190000000
1!
1'
1/
#480200000000
0!
0'
0/
#480210000000
1!
1'
1/
#480220000000
0!
0'
0/
#480230000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#480240000000
0!
0'
0/
#480250000000
1!
1'
1/
#480260000000
0!
0'
0/
#480270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#480280000000
0!
0'
0/
#480290000000
1!
1'
1/
#480300000000
0!
0'
0/
#480310000000
#480320000000
1!
1'
1/
#480330000000
0!
0'
0/
#480340000000
1!
1'
1/
#480350000000
0!
1"
0'
1(
0/
10
#480360000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#480370000000
0!
0'
0/
#480380000000
1!
1'
1/
#480390000000
0!
0'
0/
#480400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#480410000000
0!
0'
0/
#480420000000
1!
1'
1/
#480430000000
0!
1"
0'
1(
0/
10
#480440000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#480450000000
0!
1$
0'
1+
0/
#480460000000
1!
1'
1/
#480470000000
0!
0'
0/
#480480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#480490000000
0!
0'
0/
#480500000000
1!
1'
1/
#480510000000
0!
0'
0/
#480520000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#480530000000
0!
0'
0/
#480540000000
1!
1'
1/
#480550000000
0!
0'
0/
#480560000000
1!
1'
1/
#480570000000
0!
0'
0/
#480580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#480590000000
0!
0'
0/
#480600000000
1!
1'
1/
#480610000000
0!
0'
0/
#480620000000
1!
1'
1/
#480630000000
0!
0'
0/
#480640000000
1!
1'
1/
#480650000000
0!
0'
0/
#480660000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#480670000000
0!
0'
0/
#480680000000
1!
1'
1/
#480690000000
0!
0'
0/
#480700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#480710000000
0!
0'
0/
#480720000000
1!
1'
1/
#480730000000
0!
0'
0/
#480740000000
#480750000000
1!
1'
1/
#480760000000
0!
0'
0/
#480770000000
1!
1'
1/
#480780000000
0!
1"
0'
1(
0/
10
#480790000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#480800000000
0!
0'
0/
#480810000000
1!
1'
1/
#480820000000
0!
0'
0/
#480830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#480840000000
0!
0'
0/
#480850000000
1!
1'
1/
#480860000000
0!
1"
0'
1(
0/
10
#480870000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#480880000000
0!
1$
0'
1+
0/
#480890000000
1!
1'
1/
#480900000000
0!
0'
0/
#480910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#480920000000
0!
0'
0/
#480930000000
1!
1'
1/
#480940000000
0!
0'
0/
#480950000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#480960000000
0!
0'
0/
#480970000000
1!
1'
1/
#480980000000
0!
0'
0/
#480990000000
1!
1'
1/
#481000000000
0!
0'
0/
#481010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#481020000000
0!
0'
0/
#481030000000
1!
1'
1/
#481040000000
0!
0'
0/
#481050000000
1!
1'
1/
#481060000000
0!
0'
0/
#481070000000
1!
1'
1/
#481080000000
0!
0'
0/
#481090000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#481100000000
0!
0'
0/
#481110000000
1!
1'
1/
#481120000000
0!
0'
0/
#481130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#481140000000
0!
0'
0/
#481150000000
1!
1'
1/
#481160000000
0!
0'
0/
#481170000000
#481180000000
1!
1'
1/
#481190000000
0!
0'
0/
#481200000000
1!
1'
1/
#481210000000
0!
1"
0'
1(
0/
10
#481220000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#481230000000
0!
0'
0/
#481240000000
1!
1'
1/
#481250000000
0!
0'
0/
#481260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#481270000000
0!
0'
0/
#481280000000
1!
1'
1/
#481290000000
0!
1"
0'
1(
0/
10
#481300000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#481310000000
0!
1$
0'
1+
0/
#481320000000
1!
1'
1/
#481330000000
0!
0'
0/
#481340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#481350000000
0!
0'
0/
#481360000000
1!
1'
1/
#481370000000
0!
0'
0/
#481380000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#481390000000
0!
0'
0/
#481400000000
1!
1'
1/
#481410000000
0!
0'
0/
#481420000000
1!
1'
1/
#481430000000
0!
0'
0/
#481440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#481450000000
0!
0'
0/
#481460000000
1!
1'
1/
#481470000000
0!
0'
0/
#481480000000
1!
1'
1/
#481490000000
0!
0'
0/
#481500000000
1!
1'
1/
#481510000000
0!
0'
0/
#481520000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#481530000000
0!
0'
0/
#481540000000
1!
1'
1/
#481550000000
0!
0'
0/
#481560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#481570000000
0!
0'
0/
#481580000000
1!
1'
1/
#481590000000
0!
0'
0/
#481600000000
#481610000000
1!
1'
1/
#481620000000
0!
0'
0/
#481630000000
1!
1'
1/
#481640000000
0!
1"
0'
1(
0/
10
#481650000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#481660000000
0!
0'
0/
#481670000000
1!
1'
1/
#481680000000
0!
0'
0/
#481690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#481700000000
0!
0'
0/
#481710000000
1!
1'
1/
#481720000000
0!
1"
0'
1(
0/
10
#481730000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#481740000000
0!
1$
0'
1+
0/
#481750000000
1!
1'
1/
#481760000000
0!
0'
0/
#481770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#481780000000
0!
0'
0/
#481790000000
1!
1'
1/
#481800000000
0!
0'
0/
#481810000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#481820000000
0!
0'
0/
#481830000000
1!
1'
1/
#481840000000
0!
0'
0/
#481850000000
1!
1'
1/
#481860000000
0!
0'
0/
#481870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#481880000000
0!
0'
0/
#481890000000
1!
1'
1/
#481900000000
0!
0'
0/
#481910000000
1!
1'
1/
#481920000000
0!
0'
0/
#481930000000
1!
1'
1/
#481940000000
0!
0'
0/
#481950000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#481960000000
0!
0'
0/
#481970000000
1!
1'
1/
#481980000000
0!
0'
0/
#481990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#482000000000
0!
0'
0/
#482010000000
1!
1'
1/
#482020000000
0!
0'
0/
#482030000000
#482040000000
1!
1'
1/
#482050000000
0!
0'
0/
#482060000000
1!
1'
1/
#482070000000
0!
1"
0'
1(
0/
10
#482080000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#482090000000
0!
0'
0/
#482100000000
1!
1'
1/
#482110000000
0!
0'
0/
#482120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#482130000000
0!
0'
0/
#482140000000
1!
1'
1/
#482150000000
0!
1"
0'
1(
0/
10
#482160000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#482170000000
0!
1$
0'
1+
0/
#482180000000
1!
1'
1/
#482190000000
0!
0'
0/
#482200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#482210000000
0!
0'
0/
#482220000000
1!
1'
1/
#482230000000
0!
0'
0/
#482240000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#482250000000
0!
0'
0/
#482260000000
1!
1'
1/
#482270000000
0!
0'
0/
#482280000000
1!
1'
1/
#482290000000
0!
0'
0/
#482300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#482310000000
0!
0'
0/
#482320000000
1!
1'
1/
#482330000000
0!
0'
0/
#482340000000
1!
1'
1/
#482350000000
0!
0'
0/
#482360000000
1!
1'
1/
#482370000000
0!
0'
0/
#482380000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#482390000000
0!
0'
0/
#482400000000
1!
1'
1/
#482410000000
0!
0'
0/
#482420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#482430000000
0!
0'
0/
#482440000000
1!
1'
1/
#482450000000
0!
0'
0/
#482460000000
#482470000000
1!
1'
1/
#482480000000
0!
0'
0/
#482490000000
1!
1'
1/
#482500000000
0!
1"
0'
1(
0/
10
#482510000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#482520000000
0!
0'
0/
#482530000000
1!
1'
1/
#482540000000
0!
0'
0/
#482550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#482560000000
0!
0'
0/
#482570000000
1!
1'
1/
#482580000000
0!
1"
0'
1(
0/
10
#482590000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#482600000000
0!
1$
0'
1+
0/
#482610000000
1!
1'
1/
#482620000000
0!
0'
0/
#482630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#482640000000
0!
0'
0/
#482650000000
1!
1'
1/
#482660000000
0!
0'
0/
#482670000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#482680000000
0!
0'
0/
#482690000000
1!
1'
1/
#482700000000
0!
0'
0/
#482710000000
1!
1'
1/
#482720000000
0!
0'
0/
#482730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#482740000000
0!
0'
0/
#482750000000
1!
1'
1/
#482760000000
0!
0'
0/
#482770000000
1!
1'
1/
#482780000000
0!
0'
0/
#482790000000
1!
1'
1/
#482800000000
0!
0'
0/
#482810000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#482820000000
0!
0'
0/
#482830000000
1!
1'
1/
#482840000000
0!
0'
0/
#482850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#482860000000
0!
0'
0/
#482870000000
1!
1'
1/
#482880000000
0!
0'
0/
#482890000000
#482900000000
1!
1'
1/
#482910000000
0!
0'
0/
#482920000000
1!
1'
1/
#482930000000
0!
1"
0'
1(
0/
10
#482940000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#482950000000
0!
0'
0/
#482960000000
1!
1'
1/
#482970000000
0!
0'
0/
#482980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#482990000000
0!
0'
0/
#483000000000
1!
1'
1/
#483010000000
0!
1"
0'
1(
0/
10
#483020000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#483030000000
0!
1$
0'
1+
0/
#483040000000
1!
1'
1/
#483050000000
0!
0'
0/
#483060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#483070000000
0!
0'
0/
#483080000000
1!
1'
1/
#483090000000
0!
0'
0/
#483100000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#483110000000
0!
0'
0/
#483120000000
1!
1'
1/
#483130000000
0!
0'
0/
#483140000000
1!
1'
1/
#483150000000
0!
0'
0/
#483160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#483170000000
0!
0'
0/
#483180000000
1!
1'
1/
#483190000000
0!
0'
0/
#483200000000
1!
1'
1/
#483210000000
0!
0'
0/
#483220000000
1!
1'
1/
#483230000000
0!
0'
0/
#483240000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#483250000000
0!
0'
0/
#483260000000
1!
1'
1/
#483270000000
0!
0'
0/
#483280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#483290000000
0!
0'
0/
#483300000000
1!
1'
1/
#483310000000
0!
0'
0/
#483320000000
#483330000000
1!
1'
1/
#483340000000
0!
0'
0/
#483350000000
1!
1'
1/
#483360000000
0!
1"
0'
1(
0/
10
#483370000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#483380000000
0!
0'
0/
#483390000000
1!
1'
1/
#483400000000
0!
0'
0/
#483410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#483420000000
0!
0'
0/
#483430000000
1!
1'
1/
#483440000000
0!
1"
0'
1(
0/
10
#483450000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#483460000000
0!
1$
0'
1+
0/
#483470000000
1!
1'
1/
#483480000000
0!
0'
0/
#483490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#483500000000
0!
0'
0/
#483510000000
1!
1'
1/
#483520000000
0!
0'
0/
#483530000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#483540000000
0!
0'
0/
#483550000000
1!
1'
1/
#483560000000
0!
0'
0/
#483570000000
1!
1'
1/
#483580000000
0!
0'
0/
#483590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#483600000000
0!
0'
0/
#483610000000
1!
1'
1/
#483620000000
0!
0'
0/
#483630000000
1!
1'
1/
#483640000000
0!
0'
0/
#483650000000
1!
1'
1/
#483660000000
0!
0'
0/
#483670000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#483680000000
0!
0'
0/
#483690000000
1!
1'
1/
#483700000000
0!
0'
0/
#483710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#483720000000
0!
0'
0/
#483730000000
1!
1'
1/
#483740000000
0!
0'
0/
#483750000000
#483760000000
1!
1'
1/
#483770000000
0!
0'
0/
#483780000000
1!
1'
1/
#483790000000
0!
1"
0'
1(
0/
10
#483800000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#483810000000
0!
0'
0/
#483820000000
1!
1'
1/
#483830000000
0!
0'
0/
#483840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#483850000000
0!
0'
0/
#483860000000
1!
1'
1/
#483870000000
0!
1"
0'
1(
0/
10
#483880000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#483890000000
0!
1$
0'
1+
0/
#483900000000
1!
1'
1/
#483910000000
0!
0'
0/
#483920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#483930000000
0!
0'
0/
#483940000000
1!
1'
1/
#483950000000
0!
0'
0/
#483960000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#483970000000
0!
0'
0/
#483980000000
1!
1'
1/
#483990000000
0!
0'
0/
#484000000000
1!
1'
1/
#484010000000
0!
0'
0/
#484020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#484030000000
0!
0'
0/
#484040000000
1!
1'
1/
#484050000000
0!
0'
0/
#484060000000
1!
1'
1/
#484070000000
0!
0'
0/
#484080000000
1!
1'
1/
#484090000000
0!
0'
0/
#484100000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#484110000000
0!
0'
0/
#484120000000
1!
1'
1/
#484130000000
0!
0'
0/
#484140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#484150000000
0!
0'
0/
#484160000000
1!
1'
1/
#484170000000
0!
0'
0/
#484180000000
#484190000000
1!
1'
1/
#484200000000
0!
0'
0/
#484210000000
1!
1'
1/
#484220000000
0!
1"
0'
1(
0/
10
#484230000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#484240000000
0!
0'
0/
#484250000000
1!
1'
1/
#484260000000
0!
0'
0/
#484270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#484280000000
0!
0'
0/
#484290000000
1!
1'
1/
#484300000000
0!
1"
0'
1(
0/
10
#484310000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#484320000000
0!
1$
0'
1+
0/
#484330000000
1!
1'
1/
#484340000000
0!
0'
0/
#484350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#484360000000
0!
0'
0/
#484370000000
1!
1'
1/
#484380000000
0!
0'
0/
#484390000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#484400000000
0!
0'
0/
#484410000000
1!
1'
1/
#484420000000
0!
0'
0/
#484430000000
1!
1'
1/
#484440000000
0!
0'
0/
#484450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#484460000000
0!
0'
0/
#484470000000
1!
1'
1/
#484480000000
0!
0'
0/
#484490000000
1!
1'
1/
#484500000000
0!
0'
0/
#484510000000
1!
1'
1/
#484520000000
0!
0'
0/
#484530000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#484540000000
0!
0'
0/
#484550000000
1!
1'
1/
#484560000000
0!
0'
0/
#484570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#484580000000
0!
0'
0/
#484590000000
1!
1'
1/
#484600000000
0!
0'
0/
#484610000000
#484620000000
1!
1'
1/
#484630000000
0!
0'
0/
#484640000000
1!
1'
1/
#484650000000
0!
1"
0'
1(
0/
10
#484660000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#484670000000
0!
0'
0/
#484680000000
1!
1'
1/
#484690000000
0!
0'
0/
#484700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#484710000000
0!
0'
0/
#484720000000
1!
1'
1/
#484730000000
0!
1"
0'
1(
0/
10
#484740000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#484750000000
0!
1$
0'
1+
0/
#484760000000
1!
1'
1/
#484770000000
0!
0'
0/
#484780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#484790000000
0!
0'
0/
#484800000000
1!
1'
1/
#484810000000
0!
0'
0/
#484820000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#484830000000
0!
0'
0/
#484840000000
1!
1'
1/
#484850000000
0!
0'
0/
#484860000000
1!
1'
1/
#484870000000
0!
0'
0/
#484880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#484890000000
0!
0'
0/
#484900000000
1!
1'
1/
#484910000000
0!
0'
0/
#484920000000
1!
1'
1/
#484930000000
0!
0'
0/
#484940000000
1!
1'
1/
#484950000000
0!
0'
0/
#484960000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#484970000000
0!
0'
0/
#484980000000
1!
1'
1/
#484990000000
0!
0'
0/
#485000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#485010000000
0!
0'
0/
#485020000000
1!
1'
1/
#485030000000
0!
0'
0/
#485040000000
#485050000000
1!
1'
1/
#485060000000
0!
0'
0/
#485070000000
1!
1'
1/
#485080000000
0!
1"
0'
1(
0/
10
#485090000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#485100000000
0!
0'
0/
#485110000000
1!
1'
1/
#485120000000
0!
0'
0/
#485130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#485140000000
0!
0'
0/
#485150000000
1!
1'
1/
#485160000000
0!
1"
0'
1(
0/
10
#485170000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#485180000000
0!
1$
0'
1+
0/
#485190000000
1!
1'
1/
#485200000000
0!
0'
0/
#485210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#485220000000
0!
0'
0/
#485230000000
1!
1'
1/
#485240000000
0!
0'
0/
#485250000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#485260000000
0!
0'
0/
#485270000000
1!
1'
1/
#485280000000
0!
0'
0/
#485290000000
1!
1'
1/
#485300000000
0!
0'
0/
#485310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#485320000000
0!
0'
0/
#485330000000
1!
1'
1/
#485340000000
0!
0'
0/
#485350000000
1!
1'
1/
#485360000000
0!
0'
0/
#485370000000
1!
1'
1/
#485380000000
0!
0'
0/
#485390000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#485400000000
0!
0'
0/
#485410000000
1!
1'
1/
#485420000000
0!
0'
0/
#485430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#485440000000
0!
0'
0/
#485450000000
1!
1'
1/
#485460000000
0!
0'
0/
#485470000000
#485480000000
1!
1'
1/
#485490000000
0!
0'
0/
#485500000000
1!
1'
1/
#485510000000
0!
1"
0'
1(
0/
10
#485520000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#485530000000
0!
0'
0/
#485540000000
1!
1'
1/
#485550000000
0!
0'
0/
#485560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#485570000000
0!
0'
0/
#485580000000
1!
1'
1/
#485590000000
0!
1"
0'
1(
0/
10
#485600000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#485610000000
0!
1$
0'
1+
0/
#485620000000
1!
1'
1/
#485630000000
0!
0'
0/
#485640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#485650000000
0!
0'
0/
#485660000000
1!
1'
1/
#485670000000
0!
0'
0/
#485680000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#485690000000
0!
0'
0/
#485700000000
1!
1'
1/
#485710000000
0!
0'
0/
#485720000000
1!
1'
1/
#485730000000
0!
0'
0/
#485740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#485750000000
0!
0'
0/
#485760000000
1!
1'
1/
#485770000000
0!
0'
0/
#485780000000
1!
1'
1/
#485790000000
0!
0'
0/
#485800000000
1!
1'
1/
#485810000000
0!
0'
0/
#485820000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#485830000000
0!
0'
0/
#485840000000
1!
1'
1/
#485850000000
0!
0'
0/
#485860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#485870000000
0!
0'
0/
#485880000000
1!
1'
1/
#485890000000
0!
0'
0/
#485900000000
#485910000000
1!
1'
1/
#485920000000
0!
0'
0/
#485930000000
1!
1'
1/
#485940000000
0!
1"
0'
1(
0/
10
#485950000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#485960000000
0!
0'
0/
#485970000000
1!
1'
1/
#485980000000
0!
0'
0/
#485990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#486000000000
0!
0'
0/
#486010000000
1!
1'
1/
#486020000000
0!
1"
0'
1(
0/
10
#486030000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#486040000000
0!
1$
0'
1+
0/
#486050000000
1!
1'
1/
#486060000000
0!
0'
0/
#486070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#486080000000
0!
0'
0/
#486090000000
1!
1'
1/
#486100000000
0!
0'
0/
#486110000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#486120000000
0!
0'
0/
#486130000000
1!
1'
1/
#486140000000
0!
0'
0/
#486150000000
1!
1'
1/
#486160000000
0!
0'
0/
#486170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#486180000000
0!
0'
0/
#486190000000
1!
1'
1/
#486200000000
0!
0'
0/
#486210000000
1!
1'
1/
#486220000000
0!
0'
0/
#486230000000
1!
1'
1/
#486240000000
0!
0'
0/
#486250000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#486260000000
0!
0'
0/
#486270000000
1!
1'
1/
#486280000000
0!
0'
0/
#486290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#486300000000
0!
0'
0/
#486310000000
1!
1'
1/
#486320000000
0!
0'
0/
#486330000000
#486340000000
1!
1'
1/
#486350000000
0!
0'
0/
#486360000000
1!
1'
1/
#486370000000
0!
1"
0'
1(
0/
10
#486380000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#486390000000
0!
0'
0/
#486400000000
1!
1'
1/
#486410000000
0!
0'
0/
#486420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#486430000000
0!
0'
0/
#486440000000
1!
1'
1/
#486450000000
0!
1"
0'
1(
0/
10
#486460000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#486470000000
0!
1$
0'
1+
0/
#486480000000
1!
1'
1/
#486490000000
0!
0'
0/
#486500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#486510000000
0!
0'
0/
#486520000000
1!
1'
1/
#486530000000
0!
0'
0/
#486540000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#486550000000
0!
0'
0/
#486560000000
1!
1'
1/
#486570000000
0!
0'
0/
#486580000000
1!
1'
1/
#486590000000
0!
0'
0/
#486600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#486610000000
0!
0'
0/
#486620000000
1!
1'
1/
#486630000000
0!
0'
0/
#486640000000
1!
1'
1/
#486650000000
0!
0'
0/
#486660000000
1!
1'
1/
#486670000000
0!
0'
0/
#486680000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#486690000000
0!
0'
0/
#486700000000
1!
1'
1/
#486710000000
0!
0'
0/
#486720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#486730000000
0!
0'
0/
#486740000000
1!
1'
1/
#486750000000
0!
0'
0/
#486760000000
#486770000000
1!
1'
1/
#486780000000
0!
0'
0/
#486790000000
1!
1'
1/
#486800000000
0!
1"
0'
1(
0/
10
#486810000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#486820000000
0!
0'
0/
#486830000000
1!
1'
1/
#486840000000
0!
0'
0/
#486850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#486860000000
0!
0'
0/
#486870000000
1!
1'
1/
#486880000000
0!
1"
0'
1(
0/
10
#486890000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#486900000000
0!
1$
0'
1+
0/
#486910000000
1!
1'
1/
#486920000000
0!
0'
0/
#486930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#486940000000
0!
0'
0/
#486950000000
1!
1'
1/
#486960000000
0!
0'
0/
#486970000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#486980000000
0!
0'
0/
#486990000000
1!
1'
1/
#487000000000
0!
0'
0/
#487010000000
1!
1'
1/
#487020000000
0!
0'
0/
#487030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#487040000000
0!
0'
0/
#487050000000
1!
1'
1/
#487060000000
0!
0'
0/
#487070000000
1!
1'
1/
#487080000000
0!
0'
0/
#487090000000
1!
1'
1/
#487100000000
0!
0'
0/
#487110000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#487120000000
0!
0'
0/
#487130000000
1!
1'
1/
#487140000000
0!
0'
0/
#487150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#487160000000
0!
0'
0/
#487170000000
1!
1'
1/
#487180000000
0!
0'
0/
#487190000000
#487200000000
1!
1'
1/
#487210000000
0!
0'
0/
#487220000000
1!
1'
1/
#487230000000
0!
1"
0'
1(
0/
10
#487240000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#487250000000
0!
0'
0/
#487260000000
1!
1'
1/
#487270000000
0!
0'
0/
#487280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#487290000000
0!
0'
0/
#487300000000
1!
1'
1/
#487310000000
0!
1"
0'
1(
0/
10
#487320000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#487330000000
0!
1$
0'
1+
0/
#487340000000
1!
1'
1/
#487350000000
0!
0'
0/
#487360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#487370000000
0!
0'
0/
#487380000000
1!
1'
1/
#487390000000
0!
0'
0/
#487400000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#487410000000
0!
0'
0/
#487420000000
1!
1'
1/
#487430000000
0!
0'
0/
#487440000000
1!
1'
1/
#487450000000
0!
0'
0/
#487460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#487470000000
0!
0'
0/
#487480000000
1!
1'
1/
#487490000000
0!
0'
0/
#487500000000
1!
1'
1/
#487510000000
0!
0'
0/
#487520000000
1!
1'
1/
#487530000000
0!
0'
0/
#487540000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#487550000000
0!
0'
0/
#487560000000
1!
1'
1/
#487570000000
0!
0'
0/
#487580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#487590000000
0!
0'
0/
#487600000000
1!
1'
1/
#487610000000
0!
0'
0/
#487620000000
#487630000000
1!
1'
1/
#487640000000
0!
0'
0/
#487650000000
1!
1'
1/
#487660000000
0!
1"
0'
1(
0/
10
#487670000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#487680000000
0!
0'
0/
#487690000000
1!
1'
1/
#487700000000
0!
0'
0/
#487710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#487720000000
0!
0'
0/
#487730000000
1!
1'
1/
#487740000000
0!
1"
0'
1(
0/
10
#487750000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#487760000000
0!
1$
0'
1+
0/
#487770000000
1!
1'
1/
#487780000000
0!
0'
0/
#487790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#487800000000
0!
0'
0/
#487810000000
1!
1'
1/
#487820000000
0!
0'
0/
#487830000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#487840000000
0!
0'
0/
#487850000000
1!
1'
1/
#487860000000
0!
0'
0/
#487870000000
1!
1'
1/
#487880000000
0!
0'
0/
#487890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#487900000000
0!
0'
0/
#487910000000
1!
1'
1/
#487920000000
0!
0'
0/
#487930000000
1!
1'
1/
#487940000000
0!
0'
0/
#487950000000
1!
1'
1/
#487960000000
0!
0'
0/
#487970000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#487980000000
0!
0'
0/
#487990000000
1!
1'
1/
#488000000000
0!
0'
0/
#488010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#488020000000
0!
0'
0/
#488030000000
1!
1'
1/
#488040000000
0!
0'
0/
#488050000000
#488060000000
1!
1'
1/
#488070000000
0!
0'
0/
#488080000000
1!
1'
1/
#488090000000
0!
1"
0'
1(
0/
10
#488100000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#488110000000
0!
0'
0/
#488120000000
1!
1'
1/
#488130000000
0!
0'
0/
#488140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#488150000000
0!
0'
0/
#488160000000
1!
1'
1/
#488170000000
0!
1"
0'
1(
0/
10
#488180000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#488190000000
0!
1$
0'
1+
0/
#488200000000
1!
1'
1/
#488210000000
0!
0'
0/
#488220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#488230000000
0!
0'
0/
#488240000000
1!
1'
1/
#488250000000
0!
0'
0/
#488260000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#488270000000
0!
0'
0/
#488280000000
1!
1'
1/
#488290000000
0!
0'
0/
#488300000000
1!
1'
1/
#488310000000
0!
0'
0/
#488320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#488330000000
0!
0'
0/
#488340000000
1!
1'
1/
#488350000000
0!
0'
0/
#488360000000
1!
1'
1/
#488370000000
0!
0'
0/
#488380000000
1!
1'
1/
#488390000000
0!
0'
0/
#488400000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#488410000000
0!
0'
0/
#488420000000
1!
1'
1/
#488430000000
0!
0'
0/
#488440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#488450000000
0!
0'
0/
#488460000000
1!
1'
1/
#488470000000
0!
0'
0/
#488480000000
#488490000000
1!
1'
1/
#488500000000
0!
0'
0/
#488510000000
1!
1'
1/
#488520000000
0!
1"
0'
1(
0/
10
#488530000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#488540000000
0!
0'
0/
#488550000000
1!
1'
1/
#488560000000
0!
0'
0/
#488570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#488580000000
0!
0'
0/
#488590000000
1!
1'
1/
#488600000000
0!
1"
0'
1(
0/
10
#488610000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#488620000000
0!
1$
0'
1+
0/
#488630000000
1!
1'
1/
#488640000000
0!
0'
0/
#488650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#488660000000
0!
0'
0/
#488670000000
1!
1'
1/
#488680000000
0!
0'
0/
#488690000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#488700000000
0!
0'
0/
#488710000000
1!
1'
1/
#488720000000
0!
0'
0/
#488730000000
1!
1'
1/
#488740000000
0!
0'
0/
#488750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#488760000000
0!
0'
0/
#488770000000
1!
1'
1/
#488780000000
0!
0'
0/
#488790000000
1!
1'
1/
#488800000000
0!
0'
0/
#488810000000
1!
1'
1/
#488820000000
0!
0'
0/
#488830000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#488840000000
0!
0'
0/
#488850000000
1!
1'
1/
#488860000000
0!
0'
0/
#488870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#488880000000
0!
0'
0/
#488890000000
1!
1'
1/
#488900000000
0!
0'
0/
#488910000000
#488920000000
1!
1'
1/
#488930000000
0!
0'
0/
#488940000000
1!
1'
1/
#488950000000
0!
1"
0'
1(
0/
10
#488960000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#488970000000
0!
0'
0/
#488980000000
1!
1'
1/
#488990000000
0!
0'
0/
#489000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#489010000000
0!
0'
0/
#489020000000
1!
1'
1/
#489030000000
0!
1"
0'
1(
0/
10
#489040000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#489050000000
0!
1$
0'
1+
0/
#489060000000
1!
1'
1/
#489070000000
0!
0'
0/
#489080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#489090000000
0!
0'
0/
#489100000000
1!
1'
1/
#489110000000
0!
0'
0/
#489120000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#489130000000
0!
0'
0/
#489140000000
1!
1'
1/
#489150000000
0!
0'
0/
#489160000000
1!
1'
1/
#489170000000
0!
0'
0/
#489180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#489190000000
0!
0'
0/
#489200000000
1!
1'
1/
#489210000000
0!
0'
0/
#489220000000
1!
1'
1/
#489230000000
0!
0'
0/
#489240000000
1!
1'
1/
#489250000000
0!
0'
0/
#489260000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#489270000000
0!
0'
0/
#489280000000
1!
1'
1/
#489290000000
0!
0'
0/
#489300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#489310000000
0!
0'
0/
#489320000000
1!
1'
1/
#489330000000
0!
0'
0/
#489340000000
#489350000000
1!
1'
1/
#489360000000
0!
0'
0/
#489370000000
1!
1'
1/
#489380000000
0!
1"
0'
1(
0/
10
#489390000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#489400000000
0!
0'
0/
#489410000000
1!
1'
1/
#489420000000
0!
0'
0/
#489430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#489440000000
0!
0'
0/
#489450000000
1!
1'
1/
#489460000000
0!
1"
0'
1(
0/
10
#489470000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#489480000000
0!
1$
0'
1+
0/
#489490000000
1!
1'
1/
#489500000000
0!
0'
0/
#489510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#489520000000
0!
0'
0/
#489530000000
1!
1'
1/
#489540000000
0!
0'
0/
#489550000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#489560000000
0!
0'
0/
#489570000000
1!
1'
1/
#489580000000
0!
0'
0/
#489590000000
1!
1'
1/
#489600000000
0!
0'
0/
#489610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#489620000000
0!
0'
0/
#489630000000
1!
1'
1/
#489640000000
0!
0'
0/
#489650000000
1!
1'
1/
#489660000000
0!
0'
0/
#489670000000
1!
1'
1/
#489680000000
0!
0'
0/
#489690000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#489700000000
0!
0'
0/
#489710000000
1!
1'
1/
#489720000000
0!
0'
0/
#489730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#489740000000
0!
0'
0/
#489750000000
1!
1'
1/
#489760000000
0!
0'
0/
#489770000000
#489780000000
1!
1'
1/
#489790000000
0!
0'
0/
#489800000000
1!
1'
1/
#489810000000
0!
1"
0'
1(
0/
10
#489820000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#489830000000
0!
0'
0/
#489840000000
1!
1'
1/
#489850000000
0!
0'
0/
#489860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#489870000000
0!
0'
0/
#489880000000
1!
1'
1/
#489890000000
0!
1"
0'
1(
0/
10
#489900000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#489910000000
0!
1$
0'
1+
0/
#489920000000
1!
1'
1/
#489930000000
0!
0'
0/
#489940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#489950000000
0!
0'
0/
#489960000000
1!
1'
1/
#489970000000
0!
0'
0/
#489980000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#489990000000
0!
0'
0/
#490000000000
1!
1'
1/
#490010000000
0!
0'
0/
#490020000000
1!
1'
1/
#490030000000
0!
0'
0/
#490040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#490050000000
0!
0'
0/
#490060000000
1!
1'
1/
#490070000000
0!
0'
0/
#490080000000
1!
1'
1/
#490090000000
0!
0'
0/
#490100000000
1!
1'
1/
#490110000000
0!
0'
0/
#490120000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#490130000000
0!
0'
0/
#490140000000
1!
1'
1/
#490150000000
0!
0'
0/
#490160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#490170000000
0!
0'
0/
#490180000000
1!
1'
1/
#490190000000
0!
0'
0/
#490200000000
#490210000000
1!
1'
1/
#490220000000
0!
0'
0/
#490230000000
1!
1'
1/
#490240000000
0!
1"
0'
1(
0/
10
#490250000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#490260000000
0!
0'
0/
#490270000000
1!
1'
1/
#490280000000
0!
0'
0/
#490290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#490300000000
0!
0'
0/
#490310000000
1!
1'
1/
#490320000000
0!
1"
0'
1(
0/
10
#490330000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#490340000000
0!
1$
0'
1+
0/
#490350000000
1!
1'
1/
#490360000000
0!
0'
0/
#490370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#490380000000
0!
0'
0/
#490390000000
1!
1'
1/
#490400000000
0!
0'
0/
#490410000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#490420000000
0!
0'
0/
#490430000000
1!
1'
1/
#490440000000
0!
0'
0/
#490450000000
1!
1'
1/
#490460000000
0!
0'
0/
#490470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#490480000000
0!
0'
0/
#490490000000
1!
1'
1/
#490500000000
0!
0'
0/
#490510000000
1!
1'
1/
#490520000000
0!
0'
0/
#490530000000
1!
1'
1/
#490540000000
0!
0'
0/
#490550000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#490560000000
0!
0'
0/
#490570000000
1!
1'
1/
#490580000000
0!
0'
0/
#490590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#490600000000
0!
0'
0/
#490610000000
1!
1'
1/
#490620000000
0!
0'
0/
#490630000000
#490640000000
1!
1'
1/
#490650000000
0!
0'
0/
#490660000000
1!
1'
1/
#490670000000
0!
1"
0'
1(
0/
10
#490680000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#490690000000
0!
0'
0/
#490700000000
1!
1'
1/
#490710000000
0!
0'
0/
#490720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#490730000000
0!
0'
0/
#490740000000
1!
1'
1/
#490750000000
0!
1"
0'
1(
0/
10
#490760000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#490770000000
0!
1$
0'
1+
0/
#490780000000
1!
1'
1/
#490790000000
0!
0'
0/
#490800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#490810000000
0!
0'
0/
#490820000000
1!
1'
1/
#490830000000
0!
0'
0/
#490840000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#490850000000
0!
0'
0/
#490860000000
1!
1'
1/
#490870000000
0!
0'
0/
#490880000000
1!
1'
1/
#490890000000
0!
0'
0/
#490900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#490910000000
0!
0'
0/
#490920000000
1!
1'
1/
#490930000000
0!
0'
0/
#490940000000
1!
1'
1/
#490950000000
0!
0'
0/
#490960000000
1!
1'
1/
#490970000000
0!
0'
0/
#490980000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#490990000000
0!
0'
0/
#491000000000
1!
1'
1/
#491010000000
0!
0'
0/
#491020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#491030000000
0!
0'
0/
#491040000000
1!
1'
1/
#491050000000
0!
0'
0/
#491060000000
#491070000000
1!
1'
1/
#491080000000
0!
0'
0/
#491090000000
1!
1'
1/
#491100000000
0!
1"
0'
1(
0/
10
#491110000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#491120000000
0!
0'
0/
#491130000000
1!
1'
1/
#491140000000
0!
0'
0/
#491150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#491160000000
0!
0'
0/
#491170000000
1!
1'
1/
#491180000000
0!
1"
0'
1(
0/
10
#491190000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#491200000000
0!
1$
0'
1+
0/
#491210000000
1!
1'
1/
#491220000000
0!
0'
0/
#491230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#491240000000
0!
0'
0/
#491250000000
1!
1'
1/
#491260000000
0!
0'
0/
#491270000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#491280000000
0!
0'
0/
#491290000000
1!
1'
1/
#491300000000
0!
0'
0/
#491310000000
1!
1'
1/
#491320000000
0!
0'
0/
#491330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#491340000000
0!
0'
0/
#491350000000
1!
1'
1/
#491360000000
0!
0'
0/
#491370000000
1!
1'
1/
#491380000000
0!
0'
0/
#491390000000
1!
1'
1/
#491400000000
0!
0'
0/
#491410000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#491420000000
0!
0'
0/
#491430000000
1!
1'
1/
#491440000000
0!
0'
0/
#491450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#491460000000
0!
0'
0/
#491470000000
1!
1'
1/
#491480000000
0!
0'
0/
#491490000000
#491500000000
1!
1'
1/
#491510000000
0!
0'
0/
#491520000000
1!
1'
1/
#491530000000
0!
1"
0'
1(
0/
10
#491540000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#491550000000
0!
0'
0/
#491560000000
1!
1'
1/
#491570000000
0!
0'
0/
#491580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#491590000000
0!
0'
0/
#491600000000
1!
1'
1/
#491610000000
0!
1"
0'
1(
0/
10
#491620000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#491630000000
0!
1$
0'
1+
0/
#491640000000
1!
1'
1/
#491650000000
0!
0'
0/
#491660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#491670000000
0!
0'
0/
#491680000000
1!
1'
1/
#491690000000
0!
0'
0/
#491700000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#491710000000
0!
0'
0/
#491720000000
1!
1'
1/
#491730000000
0!
0'
0/
#491740000000
1!
1'
1/
#491750000000
0!
0'
0/
#491760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#491770000000
0!
0'
0/
#491780000000
1!
1'
1/
#491790000000
0!
0'
0/
#491800000000
1!
1'
1/
#491810000000
0!
0'
0/
#491820000000
1!
1'
1/
#491830000000
0!
0'
0/
#491840000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#491850000000
0!
0'
0/
#491860000000
1!
1'
1/
#491870000000
0!
0'
0/
#491880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#491890000000
0!
0'
0/
#491900000000
1!
1'
1/
#491910000000
0!
0'
0/
#491920000000
#491930000000
1!
1'
1/
#491940000000
0!
0'
0/
#491950000000
1!
1'
1/
#491960000000
0!
1"
0'
1(
0/
10
#491970000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#491980000000
0!
0'
0/
#491990000000
1!
1'
1/
#492000000000
0!
0'
0/
#492010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#492020000000
0!
0'
0/
#492030000000
1!
1'
1/
#492040000000
0!
1"
0'
1(
0/
10
#492050000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#492060000000
0!
1$
0'
1+
0/
#492070000000
1!
1'
1/
#492080000000
0!
0'
0/
#492090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#492100000000
0!
0'
0/
#492110000000
1!
1'
1/
#492120000000
0!
0'
0/
#492130000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#492140000000
0!
0'
0/
#492150000000
1!
1'
1/
#492160000000
0!
0'
0/
#492170000000
1!
1'
1/
#492180000000
0!
0'
0/
#492190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#492200000000
0!
0'
0/
#492210000000
1!
1'
1/
#492220000000
0!
0'
0/
#492230000000
1!
1'
1/
#492240000000
0!
0'
0/
#492250000000
1!
1'
1/
#492260000000
0!
0'
0/
#492270000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#492280000000
0!
0'
0/
#492290000000
1!
1'
1/
#492300000000
0!
0'
0/
#492310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#492320000000
0!
0'
0/
#492330000000
1!
1'
1/
#492340000000
0!
0'
0/
#492350000000
#492360000000
1!
1'
1/
#492370000000
0!
0'
0/
#492380000000
1!
1'
1/
#492390000000
0!
1"
0'
1(
0/
10
#492400000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#492410000000
0!
0'
0/
#492420000000
1!
1'
1/
#492430000000
0!
0'
0/
#492440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#492450000000
0!
0'
0/
#492460000000
1!
1'
1/
#492470000000
0!
1"
0'
1(
0/
10
#492480000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#492490000000
0!
1$
0'
1+
0/
#492500000000
1!
1'
1/
#492510000000
0!
0'
0/
#492520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#492530000000
0!
0'
0/
#492540000000
1!
1'
1/
#492550000000
0!
0'
0/
#492560000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#492570000000
0!
0'
0/
#492580000000
1!
1'
1/
#492590000000
0!
0'
0/
#492600000000
1!
1'
1/
#492610000000
0!
0'
0/
#492620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#492630000000
0!
0'
0/
#492640000000
1!
1'
1/
#492650000000
0!
0'
0/
#492660000000
1!
1'
1/
#492670000000
0!
0'
0/
#492680000000
1!
1'
1/
#492690000000
0!
0'
0/
#492700000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#492710000000
0!
0'
0/
#492720000000
1!
1'
1/
#492730000000
0!
0'
0/
#492740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#492750000000
0!
0'
0/
#492760000000
1!
1'
1/
#492770000000
0!
0'
0/
#492780000000
#492790000000
1!
1'
1/
#492800000000
0!
0'
0/
#492810000000
1!
1'
1/
#492820000000
0!
1"
0'
1(
0/
10
#492830000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#492840000000
0!
0'
0/
#492850000000
1!
1'
1/
#492860000000
0!
0'
0/
#492870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#492880000000
0!
0'
0/
#492890000000
1!
1'
1/
#492900000000
0!
1"
0'
1(
0/
10
#492910000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#492920000000
0!
1$
0'
1+
0/
#492930000000
1!
1'
1/
#492940000000
0!
0'
0/
#492950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#492960000000
0!
0'
0/
#492970000000
1!
1'
1/
#492980000000
0!
0'
0/
#492990000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#493000000000
0!
0'
0/
#493010000000
1!
1'
1/
#493020000000
0!
0'
0/
#493030000000
1!
1'
1/
#493040000000
0!
0'
0/
#493050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#493060000000
0!
0'
0/
#493070000000
1!
1'
1/
#493080000000
0!
0'
0/
#493090000000
1!
1'
1/
#493100000000
0!
0'
0/
#493110000000
1!
1'
1/
#493120000000
0!
0'
0/
#493130000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#493140000000
0!
0'
0/
#493150000000
1!
1'
1/
#493160000000
0!
0'
0/
#493170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#493180000000
0!
0'
0/
#493190000000
1!
1'
1/
#493200000000
0!
0'
0/
#493210000000
#493220000000
1!
1'
1/
#493230000000
0!
0'
0/
#493240000000
1!
1'
1/
#493250000000
0!
1"
0'
1(
0/
10
#493260000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#493270000000
0!
0'
0/
#493280000000
1!
1'
1/
#493290000000
0!
0'
0/
#493300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#493310000000
0!
0'
0/
#493320000000
1!
1'
1/
#493330000000
0!
1"
0'
1(
0/
10
#493340000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#493350000000
0!
1$
0'
1+
0/
#493360000000
1!
1'
1/
#493370000000
0!
0'
0/
#493380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#493390000000
0!
0'
0/
#493400000000
1!
1'
1/
#493410000000
0!
0'
0/
#493420000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#493430000000
0!
0'
0/
#493440000000
1!
1'
1/
#493450000000
0!
0'
0/
#493460000000
1!
1'
1/
#493470000000
0!
0'
0/
#493480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#493490000000
0!
0'
0/
#493500000000
1!
1'
1/
#493510000000
0!
0'
0/
#493520000000
1!
1'
1/
#493530000000
0!
0'
0/
#493540000000
1!
1'
1/
#493550000000
0!
0'
0/
#493560000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#493570000000
0!
0'
0/
#493580000000
1!
1'
1/
#493590000000
0!
0'
0/
#493600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#493610000000
0!
0'
0/
#493620000000
1!
1'
1/
#493630000000
0!
0'
0/
#493640000000
#493650000000
1!
1'
1/
#493660000000
0!
0'
0/
#493670000000
1!
1'
1/
#493680000000
0!
1"
0'
1(
0/
10
#493690000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#493700000000
0!
0'
0/
#493710000000
1!
1'
1/
#493720000000
0!
0'
0/
#493730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#493740000000
0!
0'
0/
#493750000000
1!
1'
1/
#493760000000
0!
1"
0'
1(
0/
10
#493770000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#493780000000
0!
1$
0'
1+
0/
#493790000000
1!
1'
1/
#493800000000
0!
0'
0/
#493810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#493820000000
0!
0'
0/
#493830000000
1!
1'
1/
#493840000000
0!
0'
0/
#493850000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#493860000000
0!
0'
0/
#493870000000
1!
1'
1/
#493880000000
0!
0'
0/
#493890000000
1!
1'
1/
#493900000000
0!
0'
0/
#493910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#493920000000
0!
0'
0/
#493930000000
1!
1'
1/
#493940000000
0!
0'
0/
#493950000000
1!
1'
1/
#493960000000
0!
0'
0/
#493970000000
1!
1'
1/
#493980000000
0!
0'
0/
#493990000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#494000000000
0!
0'
0/
#494010000000
1!
1'
1/
#494020000000
0!
0'
0/
#494030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#494040000000
0!
0'
0/
#494050000000
1!
1'
1/
#494060000000
0!
0'
0/
#494070000000
#494080000000
1!
1'
1/
#494090000000
0!
0'
0/
#494100000000
1!
1'
1/
#494110000000
0!
1"
0'
1(
0/
10
#494120000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#494130000000
0!
0'
0/
#494140000000
1!
1'
1/
#494150000000
0!
0'
0/
#494160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#494170000000
0!
0'
0/
#494180000000
1!
1'
1/
#494190000000
0!
1"
0'
1(
0/
10
#494200000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#494210000000
0!
1$
0'
1+
0/
#494220000000
1!
1'
1/
#494230000000
0!
0'
0/
#494240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#494250000000
0!
0'
0/
#494260000000
1!
1'
1/
#494270000000
0!
0'
0/
#494280000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#494290000000
0!
0'
0/
#494300000000
1!
1'
1/
#494310000000
0!
0'
0/
#494320000000
1!
1'
1/
#494330000000
0!
0'
0/
#494340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#494350000000
0!
0'
0/
#494360000000
1!
1'
1/
#494370000000
0!
0'
0/
#494380000000
1!
1'
1/
#494390000000
0!
0'
0/
#494400000000
1!
1'
1/
#494410000000
0!
0'
0/
#494420000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#494430000000
0!
0'
0/
#494440000000
1!
1'
1/
#494450000000
0!
0'
0/
#494460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#494470000000
0!
0'
0/
#494480000000
1!
1'
1/
#494490000000
0!
0'
0/
#494500000000
#494510000000
1!
1'
1/
#494520000000
0!
0'
0/
#494530000000
1!
1'
1/
#494540000000
0!
1"
0'
1(
0/
10
#494550000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#494560000000
0!
0'
0/
#494570000000
1!
1'
1/
#494580000000
0!
0'
0/
#494590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#494600000000
0!
0'
0/
#494610000000
1!
1'
1/
#494620000000
0!
1"
0'
1(
0/
10
#494630000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#494640000000
0!
1$
0'
1+
0/
#494650000000
1!
1'
1/
#494660000000
0!
0'
0/
#494670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#494680000000
0!
0'
0/
#494690000000
1!
1'
1/
#494700000000
0!
0'
0/
#494710000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#494720000000
0!
0'
0/
#494730000000
1!
1'
1/
#494740000000
0!
0'
0/
#494750000000
1!
1'
1/
#494760000000
0!
0'
0/
#494770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#494780000000
0!
0'
0/
#494790000000
1!
1'
1/
#494800000000
0!
0'
0/
#494810000000
1!
1'
1/
#494820000000
0!
0'
0/
#494830000000
1!
1'
1/
#494840000000
0!
0'
0/
#494850000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#494860000000
0!
0'
0/
#494870000000
1!
1'
1/
#494880000000
0!
0'
0/
#494890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#494900000000
0!
0'
0/
#494910000000
1!
1'
1/
#494920000000
0!
0'
0/
#494930000000
#494940000000
1!
1'
1/
#494950000000
0!
0'
0/
#494960000000
1!
1'
1/
#494970000000
0!
1"
0'
1(
0/
10
#494980000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#494990000000
0!
0'
0/
#495000000000
1!
1'
1/
#495010000000
0!
0'
0/
#495020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#495030000000
0!
0'
0/
#495040000000
1!
1'
1/
#495050000000
0!
1"
0'
1(
0/
10
#495060000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#495070000000
0!
1$
0'
1+
0/
#495080000000
1!
1'
1/
#495090000000
0!
0'
0/
#495100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#495110000000
0!
0'
0/
#495120000000
1!
1'
1/
#495130000000
0!
0'
0/
#495140000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#495150000000
0!
0'
0/
#495160000000
1!
1'
1/
#495170000000
0!
0'
0/
#495180000000
1!
1'
1/
#495190000000
0!
0'
0/
#495200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#495210000000
0!
0'
0/
#495220000000
1!
1'
1/
#495230000000
0!
0'
0/
#495240000000
1!
1'
1/
#495250000000
0!
0'
0/
#495260000000
1!
1'
1/
#495270000000
0!
0'
0/
#495280000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#495290000000
0!
0'
0/
#495300000000
1!
1'
1/
#495310000000
0!
0'
0/
#495320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#495330000000
0!
0'
0/
#495340000000
1!
1'
1/
#495350000000
0!
0'
0/
#495360000000
#495370000000
1!
1'
1/
#495380000000
0!
0'
0/
#495390000000
1!
1'
1/
#495400000000
0!
1"
0'
1(
0/
10
#495410000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#495420000000
0!
0'
0/
#495430000000
1!
1'
1/
#495440000000
0!
0'
0/
#495450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#495460000000
0!
0'
0/
#495470000000
1!
1'
1/
#495480000000
0!
1"
0'
1(
0/
10
#495490000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#495500000000
0!
1$
0'
1+
0/
#495510000000
1!
1'
1/
#495520000000
0!
0'
0/
#495530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#495540000000
0!
0'
0/
#495550000000
1!
1'
1/
#495560000000
0!
0'
0/
#495570000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#495580000000
0!
0'
0/
#495590000000
1!
1'
1/
#495600000000
0!
0'
0/
#495610000000
1!
1'
1/
#495620000000
0!
0'
0/
#495630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#495640000000
0!
0'
0/
#495650000000
1!
1'
1/
#495660000000
0!
0'
0/
#495670000000
1!
1'
1/
#495680000000
0!
0'
0/
#495690000000
1!
1'
1/
#495700000000
0!
0'
0/
#495710000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#495720000000
0!
0'
0/
#495730000000
1!
1'
1/
#495740000000
0!
0'
0/
#495750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#495760000000
0!
0'
0/
#495770000000
1!
1'
1/
#495780000000
0!
0'
0/
#495790000000
#495800000000
1!
1'
1/
#495810000000
0!
0'
0/
#495820000000
1!
1'
1/
#495830000000
0!
1"
0'
1(
0/
10
#495840000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#495850000000
0!
0'
0/
#495860000000
1!
1'
1/
#495870000000
0!
0'
0/
#495880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#495890000000
0!
0'
0/
#495900000000
1!
1'
1/
#495910000000
0!
1"
0'
1(
0/
10
#495920000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#495930000000
0!
1$
0'
1+
0/
#495940000000
1!
1'
1/
#495950000000
0!
0'
0/
#495960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#495970000000
0!
0'
0/
#495980000000
1!
1'
1/
#495990000000
0!
0'
0/
#496000000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#496010000000
0!
0'
0/
#496020000000
1!
1'
1/
#496030000000
0!
0'
0/
#496040000000
1!
1'
1/
#496050000000
0!
0'
0/
#496060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#496070000000
0!
0'
0/
#496080000000
1!
1'
1/
#496090000000
0!
0'
0/
#496100000000
1!
1'
1/
#496110000000
0!
0'
0/
#496120000000
1!
1'
1/
#496130000000
0!
0'
0/
#496140000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#496150000000
0!
0'
0/
#496160000000
1!
1'
1/
#496170000000
0!
0'
0/
#496180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#496190000000
0!
0'
0/
#496200000000
1!
1'
1/
#496210000000
0!
0'
0/
#496220000000
#496230000000
1!
1'
1/
#496240000000
0!
0'
0/
#496250000000
1!
1'
1/
#496260000000
0!
1"
0'
1(
0/
10
#496270000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#496280000000
0!
0'
0/
#496290000000
1!
1'
1/
#496300000000
0!
0'
0/
#496310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#496320000000
0!
0'
0/
#496330000000
1!
1'
1/
#496340000000
0!
1"
0'
1(
0/
10
#496350000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#496360000000
0!
1$
0'
1+
0/
#496370000000
1!
1'
1/
#496380000000
0!
0'
0/
#496390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#496400000000
0!
0'
0/
#496410000000
1!
1'
1/
#496420000000
0!
0'
0/
#496430000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#496440000000
0!
0'
0/
#496450000000
1!
1'
1/
#496460000000
0!
0'
0/
#496470000000
1!
1'
1/
#496480000000
0!
0'
0/
#496490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#496500000000
0!
0'
0/
#496510000000
1!
1'
1/
#496520000000
0!
0'
0/
#496530000000
1!
1'
1/
#496540000000
0!
0'
0/
#496550000000
1!
1'
1/
#496560000000
0!
0'
0/
#496570000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#496580000000
0!
0'
0/
#496590000000
1!
1'
1/
#496600000000
0!
0'
0/
#496610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#496620000000
0!
0'
0/
#496630000000
1!
1'
1/
#496640000000
0!
0'
0/
#496650000000
#496660000000
1!
1'
1/
#496670000000
0!
0'
0/
#496680000000
1!
1'
1/
#496690000000
0!
1"
0'
1(
0/
10
#496700000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#496710000000
0!
0'
0/
#496720000000
1!
1'
1/
#496730000000
0!
0'
0/
#496740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#496750000000
0!
0'
0/
#496760000000
1!
1'
1/
#496770000000
0!
1"
0'
1(
0/
10
#496780000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#496790000000
0!
1$
0'
1+
0/
#496800000000
1!
1'
1/
#496810000000
0!
0'
0/
#496820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#496830000000
0!
0'
0/
#496840000000
1!
1'
1/
#496850000000
0!
0'
0/
#496860000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#496870000000
0!
0'
0/
#496880000000
1!
1'
1/
#496890000000
0!
0'
0/
#496900000000
1!
1'
1/
#496910000000
0!
0'
0/
#496920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#496930000000
0!
0'
0/
#496940000000
1!
1'
1/
#496950000000
0!
0'
0/
#496960000000
1!
1'
1/
#496970000000
0!
0'
0/
#496980000000
1!
1'
1/
#496990000000
0!
0'
0/
#497000000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#497010000000
0!
0'
0/
#497020000000
1!
1'
1/
#497030000000
0!
0'
0/
#497040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#497050000000
0!
0'
0/
#497060000000
1!
1'
1/
#497070000000
0!
0'
0/
#497080000000
#497090000000
1!
1'
1/
#497100000000
0!
0'
0/
#497110000000
1!
1'
1/
#497120000000
0!
1"
0'
1(
0/
10
#497130000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#497140000000
0!
0'
0/
#497150000000
1!
1'
1/
#497160000000
0!
0'
0/
#497170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#497180000000
0!
0'
0/
#497190000000
1!
1'
1/
#497200000000
0!
1"
0'
1(
0/
10
#497210000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#497220000000
0!
1$
0'
1+
0/
#497230000000
1!
1'
1/
#497240000000
0!
0'
0/
#497250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#497260000000
0!
0'
0/
#497270000000
1!
1'
1/
#497280000000
0!
0'
0/
#497290000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#497300000000
0!
0'
0/
#497310000000
1!
1'
1/
#497320000000
0!
0'
0/
#497330000000
1!
1'
1/
#497340000000
0!
0'
0/
#497350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#497360000000
0!
0'
0/
#497370000000
1!
1'
1/
#497380000000
0!
0'
0/
#497390000000
1!
1'
1/
#497400000000
0!
0'
0/
#497410000000
1!
1'
1/
#497420000000
0!
0'
0/
#497430000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#497440000000
0!
0'
0/
#497450000000
1!
1'
1/
#497460000000
0!
0'
0/
#497470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#497480000000
0!
0'
0/
#497490000000
1!
1'
1/
#497500000000
0!
0'
0/
#497510000000
#497520000000
1!
1'
1/
#497530000000
0!
0'
0/
#497540000000
1!
1'
1/
#497550000000
0!
1"
0'
1(
0/
10
#497560000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#497570000000
0!
0'
0/
#497580000000
1!
1'
1/
#497590000000
0!
0'
0/
#497600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#497610000000
0!
0'
0/
#497620000000
1!
1'
1/
#497630000000
0!
1"
0'
1(
0/
10
#497640000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#497650000000
0!
1$
0'
1+
0/
#497660000000
1!
1'
1/
#497670000000
0!
0'
0/
#497680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#497690000000
0!
0'
0/
#497700000000
1!
1'
1/
#497710000000
0!
0'
0/
#497720000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#497730000000
0!
0'
0/
#497740000000
1!
1'
1/
#497750000000
0!
0'
0/
#497760000000
1!
1'
1/
#497770000000
0!
0'
0/
#497780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#497790000000
0!
0'
0/
#497800000000
1!
1'
1/
#497810000000
0!
0'
0/
#497820000000
1!
1'
1/
#497830000000
0!
0'
0/
#497840000000
1!
1'
1/
#497850000000
0!
0'
0/
#497860000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#497870000000
0!
0'
0/
#497880000000
1!
1'
1/
#497890000000
0!
0'
0/
#497900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#497910000000
0!
0'
0/
#497920000000
1!
1'
1/
#497930000000
0!
0'
0/
#497940000000
#497950000000
1!
1'
1/
#497960000000
0!
0'
0/
#497970000000
1!
1'
1/
#497980000000
0!
1"
0'
1(
0/
10
#497990000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#498000000000
0!
0'
0/
#498010000000
1!
1'
1/
#498020000000
0!
0'
0/
#498030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#498040000000
0!
0'
0/
#498050000000
1!
1'
1/
#498060000000
0!
1"
0'
1(
0/
10
#498070000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#498080000000
0!
1$
0'
1+
0/
#498090000000
1!
1'
1/
#498100000000
0!
0'
0/
#498110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#498120000000
0!
0'
0/
#498130000000
1!
1'
1/
#498140000000
0!
0'
0/
#498150000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#498160000000
0!
0'
0/
#498170000000
1!
1'
1/
#498180000000
0!
0'
0/
#498190000000
1!
1'
1/
#498200000000
0!
0'
0/
#498210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#498220000000
0!
0'
0/
#498230000000
1!
1'
1/
#498240000000
0!
0'
0/
#498250000000
1!
1'
1/
#498260000000
0!
0'
0/
#498270000000
1!
1'
1/
#498280000000
0!
0'
0/
#498290000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#498300000000
0!
0'
0/
#498310000000
1!
1'
1/
#498320000000
0!
0'
0/
#498330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#498340000000
0!
0'
0/
#498350000000
1!
1'
1/
#498360000000
0!
0'
0/
#498370000000
#498380000000
1!
1'
1/
#498390000000
0!
0'
0/
#498400000000
1!
1'
1/
#498410000000
0!
1"
0'
1(
0/
10
#498420000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#498430000000
0!
0'
0/
#498440000000
1!
1'
1/
#498450000000
0!
0'
0/
#498460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#498470000000
0!
0'
0/
#498480000000
1!
1'
1/
#498490000000
0!
1"
0'
1(
0/
10
#498500000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#498510000000
0!
1$
0'
1+
0/
#498520000000
1!
1'
1/
#498530000000
0!
0'
0/
#498540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#498550000000
0!
0'
0/
#498560000000
1!
1'
1/
#498570000000
0!
0'
0/
#498580000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#498590000000
0!
0'
0/
#498600000000
1!
1'
1/
#498610000000
0!
0'
0/
#498620000000
1!
1'
1/
#498630000000
0!
0'
0/
#498640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#498650000000
0!
0'
0/
#498660000000
1!
1'
1/
#498670000000
0!
0'
0/
#498680000000
1!
1'
1/
#498690000000
0!
0'
0/
#498700000000
1!
1'
1/
#498710000000
0!
0'
0/
#498720000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#498730000000
0!
0'
0/
#498740000000
1!
1'
1/
#498750000000
0!
0'
0/
#498760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#498770000000
0!
0'
0/
#498780000000
1!
1'
1/
#498790000000
0!
0'
0/
#498800000000
#498810000000
1!
1'
1/
#498820000000
0!
0'
0/
#498830000000
1!
1'
1/
#498840000000
0!
1"
0'
1(
0/
10
#498850000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#498860000000
0!
0'
0/
#498870000000
1!
1'
1/
#498880000000
0!
0'
0/
#498890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#498900000000
0!
0'
0/
#498910000000
1!
1'
1/
#498920000000
0!
1"
0'
1(
0/
10
#498930000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#498940000000
0!
1$
0'
1+
0/
#498950000000
1!
1'
1/
#498960000000
0!
0'
0/
#498970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#498980000000
0!
0'
0/
#498990000000
1!
1'
1/
#499000000000
0!
0'
0/
#499010000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#499020000000
0!
0'
0/
#499030000000
1!
1'
1/
#499040000000
0!
0'
0/
#499050000000
1!
1'
1/
#499060000000
0!
0'
0/
#499070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#499080000000
0!
0'
0/
#499090000000
1!
1'
1/
#499100000000
0!
0'
0/
#499110000000
1!
1'
1/
#499120000000
0!
0'
0/
#499130000000
1!
1'
1/
#499140000000
0!
0'
0/
#499150000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#499160000000
0!
0'
0/
#499170000000
1!
1'
1/
#499180000000
0!
0'
0/
#499190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#499200000000
0!
0'
0/
#499210000000
1!
1'
1/
#499220000000
0!
0'
0/
#499230000000
#499240000000
1!
1'
1/
#499250000000
0!
0'
0/
#499260000000
1!
1'
1/
#499270000000
0!
1"
0'
1(
0/
10
#499280000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#499290000000
0!
0'
0/
#499300000000
1!
1'
1/
#499310000000
0!
0'
0/
#499320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#499330000000
0!
0'
0/
#499340000000
1!
1'
1/
#499350000000
0!
1"
0'
1(
0/
10
#499360000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#499370000000
0!
1$
0'
1+
0/
#499380000000
1!
1'
1/
#499390000000
0!
0'
0/
#499400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#499410000000
0!
0'
0/
#499420000000
1!
1'
1/
#499430000000
0!
0'
0/
#499440000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#499450000000
0!
0'
0/
#499460000000
1!
1'
1/
#499470000000
0!
0'
0/
#499480000000
1!
1'
1/
#499490000000
0!
0'
0/
#499500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#499510000000
0!
0'
0/
#499520000000
1!
1'
1/
#499530000000
0!
0'
0/
#499540000000
1!
1'
1/
#499550000000
0!
0'
0/
#499560000000
1!
1'
1/
#499570000000
0!
0'
0/
#499580000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#499590000000
0!
0'
0/
#499600000000
1!
1'
1/
#499610000000
0!
0'
0/
#499620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#499630000000
0!
0'
0/
#499640000000
1!
1'
1/
#499650000000
0!
0'
0/
#499660000000
#499670000000
1!
1'
1/
#499680000000
0!
0'
0/
#499690000000
1!
1'
1/
#499700000000
0!
1"
0'
1(
0/
10
#499710000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#499720000000
0!
0'
0/
#499730000000
1!
1'
1/
#499740000000
0!
0'
0/
#499750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#499760000000
0!
0'
0/
#499770000000
1!
1'
1/
#499780000000
0!
1"
0'
1(
0/
10
#499790000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#499800000000
0!
1$
0'
1+
0/
#499810000000
1!
1'
1/
#499820000000
0!
0'
0/
#499830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#499840000000
0!
0'
0/
#499850000000
1!
1'
1/
#499860000000
0!
0'
0/
#499870000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#499880000000
0!
0'
0/
#499890000000
1!
1'
1/
#499900000000
0!
0'
0/
#499910000000
1!
1'
1/
#499920000000
0!
0'
0/
#499930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#499940000000
0!
0'
0/
#499950000000
1!
1'
1/
#499960000000
0!
0'
0/
#499970000000
1!
1'
1/
#499980000000
0!
0'
0/
#499990000000
1!
1'
1/
#500000000000
0!
0'
0/
#500010000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#500020000000
0!
0'
0/
#500030000000
1!
1'
1/
#500040000000
0!
0'
0/
#500050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#500060000000
0!
0'
0/
#500070000000
1!
1'
1/
#500080000000
0!
0'
0/
#500090000000
#500100000000
1!
1'
1/
#500110000000
0!
0'
0/
#500120000000
1!
1'
1/
#500130000000
0!
1"
0'
1(
0/
10
#500140000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#500150000000
0!
0'
0/
#500160000000
1!
1'
1/
#500170000000
0!
0'
0/
#500180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#500190000000
0!
0'
0/
#500200000000
1!
1'
1/
#500210000000
0!
1"
0'
1(
0/
10
#500220000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#500230000000
0!
1$
0'
1+
0/
#500240000000
1!
1'
1/
#500250000000
0!
0'
0/
#500260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#500270000000
0!
0'
0/
#500280000000
1!
1'
1/
#500290000000
0!
0'
0/
#500300000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#500310000000
0!
0'
0/
#500320000000
1!
1'
1/
#500330000000
0!
0'
0/
#500340000000
1!
1'
1/
#500350000000
0!
0'
0/
#500360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#500370000000
0!
0'
0/
#500380000000
1!
1'
1/
#500390000000
0!
0'
0/
#500400000000
1!
1'
1/
#500410000000
0!
0'
0/
#500420000000
1!
1'
1/
#500430000000
0!
0'
0/
#500440000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#500450000000
0!
0'
0/
#500460000000
1!
1'
1/
#500470000000
0!
0'
0/
#500480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#500490000000
0!
0'
0/
#500500000000
1!
1'
1/
#500510000000
0!
0'
0/
#500520000000
#500530000000
1!
1'
1/
#500540000000
0!
0'
0/
#500550000000
1!
1'
1/
#500560000000
0!
1"
0'
1(
0/
10
#500570000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#500580000000
0!
0'
0/
#500590000000
1!
1'
1/
#500600000000
0!
0'
0/
#500610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#500620000000
0!
0'
0/
#500630000000
1!
1'
1/
#500640000000
0!
1"
0'
1(
0/
10
#500650000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#500660000000
0!
1$
0'
1+
0/
#500670000000
1!
1'
1/
#500680000000
0!
0'
0/
#500690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#500700000000
0!
0'
0/
#500710000000
1!
1'
1/
#500720000000
0!
0'
0/
#500730000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#500740000000
0!
0'
0/
#500750000000
1!
1'
1/
#500760000000
0!
0'
0/
#500770000000
1!
1'
1/
#500780000000
0!
0'
0/
#500790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#500800000000
0!
0'
0/
#500810000000
1!
1'
1/
#500820000000
0!
0'
0/
#500830000000
1!
1'
1/
#500840000000
0!
0'
0/
#500850000000
1!
1'
1/
#500860000000
0!
0'
0/
#500870000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#500880000000
0!
0'
0/
#500890000000
1!
1'
1/
#500900000000
0!
0'
0/
#500910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#500920000000
0!
0'
0/
#500930000000
1!
1'
1/
#500940000000
0!
0'
0/
#500950000000
#500960000000
1!
1'
1/
#500970000000
0!
0'
0/
#500980000000
1!
1'
1/
#500990000000
0!
1"
0'
1(
0/
10
#501000000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#501010000000
0!
0'
0/
#501020000000
1!
1'
1/
#501030000000
0!
0'
0/
#501040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#501050000000
0!
0'
0/
#501060000000
1!
1'
1/
#501070000000
0!
1"
0'
1(
0/
10
#501080000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#501090000000
0!
1$
0'
1+
0/
#501100000000
1!
1'
1/
#501110000000
0!
0'
0/
#501120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#501130000000
0!
0'
0/
#501140000000
1!
1'
1/
#501150000000
0!
0'
0/
#501160000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#501170000000
0!
0'
0/
#501180000000
1!
1'
1/
#501190000000
0!
0'
0/
#501200000000
1!
1'
1/
#501210000000
0!
0'
0/
#501220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#501230000000
0!
0'
0/
#501240000000
1!
1'
1/
#501250000000
0!
0'
0/
#501260000000
1!
1'
1/
#501270000000
0!
0'
0/
#501280000000
1!
1'
1/
#501290000000
0!
0'
0/
#501300000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#501310000000
0!
0'
0/
#501320000000
1!
1'
1/
#501330000000
0!
0'
0/
#501340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#501350000000
0!
0'
0/
#501360000000
1!
1'
1/
#501370000000
0!
0'
0/
#501380000000
#501390000000
1!
1'
1/
#501400000000
0!
0'
0/
#501410000000
1!
1'
1/
#501420000000
0!
1"
0'
1(
0/
10
#501430000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#501440000000
0!
0'
0/
#501450000000
1!
1'
1/
#501460000000
0!
0'
0/
#501470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#501480000000
0!
0'
0/
#501490000000
1!
1'
1/
#501500000000
0!
1"
0'
1(
0/
10
#501510000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#501520000000
0!
1$
0'
1+
0/
#501530000000
1!
1'
1/
#501540000000
0!
0'
0/
#501550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#501560000000
0!
0'
0/
#501570000000
1!
1'
1/
#501580000000
0!
0'
0/
#501590000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#501600000000
0!
0'
0/
#501610000000
1!
1'
1/
#501620000000
0!
0'
0/
#501630000000
1!
1'
1/
#501640000000
0!
0'
0/
#501650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#501660000000
0!
0'
0/
#501670000000
1!
1'
1/
#501680000000
0!
0'
0/
#501690000000
1!
1'
1/
#501700000000
0!
0'
0/
#501710000000
1!
1'
1/
#501720000000
0!
0'
0/
#501730000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#501740000000
0!
0'
0/
#501750000000
1!
1'
1/
#501760000000
0!
0'
0/
#501770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#501780000000
0!
0'
0/
#501790000000
1!
1'
1/
#501800000000
0!
0'
0/
#501810000000
#501820000000
1!
1'
1/
#501830000000
0!
0'
0/
#501840000000
1!
1'
1/
#501850000000
0!
1"
0'
1(
0/
10
#501860000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#501870000000
0!
0'
0/
#501880000000
1!
1'
1/
#501890000000
0!
0'
0/
#501900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#501910000000
0!
0'
0/
#501920000000
1!
1'
1/
#501930000000
0!
1"
0'
1(
0/
10
#501940000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#501950000000
0!
1$
0'
1+
0/
#501960000000
1!
1'
1/
#501970000000
0!
0'
0/
#501980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#501990000000
0!
0'
0/
#502000000000
1!
1'
1/
#502010000000
0!
0'
0/
#502020000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#502030000000
0!
0'
0/
#502040000000
1!
1'
1/
#502050000000
0!
0'
0/
#502060000000
1!
1'
1/
#502070000000
0!
0'
0/
#502080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#502090000000
0!
0'
0/
#502100000000
1!
1'
1/
#502110000000
0!
0'
0/
#502120000000
1!
1'
1/
#502130000000
0!
0'
0/
#502140000000
1!
1'
1/
#502150000000
0!
0'
0/
#502160000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#502170000000
0!
0'
0/
#502180000000
1!
1'
1/
#502190000000
0!
0'
0/
#502200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#502210000000
0!
0'
0/
#502220000000
1!
1'
1/
#502230000000
0!
0'
0/
#502240000000
#502250000000
1!
1'
1/
#502260000000
0!
0'
0/
#502270000000
1!
1'
1/
#502280000000
0!
1"
0'
1(
0/
10
#502290000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#502300000000
0!
0'
0/
#502310000000
1!
1'
1/
#502320000000
0!
0'
0/
#502330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#502340000000
0!
0'
0/
#502350000000
1!
1'
1/
#502360000000
0!
1"
0'
1(
0/
10
#502370000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#502380000000
0!
1$
0'
1+
0/
#502390000000
1!
1'
1/
#502400000000
0!
0'
0/
#502410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#502420000000
0!
0'
0/
#502430000000
1!
1'
1/
#502440000000
0!
0'
0/
#502450000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#502460000000
0!
0'
0/
#502470000000
1!
1'
1/
#502480000000
0!
0'
0/
#502490000000
1!
1'
1/
#502500000000
0!
0'
0/
#502510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#502520000000
0!
0'
0/
#502530000000
1!
1'
1/
#502540000000
0!
0'
0/
#502550000000
1!
1'
1/
#502560000000
0!
0'
0/
#502570000000
1!
1'
1/
#502580000000
0!
0'
0/
#502590000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#502600000000
0!
0'
0/
#502610000000
1!
1'
1/
#502620000000
0!
0'
0/
#502630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#502640000000
0!
0'
0/
#502650000000
1!
1'
1/
#502660000000
0!
0'
0/
#502670000000
#502680000000
1!
1'
1/
#502690000000
0!
0'
0/
#502700000000
1!
1'
1/
#502710000000
0!
1"
0'
1(
0/
10
#502720000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#502730000000
0!
0'
0/
#502740000000
1!
1'
1/
#502750000000
0!
0'
0/
#502760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#502770000000
0!
0'
0/
#502780000000
1!
1'
1/
#502790000000
0!
1"
0'
1(
0/
10
#502800000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#502810000000
0!
1$
0'
1+
0/
#502820000000
1!
1'
1/
#502830000000
0!
0'
0/
#502840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#502850000000
0!
0'
0/
#502860000000
1!
1'
1/
#502870000000
0!
0'
0/
#502880000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#502890000000
0!
0'
0/
#502900000000
1!
1'
1/
#502910000000
0!
0'
0/
#502920000000
1!
1'
1/
#502930000000
0!
0'
0/
#502940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#502950000000
0!
0'
0/
#502960000000
1!
1'
1/
#502970000000
0!
0'
0/
#502980000000
1!
1'
1/
#502990000000
0!
0'
0/
#503000000000
1!
1'
1/
#503010000000
0!
0'
0/
#503020000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#503030000000
0!
0'
0/
#503040000000
1!
1'
1/
#503050000000
0!
0'
0/
#503060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#503070000000
0!
0'
0/
#503080000000
1!
1'
1/
#503090000000
0!
0'
0/
#503100000000
#503110000000
1!
1'
1/
#503120000000
0!
0'
0/
#503130000000
1!
1'
1/
#503140000000
0!
1"
0'
1(
0/
10
#503150000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#503160000000
0!
0'
0/
#503170000000
1!
1'
1/
#503180000000
0!
0'
0/
#503190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#503200000000
0!
0'
0/
#503210000000
1!
1'
1/
#503220000000
0!
1"
0'
1(
0/
10
#503230000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#503240000000
0!
1$
0'
1+
0/
#503250000000
1!
1'
1/
#503260000000
0!
0'
0/
#503270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#503280000000
0!
0'
0/
#503290000000
1!
1'
1/
#503300000000
0!
0'
0/
#503310000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#503320000000
0!
0'
0/
#503330000000
1!
1'
1/
#503340000000
0!
0'
0/
#503350000000
1!
1'
1/
#503360000000
0!
0'
0/
#503370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#503380000000
0!
0'
0/
#503390000000
1!
1'
1/
#503400000000
0!
0'
0/
#503410000000
1!
1'
1/
#503420000000
0!
0'
0/
#503430000000
1!
1'
1/
#503440000000
0!
0'
0/
#503450000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#503460000000
0!
0'
0/
#503470000000
1!
1'
1/
#503480000000
0!
0'
0/
#503490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#503500000000
0!
0'
0/
#503510000000
1!
1'
1/
#503520000000
0!
0'
0/
#503530000000
#503540000000
1!
1'
1/
#503550000000
0!
0'
0/
#503560000000
1!
1'
1/
#503570000000
0!
1"
0'
1(
0/
10
#503580000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#503590000000
0!
0'
0/
#503600000000
1!
1'
1/
#503610000000
0!
0'
0/
#503620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#503630000000
0!
0'
0/
#503640000000
1!
1'
1/
#503650000000
0!
1"
0'
1(
0/
10
#503660000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#503670000000
0!
1$
0'
1+
0/
#503680000000
1!
1'
1/
#503690000000
0!
0'
0/
#503700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#503710000000
0!
0'
0/
#503720000000
1!
1'
1/
#503730000000
0!
0'
0/
#503740000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#503750000000
0!
0'
0/
#503760000000
1!
1'
1/
#503770000000
0!
0'
0/
#503780000000
1!
1'
1/
#503790000000
0!
0'
0/
#503800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#503810000000
0!
0'
0/
#503820000000
1!
1'
1/
#503830000000
0!
0'
0/
#503840000000
1!
1'
1/
#503850000000
0!
0'
0/
#503860000000
1!
1'
1/
#503870000000
0!
0'
0/
#503880000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#503890000000
0!
0'
0/
#503900000000
1!
1'
1/
#503910000000
0!
0'
0/
#503920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#503930000000
0!
0'
0/
#503940000000
1!
1'
1/
#503950000000
0!
0'
0/
#503960000000
#503970000000
1!
1'
1/
#503980000000
0!
0'
0/
#503990000000
1!
1'
1/
#504000000000
0!
1"
0'
1(
0/
10
#504010000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#504020000000
0!
0'
0/
#504030000000
1!
1'
1/
#504040000000
0!
0'
0/
#504050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#504060000000
0!
0'
0/
#504070000000
1!
1'
1/
#504080000000
0!
1"
0'
1(
0/
10
#504090000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#504100000000
0!
1$
0'
1+
0/
#504110000000
1!
1'
1/
#504120000000
0!
0'
0/
#504130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#504140000000
0!
0'
0/
#504150000000
1!
1'
1/
#504160000000
0!
0'
0/
#504170000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#504180000000
0!
0'
0/
#504190000000
1!
1'
1/
#504200000000
0!
0'
0/
#504210000000
1!
1'
1/
#504220000000
0!
0'
0/
#504230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#504240000000
0!
0'
0/
#504250000000
1!
1'
1/
#504260000000
0!
0'
0/
#504270000000
1!
1'
1/
#504280000000
0!
0'
0/
#504290000000
1!
1'
1/
#504300000000
0!
0'
0/
#504310000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#504320000000
0!
0'
0/
#504330000000
1!
1'
1/
#504340000000
0!
0'
0/
#504350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#504360000000
0!
0'
0/
#504370000000
1!
1'
1/
#504380000000
0!
0'
0/
#504390000000
#504400000000
1!
1'
1/
#504410000000
0!
0'
0/
#504420000000
1!
1'
1/
#504430000000
0!
1"
0'
1(
0/
10
#504440000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#504450000000
0!
0'
0/
#504460000000
1!
1'
1/
#504470000000
0!
0'
0/
#504480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#504490000000
0!
0'
0/
#504500000000
1!
1'
1/
#504510000000
0!
1"
0'
1(
0/
10
#504520000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#504530000000
0!
1$
0'
1+
0/
#504540000000
1!
1'
1/
#504550000000
0!
0'
0/
#504560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#504570000000
0!
0'
0/
#504580000000
1!
1'
1/
#504590000000
0!
0'
0/
#504600000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#504610000000
0!
0'
0/
#504620000000
1!
1'
1/
#504630000000
0!
0'
0/
#504640000000
1!
1'
1/
#504650000000
0!
0'
0/
#504660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#504670000000
0!
0'
0/
#504680000000
1!
1'
1/
#504690000000
0!
0'
0/
#504700000000
1!
1'
1/
#504710000000
0!
0'
0/
#504720000000
1!
1'
1/
#504730000000
0!
0'
0/
#504740000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#504750000000
0!
0'
0/
#504760000000
1!
1'
1/
#504770000000
0!
0'
0/
#504780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#504790000000
0!
0'
0/
#504800000000
1!
1'
1/
#504810000000
0!
0'
0/
#504820000000
#504830000000
1!
1'
1/
#504840000000
0!
0'
0/
#504850000000
1!
1'
1/
#504860000000
0!
1"
0'
1(
0/
10
#504870000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#504880000000
0!
0'
0/
#504890000000
1!
1'
1/
#504900000000
0!
0'
0/
#504910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#504920000000
0!
0'
0/
#504930000000
1!
1'
1/
#504940000000
0!
1"
0'
1(
0/
10
#504950000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#504960000000
0!
1$
0'
1+
0/
#504970000000
1!
1'
1/
#504980000000
0!
0'
0/
#504990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#505000000000
0!
0'
0/
#505010000000
1!
1'
1/
#505020000000
0!
0'
0/
#505030000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#505040000000
0!
0'
0/
#505050000000
1!
1'
1/
#505060000000
0!
0'
0/
#505070000000
1!
1'
1/
#505080000000
0!
0'
0/
#505090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#505100000000
0!
0'
0/
#505110000000
1!
1'
1/
#505120000000
0!
0'
0/
#505130000000
1!
1'
1/
#505140000000
0!
0'
0/
#505150000000
1!
1'
1/
#505160000000
0!
0'
0/
#505170000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#505180000000
0!
0'
0/
#505190000000
1!
1'
1/
#505200000000
0!
0'
0/
#505210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#505220000000
0!
0'
0/
#505230000000
1!
1'
1/
#505240000000
0!
0'
0/
#505250000000
#505260000000
1!
1'
1/
#505270000000
0!
0'
0/
#505280000000
1!
1'
1/
#505290000000
0!
1"
0'
1(
0/
10
#505300000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#505310000000
0!
0'
0/
#505320000000
1!
1'
1/
#505330000000
0!
0'
0/
#505340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#505350000000
0!
0'
0/
#505360000000
1!
1'
1/
#505370000000
0!
1"
0'
1(
0/
10
#505380000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#505390000000
0!
1$
0'
1+
0/
#505400000000
1!
1'
1/
#505410000000
0!
0'
0/
#505420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#505430000000
0!
0'
0/
#505440000000
1!
1'
1/
#505450000000
0!
0'
0/
#505460000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#505470000000
0!
0'
0/
#505480000000
1!
1'
1/
#505490000000
0!
0'
0/
#505500000000
1!
1'
1/
#505510000000
0!
0'
0/
#505520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#505530000000
0!
0'
0/
#505540000000
1!
1'
1/
#505550000000
0!
0'
0/
#505560000000
1!
1'
1/
#505570000000
0!
0'
0/
#505580000000
1!
1'
1/
#505590000000
0!
0'
0/
#505600000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#505610000000
0!
0'
0/
#505620000000
1!
1'
1/
#505630000000
0!
0'
0/
#505640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#505650000000
0!
0'
0/
#505660000000
1!
1'
1/
#505670000000
0!
0'
0/
#505680000000
#505690000000
1!
1'
1/
#505700000000
0!
0'
0/
#505710000000
1!
1'
1/
#505720000000
0!
1"
0'
1(
0/
10
#505730000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#505740000000
0!
0'
0/
#505750000000
1!
1'
1/
#505760000000
0!
0'
0/
#505770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#505780000000
0!
0'
0/
#505790000000
1!
1'
1/
#505800000000
0!
1"
0'
1(
0/
10
#505810000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#505820000000
0!
1$
0'
1+
0/
#505830000000
1!
1'
1/
#505840000000
0!
0'
0/
#505850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#505860000000
0!
0'
0/
#505870000000
1!
1'
1/
#505880000000
0!
0'
0/
#505890000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#505900000000
0!
0'
0/
#505910000000
1!
1'
1/
#505920000000
0!
0'
0/
#505930000000
1!
1'
1/
#505940000000
0!
0'
0/
#505950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#505960000000
0!
0'
0/
#505970000000
1!
1'
1/
#505980000000
0!
0'
0/
#505990000000
1!
1'
1/
#506000000000
0!
0'
0/
#506010000000
1!
1'
1/
#506020000000
0!
0'
0/
#506030000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#506040000000
0!
0'
0/
#506050000000
1!
1'
1/
#506060000000
0!
0'
0/
#506070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#506080000000
0!
0'
0/
#506090000000
1!
1'
1/
#506100000000
0!
0'
0/
#506110000000
#506120000000
1!
1'
1/
#506130000000
0!
0'
0/
#506140000000
1!
1'
1/
#506150000000
0!
1"
0'
1(
0/
10
#506160000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#506170000000
0!
0'
0/
#506180000000
1!
1'
1/
#506190000000
0!
0'
0/
#506200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#506210000000
0!
0'
0/
#506220000000
1!
1'
1/
#506230000000
0!
1"
0'
1(
0/
10
#506240000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#506250000000
0!
1$
0'
1+
0/
#506260000000
1!
1'
1/
#506270000000
0!
0'
0/
#506280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#506290000000
0!
0'
0/
#506300000000
1!
1'
1/
#506310000000
0!
0'
0/
#506320000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#506330000000
0!
0'
0/
#506340000000
1!
1'
1/
#506350000000
0!
0'
0/
#506360000000
1!
1'
1/
#506370000000
0!
0'
0/
#506380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#506390000000
0!
0'
0/
#506400000000
1!
1'
1/
#506410000000
0!
0'
0/
#506420000000
1!
1'
1/
#506430000000
0!
0'
0/
#506440000000
1!
1'
1/
#506450000000
0!
0'
0/
#506460000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#506470000000
0!
0'
0/
#506480000000
1!
1'
1/
#506490000000
0!
0'
0/
#506500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#506510000000
0!
0'
0/
#506520000000
1!
1'
1/
#506530000000
0!
0'
0/
#506540000000
#506550000000
1!
1'
1/
#506560000000
0!
0'
0/
#506570000000
1!
1'
1/
#506580000000
0!
1"
0'
1(
0/
10
#506590000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#506600000000
0!
0'
0/
#506610000000
1!
1'
1/
#506620000000
0!
0'
0/
#506630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#506640000000
0!
0'
0/
#506650000000
1!
1'
1/
#506660000000
0!
1"
0'
1(
0/
10
#506670000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#506680000000
0!
1$
0'
1+
0/
#506690000000
1!
1'
1/
#506700000000
0!
0'
0/
#506710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#506720000000
0!
0'
0/
#506730000000
1!
1'
1/
#506740000000
0!
0'
0/
#506750000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#506760000000
0!
0'
0/
#506770000000
1!
1'
1/
#506780000000
0!
0'
0/
#506790000000
1!
1'
1/
#506800000000
0!
0'
0/
#506810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#506820000000
0!
0'
0/
#506830000000
1!
1'
1/
#506840000000
0!
0'
0/
#506850000000
1!
1'
1/
#506860000000
0!
0'
0/
#506870000000
1!
1'
1/
#506880000000
0!
0'
0/
#506890000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#506900000000
0!
0'
0/
#506910000000
1!
1'
1/
#506920000000
0!
0'
0/
#506930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#506940000000
0!
0'
0/
#506950000000
1!
1'
1/
#506960000000
0!
0'
0/
#506970000000
#506980000000
1!
1'
1/
#506990000000
0!
0'
0/
#507000000000
1!
1'
1/
#507010000000
0!
1"
0'
1(
0/
10
#507020000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#507030000000
0!
0'
0/
#507040000000
1!
1'
1/
#507050000000
0!
0'
0/
#507060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#507070000000
0!
0'
0/
#507080000000
1!
1'
1/
#507090000000
0!
1"
0'
1(
0/
10
#507100000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#507110000000
0!
1$
0'
1+
0/
#507120000000
1!
1'
1/
#507130000000
0!
0'
0/
#507140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#507150000000
0!
0'
0/
#507160000000
1!
1'
1/
#507170000000
0!
0'
0/
#507180000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#507190000000
0!
0'
0/
#507200000000
1!
1'
1/
#507210000000
0!
0'
0/
#507220000000
1!
1'
1/
#507230000000
0!
0'
0/
#507240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#507250000000
0!
0'
0/
#507260000000
1!
1'
1/
#507270000000
0!
0'
0/
#507280000000
1!
1'
1/
#507290000000
0!
0'
0/
#507300000000
1!
1'
1/
#507310000000
0!
0'
0/
#507320000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#507330000000
0!
0'
0/
#507340000000
1!
1'
1/
#507350000000
0!
0'
0/
#507360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#507370000000
0!
0'
0/
#507380000000
1!
1'
1/
#507390000000
0!
0'
0/
#507400000000
#507410000000
1!
1'
1/
#507420000000
0!
0'
0/
#507430000000
1!
1'
1/
#507440000000
0!
1"
0'
1(
0/
10
#507450000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#507460000000
0!
0'
0/
#507470000000
1!
1'
1/
#507480000000
0!
0'
0/
#507490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#507500000000
0!
0'
0/
#507510000000
1!
1'
1/
#507520000000
0!
1"
0'
1(
0/
10
#507530000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#507540000000
0!
1$
0'
1+
0/
#507550000000
1!
1'
1/
#507560000000
0!
0'
0/
#507570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#507580000000
0!
0'
0/
#507590000000
1!
1'
1/
#507600000000
0!
0'
0/
#507610000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#507620000000
0!
0'
0/
#507630000000
1!
1'
1/
#507640000000
0!
0'
0/
#507650000000
1!
1'
1/
#507660000000
0!
0'
0/
#507670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#507680000000
0!
0'
0/
#507690000000
1!
1'
1/
#507700000000
0!
0'
0/
#507710000000
1!
1'
1/
#507720000000
0!
0'
0/
#507730000000
1!
1'
1/
#507740000000
0!
0'
0/
#507750000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#507760000000
0!
0'
0/
#507770000000
1!
1'
1/
#507780000000
0!
0'
0/
#507790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#507800000000
0!
0'
0/
#507810000000
1!
1'
1/
#507820000000
0!
0'
0/
#507830000000
#507840000000
1!
1'
1/
#507850000000
0!
0'
0/
#507860000000
1!
1'
1/
#507870000000
0!
1"
0'
1(
0/
10
#507880000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#507890000000
0!
0'
0/
#507900000000
1!
1'
1/
#507910000000
0!
0'
0/
#507920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#507930000000
0!
0'
0/
#507940000000
1!
1'
1/
#507950000000
0!
1"
0'
1(
0/
10
#507960000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#507970000000
0!
1$
0'
1+
0/
#507980000000
1!
1'
1/
#507990000000
0!
0'
0/
#508000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#508010000000
0!
0'
0/
#508020000000
1!
1'
1/
#508030000000
0!
0'
0/
#508040000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#508050000000
0!
0'
0/
#508060000000
1!
1'
1/
#508070000000
0!
0'
0/
#508080000000
1!
1'
1/
#508090000000
0!
0'
0/
#508100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#508110000000
0!
0'
0/
#508120000000
1!
1'
1/
#508130000000
0!
0'
0/
#508140000000
1!
1'
1/
#508150000000
0!
0'
0/
#508160000000
1!
1'
1/
#508170000000
0!
0'
0/
#508180000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#508190000000
0!
0'
0/
#508200000000
1!
1'
1/
#508210000000
0!
0'
0/
#508220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#508230000000
0!
0'
0/
#508240000000
1!
1'
1/
#508250000000
0!
0'
0/
#508260000000
#508270000000
1!
1'
1/
#508280000000
0!
0'
0/
#508290000000
1!
1'
1/
#508300000000
0!
1"
0'
1(
0/
10
#508310000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#508320000000
0!
0'
0/
#508330000000
1!
1'
1/
#508340000000
0!
0'
0/
#508350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#508360000000
0!
0'
0/
#508370000000
1!
1'
1/
#508380000000
0!
1"
0'
1(
0/
10
#508390000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#508400000000
0!
1$
0'
1+
0/
#508410000000
1!
1'
1/
#508420000000
0!
0'
0/
#508430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#508440000000
0!
0'
0/
#508450000000
1!
1'
1/
#508460000000
0!
0'
0/
#508470000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#508480000000
0!
0'
0/
#508490000000
1!
1'
1/
#508500000000
0!
0'
0/
#508510000000
1!
1'
1/
#508520000000
0!
0'
0/
#508530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#508540000000
0!
0'
0/
#508550000000
1!
1'
1/
#508560000000
0!
0'
0/
#508570000000
1!
1'
1/
#508580000000
0!
0'
0/
#508590000000
1!
1'
1/
#508600000000
0!
0'
0/
#508610000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#508620000000
0!
0'
0/
#508630000000
1!
1'
1/
#508640000000
0!
0'
0/
#508650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#508660000000
0!
0'
0/
#508670000000
1!
1'
1/
#508680000000
0!
0'
0/
#508690000000
#508700000000
1!
1'
1/
#508710000000
0!
0'
0/
#508720000000
1!
1'
1/
#508730000000
0!
1"
0'
1(
0/
10
#508740000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#508750000000
0!
0'
0/
#508760000000
1!
1'
1/
#508770000000
0!
0'
0/
#508780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#508790000000
0!
0'
0/
#508800000000
1!
1'
1/
#508810000000
0!
1"
0'
1(
0/
10
#508820000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#508830000000
0!
1$
0'
1+
0/
#508840000000
1!
1'
1/
#508850000000
0!
0'
0/
#508860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#508870000000
0!
0'
0/
#508880000000
1!
1'
1/
#508890000000
0!
0'
0/
#508900000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#508910000000
0!
0'
0/
#508920000000
1!
1'
1/
#508930000000
0!
0'
0/
#508940000000
1!
1'
1/
#508950000000
0!
0'
0/
#508960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#508970000000
0!
0'
0/
#508980000000
1!
1'
1/
#508990000000
0!
0'
0/
#509000000000
1!
1'
1/
#509010000000
0!
0'
0/
#509020000000
1!
1'
1/
#509030000000
0!
0'
0/
#509040000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#509050000000
0!
0'
0/
#509060000000
1!
1'
1/
#509070000000
0!
0'
0/
#509080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#509090000000
0!
0'
0/
#509100000000
1!
1'
1/
#509110000000
0!
0'
0/
#509120000000
#509130000000
1!
1'
1/
#509140000000
0!
0'
0/
#509150000000
1!
1'
1/
#509160000000
0!
1"
0'
1(
0/
10
#509170000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#509180000000
0!
0'
0/
#509190000000
1!
1'
1/
#509200000000
0!
0'
0/
#509210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#509220000000
0!
0'
0/
#509230000000
1!
1'
1/
#509240000000
0!
1"
0'
1(
0/
10
#509250000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#509260000000
0!
1$
0'
1+
0/
#509270000000
1!
1'
1/
#509280000000
0!
0'
0/
#509290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#509300000000
0!
0'
0/
#509310000000
1!
1'
1/
#509320000000
0!
0'
0/
#509330000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#509340000000
0!
0'
0/
#509350000000
1!
1'
1/
#509360000000
0!
0'
0/
#509370000000
1!
1'
1/
#509380000000
0!
0'
0/
#509390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#509400000000
0!
0'
0/
#509410000000
1!
1'
1/
#509420000000
0!
0'
0/
#509430000000
1!
1'
1/
#509440000000
0!
0'
0/
#509450000000
1!
1'
1/
#509460000000
0!
0'
0/
#509470000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#509480000000
0!
0'
0/
#509490000000
1!
1'
1/
#509500000000
0!
0'
0/
#509510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#509520000000
0!
0'
0/
#509530000000
1!
1'
1/
#509540000000
0!
0'
0/
#509550000000
#509560000000
1!
1'
1/
#509570000000
0!
0'
0/
#509580000000
1!
1'
1/
#509590000000
0!
1"
0'
1(
0/
10
#509600000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#509610000000
0!
0'
0/
#509620000000
1!
1'
1/
#509630000000
0!
0'
0/
#509640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#509650000000
0!
0'
0/
#509660000000
1!
1'
1/
#509670000000
0!
1"
0'
1(
0/
10
#509680000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#509690000000
0!
1$
0'
1+
0/
#509700000000
1!
1'
1/
#509710000000
0!
0'
0/
#509720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#509730000000
0!
0'
0/
#509740000000
1!
1'
1/
#509750000000
0!
0'
0/
#509760000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#509770000000
0!
0'
0/
#509780000000
1!
1'
1/
#509790000000
0!
0'
0/
#509800000000
1!
1'
1/
#509810000000
0!
0'
0/
#509820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#509830000000
0!
0'
0/
#509840000000
1!
1'
1/
#509850000000
0!
0'
0/
#509860000000
1!
1'
1/
#509870000000
0!
0'
0/
#509880000000
1!
1'
1/
#509890000000
0!
0'
0/
#509900000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#509910000000
0!
0'
0/
#509920000000
1!
1'
1/
#509930000000
0!
0'
0/
#509940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#509950000000
0!
0'
0/
#509960000000
1!
1'
1/
#509970000000
0!
0'
0/
#509980000000
#509990000000
1!
1'
1/
#510000000000
0!
0'
0/
#510010000000
1!
1'
1/
#510020000000
0!
1"
0'
1(
0/
10
#510030000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#510040000000
0!
0'
0/
#510050000000
1!
1'
1/
#510060000000
0!
0'
0/
#510070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#510080000000
0!
0'
0/
#510090000000
1!
1'
1/
#510100000000
0!
1"
0'
1(
0/
10
#510110000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#510120000000
0!
1$
0'
1+
0/
#510130000000
1!
1'
1/
#510140000000
0!
0'
0/
#510150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#510160000000
0!
0'
0/
#510170000000
1!
1'
1/
#510180000000
0!
0'
0/
#510190000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#510200000000
0!
0'
0/
#510210000000
1!
1'
1/
#510220000000
0!
0'
0/
#510230000000
1!
1'
1/
#510240000000
0!
0'
0/
#510250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#510260000000
0!
0'
0/
#510270000000
1!
1'
1/
#510280000000
0!
0'
0/
#510290000000
1!
1'
1/
#510300000000
0!
0'
0/
#510310000000
1!
1'
1/
#510320000000
0!
0'
0/
#510330000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#510340000000
0!
0'
0/
#510350000000
1!
1'
1/
#510360000000
0!
0'
0/
#510370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#510380000000
0!
0'
0/
#510390000000
1!
1'
1/
#510400000000
0!
0'
0/
#510410000000
#510420000000
1!
1'
1/
#510430000000
0!
0'
0/
#510440000000
1!
1'
1/
#510450000000
0!
1"
0'
1(
0/
10
#510460000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#510470000000
0!
0'
0/
#510480000000
1!
1'
1/
#510490000000
0!
0'
0/
#510500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#510510000000
0!
0'
0/
#510520000000
1!
1'
1/
#510530000000
0!
1"
0'
1(
0/
10
#510540000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#510550000000
0!
1$
0'
1+
0/
#510560000000
1!
1'
1/
#510570000000
0!
0'
0/
#510580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#510590000000
0!
0'
0/
#510600000000
1!
1'
1/
#510610000000
0!
0'
0/
#510620000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#510630000000
0!
0'
0/
#510640000000
1!
1'
1/
#510650000000
0!
0'
0/
#510660000000
1!
1'
1/
#510670000000
0!
0'
0/
#510680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#510690000000
0!
0'
0/
#510700000000
1!
1'
1/
#510710000000
0!
0'
0/
#510720000000
1!
1'
1/
#510730000000
0!
0'
0/
#510740000000
1!
1'
1/
#510750000000
0!
0'
0/
#510760000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#510770000000
0!
0'
0/
#510780000000
1!
1'
1/
#510790000000
0!
0'
0/
#510800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#510810000000
0!
0'
0/
#510820000000
1!
1'
1/
#510830000000
0!
0'
0/
#510840000000
#510850000000
1!
1'
1/
#510860000000
0!
0'
0/
#510870000000
1!
1'
1/
#510880000000
0!
1"
0'
1(
0/
10
#510890000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#510900000000
0!
0'
0/
#510910000000
1!
1'
1/
#510920000000
0!
0'
0/
#510930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#510940000000
0!
0'
0/
#510950000000
1!
1'
1/
#510960000000
0!
1"
0'
1(
0/
10
#510970000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#510980000000
0!
1$
0'
1+
0/
#510990000000
1!
1'
1/
#511000000000
0!
0'
0/
#511010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#511020000000
0!
0'
0/
#511030000000
1!
1'
1/
#511040000000
0!
0'
0/
#511050000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#511060000000
0!
0'
0/
#511070000000
1!
1'
1/
#511080000000
0!
0'
0/
#511090000000
1!
1'
1/
#511100000000
0!
0'
0/
#511110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#511120000000
0!
0'
0/
#511130000000
1!
1'
1/
#511140000000
0!
0'
0/
#511150000000
1!
1'
1/
#511160000000
0!
0'
0/
#511170000000
1!
1'
1/
#511180000000
0!
0'
0/
#511190000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#511200000000
0!
0'
0/
#511210000000
1!
1'
1/
#511220000000
0!
0'
0/
#511230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#511240000000
0!
0'
0/
#511250000000
1!
1'
1/
#511260000000
0!
0'
0/
#511270000000
#511280000000
1!
1'
1/
#511290000000
0!
0'
0/
#511300000000
1!
1'
1/
#511310000000
0!
1"
0'
1(
0/
10
#511320000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#511330000000
0!
0'
0/
#511340000000
1!
1'
1/
#511350000000
0!
0'
0/
#511360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#511370000000
0!
0'
0/
#511380000000
1!
1'
1/
#511390000000
0!
1"
0'
1(
0/
10
#511400000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#511410000000
0!
1$
0'
1+
0/
#511420000000
1!
1'
1/
#511430000000
0!
0'
0/
#511440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#511450000000
0!
0'
0/
#511460000000
1!
1'
1/
#511470000000
0!
0'
0/
#511480000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#511490000000
0!
0'
0/
#511500000000
1!
1'
1/
#511510000000
0!
0'
0/
#511520000000
1!
1'
1/
#511530000000
0!
0'
0/
#511540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#511550000000
0!
0'
0/
#511560000000
1!
1'
1/
#511570000000
0!
0'
0/
#511580000000
1!
1'
1/
#511590000000
0!
0'
0/
#511600000000
1!
1'
1/
#511610000000
0!
0'
0/
#511620000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#511630000000
0!
0'
0/
#511640000000
1!
1'
1/
#511650000000
0!
0'
0/
#511660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#511670000000
0!
0'
0/
#511680000000
1!
1'
1/
#511690000000
0!
0'
0/
#511700000000
#511710000000
1!
1'
1/
#511720000000
0!
0'
0/
#511730000000
1!
1'
1/
#511740000000
0!
1"
0'
1(
0/
10
#511750000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#511760000000
0!
0'
0/
#511770000000
1!
1'
1/
#511780000000
0!
0'
0/
#511790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#511800000000
0!
0'
0/
#511810000000
1!
1'
1/
#511820000000
0!
1"
0'
1(
0/
10
#511830000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#511840000000
0!
1$
0'
1+
0/
#511850000000
1!
1'
1/
#511860000000
0!
0'
0/
#511870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#511880000000
0!
0'
0/
#511890000000
1!
1'
1/
#511900000000
0!
0'
0/
#511910000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#511920000000
0!
0'
0/
#511930000000
1!
1'
1/
#511940000000
0!
0'
0/
#511950000000
1!
1'
1/
#511960000000
0!
0'
0/
#511970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#511980000000
0!
0'
0/
#511990000000
1!
1'
1/
#512000000000
0!
0'
0/
#512010000000
1!
1'
1/
#512020000000
0!
0'
0/
#512030000000
1!
1'
1/
#512040000000
0!
0'
0/
#512050000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#512060000000
0!
0'
0/
#512070000000
1!
1'
1/
#512080000000
0!
0'
0/
#512090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#512100000000
0!
0'
0/
#512110000000
1!
1'
1/
#512120000000
0!
0'
0/
#512130000000
#512140000000
1!
1'
1/
#512150000000
0!
0'
0/
#512160000000
1!
1'
1/
#512170000000
0!
1"
0'
1(
0/
10
#512180000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#512190000000
0!
0'
0/
#512200000000
1!
1'
1/
#512210000000
0!
0'
0/
#512220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#512230000000
0!
0'
0/
#512240000000
1!
1'
1/
#512250000000
0!
1"
0'
1(
0/
10
#512260000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#512270000000
0!
1$
0'
1+
0/
#512280000000
1!
1'
1/
#512290000000
0!
0'
0/
#512300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#512310000000
0!
0'
0/
#512320000000
1!
1'
1/
#512330000000
0!
0'
0/
#512340000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#512350000000
0!
0'
0/
#512360000000
1!
1'
1/
#512370000000
0!
0'
0/
#512380000000
1!
1'
1/
#512390000000
0!
0'
0/
#512400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#512410000000
0!
0'
0/
#512420000000
1!
1'
1/
#512430000000
0!
0'
0/
#512440000000
1!
1'
1/
#512450000000
0!
0'
0/
#512460000000
1!
1'
1/
#512470000000
0!
0'
0/
#512480000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#512490000000
0!
0'
0/
#512500000000
1!
1'
1/
#512510000000
0!
0'
0/
#512520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#512530000000
0!
0'
0/
#512540000000
1!
1'
1/
#512550000000
0!
0'
0/
#512560000000
#512570000000
1!
1'
1/
#512580000000
0!
0'
0/
#512590000000
1!
1'
1/
#512600000000
0!
1"
0'
1(
0/
10
#512610000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#512620000000
0!
0'
0/
#512630000000
1!
1'
1/
#512640000000
0!
0'
0/
#512650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#512660000000
0!
0'
0/
#512670000000
1!
1'
1/
#512680000000
0!
1"
0'
1(
0/
10
#512690000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#512700000000
0!
1$
0'
1+
0/
#512710000000
1!
1'
1/
#512720000000
0!
0'
0/
#512730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#512740000000
0!
0'
0/
#512750000000
1!
1'
1/
#512760000000
0!
0'
0/
#512770000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#512780000000
0!
0'
0/
#512790000000
1!
1'
1/
#512800000000
0!
0'
0/
#512810000000
1!
1'
1/
#512820000000
0!
0'
0/
#512830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#512840000000
0!
0'
0/
#512850000000
1!
1'
1/
#512860000000
0!
0'
0/
#512870000000
1!
1'
1/
#512880000000
0!
0'
0/
#512890000000
1!
1'
1/
#512900000000
0!
0'
0/
#512910000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#512920000000
0!
0'
0/
#512930000000
1!
1'
1/
#512940000000
0!
0'
0/
#512950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#512960000000
0!
0'
0/
#512970000000
1!
1'
1/
#512980000000
0!
0'
0/
#512990000000
#513000000000
1!
1'
1/
#513010000000
0!
0'
0/
#513020000000
1!
1'
1/
#513030000000
0!
1"
0'
1(
0/
10
#513040000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#513050000000
0!
0'
0/
#513060000000
1!
1'
1/
#513070000000
0!
0'
0/
#513080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#513090000000
0!
0'
0/
#513100000000
1!
1'
1/
#513110000000
0!
1"
0'
1(
0/
10
#513120000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#513130000000
0!
1$
0'
1+
0/
#513140000000
1!
1'
1/
#513150000000
0!
0'
0/
#513160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#513170000000
0!
0'
0/
#513180000000
1!
1'
1/
#513190000000
0!
0'
0/
#513200000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#513210000000
0!
0'
0/
#513220000000
1!
1'
1/
#513230000000
0!
0'
0/
#513240000000
1!
1'
1/
#513250000000
0!
0'
0/
#513260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#513270000000
0!
0'
0/
#513280000000
1!
1'
1/
#513290000000
0!
0'
0/
#513300000000
1!
1'
1/
#513310000000
0!
0'
0/
#513320000000
1!
1'
1/
#513330000000
0!
0'
0/
#513340000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#513350000000
0!
0'
0/
#513360000000
1!
1'
1/
#513370000000
0!
0'
0/
#513380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#513390000000
0!
0'
0/
#513400000000
1!
1'
1/
#513410000000
0!
0'
0/
#513420000000
#513430000000
1!
1'
1/
#513440000000
0!
0'
0/
#513450000000
1!
1'
1/
#513460000000
0!
1"
0'
1(
0/
10
#513470000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#513480000000
0!
0'
0/
#513490000000
1!
1'
1/
#513500000000
0!
0'
0/
#513510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#513520000000
0!
0'
0/
#513530000000
1!
1'
1/
#513540000000
0!
1"
0'
1(
0/
10
#513550000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#513560000000
0!
1$
0'
1+
0/
#513570000000
1!
1'
1/
#513580000000
0!
0'
0/
#513590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#513600000000
0!
0'
0/
#513610000000
1!
1'
1/
#513620000000
0!
0'
0/
#513630000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#513640000000
0!
0'
0/
#513650000000
1!
1'
1/
#513660000000
0!
0'
0/
#513670000000
1!
1'
1/
#513680000000
0!
0'
0/
#513690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#513700000000
0!
0'
0/
#513710000000
1!
1'
1/
#513720000000
0!
0'
0/
#513730000000
1!
1'
1/
#513740000000
0!
0'
0/
#513750000000
1!
1'
1/
#513760000000
0!
0'
0/
#513770000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#513780000000
0!
0'
0/
#513790000000
1!
1'
1/
#513800000000
0!
0'
0/
#513810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#513820000000
0!
0'
0/
#513830000000
1!
1'
1/
#513840000000
0!
0'
0/
#513850000000
#513860000000
1!
1'
1/
#513870000000
0!
0'
0/
#513880000000
1!
1'
1/
#513890000000
0!
1"
0'
1(
0/
10
#513900000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#513910000000
0!
0'
0/
#513920000000
1!
1'
1/
#513930000000
0!
0'
0/
#513940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#513950000000
0!
0'
0/
#513960000000
1!
1'
1/
#513970000000
0!
1"
0'
1(
0/
10
#513980000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#513990000000
0!
1$
0'
1+
0/
#514000000000
1!
1'
1/
#514010000000
0!
0'
0/
#514020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#514030000000
0!
0'
0/
#514040000000
1!
1'
1/
#514050000000
0!
0'
0/
#514060000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#514070000000
0!
0'
0/
#514080000000
1!
1'
1/
#514090000000
0!
0'
0/
#514100000000
1!
1'
1/
#514110000000
0!
0'
0/
#514120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#514130000000
0!
0'
0/
#514140000000
1!
1'
1/
#514150000000
0!
0'
0/
#514160000000
1!
1'
1/
#514170000000
0!
0'
0/
#514180000000
1!
1'
1/
#514190000000
0!
0'
0/
#514200000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#514210000000
0!
0'
0/
#514220000000
1!
1'
1/
#514230000000
0!
0'
0/
#514240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#514250000000
0!
0'
0/
#514260000000
1!
1'
1/
#514270000000
0!
0'
0/
#514280000000
#514290000000
1!
1'
1/
#514300000000
0!
0'
0/
#514310000000
1!
1'
1/
#514320000000
0!
1"
0'
1(
0/
10
#514330000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#514340000000
0!
0'
0/
#514350000000
1!
1'
1/
#514360000000
0!
0'
0/
#514370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#514380000000
0!
0'
0/
#514390000000
1!
1'
1/
#514400000000
0!
1"
0'
1(
0/
10
#514410000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#514420000000
0!
1$
0'
1+
0/
#514430000000
1!
1'
1/
#514440000000
0!
0'
0/
#514450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#514460000000
0!
0'
0/
#514470000000
1!
1'
1/
#514480000000
0!
0'
0/
#514490000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#514500000000
0!
0'
0/
#514510000000
1!
1'
1/
#514520000000
0!
0'
0/
#514530000000
1!
1'
1/
#514540000000
0!
0'
0/
#514550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#514560000000
0!
0'
0/
#514570000000
1!
1'
1/
#514580000000
0!
0'
0/
#514590000000
1!
1'
1/
#514600000000
0!
0'
0/
#514610000000
1!
1'
1/
#514620000000
0!
0'
0/
#514630000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#514640000000
0!
0'
0/
#514650000000
1!
1'
1/
#514660000000
0!
0'
0/
#514670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#514680000000
0!
0'
0/
#514690000000
1!
1'
1/
#514700000000
0!
0'
0/
#514710000000
#514720000000
1!
1'
1/
#514730000000
0!
0'
0/
#514740000000
1!
1'
1/
#514750000000
0!
1"
0'
1(
0/
10
#514760000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#514770000000
0!
0'
0/
#514780000000
1!
1'
1/
#514790000000
0!
0'
0/
#514800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#514810000000
0!
0'
0/
#514820000000
1!
1'
1/
#514830000000
0!
1"
0'
1(
0/
10
#514840000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#514850000000
0!
1$
0'
1+
0/
#514860000000
1!
1'
1/
#514870000000
0!
0'
0/
#514880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#514890000000
0!
0'
0/
#514900000000
1!
1'
1/
#514910000000
0!
0'
0/
#514920000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#514930000000
0!
0'
0/
#514940000000
1!
1'
1/
#514950000000
0!
0'
0/
#514960000000
1!
1'
1/
#514970000000
0!
0'
0/
#514980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#514990000000
0!
0'
0/
#515000000000
1!
1'
1/
#515010000000
0!
0'
0/
#515020000000
1!
1'
1/
#515030000000
0!
0'
0/
#515040000000
1!
1'
1/
#515050000000
0!
0'
0/
#515060000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#515070000000
0!
0'
0/
#515080000000
1!
1'
1/
#515090000000
0!
0'
0/
#515100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#515110000000
0!
0'
0/
#515120000000
1!
1'
1/
#515130000000
0!
0'
0/
#515140000000
#515150000000
1!
1'
1/
#515160000000
0!
0'
0/
#515170000000
1!
1'
1/
#515180000000
0!
1"
0'
1(
0/
10
#515190000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#515200000000
0!
0'
0/
#515210000000
1!
1'
1/
#515220000000
0!
0'
0/
#515230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#515240000000
0!
0'
0/
#515250000000
1!
1'
1/
#515260000000
0!
1"
0'
1(
0/
10
#515270000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#515280000000
0!
1$
0'
1+
0/
#515290000000
1!
1'
1/
#515300000000
0!
0'
0/
#515310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#515320000000
0!
0'
0/
#515330000000
1!
1'
1/
#515340000000
0!
0'
0/
#515350000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#515360000000
0!
0'
0/
#515370000000
1!
1'
1/
#515380000000
0!
0'
0/
#515390000000
1!
1'
1/
#515400000000
0!
0'
0/
#515410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#515420000000
0!
0'
0/
#515430000000
1!
1'
1/
#515440000000
0!
0'
0/
#515450000000
1!
1'
1/
#515460000000
0!
0'
0/
#515470000000
1!
1'
1/
#515480000000
0!
0'
0/
#515490000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#515500000000
0!
0'
0/
#515510000000
1!
1'
1/
#515520000000
0!
0'
0/
#515530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#515540000000
0!
0'
0/
#515550000000
1!
1'
1/
#515560000000
0!
0'
0/
#515570000000
#515580000000
1!
1'
1/
#515590000000
0!
0'
0/
#515600000000
1!
1'
1/
#515610000000
0!
1"
0'
1(
0/
10
#515620000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#515630000000
0!
0'
0/
#515640000000
1!
1'
1/
#515650000000
0!
0'
0/
#515660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#515670000000
0!
0'
0/
#515680000000
1!
1'
1/
#515690000000
0!
1"
0'
1(
0/
10
#515700000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#515710000000
0!
1$
0'
1+
0/
#515720000000
1!
1'
1/
#515730000000
0!
0'
0/
#515740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#515750000000
0!
0'
0/
#515760000000
1!
1'
1/
#515770000000
0!
0'
0/
#515780000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#515790000000
0!
0'
0/
#515800000000
1!
1'
1/
#515810000000
0!
0'
0/
#515820000000
1!
1'
1/
#515830000000
0!
0'
0/
#515840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#515850000000
0!
0'
0/
#515860000000
1!
1'
1/
#515870000000
0!
0'
0/
#515880000000
1!
1'
1/
#515890000000
0!
0'
0/
#515900000000
1!
1'
1/
#515910000000
0!
0'
0/
#515920000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#515930000000
0!
0'
0/
#515940000000
1!
1'
1/
#515950000000
0!
0'
0/
#515960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#515970000000
0!
0'
0/
#515980000000
1!
1'
1/
#515990000000
0!
0'
0/
#516000000000
#516010000000
1!
1'
1/
#516020000000
0!
0'
0/
#516030000000
1!
1'
1/
#516040000000
0!
1"
0'
1(
0/
10
#516050000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#516060000000
0!
0'
0/
#516070000000
1!
1'
1/
#516080000000
0!
0'
0/
#516090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#516100000000
0!
0'
0/
#516110000000
1!
1'
1/
#516120000000
0!
1"
0'
1(
0/
10
#516130000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#516140000000
0!
1$
0'
1+
0/
#516150000000
1!
1'
1/
#516160000000
0!
0'
0/
#516170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#516180000000
0!
0'
0/
#516190000000
1!
1'
1/
#516200000000
0!
0'
0/
#516210000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#516220000000
0!
0'
0/
#516230000000
1!
1'
1/
#516240000000
0!
0'
0/
#516250000000
1!
1'
1/
#516260000000
0!
0'
0/
#516270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#516280000000
0!
0'
0/
#516290000000
1!
1'
1/
#516300000000
0!
0'
0/
#516310000000
1!
1'
1/
#516320000000
0!
0'
0/
#516330000000
1!
1'
1/
#516340000000
0!
0'
0/
#516350000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#516360000000
0!
0'
0/
#516370000000
1!
1'
1/
#516380000000
0!
0'
0/
#516390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#516400000000
0!
0'
0/
#516410000000
1!
1'
1/
#516420000000
0!
0'
0/
#516430000000
#516440000000
1!
1'
1/
#516450000000
0!
0'
0/
#516460000000
1!
1'
1/
#516470000000
0!
1"
0'
1(
0/
10
#516480000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#516490000000
0!
0'
0/
#516500000000
1!
1'
1/
#516510000000
0!
0'
0/
#516520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#516530000000
0!
0'
0/
#516540000000
1!
1'
1/
#516550000000
0!
1"
0'
1(
0/
10
#516560000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#516570000000
0!
1$
0'
1+
0/
#516580000000
1!
1'
1/
#516590000000
0!
0'
0/
#516600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#516610000000
0!
0'
0/
#516620000000
1!
1'
1/
#516630000000
0!
0'
0/
#516640000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#516650000000
0!
0'
0/
#516660000000
1!
1'
1/
#516670000000
0!
0'
0/
#516680000000
1!
1'
1/
#516690000000
0!
0'
0/
#516700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#516710000000
0!
0'
0/
#516720000000
1!
1'
1/
#516730000000
0!
0'
0/
#516740000000
1!
1'
1/
#516750000000
0!
0'
0/
#516760000000
1!
1'
1/
#516770000000
0!
0'
0/
#516780000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#516790000000
0!
0'
0/
#516800000000
1!
1'
1/
#516810000000
0!
0'
0/
#516820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#516830000000
0!
0'
0/
#516840000000
1!
1'
1/
#516850000000
0!
0'
0/
#516860000000
#516870000000
1!
1'
1/
#516880000000
0!
0'
0/
#516890000000
1!
1'
1/
#516900000000
0!
1"
0'
1(
0/
10
#516910000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#516920000000
0!
0'
0/
#516930000000
1!
1'
1/
#516940000000
0!
0'
0/
#516950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#516960000000
0!
0'
0/
#516970000000
1!
1'
1/
#516980000000
0!
1"
0'
1(
0/
10
#516990000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#517000000000
0!
1$
0'
1+
0/
#517010000000
1!
1'
1/
#517020000000
0!
0'
0/
#517030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#517040000000
0!
0'
0/
#517050000000
1!
1'
1/
#517060000000
0!
0'
0/
#517070000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#517080000000
0!
0'
0/
#517090000000
1!
1'
1/
#517100000000
0!
0'
0/
#517110000000
1!
1'
1/
#517120000000
0!
0'
0/
#517130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#517140000000
0!
0'
0/
#517150000000
1!
1'
1/
#517160000000
0!
0'
0/
#517170000000
1!
1'
1/
#517180000000
0!
0'
0/
#517190000000
1!
1'
1/
#517200000000
0!
0'
0/
#517210000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#517220000000
0!
0'
0/
#517230000000
1!
1'
1/
#517240000000
0!
0'
0/
#517250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#517260000000
0!
0'
0/
#517270000000
1!
1'
1/
#517280000000
0!
0'
0/
#517290000000
#517300000000
1!
1'
1/
#517310000000
0!
0'
0/
#517320000000
1!
1'
1/
#517330000000
0!
1"
0'
1(
0/
10
#517340000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#517350000000
0!
0'
0/
#517360000000
1!
1'
1/
#517370000000
0!
0'
0/
#517380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#517390000000
0!
0'
0/
#517400000000
1!
1'
1/
#517410000000
0!
1"
0'
1(
0/
10
#517420000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#517430000000
0!
1$
0'
1+
0/
#517440000000
1!
1'
1/
#517450000000
0!
0'
0/
#517460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#517470000000
0!
0'
0/
#517480000000
1!
1'
1/
#517490000000
0!
0'
0/
#517500000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#517510000000
0!
0'
0/
#517520000000
1!
1'
1/
#517530000000
0!
0'
0/
#517540000000
1!
1'
1/
#517550000000
0!
0'
0/
#517560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#517570000000
0!
0'
0/
#517580000000
1!
1'
1/
#517590000000
0!
0'
0/
#517600000000
1!
1'
1/
#517610000000
0!
0'
0/
#517620000000
1!
1'
1/
#517630000000
0!
0'
0/
#517640000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#517650000000
0!
0'
0/
#517660000000
1!
1'
1/
#517670000000
0!
0'
0/
#517680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#517690000000
0!
0'
0/
#517700000000
1!
1'
1/
#517710000000
0!
0'
0/
#517720000000
#517730000000
1!
1'
1/
#517740000000
0!
0'
0/
#517750000000
1!
1'
1/
#517760000000
0!
1"
0'
1(
0/
10
#517770000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#517780000000
0!
0'
0/
#517790000000
1!
1'
1/
#517800000000
0!
0'
0/
#517810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#517820000000
0!
0'
0/
#517830000000
1!
1'
1/
#517840000000
0!
1"
0'
1(
0/
10
#517850000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#517860000000
0!
1$
0'
1+
0/
#517870000000
1!
1'
1/
#517880000000
0!
0'
0/
#517890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#517900000000
0!
0'
0/
#517910000000
1!
1'
1/
#517920000000
0!
0'
0/
#517930000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#517940000000
0!
0'
0/
#517950000000
1!
1'
1/
#517960000000
0!
0'
0/
#517970000000
1!
1'
1/
#517980000000
0!
0'
0/
#517990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#518000000000
0!
0'
0/
#518010000000
1!
1'
1/
#518020000000
0!
0'
0/
#518030000000
1!
1'
1/
#518040000000
0!
0'
0/
#518050000000
1!
1'
1/
#518060000000
0!
0'
0/
#518070000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#518080000000
0!
0'
0/
#518090000000
1!
1'
1/
#518100000000
0!
0'
0/
#518110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#518120000000
0!
0'
0/
#518130000000
1!
1'
1/
#518140000000
0!
0'
0/
#518150000000
#518160000000
1!
1'
1/
#518170000000
0!
0'
0/
#518180000000
1!
1'
1/
#518190000000
0!
1"
0'
1(
0/
10
#518200000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#518210000000
0!
0'
0/
#518220000000
1!
1'
1/
#518230000000
0!
0'
0/
#518240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#518250000000
0!
0'
0/
#518260000000
1!
1'
1/
#518270000000
0!
1"
0'
1(
0/
10
#518280000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#518290000000
0!
1$
0'
1+
0/
#518300000000
1!
1'
1/
#518310000000
0!
0'
0/
#518320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#518330000000
0!
0'
0/
#518340000000
1!
1'
1/
#518350000000
0!
0'
0/
#518360000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#518370000000
0!
0'
0/
#518380000000
1!
1'
1/
#518390000000
0!
0'
0/
#518400000000
1!
1'
1/
#518410000000
0!
0'
0/
#518420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#518430000000
0!
0'
0/
#518440000000
1!
1'
1/
#518450000000
0!
0'
0/
#518460000000
1!
1'
1/
#518470000000
0!
0'
0/
#518480000000
1!
1'
1/
#518490000000
0!
0'
0/
#518500000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#518510000000
0!
0'
0/
#518520000000
1!
1'
1/
#518530000000
0!
0'
0/
#518540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#518550000000
0!
0'
0/
#518560000000
1!
1'
1/
#518570000000
0!
0'
0/
#518580000000
#518590000000
1!
1'
1/
#518600000000
0!
0'
0/
#518610000000
1!
1'
1/
#518620000000
0!
1"
0'
1(
0/
10
#518630000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#518640000000
0!
0'
0/
#518650000000
1!
1'
1/
#518660000000
0!
0'
0/
#518670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#518680000000
0!
0'
0/
#518690000000
1!
1'
1/
#518700000000
0!
1"
0'
1(
0/
10
#518710000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#518720000000
0!
1$
0'
1+
0/
#518730000000
1!
1'
1/
#518740000000
0!
0'
0/
#518750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#518760000000
0!
0'
0/
#518770000000
1!
1'
1/
#518780000000
0!
0'
0/
#518790000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#518800000000
0!
0'
0/
#518810000000
1!
1'
1/
#518820000000
0!
0'
0/
#518830000000
1!
1'
1/
#518840000000
0!
0'
0/
#518850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#518860000000
0!
0'
0/
#518870000000
1!
1'
1/
#518880000000
0!
0'
0/
#518890000000
1!
1'
1/
#518900000000
0!
0'
0/
#518910000000
1!
1'
1/
#518920000000
0!
0'
0/
#518930000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#518940000000
0!
0'
0/
#518950000000
1!
1'
1/
#518960000000
0!
0'
0/
#518970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#518980000000
0!
0'
0/
#518990000000
1!
1'
1/
#519000000000
0!
0'
0/
#519010000000
#519020000000
1!
1'
1/
#519030000000
0!
0'
0/
#519040000000
1!
1'
1/
#519050000000
0!
1"
0'
1(
0/
10
#519060000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#519070000000
0!
0'
0/
#519080000000
1!
1'
1/
#519090000000
0!
0'
0/
#519100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#519110000000
0!
0'
0/
#519120000000
1!
1'
1/
#519130000000
0!
1"
0'
1(
0/
10
#519140000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#519150000000
0!
1$
0'
1+
0/
#519160000000
1!
1'
1/
#519170000000
0!
0'
0/
#519180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#519190000000
0!
0'
0/
#519200000000
1!
1'
1/
#519210000000
0!
0'
0/
#519220000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#519230000000
0!
0'
0/
#519240000000
1!
1'
1/
#519250000000
0!
0'
0/
#519260000000
1!
1'
1/
#519270000000
0!
0'
0/
#519280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#519290000000
0!
0'
0/
#519300000000
1!
1'
1/
#519310000000
0!
0'
0/
#519320000000
1!
1'
1/
#519330000000
0!
0'
0/
#519340000000
1!
1'
1/
#519350000000
0!
0'
0/
#519360000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#519370000000
0!
0'
0/
#519380000000
1!
1'
1/
#519390000000
0!
0'
0/
#519400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#519410000000
0!
0'
0/
#519420000000
1!
1'
1/
#519430000000
0!
0'
0/
#519440000000
#519450000000
1!
1'
1/
#519460000000
0!
0'
0/
#519470000000
1!
1'
1/
#519480000000
0!
1"
0'
1(
0/
10
#519490000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#519500000000
0!
0'
0/
#519510000000
1!
1'
1/
#519520000000
0!
0'
0/
#519530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#519540000000
0!
0'
0/
#519550000000
1!
1'
1/
#519560000000
0!
1"
0'
1(
0/
10
#519570000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#519580000000
0!
1$
0'
1+
0/
#519590000000
1!
1'
1/
#519600000000
0!
0'
0/
#519610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#519620000000
0!
0'
0/
#519630000000
1!
1'
1/
#519640000000
0!
0'
0/
#519650000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#519660000000
0!
0'
0/
#519670000000
1!
1'
1/
#519680000000
0!
0'
0/
#519690000000
1!
1'
1/
#519700000000
0!
0'
0/
#519710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#519720000000
0!
0'
0/
#519730000000
1!
1'
1/
#519740000000
0!
0'
0/
#519750000000
1!
1'
1/
#519760000000
0!
0'
0/
#519770000000
1!
1'
1/
#519780000000
0!
0'
0/
#519790000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#519800000000
0!
0'
0/
#519810000000
1!
1'
1/
#519820000000
0!
0'
0/
#519830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#519840000000
0!
0'
0/
#519850000000
1!
1'
1/
#519860000000
0!
0'
0/
#519870000000
#519880000000
1!
1'
1/
#519890000000
0!
0'
0/
#519900000000
1!
1'
1/
#519910000000
0!
1"
0'
1(
0/
10
#519920000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#519930000000
0!
0'
0/
#519940000000
1!
1'
1/
#519950000000
0!
0'
0/
#519960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#519970000000
0!
0'
0/
#519980000000
1!
1'
1/
#519990000000
0!
1"
0'
1(
0/
10
#520000000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#520010000000
0!
1$
0'
1+
0/
#520020000000
1!
1'
1/
#520030000000
0!
0'
0/
#520040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#520050000000
0!
0'
0/
#520060000000
1!
1'
1/
#520070000000
0!
0'
0/
#520080000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#520090000000
0!
0'
0/
#520100000000
1!
1'
1/
#520110000000
0!
0'
0/
#520120000000
1!
1'
1/
#520130000000
0!
0'
0/
#520140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#520150000000
0!
0'
0/
#520160000000
1!
1'
1/
#520170000000
0!
0'
0/
#520180000000
1!
1'
1/
#520190000000
0!
0'
0/
#520200000000
1!
1'
1/
#520210000000
0!
0'
0/
#520220000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#520230000000
0!
0'
0/
#520240000000
1!
1'
1/
#520250000000
0!
0'
0/
#520260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#520270000000
0!
0'
0/
#520280000000
1!
1'
1/
#520290000000
0!
0'
0/
#520300000000
#520310000000
1!
1'
1/
#520320000000
0!
0'
0/
#520330000000
1!
1'
1/
#520340000000
0!
1"
0'
1(
0/
10
#520350000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#520360000000
0!
0'
0/
#520370000000
1!
1'
1/
#520380000000
0!
0'
0/
#520390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#520400000000
0!
0'
0/
#520410000000
1!
1'
1/
#520420000000
0!
1"
0'
1(
0/
10
#520430000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#520440000000
0!
1$
0'
1+
0/
#520450000000
1!
1'
1/
#520460000000
0!
0'
0/
#520470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#520480000000
0!
0'
0/
#520490000000
1!
1'
1/
#520500000000
0!
0'
0/
#520510000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#520520000000
0!
0'
0/
#520530000000
1!
1'
1/
#520540000000
0!
0'
0/
#520550000000
1!
1'
1/
#520560000000
0!
0'
0/
#520570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#520580000000
0!
0'
0/
#520590000000
1!
1'
1/
#520600000000
0!
0'
0/
#520610000000
1!
1'
1/
#520620000000
0!
0'
0/
#520630000000
1!
1'
1/
#520640000000
0!
0'
0/
#520650000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#520660000000
0!
0'
0/
#520670000000
1!
1'
1/
#520680000000
0!
0'
0/
#520690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#520700000000
0!
0'
0/
#520710000000
1!
1'
1/
#520720000000
0!
0'
0/
#520730000000
#520740000000
1!
1'
1/
#520750000000
0!
0'
0/
#520760000000
1!
1'
1/
#520770000000
0!
1"
0'
1(
0/
10
#520780000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#520790000000
0!
0'
0/
#520800000000
1!
1'
1/
#520810000000
0!
0'
0/
#520820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#520830000000
0!
0'
0/
#520840000000
1!
1'
1/
#520850000000
0!
1"
0'
1(
0/
10
#520860000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#520870000000
0!
1$
0'
1+
0/
#520880000000
1!
1'
1/
#520890000000
0!
0'
0/
#520900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#520910000000
0!
0'
0/
#520920000000
1!
1'
1/
#520930000000
0!
0'
0/
#520940000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#520950000000
0!
0'
0/
#520960000000
1!
1'
1/
#520970000000
0!
0'
0/
#520980000000
1!
1'
1/
#520990000000
0!
0'
0/
#521000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#521010000000
0!
0'
0/
#521020000000
1!
1'
1/
#521030000000
0!
0'
0/
#521040000000
1!
1'
1/
#521050000000
0!
0'
0/
#521060000000
1!
1'
1/
#521070000000
0!
0'
0/
#521080000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#521090000000
0!
0'
0/
#521100000000
1!
1'
1/
#521110000000
0!
0'
0/
#521120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#521130000000
0!
0'
0/
#521140000000
1!
1'
1/
#521150000000
0!
0'
0/
#521160000000
#521170000000
1!
1'
1/
#521180000000
0!
0'
0/
#521190000000
1!
1'
1/
#521200000000
0!
1"
0'
1(
0/
10
#521210000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#521220000000
0!
0'
0/
#521230000000
1!
1'
1/
#521240000000
0!
0'
0/
#521250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#521260000000
0!
0'
0/
#521270000000
1!
1'
1/
#521280000000
0!
1"
0'
1(
0/
10
#521290000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#521300000000
0!
1$
0'
1+
0/
#521310000000
1!
1'
1/
#521320000000
0!
0'
0/
#521330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#521340000000
0!
0'
0/
#521350000000
1!
1'
1/
#521360000000
0!
0'
0/
#521370000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#521380000000
0!
0'
0/
#521390000000
1!
1'
1/
#521400000000
0!
0'
0/
#521410000000
1!
1'
1/
#521420000000
0!
0'
0/
#521430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#521440000000
0!
0'
0/
#521450000000
1!
1'
1/
#521460000000
0!
0'
0/
#521470000000
1!
1'
1/
#521480000000
0!
0'
0/
#521490000000
1!
1'
1/
#521500000000
0!
0'
0/
#521510000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#521520000000
0!
0'
0/
#521530000000
1!
1'
1/
#521540000000
0!
0'
0/
#521550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#521560000000
0!
0'
0/
#521570000000
1!
1'
1/
#521580000000
0!
0'
0/
#521590000000
#521600000000
1!
1'
1/
#521610000000
0!
0'
0/
#521620000000
1!
1'
1/
#521630000000
0!
1"
0'
1(
0/
10
#521640000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#521650000000
0!
0'
0/
#521660000000
1!
1'
1/
#521670000000
0!
0'
0/
#521680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#521690000000
0!
0'
0/
#521700000000
1!
1'
1/
#521710000000
0!
1"
0'
1(
0/
10
#521720000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#521730000000
0!
1$
0'
1+
0/
#521740000000
1!
1'
1/
#521750000000
0!
0'
0/
#521760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#521770000000
0!
0'
0/
#521780000000
1!
1'
1/
#521790000000
0!
0'
0/
#521800000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#521810000000
0!
0'
0/
#521820000000
1!
1'
1/
#521830000000
0!
0'
0/
#521840000000
1!
1'
1/
#521850000000
0!
0'
0/
#521860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#521870000000
0!
0'
0/
#521880000000
1!
1'
1/
#521890000000
0!
0'
0/
#521900000000
1!
1'
1/
#521910000000
0!
0'
0/
#521920000000
1!
1'
1/
#521930000000
0!
0'
0/
#521940000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#521950000000
0!
0'
0/
#521960000000
1!
1'
1/
#521970000000
0!
0'
0/
#521980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#521990000000
0!
0'
0/
#522000000000
1!
1'
1/
#522010000000
0!
0'
0/
#522020000000
#522030000000
1!
1'
1/
#522040000000
0!
0'
0/
#522050000000
1!
1'
1/
#522060000000
0!
1"
0'
1(
0/
10
#522070000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#522080000000
0!
0'
0/
#522090000000
1!
1'
1/
#522100000000
0!
0'
0/
#522110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#522120000000
0!
0'
0/
#522130000000
1!
1'
1/
#522140000000
0!
1"
0'
1(
0/
10
#522150000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#522160000000
0!
1$
0'
1+
0/
#522170000000
1!
1'
1/
#522180000000
0!
0'
0/
#522190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#522200000000
0!
0'
0/
#522210000000
1!
1'
1/
#522220000000
0!
0'
0/
#522230000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#522240000000
0!
0'
0/
#522250000000
1!
1'
1/
#522260000000
0!
0'
0/
#522270000000
1!
1'
1/
#522280000000
0!
0'
0/
#522290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#522300000000
0!
0'
0/
#522310000000
1!
1'
1/
#522320000000
0!
0'
0/
#522330000000
1!
1'
1/
#522340000000
0!
0'
0/
#522350000000
1!
1'
1/
#522360000000
0!
0'
0/
#522370000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#522380000000
0!
0'
0/
#522390000000
1!
1'
1/
#522400000000
0!
0'
0/
#522410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#522420000000
0!
0'
0/
#522430000000
1!
1'
1/
#522440000000
0!
0'
0/
#522450000000
#522460000000
1!
1'
1/
#522470000000
0!
0'
0/
#522480000000
1!
1'
1/
#522490000000
0!
1"
0'
1(
0/
10
#522500000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#522510000000
0!
0'
0/
#522520000000
1!
1'
1/
#522530000000
0!
0'
0/
#522540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#522550000000
0!
0'
0/
#522560000000
1!
1'
1/
#522570000000
0!
1"
0'
1(
0/
10
#522580000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#522590000000
0!
1$
0'
1+
0/
#522600000000
1!
1'
1/
#522610000000
0!
0'
0/
#522620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#522630000000
0!
0'
0/
#522640000000
1!
1'
1/
#522650000000
0!
0'
0/
#522660000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#522670000000
0!
0'
0/
#522680000000
1!
1'
1/
#522690000000
0!
0'
0/
#522700000000
1!
1'
1/
#522710000000
0!
0'
0/
#522720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#522730000000
0!
0'
0/
#522740000000
1!
1'
1/
#522750000000
0!
0'
0/
#522760000000
1!
1'
1/
#522770000000
0!
0'
0/
#522780000000
1!
1'
1/
#522790000000
0!
0'
0/
#522800000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#522810000000
0!
0'
0/
#522820000000
1!
1'
1/
#522830000000
0!
0'
0/
#522840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#522850000000
0!
0'
0/
#522860000000
1!
1'
1/
#522870000000
0!
0'
0/
#522880000000
#522890000000
1!
1'
1/
#522900000000
0!
0'
0/
#522910000000
1!
1'
1/
#522920000000
0!
1"
0'
1(
0/
10
#522930000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#522940000000
0!
0'
0/
#522950000000
1!
1'
1/
#522960000000
0!
0'
0/
#522970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#522980000000
0!
0'
0/
#522990000000
1!
1'
1/
#523000000000
0!
1"
0'
1(
0/
10
#523010000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#523020000000
0!
1$
0'
1+
0/
#523030000000
1!
1'
1/
#523040000000
0!
0'
0/
#523050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#523060000000
0!
0'
0/
#523070000000
1!
1'
1/
#523080000000
0!
0'
0/
#523090000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#523100000000
0!
0'
0/
#523110000000
1!
1'
1/
#523120000000
0!
0'
0/
#523130000000
1!
1'
1/
#523140000000
0!
0'
0/
#523150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#523160000000
0!
0'
0/
#523170000000
1!
1'
1/
#523180000000
0!
0'
0/
#523190000000
1!
1'
1/
#523200000000
0!
0'
0/
#523210000000
1!
1'
1/
#523220000000
0!
0'
0/
#523230000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#523240000000
0!
0'
0/
#523250000000
1!
1'
1/
#523260000000
0!
0'
0/
#523270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#523280000000
0!
0'
0/
#523290000000
1!
1'
1/
#523300000000
0!
0'
0/
#523310000000
#523320000000
1!
1'
1/
#523330000000
0!
0'
0/
#523340000000
1!
1'
1/
#523350000000
0!
1"
0'
1(
0/
10
#523360000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#523370000000
0!
0'
0/
#523380000000
1!
1'
1/
#523390000000
0!
0'
0/
#523400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#523410000000
0!
0'
0/
#523420000000
1!
1'
1/
#523430000000
0!
1"
0'
1(
0/
10
#523440000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#523450000000
0!
1$
0'
1+
0/
#523460000000
1!
1'
1/
#523470000000
0!
0'
0/
#523480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#523490000000
0!
0'
0/
#523500000000
1!
1'
1/
#523510000000
0!
0'
0/
#523520000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#523530000000
0!
0'
0/
#523540000000
1!
1'
1/
#523550000000
0!
0'
0/
#523560000000
1!
1'
1/
#523570000000
0!
0'
0/
#523580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#523590000000
0!
0'
0/
#523600000000
1!
1'
1/
#523610000000
0!
0'
0/
#523620000000
1!
1'
1/
#523630000000
0!
0'
0/
#523640000000
1!
1'
1/
#523650000000
0!
0'
0/
#523660000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#523670000000
0!
0'
0/
#523680000000
1!
1'
1/
#523690000000
0!
0'
0/
#523700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#523710000000
0!
0'
0/
#523720000000
1!
1'
1/
#523730000000
0!
0'
0/
#523740000000
#523750000000
1!
1'
1/
#523760000000
0!
0'
0/
#523770000000
1!
1'
1/
#523780000000
0!
1"
0'
1(
0/
10
#523790000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#523800000000
0!
0'
0/
#523810000000
1!
1'
1/
#523820000000
0!
0'
0/
#523830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#523840000000
0!
0'
0/
#523850000000
1!
1'
1/
#523860000000
0!
1"
0'
1(
0/
10
#523870000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#523880000000
0!
1$
0'
1+
0/
#523890000000
1!
1'
1/
#523900000000
0!
0'
0/
#523910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#523920000000
0!
0'
0/
#523930000000
1!
1'
1/
#523940000000
0!
0'
0/
#523950000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#523960000000
0!
0'
0/
#523970000000
1!
1'
1/
#523980000000
0!
0'
0/
#523990000000
1!
1'
1/
#524000000000
0!
0'
0/
#524010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#524020000000
0!
0'
0/
#524030000000
1!
1'
1/
#524040000000
0!
0'
0/
#524050000000
1!
1'
1/
#524060000000
0!
0'
0/
#524070000000
1!
1'
1/
#524080000000
0!
0'
0/
#524090000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#524100000000
0!
0'
0/
#524110000000
1!
1'
1/
#524120000000
0!
0'
0/
#524130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#524140000000
0!
0'
0/
#524150000000
1!
1'
1/
#524160000000
0!
0'
0/
#524170000000
#524180000000
1!
1'
1/
#524190000000
0!
0'
0/
#524200000000
1!
1'
1/
#524210000000
0!
1"
0'
1(
0/
10
#524220000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#524230000000
0!
0'
0/
#524240000000
1!
1'
1/
#524250000000
0!
0'
0/
#524260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#524270000000
0!
0'
0/
#524280000000
1!
1'
1/
#524290000000
0!
1"
0'
1(
0/
10
#524300000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#524310000000
0!
1$
0'
1+
0/
#524320000000
1!
1'
1/
#524330000000
0!
0'
0/
#524340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#524350000000
0!
0'
0/
#524360000000
1!
1'
1/
#524370000000
0!
0'
0/
#524380000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#524390000000
0!
0'
0/
#524400000000
1!
1'
1/
#524410000000
0!
0'
0/
#524420000000
1!
1'
1/
#524430000000
0!
0'
0/
#524440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#524450000000
0!
0'
0/
#524460000000
1!
1'
1/
#524470000000
0!
0'
0/
#524480000000
1!
1'
1/
#524490000000
0!
0'
0/
#524500000000
1!
1'
1/
#524510000000
0!
0'
0/
#524520000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#524530000000
0!
0'
0/
#524540000000
1!
1'
1/
#524550000000
0!
0'
0/
#524560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#524570000000
0!
0'
0/
#524580000000
1!
1'
1/
#524590000000
0!
0'
0/
#524600000000
#524610000000
1!
1'
1/
#524620000000
0!
0'
0/
#524630000000
1!
1'
1/
#524640000000
0!
1"
0'
1(
0/
10
#524650000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#524660000000
0!
0'
0/
#524670000000
1!
1'
1/
#524680000000
0!
0'
0/
#524690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#524700000000
0!
0'
0/
#524710000000
1!
1'
1/
#524720000000
0!
1"
0'
1(
0/
10
#524730000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#524740000000
0!
1$
0'
1+
0/
#524750000000
1!
1'
1/
#524760000000
0!
0'
0/
#524770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#524780000000
0!
0'
0/
#524790000000
1!
1'
1/
#524800000000
0!
0'
0/
#524810000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#524820000000
0!
0'
0/
#524830000000
1!
1'
1/
#524840000000
0!
0'
0/
#524850000000
1!
1'
1/
#524860000000
0!
0'
0/
#524870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#524880000000
0!
0'
0/
#524890000000
1!
1'
1/
#524900000000
0!
0'
0/
#524910000000
1!
1'
1/
#524920000000
0!
0'
0/
#524930000000
1!
1'
1/
#524940000000
0!
0'
0/
#524950000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#524960000000
0!
0'
0/
#524970000000
1!
1'
1/
#524980000000
0!
0'
0/
#524990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#525000000000
0!
0'
0/
#525010000000
1!
1'
1/
#525020000000
0!
0'
0/
#525030000000
#525040000000
1!
1'
1/
#525050000000
0!
0'
0/
#525060000000
1!
1'
1/
#525070000000
0!
1"
0'
1(
0/
10
#525080000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#525090000000
0!
0'
0/
#525100000000
1!
1'
1/
#525110000000
0!
0'
0/
#525120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#525130000000
0!
0'
0/
#525140000000
1!
1'
1/
#525150000000
0!
1"
0'
1(
0/
10
#525160000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#525170000000
0!
1$
0'
1+
0/
#525180000000
1!
1'
1/
#525190000000
0!
0'
0/
#525200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#525210000000
0!
0'
0/
#525220000000
1!
1'
1/
#525230000000
0!
0'
0/
#525240000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#525250000000
0!
0'
0/
#525260000000
1!
1'
1/
#525270000000
0!
0'
0/
#525280000000
1!
1'
1/
#525290000000
0!
0'
0/
#525300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#525310000000
0!
0'
0/
#525320000000
1!
1'
1/
#525330000000
0!
0'
0/
#525340000000
1!
1'
1/
#525350000000
0!
0'
0/
#525360000000
1!
1'
1/
#525370000000
0!
0'
0/
#525380000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#525390000000
0!
0'
0/
#525400000000
1!
1'
1/
#525410000000
0!
0'
0/
#525420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#525430000000
0!
0'
0/
#525440000000
1!
1'
1/
#525450000000
0!
0'
0/
#525460000000
#525470000000
1!
1'
1/
#525480000000
0!
0'
0/
#525490000000
1!
1'
1/
#525500000000
0!
1"
0'
1(
0/
10
#525510000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#525520000000
0!
0'
0/
#525530000000
1!
1'
1/
#525540000000
0!
0'
0/
#525550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#525560000000
0!
0'
0/
#525570000000
1!
1'
1/
#525580000000
0!
1"
0'
1(
0/
10
#525590000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#525600000000
0!
1$
0'
1+
0/
#525610000000
1!
1'
1/
#525620000000
0!
0'
0/
#525630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#525640000000
0!
0'
0/
#525650000000
1!
1'
1/
#525660000000
0!
0'
0/
#525670000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#525680000000
0!
0'
0/
#525690000000
1!
1'
1/
#525700000000
0!
0'
0/
#525710000000
1!
1'
1/
#525720000000
0!
0'
0/
#525730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#525740000000
0!
0'
0/
#525750000000
1!
1'
1/
#525760000000
0!
0'
0/
#525770000000
1!
1'
1/
#525780000000
0!
0'
0/
#525790000000
1!
1'
1/
#525800000000
0!
0'
0/
#525810000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#525820000000
0!
0'
0/
#525830000000
1!
1'
1/
#525840000000
0!
0'
0/
#525850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#525860000000
0!
0'
0/
#525870000000
1!
1'
1/
#525880000000
0!
0'
0/
#525890000000
#525900000000
1!
1'
1/
#525910000000
0!
0'
0/
#525920000000
1!
1'
1/
#525930000000
0!
1"
0'
1(
0/
10
#525940000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#525950000000
0!
0'
0/
#525960000000
1!
1'
1/
#525970000000
0!
0'
0/
#525980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#525990000000
0!
0'
0/
#526000000000
1!
1'
1/
#526010000000
0!
1"
0'
1(
0/
10
#526020000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#526030000000
0!
1$
0'
1+
0/
#526040000000
1!
1'
1/
#526050000000
0!
0'
0/
#526060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#526070000000
0!
0'
0/
#526080000000
1!
1'
1/
#526090000000
0!
0'
0/
#526100000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#526110000000
0!
0'
0/
#526120000000
1!
1'
1/
#526130000000
0!
0'
0/
#526140000000
1!
1'
1/
#526150000000
0!
0'
0/
#526160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#526170000000
0!
0'
0/
#526180000000
1!
1'
1/
#526190000000
0!
0'
0/
#526200000000
1!
1'
1/
#526210000000
0!
0'
0/
#526220000000
1!
1'
1/
#526230000000
0!
0'
0/
#526240000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#526250000000
0!
0'
0/
#526260000000
1!
1'
1/
#526270000000
0!
0'
0/
#526280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#526290000000
0!
0'
0/
#526300000000
1!
1'
1/
#526310000000
0!
0'
0/
#526320000000
#526330000000
1!
1'
1/
#526340000000
0!
0'
0/
#526350000000
1!
1'
1/
#526360000000
0!
1"
0'
1(
0/
10
#526370000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#526380000000
0!
0'
0/
#526390000000
1!
1'
1/
#526400000000
0!
0'
0/
#526410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#526420000000
0!
0'
0/
#526430000000
1!
1'
1/
#526440000000
0!
1"
0'
1(
0/
10
#526450000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#526460000000
0!
1$
0'
1+
0/
#526470000000
1!
1'
1/
#526480000000
0!
0'
0/
#526490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#526500000000
0!
0'
0/
#526510000000
1!
1'
1/
#526520000000
0!
0'
0/
#526530000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#526540000000
0!
0'
0/
#526550000000
1!
1'
1/
#526560000000
0!
0'
0/
#526570000000
1!
1'
1/
#526580000000
0!
0'
0/
#526590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#526600000000
0!
0'
0/
#526610000000
1!
1'
1/
#526620000000
0!
0'
0/
#526630000000
1!
1'
1/
#526640000000
0!
0'
0/
#526650000000
1!
1'
1/
#526660000000
0!
0'
0/
#526670000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#526680000000
0!
0'
0/
#526690000000
1!
1'
1/
#526700000000
0!
0'
0/
#526710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#526720000000
0!
0'
0/
#526730000000
1!
1'
1/
#526740000000
0!
0'
0/
#526750000000
#526760000000
1!
1'
1/
#526770000000
0!
0'
0/
#526780000000
1!
1'
1/
#526790000000
0!
1"
0'
1(
0/
10
#526800000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#526810000000
0!
0'
0/
#526820000000
1!
1'
1/
#526830000000
0!
0'
0/
#526840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#526850000000
0!
0'
0/
#526860000000
1!
1'
1/
#526870000000
0!
1"
0'
1(
0/
10
#526880000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#526890000000
0!
1$
0'
1+
0/
#526900000000
1!
1'
1/
#526910000000
0!
0'
0/
#526920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#526930000000
0!
0'
0/
#526940000000
1!
1'
1/
#526950000000
0!
0'
0/
#526960000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#526970000000
0!
0'
0/
#526980000000
1!
1'
1/
#526990000000
0!
0'
0/
#527000000000
1!
1'
1/
#527010000000
0!
0'
0/
#527020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#527030000000
0!
0'
0/
#527040000000
1!
1'
1/
#527050000000
0!
0'
0/
#527060000000
1!
1'
1/
#527070000000
0!
0'
0/
#527080000000
1!
1'
1/
#527090000000
0!
0'
0/
#527100000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#527110000000
0!
0'
0/
#527120000000
1!
1'
1/
#527130000000
0!
0'
0/
#527140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#527150000000
0!
0'
0/
#527160000000
1!
1'
1/
#527170000000
0!
0'
0/
#527180000000
#527190000000
1!
1'
1/
#527200000000
0!
0'
0/
#527210000000
1!
1'
1/
#527220000000
0!
1"
0'
1(
0/
10
#527230000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#527240000000
0!
0'
0/
#527250000000
1!
1'
1/
#527260000000
0!
0'
0/
#527270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#527280000000
0!
0'
0/
#527290000000
1!
1'
1/
#527300000000
0!
1"
0'
1(
0/
10
#527310000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#527320000000
0!
1$
0'
1+
0/
#527330000000
1!
1'
1/
#527340000000
0!
0'
0/
#527350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#527360000000
0!
0'
0/
#527370000000
1!
1'
1/
#527380000000
0!
0'
0/
#527390000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#527400000000
0!
0'
0/
#527410000000
1!
1'
1/
#527420000000
0!
0'
0/
#527430000000
1!
1'
1/
#527440000000
0!
0'
0/
#527450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#527460000000
0!
0'
0/
#527470000000
1!
1'
1/
#527480000000
0!
0'
0/
#527490000000
1!
1'
1/
#527500000000
0!
0'
0/
#527510000000
1!
1'
1/
#527520000000
0!
0'
0/
#527530000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#527540000000
0!
0'
0/
#527550000000
1!
1'
1/
#527560000000
0!
0'
0/
#527570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#527580000000
0!
0'
0/
#527590000000
1!
1'
1/
#527600000000
0!
0'
0/
#527610000000
#527620000000
1!
1'
1/
#527630000000
0!
0'
0/
#527640000000
1!
1'
1/
#527650000000
0!
1"
0'
1(
0/
10
#527660000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#527670000000
0!
0'
0/
#527680000000
1!
1'
1/
#527690000000
0!
0'
0/
#527700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#527710000000
0!
0'
0/
#527720000000
1!
1'
1/
#527730000000
0!
1"
0'
1(
0/
10
#527740000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#527750000000
0!
1$
0'
1+
0/
#527760000000
1!
1'
1/
#527770000000
0!
0'
0/
#527780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#527790000000
0!
0'
0/
#527800000000
1!
1'
1/
#527810000000
0!
0'
0/
#527820000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#527830000000
0!
0'
0/
#527840000000
1!
1'
1/
#527850000000
0!
0'
0/
#527860000000
1!
1'
1/
#527870000000
0!
0'
0/
#527880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#527890000000
0!
0'
0/
#527900000000
1!
1'
1/
#527910000000
0!
0'
0/
#527920000000
1!
1'
1/
#527930000000
0!
0'
0/
#527940000000
1!
1'
1/
#527950000000
0!
0'
0/
#527960000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#527970000000
0!
0'
0/
#527980000000
1!
1'
1/
#527990000000
0!
0'
0/
#528000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#528010000000
0!
0'
0/
#528020000000
1!
1'
1/
#528030000000
0!
0'
0/
#528040000000
#528050000000
1!
1'
1/
#528060000000
0!
0'
0/
#528070000000
1!
1'
1/
#528080000000
0!
1"
0'
1(
0/
10
#528090000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#528100000000
0!
0'
0/
#528110000000
1!
1'
1/
#528120000000
0!
0'
0/
#528130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#528140000000
0!
0'
0/
#528150000000
1!
1'
1/
#528160000000
0!
1"
0'
1(
0/
10
#528170000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#528180000000
0!
1$
0'
1+
0/
#528190000000
1!
1'
1/
#528200000000
0!
0'
0/
#528210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#528220000000
0!
0'
0/
#528230000000
1!
1'
1/
#528240000000
0!
0'
0/
#528250000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#528260000000
0!
0'
0/
#528270000000
1!
1'
1/
#528280000000
0!
0'
0/
#528290000000
1!
1'
1/
#528300000000
0!
0'
0/
#528310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#528320000000
0!
0'
0/
#528330000000
1!
1'
1/
#528340000000
0!
0'
0/
#528350000000
1!
1'
1/
#528360000000
0!
0'
0/
#528370000000
1!
1'
1/
#528380000000
0!
0'
0/
#528390000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#528400000000
0!
0'
0/
#528410000000
1!
1'
1/
#528420000000
0!
0'
0/
#528430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#528440000000
0!
0'
0/
#528450000000
1!
1'
1/
#528460000000
0!
0'
0/
#528470000000
#528480000000
1!
1'
1/
#528490000000
0!
0'
0/
#528500000000
1!
1'
1/
#528510000000
0!
1"
0'
1(
0/
10
#528520000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#528530000000
0!
0'
0/
#528540000000
1!
1'
1/
#528550000000
0!
0'
0/
#528560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#528570000000
0!
0'
0/
#528580000000
1!
1'
1/
#528590000000
0!
1"
0'
1(
0/
10
#528600000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#528610000000
0!
1$
0'
1+
0/
#528620000000
1!
1'
1/
#528630000000
0!
0'
0/
#528640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#528650000000
0!
0'
0/
#528660000000
1!
1'
1/
#528670000000
0!
0'
0/
#528680000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#528690000000
0!
0'
0/
#528700000000
1!
1'
1/
#528710000000
0!
0'
0/
#528720000000
1!
1'
1/
#528730000000
0!
0'
0/
#528740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#528750000000
0!
0'
0/
#528760000000
1!
1'
1/
#528770000000
0!
0'
0/
#528780000000
1!
1'
1/
#528790000000
0!
0'
0/
#528800000000
1!
1'
1/
#528810000000
0!
0'
0/
#528820000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#528830000000
0!
0'
0/
#528840000000
1!
1'
1/
#528850000000
0!
0'
0/
#528860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#528870000000
0!
0'
0/
#528880000000
1!
1'
1/
#528890000000
0!
0'
0/
#528900000000
#528910000000
1!
1'
1/
#528920000000
0!
0'
0/
#528930000000
1!
1'
1/
#528940000000
0!
1"
0'
1(
0/
10
#528950000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#528960000000
0!
0'
0/
#528970000000
1!
1'
1/
#528980000000
0!
0'
0/
#528990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#529000000000
0!
0'
0/
#529010000000
1!
1'
1/
#529020000000
0!
1"
0'
1(
0/
10
#529030000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#529040000000
0!
1$
0'
1+
0/
#529050000000
1!
1'
1/
#529060000000
0!
0'
0/
#529070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#529080000000
0!
0'
0/
#529090000000
1!
1'
1/
#529100000000
0!
0'
0/
#529110000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#529120000000
0!
0'
0/
#529130000000
1!
1'
1/
#529140000000
0!
0'
0/
#529150000000
1!
1'
1/
#529160000000
0!
0'
0/
#529170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#529180000000
0!
0'
0/
#529190000000
1!
1'
1/
#529200000000
0!
0'
0/
#529210000000
1!
1'
1/
#529220000000
0!
0'
0/
#529230000000
1!
1'
1/
#529240000000
0!
0'
0/
#529250000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#529260000000
0!
0'
0/
#529270000000
1!
1'
1/
#529280000000
0!
0'
0/
#529290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#529300000000
0!
0'
0/
#529310000000
1!
1'
1/
#529320000000
0!
0'
0/
#529330000000
#529340000000
1!
1'
1/
#529350000000
0!
0'
0/
#529360000000
1!
1'
1/
#529370000000
0!
1"
0'
1(
0/
10
#529380000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#529390000000
0!
0'
0/
#529400000000
1!
1'
1/
#529410000000
0!
0'
0/
#529420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#529430000000
0!
0'
0/
#529440000000
1!
1'
1/
#529450000000
0!
1"
0'
1(
0/
10
#529460000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#529470000000
0!
1$
0'
1+
0/
#529480000000
1!
1'
1/
#529490000000
0!
0'
0/
#529500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#529510000000
0!
0'
0/
#529520000000
1!
1'
1/
#529530000000
0!
0'
0/
#529540000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#529550000000
0!
0'
0/
#529560000000
1!
1'
1/
#529570000000
0!
0'
0/
#529580000000
1!
1'
1/
#529590000000
0!
0'
0/
#529600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#529610000000
0!
0'
0/
#529620000000
1!
1'
1/
#529630000000
0!
0'
0/
#529640000000
1!
1'
1/
#529650000000
0!
0'
0/
#529660000000
1!
1'
1/
#529670000000
0!
0'
0/
#529680000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#529690000000
0!
0'
0/
#529700000000
1!
1'
1/
#529710000000
0!
0'
0/
#529720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#529730000000
0!
0'
0/
#529740000000
1!
1'
1/
#529750000000
0!
0'
0/
#529760000000
#529770000000
1!
1'
1/
#529780000000
0!
0'
0/
#529790000000
1!
1'
1/
#529800000000
0!
1"
0'
1(
0/
10
#529810000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#529820000000
0!
0'
0/
#529830000000
1!
1'
1/
#529840000000
0!
0'
0/
#529850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#529860000000
0!
0'
0/
#529870000000
1!
1'
1/
#529880000000
0!
1"
0'
1(
0/
10
#529890000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#529900000000
0!
1$
0'
1+
0/
#529910000000
1!
1'
1/
#529920000000
0!
0'
0/
#529930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#529940000000
0!
0'
0/
#529950000000
1!
1'
1/
#529960000000
0!
0'
0/
#529970000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#529980000000
0!
0'
0/
#529990000000
1!
1'
1/
#530000000000
0!
0'
0/
#530010000000
1!
1'
1/
#530020000000
0!
0'
0/
#530030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#530040000000
0!
0'
0/
#530050000000
1!
1'
1/
#530060000000
0!
0'
0/
#530070000000
1!
1'
1/
#530080000000
0!
0'
0/
#530090000000
1!
1'
1/
#530100000000
0!
0'
0/
#530110000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#530120000000
0!
0'
0/
#530130000000
1!
1'
1/
#530140000000
0!
0'
0/
#530150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#530160000000
0!
0'
0/
#530170000000
1!
1'
1/
#530180000000
0!
0'
0/
#530190000000
#530200000000
1!
1'
1/
#530210000000
0!
0'
0/
#530220000000
1!
1'
1/
#530230000000
0!
1"
0'
1(
0/
10
#530240000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#530250000000
0!
0'
0/
#530260000000
1!
1'
1/
#530270000000
0!
0'
0/
#530280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#530290000000
0!
0'
0/
#530300000000
1!
1'
1/
#530310000000
0!
1"
0'
1(
0/
10
#530320000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#530330000000
0!
1$
0'
1+
0/
#530340000000
1!
1'
1/
#530350000000
0!
0'
0/
#530360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#530370000000
0!
0'
0/
#530380000000
1!
1'
1/
#530390000000
0!
0'
0/
#530400000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#530410000000
0!
0'
0/
#530420000000
1!
1'
1/
#530430000000
0!
0'
0/
#530440000000
1!
1'
1/
#530450000000
0!
0'
0/
#530460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#530470000000
0!
0'
0/
#530480000000
1!
1'
1/
#530490000000
0!
0'
0/
#530500000000
1!
1'
1/
#530510000000
0!
0'
0/
#530520000000
1!
1'
1/
#530530000000
0!
0'
0/
#530540000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#530550000000
0!
0'
0/
#530560000000
1!
1'
1/
#530570000000
0!
0'
0/
#530580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#530590000000
0!
0'
0/
#530600000000
1!
1'
1/
#530610000000
0!
0'
0/
#530620000000
#530630000000
1!
1'
1/
#530640000000
0!
0'
0/
#530650000000
1!
1'
1/
#530660000000
0!
1"
0'
1(
0/
10
#530670000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#530680000000
0!
0'
0/
#530690000000
1!
1'
1/
#530700000000
0!
0'
0/
#530710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#530720000000
0!
0'
0/
#530730000000
1!
1'
1/
#530740000000
0!
1"
0'
1(
0/
10
#530750000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#530760000000
0!
1$
0'
1+
0/
#530770000000
1!
1'
1/
#530780000000
0!
0'
0/
#530790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#530800000000
0!
0'
0/
#530810000000
1!
1'
1/
#530820000000
0!
0'
0/
#530830000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#530840000000
0!
0'
0/
#530850000000
1!
1'
1/
#530860000000
0!
0'
0/
#530870000000
1!
1'
1/
#530880000000
0!
0'
0/
#530890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#530900000000
0!
0'
0/
#530910000000
1!
1'
1/
#530920000000
0!
0'
0/
#530930000000
1!
1'
1/
#530940000000
0!
0'
0/
#530950000000
1!
1'
1/
#530960000000
0!
0'
0/
#530970000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#530980000000
0!
0'
0/
#530990000000
1!
1'
1/
#531000000000
0!
0'
0/
#531010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#531020000000
0!
0'
0/
#531030000000
1!
1'
1/
#531040000000
0!
0'
0/
#531050000000
#531060000000
1!
1'
1/
#531070000000
0!
0'
0/
#531080000000
1!
1'
1/
#531090000000
0!
1"
0'
1(
0/
10
#531100000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#531110000000
0!
0'
0/
#531120000000
1!
1'
1/
#531130000000
0!
0'
0/
#531140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#531150000000
0!
0'
0/
#531160000000
1!
1'
1/
#531170000000
0!
1"
0'
1(
0/
10
#531180000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#531190000000
0!
1$
0'
1+
0/
#531200000000
1!
1'
1/
#531210000000
0!
0'
0/
#531220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#531230000000
0!
0'
0/
#531240000000
1!
1'
1/
#531250000000
0!
0'
0/
#531260000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#531270000000
0!
0'
0/
#531280000000
1!
1'
1/
#531290000000
0!
0'
0/
#531300000000
1!
1'
1/
#531310000000
0!
0'
0/
#531320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#531330000000
0!
0'
0/
#531340000000
1!
1'
1/
#531350000000
0!
0'
0/
#531360000000
1!
1'
1/
#531370000000
0!
0'
0/
#531380000000
1!
1'
1/
#531390000000
0!
0'
0/
#531400000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#531410000000
0!
0'
0/
#531420000000
1!
1'
1/
#531430000000
0!
0'
0/
#531440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#531450000000
0!
0'
0/
#531460000000
1!
1'
1/
#531470000000
0!
0'
0/
#531480000000
#531490000000
1!
1'
1/
#531500000000
0!
0'
0/
#531510000000
1!
1'
1/
#531520000000
0!
1"
0'
1(
0/
10
#531530000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#531540000000
0!
0'
0/
#531550000000
1!
1'
1/
#531560000000
0!
0'
0/
#531570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#531580000000
0!
0'
0/
#531590000000
1!
1'
1/
#531600000000
0!
1"
0'
1(
0/
10
#531610000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#531620000000
0!
1$
0'
1+
0/
#531630000000
1!
1'
1/
#531640000000
0!
0'
0/
#531650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#531660000000
0!
0'
0/
#531670000000
1!
1'
1/
#531680000000
0!
0'
0/
#531690000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#531700000000
0!
0'
0/
#531710000000
1!
1'
1/
#531720000000
0!
0'
0/
#531730000000
1!
1'
1/
#531740000000
0!
0'
0/
#531750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#531760000000
0!
0'
0/
#531770000000
1!
1'
1/
#531780000000
0!
0'
0/
#531790000000
1!
1'
1/
#531800000000
0!
0'
0/
#531810000000
1!
1'
1/
#531820000000
0!
0'
0/
#531830000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#531840000000
0!
0'
0/
#531850000000
1!
1'
1/
#531860000000
0!
0'
0/
#531870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#531880000000
0!
0'
0/
#531890000000
1!
1'
1/
#531900000000
0!
0'
0/
#531910000000
#531920000000
1!
1'
1/
#531930000000
0!
0'
0/
#531940000000
1!
1'
1/
#531950000000
0!
1"
0'
1(
0/
10
#531960000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#531970000000
0!
0'
0/
#531980000000
1!
1'
1/
#531990000000
0!
0'
0/
#532000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#532010000000
0!
0'
0/
#532020000000
1!
1'
1/
#532030000000
0!
1"
0'
1(
0/
10
#532040000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#532050000000
0!
1$
0'
1+
0/
#532060000000
1!
1'
1/
#532070000000
0!
0'
0/
#532080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#532090000000
0!
0'
0/
#532100000000
1!
1'
1/
#532110000000
0!
0'
0/
#532120000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#532130000000
0!
0'
0/
#532140000000
1!
1'
1/
#532150000000
0!
0'
0/
#532160000000
1!
1'
1/
#532170000000
0!
0'
0/
#532180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#532190000000
0!
0'
0/
#532200000000
1!
1'
1/
#532210000000
0!
0'
0/
#532220000000
1!
1'
1/
#532230000000
0!
0'
0/
#532240000000
1!
1'
1/
#532250000000
0!
0'
0/
#532260000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#532270000000
0!
0'
0/
#532280000000
1!
1'
1/
#532290000000
0!
0'
0/
#532300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#532310000000
0!
0'
0/
#532320000000
1!
1'
1/
#532330000000
0!
0'
0/
#532340000000
#532350000000
1!
1'
1/
#532360000000
0!
0'
0/
#532370000000
1!
1'
1/
#532380000000
0!
1"
0'
1(
0/
10
#532390000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#532400000000
0!
0'
0/
#532410000000
1!
1'
1/
#532420000000
0!
0'
0/
#532430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#532440000000
0!
0'
0/
#532450000000
1!
1'
1/
#532460000000
0!
1"
0'
1(
0/
10
#532470000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#532480000000
0!
1$
0'
1+
0/
#532490000000
1!
1'
1/
#532500000000
0!
0'
0/
#532510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#532520000000
0!
0'
0/
#532530000000
1!
1'
1/
#532540000000
0!
0'
0/
#532550000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#532560000000
0!
0'
0/
#532570000000
1!
1'
1/
#532580000000
0!
0'
0/
#532590000000
1!
1'
1/
#532600000000
0!
0'
0/
#532610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#532620000000
0!
0'
0/
#532630000000
1!
1'
1/
#532640000000
0!
0'
0/
#532650000000
1!
1'
1/
#532660000000
0!
0'
0/
#532670000000
1!
1'
1/
#532680000000
0!
0'
0/
#532690000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#532700000000
0!
0'
0/
#532710000000
1!
1'
1/
#532720000000
0!
0'
0/
#532730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#532740000000
0!
0'
0/
#532750000000
1!
1'
1/
#532760000000
0!
0'
0/
#532770000000
#532780000000
1!
1'
1/
#532790000000
0!
0'
0/
#532800000000
1!
1'
1/
#532810000000
0!
1"
0'
1(
0/
10
#532820000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#532830000000
0!
0'
0/
#532840000000
1!
1'
1/
#532850000000
0!
0'
0/
#532860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#532870000000
0!
0'
0/
#532880000000
1!
1'
1/
#532890000000
0!
1"
0'
1(
0/
10
#532900000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#532910000000
0!
1$
0'
1+
0/
#532920000000
1!
1'
1/
#532930000000
0!
0'
0/
#532940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#532950000000
0!
0'
0/
#532960000000
1!
1'
1/
#532970000000
0!
0'
0/
#532980000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#532990000000
0!
0'
0/
#533000000000
1!
1'
1/
#533010000000
0!
0'
0/
#533020000000
1!
1'
1/
#533030000000
0!
0'
0/
#533040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#533050000000
0!
0'
0/
#533060000000
1!
1'
1/
#533070000000
0!
0'
0/
#533080000000
1!
1'
1/
#533090000000
0!
0'
0/
#533100000000
1!
1'
1/
#533110000000
0!
0'
0/
#533120000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#533130000000
0!
0'
0/
#533140000000
1!
1'
1/
#533150000000
0!
0'
0/
#533160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#533170000000
0!
0'
0/
#533180000000
1!
1'
1/
#533190000000
0!
0'
0/
#533200000000
#533210000000
1!
1'
1/
#533220000000
0!
0'
0/
#533230000000
1!
1'
1/
#533240000000
0!
1"
0'
1(
0/
10
#533250000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#533260000000
0!
0'
0/
#533270000000
1!
1'
1/
#533280000000
0!
0'
0/
#533290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#533300000000
0!
0'
0/
#533310000000
1!
1'
1/
#533320000000
0!
1"
0'
1(
0/
10
#533330000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#533340000000
0!
1$
0'
1+
0/
#533350000000
1!
1'
1/
#533360000000
0!
0'
0/
#533370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#533380000000
0!
0'
0/
#533390000000
1!
1'
1/
#533400000000
0!
0'
0/
#533410000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#533420000000
0!
0'
0/
#533430000000
1!
1'
1/
#533440000000
0!
0'
0/
#533450000000
1!
1'
1/
#533460000000
0!
0'
0/
#533470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#533480000000
0!
0'
0/
#533490000000
1!
1'
1/
#533500000000
0!
0'
0/
#533510000000
1!
1'
1/
#533520000000
0!
0'
0/
#533530000000
1!
1'
1/
#533540000000
0!
0'
0/
#533550000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#533560000000
0!
0'
0/
#533570000000
1!
1'
1/
#533580000000
0!
0'
0/
#533590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#533600000000
0!
0'
0/
#533610000000
1!
1'
1/
#533620000000
0!
0'
0/
#533630000000
#533640000000
1!
1'
1/
#533650000000
0!
0'
0/
#533660000000
1!
1'
1/
#533670000000
0!
1"
0'
1(
0/
10
#533680000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#533690000000
0!
0'
0/
#533700000000
1!
1'
1/
#533710000000
0!
0'
0/
#533720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#533730000000
0!
0'
0/
#533740000000
1!
1'
1/
#533750000000
0!
1"
0'
1(
0/
10
#533760000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#533770000000
0!
1$
0'
1+
0/
#533780000000
1!
1'
1/
#533790000000
0!
0'
0/
#533800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#533810000000
0!
0'
0/
#533820000000
1!
1'
1/
#533830000000
0!
0'
0/
#533840000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#533850000000
0!
0'
0/
#533860000000
1!
1'
1/
#533870000000
0!
0'
0/
#533880000000
1!
1'
1/
#533890000000
0!
0'
0/
#533900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#533910000000
0!
0'
0/
#533920000000
1!
1'
1/
#533930000000
0!
0'
0/
#533940000000
1!
1'
1/
#533950000000
0!
0'
0/
#533960000000
1!
1'
1/
#533970000000
0!
0'
0/
#533980000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#533990000000
0!
0'
0/
#534000000000
1!
1'
1/
#534010000000
0!
0'
0/
#534020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#534030000000
0!
0'
0/
#534040000000
1!
1'
1/
#534050000000
0!
0'
0/
#534060000000
#534070000000
1!
1'
1/
#534080000000
0!
0'
0/
#534090000000
1!
1'
1/
#534100000000
0!
1"
0'
1(
0/
10
#534110000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#534120000000
0!
0'
0/
#534130000000
1!
1'
1/
#534140000000
0!
0'
0/
#534150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#534160000000
0!
0'
0/
#534170000000
1!
1'
1/
#534180000000
0!
1"
0'
1(
0/
10
#534190000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#534200000000
0!
1$
0'
1+
0/
#534210000000
1!
1'
1/
#534220000000
0!
0'
0/
#534230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#534240000000
0!
0'
0/
#534250000000
1!
1'
1/
#534260000000
0!
0'
0/
#534270000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#534280000000
0!
0'
0/
#534290000000
1!
1'
1/
#534300000000
0!
0'
0/
#534310000000
1!
1'
1/
#534320000000
0!
0'
0/
#534330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#534340000000
0!
0'
0/
#534350000000
1!
1'
1/
#534360000000
0!
0'
0/
#534370000000
1!
1'
1/
#534380000000
0!
0'
0/
#534390000000
1!
1'
1/
#534400000000
0!
0'
0/
#534410000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#534420000000
0!
0'
0/
#534430000000
1!
1'
1/
#534440000000
0!
0'
0/
#534450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#534460000000
0!
0'
0/
#534470000000
1!
1'
1/
#534480000000
0!
0'
0/
#534490000000
#534500000000
1!
1'
1/
#534510000000
0!
0'
0/
#534520000000
1!
1'
1/
#534530000000
0!
1"
0'
1(
0/
10
#534540000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#534550000000
0!
0'
0/
#534560000000
1!
1'
1/
#534570000000
0!
0'
0/
#534580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#534590000000
0!
0'
0/
#534600000000
1!
1'
1/
#534610000000
0!
1"
0'
1(
0/
10
#534620000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#534630000000
0!
1$
0'
1+
0/
#534640000000
1!
1'
1/
#534650000000
0!
0'
0/
#534660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#534670000000
0!
0'
0/
#534680000000
1!
1'
1/
#534690000000
0!
0'
0/
#534700000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#534710000000
0!
0'
0/
#534720000000
1!
1'
1/
#534730000000
0!
0'
0/
#534740000000
1!
1'
1/
#534750000000
0!
0'
0/
#534760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#534770000000
0!
0'
0/
#534780000000
1!
1'
1/
#534790000000
0!
0'
0/
#534800000000
1!
1'
1/
#534810000000
0!
0'
0/
#534820000000
1!
1'
1/
#534830000000
0!
0'
0/
#534840000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#534850000000
0!
0'
0/
#534860000000
1!
1'
1/
#534870000000
0!
0'
0/
#534880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#534890000000
0!
0'
0/
#534900000000
1!
1'
1/
#534910000000
0!
0'
0/
#534920000000
#534930000000
1!
1'
1/
#534940000000
0!
0'
0/
#534950000000
1!
1'
1/
#534960000000
0!
1"
0'
1(
0/
10
#534970000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#534980000000
0!
0'
0/
#534990000000
1!
1'
1/
#535000000000
0!
0'
0/
#535010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#535020000000
0!
0'
0/
#535030000000
1!
1'
1/
#535040000000
0!
1"
0'
1(
0/
10
#535050000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#535060000000
0!
1$
0'
1+
0/
#535070000000
1!
1'
1/
#535080000000
0!
0'
0/
#535090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#535100000000
0!
0'
0/
#535110000000
1!
1'
1/
#535120000000
0!
0'
0/
#535130000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#535140000000
0!
0'
0/
#535150000000
1!
1'
1/
#535160000000
0!
0'
0/
#535170000000
1!
1'
1/
#535180000000
0!
0'
0/
#535190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#535200000000
0!
0'
0/
#535210000000
1!
1'
1/
#535220000000
0!
0'
0/
#535230000000
1!
1'
1/
#535240000000
0!
0'
0/
#535250000000
1!
1'
1/
#535260000000
0!
0'
0/
#535270000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#535280000000
0!
0'
0/
#535290000000
1!
1'
1/
#535300000000
0!
0'
0/
#535310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#535320000000
0!
0'
0/
#535330000000
1!
1'
1/
#535340000000
0!
0'
0/
#535350000000
#535360000000
1!
1'
1/
#535370000000
0!
0'
0/
#535380000000
1!
1'
1/
#535390000000
0!
1"
0'
1(
0/
10
#535400000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#535410000000
0!
0'
0/
#535420000000
1!
1'
1/
#535430000000
0!
0'
0/
#535440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#535450000000
0!
0'
0/
#535460000000
1!
1'
1/
#535470000000
0!
1"
0'
1(
0/
10
#535480000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#535490000000
0!
1$
0'
1+
0/
#535500000000
1!
1'
1/
#535510000000
0!
0'
0/
#535520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#535530000000
0!
0'
0/
#535540000000
1!
1'
1/
#535550000000
0!
0'
0/
#535560000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#535570000000
0!
0'
0/
#535580000000
1!
1'
1/
#535590000000
0!
0'
0/
#535600000000
1!
1'
1/
#535610000000
0!
0'
0/
#535620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#535630000000
0!
0'
0/
#535640000000
1!
1'
1/
#535650000000
0!
0'
0/
#535660000000
1!
1'
1/
#535670000000
0!
0'
0/
#535680000000
1!
1'
1/
#535690000000
0!
0'
0/
#535700000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#535710000000
0!
0'
0/
#535720000000
1!
1'
1/
#535730000000
0!
0'
0/
#535740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#535750000000
0!
0'
0/
#535760000000
1!
1'
1/
#535770000000
0!
0'
0/
#535780000000
#535790000000
1!
1'
1/
#535800000000
0!
0'
0/
#535810000000
1!
1'
1/
#535820000000
0!
1"
0'
1(
0/
10
#535830000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#535840000000
0!
0'
0/
#535850000000
1!
1'
1/
#535860000000
0!
0'
0/
#535870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#535880000000
0!
0'
0/
#535890000000
1!
1'
1/
#535900000000
0!
1"
0'
1(
0/
10
#535910000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#535920000000
0!
1$
0'
1+
0/
#535930000000
1!
1'
1/
#535940000000
0!
0'
0/
#535950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#535960000000
0!
0'
0/
#535970000000
1!
1'
1/
#535980000000
0!
0'
0/
#535990000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#536000000000
0!
0'
0/
#536010000000
1!
1'
1/
#536020000000
0!
0'
0/
#536030000000
1!
1'
1/
#536040000000
0!
0'
0/
#536050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#536060000000
0!
0'
0/
#536070000000
1!
1'
1/
#536080000000
0!
0'
0/
#536090000000
1!
1'
1/
#536100000000
0!
0'
0/
#536110000000
1!
1'
1/
#536120000000
0!
0'
0/
#536130000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#536140000000
0!
0'
0/
#536150000000
1!
1'
1/
#536160000000
0!
0'
0/
#536170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#536180000000
0!
0'
0/
#536190000000
1!
1'
1/
#536200000000
0!
0'
0/
#536210000000
#536220000000
1!
1'
1/
#536230000000
0!
0'
0/
#536240000000
1!
1'
1/
#536250000000
0!
1"
0'
1(
0/
10
#536260000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#536270000000
0!
0'
0/
#536280000000
1!
1'
1/
#536290000000
0!
0'
0/
#536300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#536310000000
0!
0'
0/
#536320000000
1!
1'
1/
#536330000000
0!
1"
0'
1(
0/
10
#536340000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#536350000000
0!
1$
0'
1+
0/
#536360000000
1!
1'
1/
#536370000000
0!
0'
0/
#536380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#536390000000
0!
0'
0/
#536400000000
1!
1'
1/
#536410000000
0!
0'
0/
#536420000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#536430000000
0!
0'
0/
#536440000000
1!
1'
1/
#536450000000
0!
0'
0/
#536460000000
1!
1'
1/
#536470000000
0!
0'
0/
#536480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#536490000000
0!
0'
0/
#536500000000
1!
1'
1/
#536510000000
0!
0'
0/
#536520000000
1!
1'
1/
#536530000000
0!
0'
0/
#536540000000
1!
1'
1/
#536550000000
0!
0'
0/
#536560000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#536570000000
0!
0'
0/
#536580000000
1!
1'
1/
#536590000000
0!
0'
0/
#536600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#536610000000
0!
0'
0/
#536620000000
1!
1'
1/
#536630000000
0!
0'
0/
#536640000000
#536650000000
1!
1'
1/
#536660000000
0!
0'
0/
#536670000000
1!
1'
1/
#536680000000
0!
1"
0'
1(
0/
10
#536690000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#536700000000
0!
0'
0/
#536710000000
1!
1'
1/
#536720000000
0!
0'
0/
#536730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#536740000000
0!
0'
0/
#536750000000
1!
1'
1/
#536760000000
0!
1"
0'
1(
0/
10
#536770000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#536780000000
0!
1$
0'
1+
0/
#536790000000
1!
1'
1/
#536800000000
0!
0'
0/
#536810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#536820000000
0!
0'
0/
#536830000000
1!
1'
1/
#536840000000
0!
0'
0/
#536850000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#536860000000
0!
0'
0/
#536870000000
1!
1'
1/
#536880000000
0!
0'
0/
#536890000000
1!
1'
1/
#536900000000
0!
0'
0/
#536910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#536920000000
0!
0'
0/
#536930000000
1!
1'
1/
#536940000000
0!
0'
0/
#536950000000
1!
1'
1/
#536960000000
0!
0'
0/
#536970000000
1!
1'
1/
#536980000000
0!
0'
0/
#536990000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#537000000000
0!
0'
0/
#537010000000
1!
1'
1/
#537020000000
0!
0'
0/
#537030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#537040000000
0!
0'
0/
#537050000000
1!
1'
1/
#537060000000
0!
0'
0/
#537070000000
#537080000000
1!
1'
1/
#537090000000
0!
0'
0/
#537100000000
1!
1'
1/
#537110000000
0!
1"
0'
1(
0/
10
#537120000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#537130000000
0!
0'
0/
#537140000000
1!
1'
1/
#537150000000
0!
0'
0/
#537160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#537170000000
0!
0'
0/
#537180000000
1!
1'
1/
#537190000000
0!
1"
0'
1(
0/
10
#537200000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#537210000000
0!
1$
0'
1+
0/
#537220000000
1!
1'
1/
#537230000000
0!
0'
0/
#537240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#537250000000
0!
0'
0/
#537260000000
1!
1'
1/
#537270000000
0!
0'
0/
#537280000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#537290000000
0!
0'
0/
#537300000000
1!
1'
1/
#537310000000
0!
0'
0/
#537320000000
1!
1'
1/
#537330000000
0!
0'
0/
#537340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#537350000000
0!
0'
0/
#537360000000
1!
1'
1/
#537370000000
0!
0'
0/
#537380000000
1!
1'
1/
#537390000000
0!
0'
0/
#537400000000
1!
1'
1/
#537410000000
0!
0'
0/
#537420000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#537430000000
0!
0'
0/
#537440000000
1!
1'
1/
#537450000000
0!
0'
0/
#537460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#537470000000
0!
0'
0/
#537480000000
1!
1'
1/
#537490000000
0!
0'
0/
#537500000000
#537510000000
1!
1'
1/
#537520000000
0!
0'
0/
#537530000000
1!
1'
1/
#537540000000
0!
1"
0'
1(
0/
10
#537550000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#537560000000
0!
0'
0/
#537570000000
1!
1'
1/
#537580000000
0!
0'
0/
#537590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#537600000000
0!
0'
0/
#537610000000
1!
1'
1/
#537620000000
0!
1"
0'
1(
0/
10
#537630000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#537640000000
0!
1$
0'
1+
0/
#537650000000
1!
1'
1/
#537660000000
0!
0'
0/
#537670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#537680000000
0!
0'
0/
#537690000000
1!
1'
1/
#537700000000
0!
0'
0/
#537710000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#537720000000
0!
0'
0/
#537730000000
1!
1'
1/
#537740000000
0!
0'
0/
#537750000000
1!
1'
1/
#537760000000
0!
0'
0/
#537770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#537780000000
0!
0'
0/
#537790000000
1!
1'
1/
#537800000000
0!
0'
0/
#537810000000
1!
1'
1/
#537820000000
0!
0'
0/
#537830000000
1!
1'
1/
#537840000000
0!
0'
0/
#537850000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#537860000000
0!
0'
0/
#537870000000
1!
1'
1/
#537880000000
0!
0'
0/
#537890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#537900000000
0!
0'
0/
#537910000000
1!
1'
1/
#537920000000
0!
0'
0/
#537930000000
#537940000000
1!
1'
1/
#537950000000
0!
0'
0/
#537960000000
1!
1'
1/
#537970000000
0!
1"
0'
1(
0/
10
#537980000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#537990000000
0!
0'
0/
#538000000000
1!
1'
1/
#538010000000
0!
0'
0/
#538020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#538030000000
0!
0'
0/
#538040000000
1!
1'
1/
#538050000000
0!
1"
0'
1(
0/
10
#538060000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#538070000000
0!
1$
0'
1+
0/
#538080000000
1!
1'
1/
#538090000000
0!
0'
0/
#538100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#538110000000
0!
0'
0/
#538120000000
1!
1'
1/
#538130000000
0!
0'
0/
#538140000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#538150000000
0!
0'
0/
#538160000000
1!
1'
1/
#538170000000
0!
0'
0/
#538180000000
1!
1'
1/
#538190000000
0!
0'
0/
#538200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#538210000000
0!
0'
0/
#538220000000
1!
1'
1/
#538230000000
0!
0'
0/
#538240000000
1!
1'
1/
#538250000000
0!
0'
0/
#538260000000
1!
1'
1/
#538270000000
0!
0'
0/
#538280000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#538290000000
0!
0'
0/
#538300000000
1!
1'
1/
#538310000000
0!
0'
0/
#538320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#538330000000
0!
0'
0/
#538340000000
1!
1'
1/
#538350000000
0!
0'
0/
#538360000000
#538370000000
1!
1'
1/
#538380000000
0!
0'
0/
#538390000000
1!
1'
1/
#538400000000
0!
1"
0'
1(
0/
10
#538410000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#538420000000
0!
0'
0/
#538430000000
1!
1'
1/
#538440000000
0!
0'
0/
#538450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#538460000000
0!
0'
0/
#538470000000
1!
1'
1/
#538480000000
0!
1"
0'
1(
0/
10
#538490000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#538500000000
0!
1$
0'
1+
0/
#538510000000
1!
1'
1/
#538520000000
0!
0'
0/
#538530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#538540000000
0!
0'
0/
#538550000000
1!
1'
1/
#538560000000
0!
0'
0/
#538570000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#538580000000
0!
0'
0/
#538590000000
1!
1'
1/
#538600000000
0!
0'
0/
#538610000000
1!
1'
1/
#538620000000
0!
0'
0/
#538630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#538640000000
0!
0'
0/
#538650000000
1!
1'
1/
#538660000000
0!
0'
0/
#538670000000
1!
1'
1/
#538680000000
0!
0'
0/
#538690000000
1!
1'
1/
#538700000000
0!
0'
0/
#538710000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#538720000000
0!
0'
0/
#538730000000
1!
1'
1/
#538740000000
0!
0'
0/
#538750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#538760000000
0!
0'
0/
#538770000000
1!
1'
1/
#538780000000
0!
0'
0/
#538790000000
#538800000000
1!
1'
1/
#538810000000
0!
0'
0/
#538820000000
1!
1'
1/
#538830000000
0!
1"
0'
1(
0/
10
#538840000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#538850000000
0!
0'
0/
#538860000000
1!
1'
1/
#538870000000
0!
0'
0/
#538880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#538890000000
0!
0'
0/
#538900000000
1!
1'
1/
#538910000000
0!
1"
0'
1(
0/
10
#538920000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#538930000000
0!
1$
0'
1+
0/
#538940000000
1!
1'
1/
#538950000000
0!
0'
0/
#538960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#538970000000
0!
0'
0/
#538980000000
1!
1'
1/
#538990000000
0!
0'
0/
#539000000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#539010000000
0!
0'
0/
#539020000000
1!
1'
1/
#539030000000
0!
0'
0/
#539040000000
1!
1'
1/
#539050000000
0!
0'
0/
#539060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#539070000000
0!
0'
0/
#539080000000
1!
1'
1/
#539090000000
0!
0'
0/
#539100000000
1!
1'
1/
#539110000000
0!
0'
0/
#539120000000
1!
1'
1/
#539130000000
0!
0'
0/
#539140000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#539150000000
0!
0'
0/
#539160000000
1!
1'
1/
#539170000000
0!
0'
0/
#539180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#539190000000
0!
0'
0/
#539200000000
1!
1'
1/
#539210000000
0!
0'
0/
#539220000000
#539230000000
1!
1'
1/
#539240000000
0!
0'
0/
#539250000000
1!
1'
1/
#539260000000
0!
1"
0'
1(
0/
10
#539270000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#539280000000
0!
0'
0/
#539290000000
1!
1'
1/
#539300000000
0!
0'
0/
#539310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#539320000000
0!
0'
0/
#539330000000
1!
1'
1/
#539340000000
0!
1"
0'
1(
0/
10
#539350000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#539360000000
0!
1$
0'
1+
0/
#539370000000
1!
1'
1/
#539380000000
0!
0'
0/
#539390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#539400000000
0!
0'
0/
#539410000000
1!
1'
1/
#539420000000
0!
0'
0/
#539430000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#539440000000
0!
0'
0/
#539450000000
1!
1'
1/
#539460000000
0!
0'
0/
#539470000000
1!
1'
1/
#539480000000
0!
0'
0/
#539490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#539500000000
0!
0'
0/
#539510000000
1!
1'
1/
#539520000000
0!
0'
0/
#539530000000
1!
1'
1/
#539540000000
0!
0'
0/
#539550000000
1!
1'
1/
#539560000000
0!
0'
0/
#539570000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#539580000000
0!
0'
0/
#539590000000
1!
1'
1/
#539600000000
0!
0'
0/
#539610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#539620000000
0!
0'
0/
#539630000000
1!
1'
1/
#539640000000
0!
0'
0/
#539650000000
#539660000000
1!
1'
1/
#539670000000
0!
0'
0/
#539680000000
1!
1'
1/
#539690000000
0!
1"
0'
1(
0/
10
#539700000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#539710000000
0!
0'
0/
#539720000000
1!
1'
1/
#539730000000
0!
0'
0/
#539740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#539750000000
0!
0'
0/
#539760000000
1!
1'
1/
#539770000000
0!
1"
0'
1(
0/
10
#539780000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#539790000000
0!
1$
0'
1+
0/
#539800000000
1!
1'
1/
#539810000000
0!
0'
0/
#539820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#539830000000
0!
0'
0/
#539840000000
1!
1'
1/
#539850000000
0!
0'
0/
#539860000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#539870000000
0!
0'
0/
#539880000000
1!
1'
1/
#539890000000
0!
0'
0/
#539900000000
1!
1'
1/
#539910000000
0!
0'
0/
#539920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#539930000000
0!
0'
0/
#539940000000
1!
1'
1/
#539950000000
0!
0'
0/
#539960000000
1!
1'
1/
#539970000000
0!
0'
0/
#539980000000
1!
1'
1/
#539990000000
0!
0'
0/
#540000000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#540010000000
0!
0'
0/
#540020000000
1!
1'
1/
#540030000000
0!
0'
0/
#540040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#540050000000
0!
0'
0/
#540060000000
1!
1'
1/
#540070000000
0!
0'
0/
#540080000000
#540090000000
1!
1'
1/
#540100000000
0!
0'
0/
#540110000000
1!
1'
1/
#540120000000
0!
1"
0'
1(
0/
10
#540130000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#540140000000
0!
0'
0/
#540150000000
1!
1'
1/
#540160000000
0!
0'
0/
#540170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#540180000000
0!
0'
0/
#540190000000
1!
1'
1/
#540200000000
0!
1"
0'
1(
0/
10
#540210000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#540220000000
0!
1$
0'
1+
0/
#540230000000
1!
1'
1/
#540240000000
0!
0'
0/
#540250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#540260000000
0!
0'
0/
#540270000000
1!
1'
1/
#540280000000
0!
0'
0/
#540290000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#540300000000
0!
0'
0/
#540310000000
1!
1'
1/
#540320000000
0!
0'
0/
#540330000000
1!
1'
1/
#540340000000
0!
0'
0/
#540350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#540360000000
0!
0'
0/
#540370000000
1!
1'
1/
#540380000000
0!
0'
0/
#540390000000
1!
1'
1/
#540400000000
0!
0'
0/
#540410000000
1!
1'
1/
#540420000000
0!
0'
0/
#540430000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#540440000000
0!
0'
0/
#540450000000
1!
1'
1/
#540460000000
0!
0'
0/
#540470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#540480000000
0!
0'
0/
#540490000000
1!
1'
1/
#540500000000
0!
0'
0/
#540510000000
#540520000000
1!
1'
1/
#540530000000
0!
0'
0/
#540540000000
1!
1'
1/
#540550000000
0!
1"
0'
1(
0/
10
#540560000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#540570000000
0!
0'
0/
#540580000000
1!
1'
1/
#540590000000
0!
0'
0/
#540600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#540610000000
0!
0'
0/
#540620000000
1!
1'
1/
#540630000000
0!
1"
0'
1(
0/
10
#540640000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#540650000000
0!
1$
0'
1+
0/
#540660000000
1!
1'
1/
#540670000000
0!
0'
0/
#540680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#540690000000
0!
0'
0/
#540700000000
1!
1'
1/
#540710000000
0!
0'
0/
#540720000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#540730000000
0!
0'
0/
#540740000000
1!
1'
1/
#540750000000
0!
0'
0/
#540760000000
1!
1'
1/
#540770000000
0!
0'
0/
#540780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#540790000000
0!
0'
0/
#540800000000
1!
1'
1/
#540810000000
0!
0'
0/
#540820000000
1!
1'
1/
#540830000000
0!
0'
0/
#540840000000
1!
1'
1/
#540850000000
0!
0'
0/
#540860000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#540870000000
0!
0'
0/
#540880000000
1!
1'
1/
#540890000000
0!
0'
0/
#540900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#540910000000
0!
0'
0/
#540920000000
1!
1'
1/
#540930000000
0!
0'
0/
#540940000000
#540950000000
1!
1'
1/
#540960000000
0!
0'
0/
#540970000000
1!
1'
1/
#540980000000
0!
1"
0'
1(
0/
10
#540990000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#541000000000
0!
0'
0/
#541010000000
1!
1'
1/
#541020000000
0!
0'
0/
#541030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#541040000000
0!
0'
0/
#541050000000
1!
1'
1/
#541060000000
0!
1"
0'
1(
0/
10
#541070000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#541080000000
0!
1$
0'
1+
0/
#541090000000
1!
1'
1/
#541100000000
0!
0'
0/
#541110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#541120000000
0!
0'
0/
#541130000000
1!
1'
1/
#541140000000
0!
0'
0/
#541150000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#541160000000
0!
0'
0/
#541170000000
1!
1'
1/
#541180000000
0!
0'
0/
#541190000000
1!
1'
1/
#541200000000
0!
0'
0/
#541210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#541220000000
0!
0'
0/
#541230000000
1!
1'
1/
#541240000000
0!
0'
0/
#541250000000
1!
1'
1/
#541260000000
0!
0'
0/
#541270000000
1!
1'
1/
#541280000000
0!
0'
0/
#541290000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#541300000000
0!
0'
0/
#541310000000
1!
1'
1/
#541320000000
0!
0'
0/
#541330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#541340000000
0!
0'
0/
#541350000000
1!
1'
1/
#541360000000
0!
0'
0/
#541370000000
#541380000000
1!
1'
1/
#541390000000
0!
0'
0/
#541400000000
1!
1'
1/
#541410000000
0!
1"
0'
1(
0/
10
#541420000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#541430000000
0!
0'
0/
#541440000000
1!
1'
1/
#541450000000
0!
0'
0/
#541460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#541470000000
0!
0'
0/
#541480000000
1!
1'
1/
#541490000000
0!
1"
0'
1(
0/
10
#541500000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#541510000000
0!
1$
0'
1+
0/
#541520000000
1!
1'
1/
#541530000000
0!
0'
0/
#541540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#541550000000
0!
0'
0/
#541560000000
1!
1'
1/
#541570000000
0!
0'
0/
#541580000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#541590000000
0!
0'
0/
#541600000000
1!
1'
1/
#541610000000
0!
0'
0/
#541620000000
1!
1'
1/
#541630000000
0!
0'
0/
#541640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#541650000000
0!
0'
0/
#541660000000
1!
1'
1/
#541670000000
0!
0'
0/
#541680000000
1!
1'
1/
#541690000000
0!
0'
0/
#541700000000
1!
1'
1/
#541710000000
0!
0'
0/
#541720000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#541730000000
0!
0'
0/
#541740000000
1!
1'
1/
#541750000000
0!
0'
0/
#541760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#541770000000
0!
0'
0/
#541780000000
1!
1'
1/
#541790000000
0!
0'
0/
#541800000000
#541810000000
1!
1'
1/
#541820000000
0!
0'
0/
#541830000000
1!
1'
1/
#541840000000
0!
1"
0'
1(
0/
10
#541850000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#541860000000
0!
0'
0/
#541870000000
1!
1'
1/
#541880000000
0!
0'
0/
#541890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#541900000000
0!
0'
0/
#541910000000
1!
1'
1/
#541920000000
0!
1"
0'
1(
0/
10
#541930000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#541940000000
0!
1$
0'
1+
0/
#541950000000
1!
1'
1/
#541960000000
0!
0'
0/
#541970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#541980000000
0!
0'
0/
#541990000000
1!
1'
1/
#542000000000
0!
0'
0/
#542010000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#542020000000
0!
0'
0/
#542030000000
1!
1'
1/
#542040000000
0!
0'
0/
#542050000000
1!
1'
1/
#542060000000
0!
0'
0/
#542070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#542080000000
0!
0'
0/
#542090000000
1!
1'
1/
#542100000000
0!
0'
0/
#542110000000
1!
1'
1/
#542120000000
0!
0'
0/
#542130000000
1!
1'
1/
#542140000000
0!
0'
0/
#542150000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#542160000000
0!
0'
0/
#542170000000
1!
1'
1/
#542180000000
0!
0'
0/
#542190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#542200000000
0!
0'
0/
#542210000000
1!
1'
1/
#542220000000
0!
0'
0/
#542230000000
#542240000000
1!
1'
1/
#542250000000
0!
0'
0/
#542260000000
1!
1'
1/
#542270000000
0!
1"
0'
1(
0/
10
#542280000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#542290000000
0!
0'
0/
#542300000000
1!
1'
1/
#542310000000
0!
0'
0/
#542320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#542330000000
0!
0'
0/
#542340000000
1!
1'
1/
#542350000000
0!
1"
0'
1(
0/
10
#542360000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#542370000000
0!
1$
0'
1+
0/
#542380000000
1!
1'
1/
#542390000000
0!
0'
0/
#542400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#542410000000
0!
0'
0/
#542420000000
1!
1'
1/
#542430000000
0!
0'
0/
#542440000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#542450000000
0!
0'
0/
#542460000000
1!
1'
1/
#542470000000
0!
0'
0/
#542480000000
1!
1'
1/
#542490000000
0!
0'
0/
#542500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#542510000000
0!
0'
0/
#542520000000
1!
1'
1/
#542530000000
0!
0'
0/
#542540000000
1!
1'
1/
#542550000000
0!
0'
0/
#542560000000
1!
1'
1/
#542570000000
0!
0'
0/
#542580000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#542590000000
0!
0'
0/
#542600000000
1!
1'
1/
#542610000000
0!
0'
0/
#542620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#542630000000
0!
0'
0/
#542640000000
1!
1'
1/
#542650000000
0!
0'
0/
#542660000000
#542670000000
1!
1'
1/
#542680000000
0!
0'
0/
#542690000000
1!
1'
1/
#542700000000
0!
1"
0'
1(
0/
10
#542710000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#542720000000
0!
0'
0/
#542730000000
1!
1'
1/
#542740000000
0!
0'
0/
#542750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#542760000000
0!
0'
0/
#542770000000
1!
1'
1/
#542780000000
0!
1"
0'
1(
0/
10
#542790000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#542800000000
0!
1$
0'
1+
0/
#542810000000
1!
1'
1/
#542820000000
0!
0'
0/
#542830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#542840000000
0!
0'
0/
#542850000000
1!
1'
1/
#542860000000
0!
0'
0/
#542870000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#542880000000
0!
0'
0/
#542890000000
1!
1'
1/
#542900000000
0!
0'
0/
#542910000000
1!
1'
1/
#542920000000
0!
0'
0/
#542930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#542940000000
0!
0'
0/
#542950000000
1!
1'
1/
#542960000000
0!
0'
0/
#542970000000
1!
1'
1/
#542980000000
0!
0'
0/
#542990000000
1!
1'
1/
#543000000000
0!
0'
0/
#543010000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#543020000000
0!
0'
0/
#543030000000
1!
1'
1/
#543040000000
0!
0'
0/
#543050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#543060000000
0!
0'
0/
#543070000000
1!
1'
1/
#543080000000
0!
0'
0/
#543090000000
#543100000000
1!
1'
1/
#543110000000
0!
0'
0/
#543120000000
1!
1'
1/
#543130000000
0!
1"
0'
1(
0/
10
#543140000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#543150000000
0!
0'
0/
#543160000000
1!
1'
1/
#543170000000
0!
0'
0/
#543180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#543190000000
0!
0'
0/
#543200000000
1!
1'
1/
#543210000000
0!
1"
0'
1(
0/
10
#543220000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#543230000000
0!
1$
0'
1+
0/
#543240000000
1!
1'
1/
#543250000000
0!
0'
0/
#543260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#543270000000
0!
0'
0/
#543280000000
1!
1'
1/
#543290000000
0!
0'
0/
#543300000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#543310000000
0!
0'
0/
#543320000000
1!
1'
1/
#543330000000
0!
0'
0/
#543340000000
1!
1'
1/
#543350000000
0!
0'
0/
#543360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#543370000000
0!
0'
0/
#543380000000
1!
1'
1/
#543390000000
0!
0'
0/
#543400000000
1!
1'
1/
#543410000000
0!
0'
0/
#543420000000
1!
1'
1/
#543430000000
0!
0'
0/
#543440000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#543450000000
0!
0'
0/
#543460000000
1!
1'
1/
#543470000000
0!
0'
0/
#543480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#543490000000
0!
0'
0/
#543500000000
1!
1'
1/
#543510000000
0!
0'
0/
#543520000000
#543530000000
1!
1'
1/
#543540000000
0!
0'
0/
#543550000000
1!
1'
1/
#543560000000
0!
1"
0'
1(
0/
10
#543570000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#543580000000
0!
0'
0/
#543590000000
1!
1'
1/
#543600000000
0!
0'
0/
#543610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#543620000000
0!
0'
0/
#543630000000
1!
1'
1/
#543640000000
0!
1"
0'
1(
0/
10
#543650000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#543660000000
0!
1$
0'
1+
0/
#543670000000
1!
1'
1/
#543680000000
0!
0'
0/
#543690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#543700000000
0!
0'
0/
#543710000000
1!
1'
1/
#543720000000
0!
0'
0/
#543730000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#543740000000
0!
0'
0/
#543750000000
1!
1'
1/
#543760000000
0!
0'
0/
#543770000000
1!
1'
1/
#543780000000
0!
0'
0/
#543790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#543800000000
0!
0'
0/
#543810000000
1!
1'
1/
#543820000000
0!
0'
0/
#543830000000
1!
1'
1/
#543840000000
0!
0'
0/
#543850000000
1!
1'
1/
#543860000000
0!
0'
0/
#543870000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#543880000000
0!
0'
0/
#543890000000
1!
1'
1/
#543900000000
0!
0'
0/
#543910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#543920000000
0!
0'
0/
#543930000000
1!
1'
1/
#543940000000
0!
0'
0/
#543950000000
#543960000000
1!
1'
1/
#543970000000
0!
0'
0/
#543980000000
1!
1'
1/
#543990000000
0!
1"
0'
1(
0/
10
#544000000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#544010000000
0!
0'
0/
#544020000000
1!
1'
1/
#544030000000
0!
0'
0/
#544040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#544050000000
0!
0'
0/
#544060000000
1!
1'
1/
#544070000000
0!
1"
0'
1(
0/
10
#544080000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#544090000000
0!
1$
0'
1+
0/
#544100000000
1!
1'
1/
#544110000000
0!
0'
0/
#544120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#544130000000
0!
0'
0/
#544140000000
1!
1'
1/
#544150000000
0!
0'
0/
#544160000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#544170000000
0!
0'
0/
#544180000000
1!
1'
1/
#544190000000
0!
0'
0/
#544200000000
1!
1'
1/
#544210000000
0!
0'
0/
#544220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#544230000000
0!
0'
0/
#544240000000
1!
1'
1/
#544250000000
0!
0'
0/
#544260000000
1!
1'
1/
#544270000000
0!
0'
0/
#544280000000
1!
1'
1/
#544290000000
0!
0'
0/
#544300000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#544310000000
0!
0'
0/
#544320000000
1!
1'
1/
#544330000000
0!
0'
0/
#544340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#544350000000
0!
0'
0/
#544360000000
1!
1'
1/
#544370000000
0!
0'
0/
#544380000000
#544390000000
1!
1'
1/
#544400000000
0!
0'
0/
#544410000000
1!
1'
1/
#544420000000
0!
1"
0'
1(
0/
10
#544430000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#544440000000
0!
0'
0/
#544450000000
1!
1'
1/
#544460000000
0!
0'
0/
#544470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#544480000000
0!
0'
0/
#544490000000
1!
1'
1/
#544500000000
0!
1"
0'
1(
0/
10
#544510000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#544520000000
0!
1$
0'
1+
0/
#544530000000
1!
1'
1/
#544540000000
0!
0'
0/
#544550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#544560000000
0!
0'
0/
#544570000000
1!
1'
1/
#544580000000
0!
0'
0/
#544590000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#544600000000
0!
0'
0/
#544610000000
1!
1'
1/
#544620000000
0!
0'
0/
#544630000000
1!
1'
1/
#544640000000
0!
0'
0/
#544650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#544660000000
0!
0'
0/
#544670000000
1!
1'
1/
#544680000000
0!
0'
0/
#544690000000
1!
1'
1/
#544700000000
0!
0'
0/
#544710000000
1!
1'
1/
#544720000000
0!
0'
0/
#544730000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#544740000000
0!
0'
0/
#544750000000
1!
1'
1/
#544760000000
0!
0'
0/
#544770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#544780000000
0!
0'
0/
#544790000000
1!
1'
1/
#544800000000
0!
0'
0/
#544810000000
#544820000000
1!
1'
1/
#544830000000
0!
0'
0/
#544840000000
1!
1'
1/
#544850000000
0!
1"
0'
1(
0/
10
#544860000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#544870000000
0!
0'
0/
#544880000000
1!
1'
1/
#544890000000
0!
0'
0/
#544900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#544910000000
0!
0'
0/
#544920000000
1!
1'
1/
#544930000000
0!
1"
0'
1(
0/
10
#544940000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#544950000000
0!
1$
0'
1+
0/
#544960000000
1!
1'
1/
#544970000000
0!
0'
0/
#544980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#544990000000
0!
0'
0/
#545000000000
1!
1'
1/
#545010000000
0!
0'
0/
#545020000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#545030000000
0!
0'
0/
#545040000000
1!
1'
1/
#545050000000
0!
0'
0/
#545060000000
1!
1'
1/
#545070000000
0!
0'
0/
#545080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#545090000000
0!
0'
0/
#545100000000
1!
1'
1/
#545110000000
0!
0'
0/
#545120000000
1!
1'
1/
#545130000000
0!
0'
0/
#545140000000
1!
1'
1/
#545150000000
0!
0'
0/
#545160000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#545170000000
0!
0'
0/
#545180000000
1!
1'
1/
#545190000000
0!
0'
0/
#545200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#545210000000
0!
0'
0/
#545220000000
1!
1'
1/
#545230000000
0!
0'
0/
#545240000000
#545250000000
1!
1'
1/
#545260000000
0!
0'
0/
#545270000000
1!
1'
1/
#545280000000
0!
1"
0'
1(
0/
10
#545290000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#545300000000
0!
0'
0/
#545310000000
1!
1'
1/
#545320000000
0!
0'
0/
#545330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#545340000000
0!
0'
0/
#545350000000
1!
1'
1/
#545360000000
0!
1"
0'
1(
0/
10
#545370000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#545380000000
0!
1$
0'
1+
0/
#545390000000
1!
1'
1/
#545400000000
0!
0'
0/
#545410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#545420000000
0!
0'
0/
#545430000000
1!
1'
1/
#545440000000
0!
0'
0/
#545450000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#545460000000
0!
0'
0/
#545470000000
1!
1'
1/
#545480000000
0!
0'
0/
#545490000000
1!
1'
1/
#545500000000
0!
0'
0/
#545510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#545520000000
0!
0'
0/
#545530000000
1!
1'
1/
#545540000000
0!
0'
0/
#545550000000
1!
1'
1/
#545560000000
0!
0'
0/
#545570000000
1!
1'
1/
#545580000000
0!
0'
0/
#545590000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#545600000000
0!
0'
0/
#545610000000
1!
1'
1/
#545620000000
0!
0'
0/
#545630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#545640000000
0!
0'
0/
#545650000000
1!
1'
1/
#545660000000
0!
0'
0/
#545670000000
#545680000000
1!
1'
1/
#545690000000
0!
0'
0/
#545700000000
1!
1'
1/
#545710000000
0!
1"
0'
1(
0/
10
#545720000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#545730000000
0!
0'
0/
#545740000000
1!
1'
1/
#545750000000
0!
0'
0/
#545760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#545770000000
0!
0'
0/
#545780000000
1!
1'
1/
#545790000000
0!
1"
0'
1(
0/
10
#545800000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#545810000000
0!
1$
0'
1+
0/
#545820000000
1!
1'
1/
#545830000000
0!
0'
0/
#545840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#545850000000
0!
0'
0/
#545860000000
1!
1'
1/
#545870000000
0!
0'
0/
#545880000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#545890000000
0!
0'
0/
#545900000000
1!
1'
1/
#545910000000
0!
0'
0/
#545920000000
1!
1'
1/
#545930000000
0!
0'
0/
#545940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#545950000000
0!
0'
0/
#545960000000
1!
1'
1/
#545970000000
0!
0'
0/
#545980000000
1!
1'
1/
#545990000000
0!
0'
0/
#546000000000
1!
1'
1/
#546010000000
0!
0'
0/
#546020000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#546030000000
0!
0'
0/
#546040000000
1!
1'
1/
#546050000000
0!
0'
0/
#546060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#546070000000
0!
0'
0/
#546080000000
1!
1'
1/
#546090000000
0!
0'
0/
#546100000000
#546110000000
1!
1'
1/
#546120000000
0!
0'
0/
#546130000000
1!
1'
1/
#546140000000
0!
1"
0'
1(
0/
10
#546150000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#546160000000
0!
0'
0/
#546170000000
1!
1'
1/
#546180000000
0!
0'
0/
#546190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#546200000000
0!
0'
0/
#546210000000
1!
1'
1/
#546220000000
0!
1"
0'
1(
0/
10
#546230000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#546240000000
0!
1$
0'
1+
0/
#546250000000
1!
1'
1/
#546260000000
0!
0'
0/
#546270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#546280000000
0!
0'
0/
#546290000000
1!
1'
1/
#546300000000
0!
0'
0/
#546310000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#546320000000
0!
0'
0/
#546330000000
1!
1'
1/
#546340000000
0!
0'
0/
#546350000000
1!
1'
1/
#546360000000
0!
0'
0/
#546370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#546380000000
0!
0'
0/
#546390000000
1!
1'
1/
#546400000000
0!
0'
0/
#546410000000
1!
1'
1/
#546420000000
0!
0'
0/
#546430000000
1!
1'
1/
#546440000000
0!
0'
0/
#546450000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#546460000000
0!
0'
0/
#546470000000
1!
1'
1/
#546480000000
0!
0'
0/
#546490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#546500000000
0!
0'
0/
#546510000000
1!
1'
1/
#546520000000
0!
0'
0/
#546530000000
#546540000000
1!
1'
1/
#546550000000
0!
0'
0/
#546560000000
1!
1'
1/
#546570000000
0!
1"
0'
1(
0/
10
#546580000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#546590000000
0!
0'
0/
#546600000000
1!
1'
1/
#546610000000
0!
0'
0/
#546620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#546630000000
0!
0'
0/
#546640000000
1!
1'
1/
#546650000000
0!
1"
0'
1(
0/
10
#546660000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#546670000000
0!
1$
0'
1+
0/
#546680000000
1!
1'
1/
#546690000000
0!
0'
0/
#546700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#546710000000
0!
0'
0/
#546720000000
1!
1'
1/
#546730000000
0!
0'
0/
#546740000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#546750000000
0!
0'
0/
#546760000000
1!
1'
1/
#546770000000
0!
0'
0/
#546780000000
1!
1'
1/
#546790000000
0!
0'
0/
#546800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#546810000000
0!
0'
0/
#546820000000
1!
1'
1/
#546830000000
0!
0'
0/
#546840000000
1!
1'
1/
#546850000000
0!
0'
0/
#546860000000
1!
1'
1/
#546870000000
0!
0'
0/
#546880000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#546890000000
0!
0'
0/
#546900000000
1!
1'
1/
#546910000000
0!
0'
0/
#546920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#546930000000
0!
0'
0/
#546940000000
1!
1'
1/
#546950000000
0!
0'
0/
#546960000000
#546970000000
1!
1'
1/
#546980000000
0!
0'
0/
#546990000000
1!
1'
1/
#547000000000
0!
1"
0'
1(
0/
10
#547010000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#547020000000
0!
0'
0/
#547030000000
1!
1'
1/
#547040000000
0!
0'
0/
#547050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#547060000000
0!
0'
0/
#547070000000
1!
1'
1/
#547080000000
0!
1"
0'
1(
0/
10
#547090000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#547100000000
0!
1$
0'
1+
0/
#547110000000
1!
1'
1/
#547120000000
0!
0'
0/
#547130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#547140000000
0!
0'
0/
#547150000000
1!
1'
1/
#547160000000
0!
0'
0/
#547170000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#547180000000
0!
0'
0/
#547190000000
1!
1'
1/
#547200000000
0!
0'
0/
#547210000000
1!
1'
1/
#547220000000
0!
0'
0/
#547230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#547240000000
0!
0'
0/
#547250000000
1!
1'
1/
#547260000000
0!
0'
0/
#547270000000
1!
1'
1/
#547280000000
0!
0'
0/
#547290000000
1!
1'
1/
#547300000000
0!
0'
0/
#547310000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#547320000000
0!
0'
0/
#547330000000
1!
1'
1/
#547340000000
0!
0'
0/
#547350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#547360000000
0!
0'
0/
#547370000000
1!
1'
1/
#547380000000
0!
0'
0/
#547390000000
#547400000000
1!
1'
1/
#547410000000
0!
0'
0/
#547420000000
1!
1'
1/
#547430000000
0!
1"
0'
1(
0/
10
#547440000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#547450000000
0!
0'
0/
#547460000000
1!
1'
1/
#547470000000
0!
0'
0/
#547480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#547490000000
0!
0'
0/
#547500000000
1!
1'
1/
#547510000000
0!
1"
0'
1(
0/
10
#547520000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#547530000000
0!
1$
0'
1+
0/
#547540000000
1!
1'
1/
#547550000000
0!
0'
0/
#547560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#547570000000
0!
0'
0/
#547580000000
1!
1'
1/
#547590000000
0!
0'
0/
#547600000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#547610000000
0!
0'
0/
#547620000000
1!
1'
1/
#547630000000
0!
0'
0/
#547640000000
1!
1'
1/
#547650000000
0!
0'
0/
#547660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#547670000000
0!
0'
0/
#547680000000
1!
1'
1/
#547690000000
0!
0'
0/
#547700000000
1!
1'
1/
#547710000000
0!
0'
0/
#547720000000
1!
1'
1/
#547730000000
0!
0'
0/
#547740000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#547750000000
0!
0'
0/
#547760000000
1!
1'
1/
#547770000000
0!
0'
0/
#547780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#547790000000
0!
0'
0/
#547800000000
1!
1'
1/
#547810000000
0!
0'
0/
#547820000000
#547830000000
1!
1'
1/
#547840000000
0!
0'
0/
#547850000000
1!
1'
1/
#547860000000
0!
1"
0'
1(
0/
10
#547870000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#547880000000
0!
0'
0/
#547890000000
1!
1'
1/
#547900000000
0!
0'
0/
#547910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#547920000000
0!
0'
0/
#547930000000
1!
1'
1/
#547940000000
0!
1"
0'
1(
0/
10
#547950000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#547960000000
0!
1$
0'
1+
0/
#547970000000
1!
1'
1/
#547980000000
0!
0'
0/
#547990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#548000000000
0!
0'
0/
#548010000000
1!
1'
1/
#548020000000
0!
0'
0/
#548030000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#548040000000
0!
0'
0/
#548050000000
1!
1'
1/
#548060000000
0!
0'
0/
#548070000000
1!
1'
1/
#548080000000
0!
0'
0/
#548090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#548100000000
0!
0'
0/
#548110000000
1!
1'
1/
#548120000000
0!
0'
0/
#548130000000
1!
1'
1/
#548140000000
0!
0'
0/
#548150000000
1!
1'
1/
#548160000000
0!
0'
0/
#548170000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#548180000000
0!
0'
0/
#548190000000
1!
1'
1/
#548200000000
0!
0'
0/
#548210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#548220000000
0!
0'
0/
#548230000000
1!
1'
1/
#548240000000
0!
0'
0/
#548250000000
#548260000000
1!
1'
1/
#548270000000
0!
0'
0/
#548280000000
1!
1'
1/
#548290000000
0!
1"
0'
1(
0/
10
#548300000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#548310000000
0!
0'
0/
#548320000000
1!
1'
1/
#548330000000
0!
0'
0/
#548340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#548350000000
0!
0'
0/
#548360000000
1!
1'
1/
#548370000000
0!
1"
0'
1(
0/
10
#548380000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#548390000000
0!
1$
0'
1+
0/
#548400000000
1!
1'
1/
#548410000000
0!
0'
0/
#548420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#548430000000
0!
0'
0/
#548440000000
1!
1'
1/
#548450000000
0!
0'
0/
#548460000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#548470000000
0!
0'
0/
#548480000000
1!
1'
1/
#548490000000
0!
0'
0/
#548500000000
1!
1'
1/
#548510000000
0!
0'
0/
#548520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#548530000000
0!
0'
0/
#548540000000
1!
1'
1/
#548550000000
0!
0'
0/
#548560000000
1!
1'
1/
#548570000000
0!
0'
0/
#548580000000
1!
1'
1/
#548590000000
0!
0'
0/
#548600000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#548610000000
0!
0'
0/
#548620000000
1!
1'
1/
#548630000000
0!
0'
0/
#548640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#548650000000
0!
0'
0/
#548660000000
1!
1'
1/
#548670000000
0!
0'
0/
#548680000000
#548690000000
1!
1'
1/
#548700000000
0!
0'
0/
#548710000000
1!
1'
1/
#548720000000
0!
1"
0'
1(
0/
10
#548730000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#548740000000
0!
0'
0/
#548750000000
1!
1'
1/
#548760000000
0!
0'
0/
#548770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#548780000000
0!
0'
0/
#548790000000
1!
1'
1/
#548800000000
0!
1"
0'
1(
0/
10
#548810000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#548820000000
0!
1$
0'
1+
0/
#548830000000
1!
1'
1/
#548840000000
0!
0'
0/
#548850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#548860000000
0!
0'
0/
#548870000000
1!
1'
1/
#548880000000
0!
0'
0/
#548890000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#548900000000
0!
0'
0/
#548910000000
1!
1'
1/
#548920000000
0!
0'
0/
#548930000000
1!
1'
1/
#548940000000
0!
0'
0/
#548950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#548960000000
0!
0'
0/
#548970000000
1!
1'
1/
#548980000000
0!
0'
0/
#548990000000
1!
1'
1/
#549000000000
0!
0'
0/
#549010000000
1!
1'
1/
#549020000000
0!
0'
0/
#549030000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#549040000000
0!
0'
0/
#549050000000
1!
1'
1/
#549060000000
0!
0'
0/
#549070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#549080000000
0!
0'
0/
#549090000000
1!
1'
1/
#549100000000
0!
0'
0/
#549110000000
#549120000000
1!
1'
1/
#549130000000
0!
0'
0/
#549140000000
1!
1'
1/
#549150000000
0!
1"
0'
1(
0/
10
#549160000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#549170000000
0!
0'
0/
#549180000000
1!
1'
1/
#549190000000
0!
0'
0/
#549200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#549210000000
0!
0'
0/
#549220000000
1!
1'
1/
#549230000000
0!
1"
0'
1(
0/
10
#549240000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#549250000000
0!
1$
0'
1+
0/
#549260000000
1!
1'
1/
#549270000000
0!
0'
0/
#549280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#549290000000
0!
0'
0/
#549300000000
1!
1'
1/
#549310000000
0!
0'
0/
#549320000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#549330000000
0!
0'
0/
#549340000000
1!
1'
1/
#549350000000
0!
0'
0/
#549360000000
1!
1'
1/
#549370000000
0!
0'
0/
#549380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#549390000000
0!
0'
0/
#549400000000
1!
1'
1/
#549410000000
0!
0'
0/
#549420000000
1!
1'
1/
#549430000000
0!
0'
0/
#549440000000
1!
1'
1/
#549450000000
0!
0'
0/
#549460000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#549470000000
0!
0'
0/
#549480000000
1!
1'
1/
#549490000000
0!
0'
0/
#549500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#549510000000
0!
0'
0/
#549520000000
1!
1'
1/
#549530000000
0!
0'
0/
#549540000000
#549550000000
1!
1'
1/
#549560000000
0!
0'
0/
#549570000000
1!
1'
1/
#549580000000
0!
1"
0'
1(
0/
10
#549590000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#549600000000
0!
0'
0/
#549610000000
1!
1'
1/
#549620000000
0!
0'
0/
#549630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#549640000000
0!
0'
0/
#549650000000
1!
1'
1/
#549660000000
0!
1"
0'
1(
0/
10
#549670000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#549680000000
0!
1$
0'
1+
0/
#549690000000
1!
1'
1/
#549700000000
0!
0'
0/
#549710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#549720000000
0!
0'
0/
#549730000000
1!
1'
1/
#549740000000
0!
0'
0/
#549750000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#549760000000
0!
0'
0/
#549770000000
1!
1'
1/
#549780000000
0!
0'
0/
#549790000000
1!
1'
1/
#549800000000
0!
0'
0/
#549810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#549820000000
0!
0'
0/
#549830000000
1!
1'
1/
#549840000000
0!
0'
0/
#549850000000
1!
1'
1/
#549860000000
0!
0'
0/
#549870000000
1!
1'
1/
#549880000000
0!
0'
0/
#549890000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#549900000000
0!
0'
0/
#549910000000
1!
1'
1/
#549920000000
0!
0'
0/
#549930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#549940000000
0!
0'
0/
#549950000000
1!
1'
1/
#549960000000
0!
0'
0/
#549970000000
#549980000000
1!
1'
1/
#549990000000
0!
0'
0/
#550000000000
1!
1'
1/
#550010000000
0!
1"
0'
1(
0/
10
#550020000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#550030000000
0!
0'
0/
#550040000000
1!
1'
1/
#550050000000
0!
0'
0/
#550060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#550070000000
0!
0'
0/
#550080000000
1!
1'
1/
#550090000000
0!
1"
0'
1(
0/
10
#550100000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#550110000000
0!
1$
0'
1+
0/
#550120000000
1!
1'
1/
#550130000000
0!
0'
0/
#550140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#550150000000
0!
0'
0/
#550160000000
1!
1'
1/
#550170000000
0!
0'
0/
#550180000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#550190000000
0!
0'
0/
#550200000000
1!
1'
1/
#550210000000
0!
0'
0/
#550220000000
1!
1'
1/
#550230000000
0!
0'
0/
#550240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#550250000000
0!
0'
0/
#550260000000
1!
1'
1/
#550270000000
0!
0'
0/
#550280000000
1!
1'
1/
#550290000000
0!
0'
0/
#550300000000
1!
1'
1/
#550310000000
0!
0'
0/
#550320000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#550330000000
0!
0'
0/
#550340000000
1!
1'
1/
#550350000000
0!
0'
0/
#550360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#550370000000
0!
0'
0/
#550380000000
1!
1'
1/
#550390000000
0!
0'
0/
#550400000000
#550410000000
1!
1'
1/
#550420000000
0!
0'
0/
#550430000000
1!
1'
1/
#550440000000
0!
1"
0'
1(
0/
10
#550450000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#550460000000
0!
0'
0/
#550470000000
1!
1'
1/
#550480000000
0!
0'
0/
#550490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#550500000000
0!
0'
0/
#550510000000
1!
1'
1/
#550520000000
0!
1"
0'
1(
0/
10
#550530000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#550540000000
0!
1$
0'
1+
0/
#550550000000
1!
1'
1/
#550560000000
0!
0'
0/
#550570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#550580000000
0!
0'
0/
#550590000000
1!
1'
1/
#550600000000
0!
0'
0/
#550610000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#550620000000
0!
0'
0/
#550630000000
1!
1'
1/
#550640000000
0!
0'
0/
#550650000000
1!
1'
1/
#550660000000
0!
0'
0/
#550670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#550680000000
0!
0'
0/
#550690000000
1!
1'
1/
#550700000000
0!
0'
0/
#550710000000
1!
1'
1/
#550720000000
0!
0'
0/
#550730000000
1!
1'
1/
#550740000000
0!
0'
0/
#550750000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#550760000000
0!
0'
0/
#550770000000
1!
1'
1/
#550780000000
0!
0'
0/
#550790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#550800000000
0!
0'
0/
#550810000000
1!
1'
1/
#550820000000
0!
0'
0/
#550830000000
#550840000000
1!
1'
1/
#550850000000
0!
0'
0/
#550860000000
1!
1'
1/
#550870000000
0!
1"
0'
1(
0/
10
#550880000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#550890000000
0!
0'
0/
#550900000000
1!
1'
1/
#550910000000
0!
0'
0/
#550920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#550930000000
0!
0'
0/
#550940000000
1!
1'
1/
#550950000000
0!
1"
0'
1(
0/
10
#550960000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#550970000000
0!
1$
0'
1+
0/
#550980000000
1!
1'
1/
#550990000000
0!
0'
0/
#551000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#551010000000
0!
0'
0/
#551020000000
1!
1'
1/
#551030000000
0!
0'
0/
#551040000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#551050000000
0!
0'
0/
#551060000000
1!
1'
1/
#551070000000
0!
0'
0/
#551080000000
1!
1'
1/
#551090000000
0!
0'
0/
#551100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#551110000000
0!
0'
0/
#551120000000
1!
1'
1/
#551130000000
0!
0'
0/
#551140000000
1!
1'
1/
#551150000000
0!
0'
0/
#551160000000
1!
1'
1/
#551170000000
0!
0'
0/
#551180000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#551190000000
0!
0'
0/
#551200000000
1!
1'
1/
#551210000000
0!
0'
0/
#551220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#551230000000
0!
0'
0/
#551240000000
1!
1'
1/
#551250000000
0!
0'
0/
#551260000000
#551270000000
1!
1'
1/
#551280000000
0!
0'
0/
#551290000000
1!
1'
1/
#551300000000
0!
1"
0'
1(
0/
10
#551310000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#551320000000
0!
0'
0/
#551330000000
1!
1'
1/
#551340000000
0!
0'
0/
#551350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#551360000000
0!
0'
0/
#551370000000
1!
1'
1/
#551380000000
0!
1"
0'
1(
0/
10
#551390000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#551400000000
0!
1$
0'
1+
0/
#551410000000
1!
1'
1/
#551420000000
0!
0'
0/
#551430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#551440000000
0!
0'
0/
#551450000000
1!
1'
1/
#551460000000
0!
0'
0/
#551470000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#551480000000
0!
0'
0/
#551490000000
1!
1'
1/
#551500000000
0!
0'
0/
#551510000000
1!
1'
1/
#551520000000
0!
0'
0/
#551530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#551540000000
0!
0'
0/
#551550000000
1!
1'
1/
#551560000000
0!
0'
0/
#551570000000
1!
1'
1/
#551580000000
0!
0'
0/
#551590000000
1!
1'
1/
#551600000000
0!
0'
0/
#551610000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#551620000000
0!
0'
0/
#551630000000
1!
1'
1/
#551640000000
0!
0'
0/
#551650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#551660000000
0!
0'
0/
#551670000000
1!
1'
1/
#551680000000
0!
0'
0/
#551690000000
#551700000000
1!
1'
1/
#551710000000
0!
0'
0/
#551720000000
1!
1'
1/
#551730000000
0!
1"
0'
1(
0/
10
#551740000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#551750000000
0!
0'
0/
#551760000000
1!
1'
1/
#551770000000
0!
0'
0/
#551780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#551790000000
0!
0'
0/
#551800000000
1!
1'
1/
#551810000000
0!
1"
0'
1(
0/
10
#551820000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#551830000000
0!
1$
0'
1+
0/
#551840000000
1!
1'
1/
#551850000000
0!
0'
0/
#551860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#551870000000
0!
0'
0/
#551880000000
1!
1'
1/
#551890000000
0!
0'
0/
#551900000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#551910000000
0!
0'
0/
#551920000000
1!
1'
1/
#551930000000
0!
0'
0/
#551940000000
1!
1'
1/
#551950000000
0!
0'
0/
#551960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#551970000000
0!
0'
0/
#551980000000
1!
1'
1/
#551990000000
0!
0'
0/
#552000000000
1!
1'
1/
#552010000000
0!
0'
0/
#552020000000
1!
1'
1/
#552030000000
0!
0'
0/
#552040000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#552050000000
0!
0'
0/
#552060000000
1!
1'
1/
#552070000000
0!
0'
0/
#552080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#552090000000
0!
0'
0/
#552100000000
1!
1'
1/
#552110000000
0!
0'
0/
#552120000000
#552130000000
1!
1'
1/
#552140000000
0!
0'
0/
#552150000000
1!
1'
1/
#552160000000
0!
1"
0'
1(
0/
10
#552170000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#552180000000
0!
0'
0/
#552190000000
1!
1'
1/
#552200000000
0!
0'
0/
#552210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#552220000000
0!
0'
0/
#552230000000
1!
1'
1/
#552240000000
0!
1"
0'
1(
0/
10
#552250000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#552260000000
0!
1$
0'
1+
0/
#552270000000
1!
1'
1/
#552280000000
0!
0'
0/
#552290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#552300000000
0!
0'
0/
#552310000000
1!
1'
1/
#552320000000
0!
0'
0/
#552330000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#552340000000
0!
0'
0/
#552350000000
1!
1'
1/
#552360000000
0!
0'
0/
#552370000000
1!
1'
1/
#552380000000
0!
0'
0/
#552390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#552400000000
0!
0'
0/
#552410000000
1!
1'
1/
#552420000000
0!
0'
0/
#552430000000
1!
1'
1/
#552440000000
0!
0'
0/
#552450000000
1!
1'
1/
#552460000000
0!
0'
0/
#552470000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#552480000000
0!
0'
0/
#552490000000
1!
1'
1/
#552500000000
0!
0'
0/
#552510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#552520000000
0!
0'
0/
#552530000000
1!
1'
1/
#552540000000
0!
0'
0/
#552550000000
#552560000000
1!
1'
1/
#552570000000
0!
0'
0/
#552580000000
1!
1'
1/
#552590000000
0!
1"
0'
1(
0/
10
#552600000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#552610000000
0!
0'
0/
#552620000000
1!
1'
1/
#552630000000
0!
0'
0/
#552640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#552650000000
0!
0'
0/
#552660000000
1!
1'
1/
#552670000000
0!
1"
0'
1(
0/
10
#552680000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#552690000000
0!
1$
0'
1+
0/
#552700000000
1!
1'
1/
#552710000000
0!
0'
0/
#552720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#552730000000
0!
0'
0/
#552740000000
1!
1'
1/
#552750000000
0!
0'
0/
#552760000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#552770000000
0!
0'
0/
#552780000000
1!
1'
1/
#552790000000
0!
0'
0/
#552800000000
1!
1'
1/
#552810000000
0!
0'
0/
#552820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#552830000000
0!
0'
0/
#552840000000
1!
1'
1/
#552850000000
0!
0'
0/
#552860000000
1!
1'
1/
#552870000000
0!
0'
0/
#552880000000
1!
1'
1/
#552890000000
0!
0'
0/
#552900000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#552910000000
0!
0'
0/
#552920000000
1!
1'
1/
#552930000000
0!
0'
0/
#552940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#552950000000
0!
0'
0/
#552960000000
1!
1'
1/
#552970000000
0!
0'
0/
#552980000000
#552990000000
1!
1'
1/
#553000000000
0!
0'
0/
#553010000000
1!
1'
1/
#553020000000
0!
1"
0'
1(
0/
10
#553030000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#553040000000
0!
0'
0/
#553050000000
1!
1'
1/
#553060000000
0!
0'
0/
#553070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#553080000000
0!
0'
0/
#553090000000
1!
1'
1/
#553100000000
0!
1"
0'
1(
0/
10
#553110000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#553120000000
0!
1$
0'
1+
0/
#553130000000
1!
1'
1/
#553140000000
0!
0'
0/
#553150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#553160000000
0!
0'
0/
#553170000000
1!
1'
1/
#553180000000
0!
0'
0/
#553190000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#553200000000
0!
0'
0/
#553210000000
1!
1'
1/
#553220000000
0!
0'
0/
#553230000000
1!
1'
1/
#553240000000
0!
0'
0/
#553250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#553260000000
0!
0'
0/
#553270000000
1!
1'
1/
#553280000000
0!
0'
0/
#553290000000
1!
1'
1/
#553300000000
0!
0'
0/
#553310000000
1!
1'
1/
#553320000000
0!
0'
0/
#553330000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#553340000000
0!
0'
0/
#553350000000
1!
1'
1/
#553360000000
0!
0'
0/
#553370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#553380000000
0!
0'
0/
#553390000000
1!
1'
1/
#553400000000
0!
0'
0/
#553410000000
#553420000000
1!
1'
1/
#553430000000
0!
0'
0/
#553440000000
1!
1'
1/
#553450000000
0!
1"
0'
1(
0/
10
#553460000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#553470000000
0!
0'
0/
#553480000000
1!
1'
1/
#553490000000
0!
0'
0/
#553500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#553510000000
0!
0'
0/
#553520000000
1!
1'
1/
#553530000000
0!
1"
0'
1(
0/
10
#553540000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#553550000000
0!
1$
0'
1+
0/
#553560000000
1!
1'
1/
#553570000000
0!
0'
0/
#553580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#553590000000
0!
0'
0/
#553600000000
1!
1'
1/
#553610000000
0!
0'
0/
#553620000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#553630000000
0!
0'
0/
#553640000000
1!
1'
1/
#553650000000
0!
0'
0/
#553660000000
1!
1'
1/
#553670000000
0!
0'
0/
#553680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#553690000000
0!
0'
0/
#553700000000
1!
1'
1/
#553710000000
0!
0'
0/
#553720000000
1!
1'
1/
#553730000000
0!
0'
0/
#553740000000
1!
1'
1/
#553750000000
0!
0'
0/
#553760000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#553770000000
0!
0'
0/
#553780000000
1!
1'
1/
#553790000000
0!
0'
0/
#553800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#553810000000
0!
0'
0/
#553820000000
1!
1'
1/
#553830000000
0!
0'
0/
#553840000000
#553850000000
1!
1'
1/
#553860000000
0!
0'
0/
#553870000000
1!
1'
1/
#553880000000
0!
1"
0'
1(
0/
10
#553890000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#553900000000
0!
0'
0/
#553910000000
1!
1'
1/
#553920000000
0!
0'
0/
#553930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#553940000000
0!
0'
0/
#553950000000
1!
1'
1/
#553960000000
0!
1"
0'
1(
0/
10
#553970000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#553980000000
0!
1$
0'
1+
0/
#553990000000
1!
1'
1/
#554000000000
0!
0'
0/
#554010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#554020000000
0!
0'
0/
#554030000000
1!
1'
1/
#554040000000
0!
0'
0/
#554050000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#554060000000
0!
0'
0/
#554070000000
1!
1'
1/
#554080000000
0!
0'
0/
#554090000000
1!
1'
1/
#554100000000
0!
0'
0/
#554110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#554120000000
0!
0'
0/
#554130000000
1!
1'
1/
#554140000000
0!
0'
0/
#554150000000
1!
1'
1/
#554160000000
0!
0'
0/
#554170000000
1!
1'
1/
#554180000000
0!
0'
0/
#554190000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#554200000000
0!
0'
0/
#554210000000
1!
1'
1/
#554220000000
0!
0'
0/
#554230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#554240000000
0!
0'
0/
#554250000000
1!
1'
1/
#554260000000
0!
0'
0/
#554270000000
#554280000000
1!
1'
1/
#554290000000
0!
0'
0/
#554300000000
1!
1'
1/
#554310000000
0!
1"
0'
1(
0/
10
#554320000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#554330000000
0!
0'
0/
#554340000000
1!
1'
1/
#554350000000
0!
0'
0/
#554360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#554370000000
0!
0'
0/
#554380000000
1!
1'
1/
#554390000000
0!
1"
0'
1(
0/
10
#554400000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#554410000000
0!
1$
0'
1+
0/
#554420000000
1!
1'
1/
#554430000000
0!
0'
0/
#554440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#554450000000
0!
0'
0/
#554460000000
1!
1'
1/
#554470000000
0!
0'
0/
#554480000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#554490000000
0!
0'
0/
#554500000000
1!
1'
1/
#554510000000
0!
0'
0/
#554520000000
1!
1'
1/
#554530000000
0!
0'
0/
#554540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#554550000000
0!
0'
0/
#554560000000
1!
1'
1/
#554570000000
0!
0'
0/
#554580000000
1!
1'
1/
#554590000000
0!
0'
0/
#554600000000
1!
1'
1/
#554610000000
0!
0'
0/
#554620000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#554630000000
0!
0'
0/
#554640000000
1!
1'
1/
#554650000000
0!
0'
0/
#554660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#554670000000
0!
0'
0/
#554680000000
1!
1'
1/
#554690000000
0!
0'
0/
#554700000000
#554710000000
1!
1'
1/
#554720000000
0!
0'
0/
#554730000000
1!
1'
1/
#554740000000
0!
1"
0'
1(
0/
10
#554750000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#554760000000
0!
0'
0/
#554770000000
1!
1'
1/
#554780000000
0!
0'
0/
#554790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#554800000000
0!
0'
0/
#554810000000
1!
1'
1/
#554820000000
0!
1"
0'
1(
0/
10
#554830000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#554840000000
0!
1$
0'
1+
0/
#554850000000
1!
1'
1/
#554860000000
0!
0'
0/
#554870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#554880000000
0!
0'
0/
#554890000000
1!
1'
1/
#554900000000
0!
0'
0/
#554910000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#554920000000
0!
0'
0/
#554930000000
1!
1'
1/
#554940000000
0!
0'
0/
#554950000000
1!
1'
1/
#554960000000
0!
0'
0/
#554970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#554980000000
0!
0'
0/
#554990000000
1!
1'
1/
#555000000000
0!
0'
0/
#555010000000
1!
1'
1/
#555020000000
0!
0'
0/
#555030000000
1!
1'
1/
#555040000000
0!
0'
0/
#555050000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#555060000000
0!
0'
0/
#555070000000
1!
1'
1/
#555080000000
0!
0'
0/
#555090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#555100000000
0!
0'
0/
#555110000000
1!
1'
1/
#555120000000
0!
0'
0/
#555130000000
#555140000000
1!
1'
1/
#555150000000
0!
0'
0/
#555160000000
1!
1'
1/
#555170000000
0!
1"
0'
1(
0/
10
#555180000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#555190000000
0!
0'
0/
#555200000000
1!
1'
1/
#555210000000
0!
0'
0/
#555220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#555230000000
0!
0'
0/
#555240000000
1!
1'
1/
#555250000000
0!
1"
0'
1(
0/
10
#555260000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#555270000000
0!
1$
0'
1+
0/
#555280000000
1!
1'
1/
#555290000000
0!
0'
0/
#555300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#555310000000
0!
0'
0/
#555320000000
1!
1'
1/
#555330000000
0!
0'
0/
#555340000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#555350000000
0!
0'
0/
#555360000000
1!
1'
1/
#555370000000
0!
0'
0/
#555380000000
1!
1'
1/
#555390000000
0!
0'
0/
#555400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#555410000000
0!
0'
0/
#555420000000
1!
1'
1/
#555430000000
0!
0'
0/
#555440000000
1!
1'
1/
#555450000000
0!
0'
0/
#555460000000
1!
1'
1/
#555470000000
0!
0'
0/
#555480000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#555490000000
0!
0'
0/
#555500000000
1!
1'
1/
#555510000000
0!
0'
0/
#555520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#555530000000
0!
0'
0/
#555540000000
1!
1'
1/
#555550000000
0!
0'
0/
#555560000000
#555570000000
1!
1'
1/
#555580000000
0!
0'
0/
#555590000000
1!
1'
1/
#555600000000
0!
1"
0'
1(
0/
10
#555610000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#555620000000
0!
0'
0/
#555630000000
1!
1'
1/
#555640000000
0!
0'
0/
#555650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#555660000000
0!
0'
0/
#555670000000
1!
1'
1/
#555680000000
0!
1"
0'
1(
0/
10
#555690000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#555700000000
0!
1$
0'
1+
0/
#555710000000
1!
1'
1/
#555720000000
0!
0'
0/
#555730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#555740000000
0!
0'
0/
#555750000000
1!
1'
1/
#555760000000
0!
0'
0/
#555770000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#555780000000
0!
0'
0/
#555790000000
1!
1'
1/
#555800000000
0!
0'
0/
#555810000000
1!
1'
1/
#555820000000
0!
0'
0/
#555830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#555840000000
0!
0'
0/
#555850000000
1!
1'
1/
#555860000000
0!
0'
0/
#555870000000
1!
1'
1/
#555880000000
0!
0'
0/
#555890000000
1!
1'
1/
#555900000000
0!
0'
0/
#555910000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#555920000000
0!
0'
0/
#555930000000
1!
1'
1/
#555940000000
0!
0'
0/
#555950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#555960000000
0!
0'
0/
#555970000000
1!
1'
1/
#555980000000
0!
0'
0/
#555990000000
#556000000000
1!
1'
1/
#556010000000
0!
0'
0/
#556020000000
1!
1'
1/
#556030000000
0!
1"
0'
1(
0/
10
#556040000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#556050000000
0!
0'
0/
#556060000000
1!
1'
1/
#556070000000
0!
0'
0/
#556080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#556090000000
0!
0'
0/
#556100000000
1!
1'
1/
#556110000000
0!
1"
0'
1(
0/
10
#556120000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#556130000000
0!
1$
0'
1+
0/
#556140000000
1!
1'
1/
#556150000000
0!
0'
0/
#556160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#556170000000
0!
0'
0/
#556180000000
1!
1'
1/
#556190000000
0!
0'
0/
#556200000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#556210000000
0!
0'
0/
#556220000000
1!
1'
1/
#556230000000
0!
0'
0/
#556240000000
1!
1'
1/
#556250000000
0!
0'
0/
#556260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#556270000000
0!
0'
0/
#556280000000
1!
1'
1/
#556290000000
0!
0'
0/
#556300000000
1!
1'
1/
#556310000000
0!
0'
0/
#556320000000
1!
1'
1/
#556330000000
0!
0'
0/
#556340000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#556350000000
0!
0'
0/
#556360000000
1!
1'
1/
#556370000000
0!
0'
0/
#556380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#556390000000
0!
0'
0/
#556400000000
1!
1'
1/
#556410000000
0!
0'
0/
#556420000000
#556430000000
1!
1'
1/
#556440000000
0!
0'
0/
#556450000000
1!
1'
1/
#556460000000
0!
1"
0'
1(
0/
10
#556470000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#556480000000
0!
0'
0/
#556490000000
1!
1'
1/
#556500000000
0!
0'
0/
#556510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#556520000000
0!
0'
0/
#556530000000
1!
1'
1/
#556540000000
0!
1"
0'
1(
0/
10
#556550000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#556560000000
0!
1$
0'
1+
0/
#556570000000
1!
1'
1/
#556580000000
0!
0'
0/
#556590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#556600000000
0!
0'
0/
#556610000000
1!
1'
1/
#556620000000
0!
0'
0/
#556630000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#556640000000
0!
0'
0/
#556650000000
1!
1'
1/
#556660000000
0!
0'
0/
#556670000000
1!
1'
1/
#556680000000
0!
0'
0/
#556690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#556700000000
0!
0'
0/
#556710000000
1!
1'
1/
#556720000000
0!
0'
0/
#556730000000
1!
1'
1/
#556740000000
0!
0'
0/
#556750000000
1!
1'
1/
#556760000000
0!
0'
0/
#556770000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#556780000000
0!
0'
0/
#556790000000
1!
1'
1/
#556800000000
0!
0'
0/
#556810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#556820000000
0!
0'
0/
#556830000000
1!
1'
1/
#556840000000
0!
0'
0/
#556850000000
#556860000000
1!
1'
1/
#556870000000
0!
0'
0/
#556880000000
1!
1'
1/
#556890000000
0!
1"
0'
1(
0/
10
#556900000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#556910000000
0!
0'
0/
#556920000000
1!
1'
1/
#556930000000
0!
0'
0/
#556940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#556950000000
0!
0'
0/
#556960000000
1!
1'
1/
#556970000000
0!
1"
0'
1(
0/
10
#556980000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#556990000000
0!
1$
0'
1+
0/
#557000000000
1!
1'
1/
#557010000000
0!
0'
0/
#557020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#557030000000
0!
0'
0/
#557040000000
1!
1'
1/
#557050000000
0!
0'
0/
#557060000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#557070000000
0!
0'
0/
#557080000000
1!
1'
1/
#557090000000
0!
0'
0/
#557100000000
1!
1'
1/
#557110000000
0!
0'
0/
#557120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#557130000000
0!
0'
0/
#557140000000
1!
1'
1/
#557150000000
0!
0'
0/
#557160000000
1!
1'
1/
#557170000000
0!
0'
0/
#557180000000
1!
1'
1/
#557190000000
0!
0'
0/
#557200000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#557210000000
0!
0'
0/
#557220000000
1!
1'
1/
#557230000000
0!
0'
0/
#557240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#557250000000
0!
0'
0/
#557260000000
1!
1'
1/
#557270000000
0!
0'
0/
#557280000000
#557290000000
1!
1'
1/
#557300000000
0!
0'
0/
#557310000000
1!
1'
1/
#557320000000
0!
1"
0'
1(
0/
10
#557330000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#557340000000
0!
0'
0/
#557350000000
1!
1'
1/
#557360000000
0!
0'
0/
#557370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#557380000000
0!
0'
0/
#557390000000
1!
1'
1/
#557400000000
0!
1"
0'
1(
0/
10
#557410000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#557420000000
0!
1$
0'
1+
0/
#557430000000
1!
1'
1/
#557440000000
0!
0'
0/
#557450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#557460000000
0!
0'
0/
#557470000000
1!
1'
1/
#557480000000
0!
0'
0/
#557490000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#557500000000
0!
0'
0/
#557510000000
1!
1'
1/
#557520000000
0!
0'
0/
#557530000000
1!
1'
1/
#557540000000
0!
0'
0/
#557550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#557560000000
0!
0'
0/
#557570000000
1!
1'
1/
#557580000000
0!
0'
0/
#557590000000
1!
1'
1/
#557600000000
0!
0'
0/
#557610000000
1!
1'
1/
#557620000000
0!
0'
0/
#557630000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#557640000000
0!
0'
0/
#557650000000
1!
1'
1/
#557660000000
0!
0'
0/
#557670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#557680000000
0!
0'
0/
#557690000000
1!
1'
1/
#557700000000
0!
0'
0/
#557710000000
#557720000000
1!
1'
1/
#557730000000
0!
0'
0/
#557740000000
1!
1'
1/
#557750000000
0!
1"
0'
1(
0/
10
#557760000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#557770000000
0!
0'
0/
#557780000000
1!
1'
1/
#557790000000
0!
0'
0/
#557800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#557810000000
0!
0'
0/
#557820000000
1!
1'
1/
#557830000000
0!
1"
0'
1(
0/
10
#557840000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#557850000000
0!
1$
0'
1+
0/
#557860000000
1!
1'
1/
#557870000000
0!
0'
0/
#557880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#557890000000
0!
0'
0/
#557900000000
1!
1'
1/
#557910000000
0!
0'
0/
#557920000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#557930000000
0!
0'
0/
#557940000000
1!
1'
1/
#557950000000
0!
0'
0/
#557960000000
1!
1'
1/
#557970000000
0!
0'
0/
#557980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#557990000000
0!
0'
0/
#558000000000
1!
1'
1/
#558010000000
0!
0'
0/
#558020000000
1!
1'
1/
#558030000000
0!
0'
0/
#558040000000
1!
1'
1/
#558050000000
0!
0'
0/
#558060000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#558070000000
0!
0'
0/
#558080000000
1!
1'
1/
#558090000000
0!
0'
0/
#558100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#558110000000
0!
0'
0/
#558120000000
1!
1'
1/
#558130000000
0!
0'
0/
#558140000000
#558150000000
1!
1'
1/
#558160000000
0!
0'
0/
#558170000000
1!
1'
1/
#558180000000
0!
1"
0'
1(
0/
10
#558190000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#558200000000
0!
0'
0/
#558210000000
1!
1'
1/
#558220000000
0!
0'
0/
#558230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#558240000000
0!
0'
0/
#558250000000
1!
1'
1/
#558260000000
0!
1"
0'
1(
0/
10
#558270000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#558280000000
0!
1$
0'
1+
0/
#558290000000
1!
1'
1/
#558300000000
0!
0'
0/
#558310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#558320000000
0!
0'
0/
#558330000000
1!
1'
1/
#558340000000
0!
0'
0/
#558350000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#558360000000
0!
0'
0/
#558370000000
1!
1'
1/
#558380000000
0!
0'
0/
#558390000000
1!
1'
1/
#558400000000
0!
0'
0/
#558410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#558420000000
0!
0'
0/
#558430000000
1!
1'
1/
#558440000000
0!
0'
0/
#558450000000
1!
1'
1/
#558460000000
0!
0'
0/
#558470000000
1!
1'
1/
#558480000000
0!
0'
0/
#558490000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#558500000000
0!
0'
0/
#558510000000
1!
1'
1/
#558520000000
0!
0'
0/
#558530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#558540000000
0!
0'
0/
#558550000000
1!
1'
1/
#558560000000
0!
0'
0/
#558570000000
#558580000000
1!
1'
1/
#558590000000
0!
0'
0/
#558600000000
1!
1'
1/
#558610000000
0!
1"
0'
1(
0/
10
#558620000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#558630000000
0!
0'
0/
#558640000000
1!
1'
1/
#558650000000
0!
0'
0/
#558660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#558670000000
0!
0'
0/
#558680000000
1!
1'
1/
#558690000000
0!
1"
0'
1(
0/
10
#558700000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#558710000000
0!
1$
0'
1+
0/
#558720000000
1!
1'
1/
#558730000000
0!
0'
0/
#558740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#558750000000
0!
0'
0/
#558760000000
1!
1'
1/
#558770000000
0!
0'
0/
#558780000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#558790000000
0!
0'
0/
#558800000000
1!
1'
1/
#558810000000
0!
0'
0/
#558820000000
1!
1'
1/
#558830000000
0!
0'
0/
#558840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#558850000000
0!
0'
0/
#558860000000
1!
1'
1/
#558870000000
0!
0'
0/
#558880000000
1!
1'
1/
#558890000000
0!
0'
0/
#558900000000
1!
1'
1/
#558910000000
0!
0'
0/
#558920000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#558930000000
0!
0'
0/
#558940000000
1!
1'
1/
#558950000000
0!
0'
0/
#558960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#558970000000
0!
0'
0/
#558980000000
1!
1'
1/
#558990000000
0!
0'
0/
#559000000000
#559010000000
1!
1'
1/
#559020000000
0!
0'
0/
#559030000000
1!
1'
1/
#559040000000
0!
1"
0'
1(
0/
10
#559050000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#559060000000
0!
0'
0/
#559070000000
1!
1'
1/
#559080000000
0!
0'
0/
#559090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#559100000000
0!
0'
0/
#559110000000
1!
1'
1/
#559120000000
0!
1"
0'
1(
0/
10
#559130000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#559140000000
0!
1$
0'
1+
0/
#559150000000
1!
1'
1/
#559160000000
0!
0'
0/
#559170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#559180000000
0!
0'
0/
#559190000000
1!
1'
1/
#559200000000
0!
0'
0/
#559210000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#559220000000
0!
0'
0/
#559230000000
1!
1'
1/
#559240000000
0!
0'
0/
#559250000000
1!
1'
1/
#559260000000
0!
0'
0/
#559270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#559280000000
0!
0'
0/
#559290000000
1!
1'
1/
#559300000000
0!
0'
0/
#559310000000
1!
1'
1/
#559320000000
0!
0'
0/
#559330000000
1!
1'
1/
#559340000000
0!
0'
0/
#559350000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#559360000000
0!
0'
0/
#559370000000
1!
1'
1/
#559380000000
0!
0'
0/
#559390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#559400000000
0!
0'
0/
#559410000000
1!
1'
1/
#559420000000
0!
0'
0/
#559430000000
#559440000000
1!
1'
1/
#559450000000
0!
0'
0/
#559460000000
1!
1'
1/
#559470000000
0!
1"
0'
1(
0/
10
#559480000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#559490000000
0!
0'
0/
#559500000000
1!
1'
1/
#559510000000
0!
0'
0/
#559520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#559530000000
0!
0'
0/
#559540000000
1!
1'
1/
#559550000000
0!
1"
0'
1(
0/
10
#559560000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#559570000000
0!
1$
0'
1+
0/
#559580000000
1!
1'
1/
#559590000000
0!
0'
0/
#559600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#559610000000
0!
0'
0/
#559620000000
1!
1'
1/
#559630000000
0!
0'
0/
#559640000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#559650000000
0!
0'
0/
#559660000000
1!
1'
1/
#559670000000
0!
0'
0/
#559680000000
1!
1'
1/
#559690000000
0!
0'
0/
#559700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#559710000000
0!
0'
0/
#559720000000
1!
1'
1/
#559730000000
0!
0'
0/
#559740000000
1!
1'
1/
#559750000000
0!
0'
0/
#559760000000
1!
1'
1/
#559770000000
0!
0'
0/
#559780000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#559790000000
0!
0'
0/
#559800000000
1!
1'
1/
#559810000000
0!
0'
0/
#559820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#559830000000
0!
0'
0/
#559840000000
1!
1'
1/
#559850000000
0!
0'
0/
#559860000000
#559870000000
1!
1'
1/
#559880000000
0!
0'
0/
#559890000000
1!
1'
1/
#559900000000
0!
1"
0'
1(
0/
10
#559910000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#559920000000
0!
0'
0/
#559930000000
1!
1'
1/
#559940000000
0!
0'
0/
#559950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#559960000000
0!
0'
0/
#559970000000
1!
1'
1/
#559980000000
0!
1"
0'
1(
0/
10
#559990000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#560000000000
0!
1$
0'
1+
0/
#560010000000
1!
1'
1/
#560020000000
0!
0'
0/
#560030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#560040000000
0!
0'
0/
#560050000000
1!
1'
1/
#560060000000
0!
0'
0/
#560070000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#560080000000
0!
0'
0/
#560090000000
1!
1'
1/
#560100000000
0!
0'
0/
#560110000000
1!
1'
1/
#560120000000
0!
0'
0/
#560130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#560140000000
0!
0'
0/
#560150000000
1!
1'
1/
#560160000000
0!
0'
0/
#560170000000
1!
1'
1/
#560180000000
0!
0'
0/
#560190000000
1!
1'
1/
#560200000000
0!
0'
0/
#560210000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#560220000000
0!
0'
0/
#560230000000
1!
1'
1/
#560240000000
0!
0'
0/
#560250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#560260000000
0!
0'
0/
#560270000000
1!
1'
1/
#560280000000
0!
0'
0/
#560290000000
#560300000000
1!
1'
1/
#560310000000
0!
0'
0/
#560320000000
1!
1'
1/
#560330000000
0!
1"
0'
1(
0/
10
#560340000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#560350000000
0!
0'
0/
#560360000000
1!
1'
1/
#560370000000
0!
0'
0/
#560380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#560390000000
0!
0'
0/
#560400000000
1!
1'
1/
#560410000000
0!
1"
0'
1(
0/
10
#560420000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#560430000000
0!
1$
0'
1+
0/
#560440000000
1!
1'
1/
#560450000000
0!
0'
0/
#560460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#560470000000
0!
0'
0/
#560480000000
1!
1'
1/
#560490000000
0!
0'
0/
#560500000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#560510000000
0!
0'
0/
#560520000000
1!
1'
1/
#560530000000
0!
0'
0/
#560540000000
1!
1'
1/
#560550000000
0!
0'
0/
#560560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#560570000000
0!
0'
0/
#560580000000
1!
1'
1/
#560590000000
0!
0'
0/
#560600000000
1!
1'
1/
#560610000000
0!
0'
0/
#560620000000
1!
1'
1/
#560630000000
0!
0'
0/
#560640000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#560650000000
0!
0'
0/
#560660000000
1!
1'
1/
#560670000000
0!
0'
0/
#560680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#560690000000
0!
0'
0/
#560700000000
1!
1'
1/
#560710000000
0!
0'
0/
#560720000000
#560730000000
1!
1'
1/
#560740000000
0!
0'
0/
#560750000000
1!
1'
1/
#560760000000
0!
1"
0'
1(
0/
10
#560770000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#560780000000
0!
0'
0/
#560790000000
1!
1'
1/
#560800000000
0!
0'
0/
#560810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#560820000000
0!
0'
0/
#560830000000
1!
1'
1/
#560840000000
0!
1"
0'
1(
0/
10
#560850000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#560860000000
0!
1$
0'
1+
0/
#560870000000
1!
1'
1/
#560880000000
0!
0'
0/
#560890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#560900000000
0!
0'
0/
#560910000000
1!
1'
1/
#560920000000
0!
0'
0/
#560930000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#560940000000
0!
0'
0/
#560950000000
1!
1'
1/
#560960000000
0!
0'
0/
#560970000000
1!
1'
1/
#560980000000
0!
0'
0/
#560990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#561000000000
0!
0'
0/
#561010000000
1!
1'
1/
#561020000000
0!
0'
0/
#561030000000
1!
1'
1/
#561040000000
0!
0'
0/
#561050000000
1!
1'
1/
#561060000000
0!
0'
0/
#561070000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#561080000000
0!
0'
0/
#561090000000
1!
1'
1/
#561100000000
0!
0'
0/
#561110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#561120000000
0!
0'
0/
#561130000000
1!
1'
1/
#561140000000
0!
0'
0/
#561150000000
#561160000000
1!
1'
1/
#561170000000
0!
0'
0/
#561180000000
1!
1'
1/
#561190000000
0!
1"
0'
1(
0/
10
#561200000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#561210000000
0!
0'
0/
#561220000000
1!
1'
1/
#561230000000
0!
0'
0/
#561240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#561250000000
0!
0'
0/
#561260000000
1!
1'
1/
#561270000000
0!
1"
0'
1(
0/
10
#561280000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#561290000000
0!
1$
0'
1+
0/
#561300000000
1!
1'
1/
#561310000000
0!
0'
0/
#561320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#561330000000
0!
0'
0/
#561340000000
1!
1'
1/
#561350000000
0!
0'
0/
#561360000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#561370000000
0!
0'
0/
#561380000000
1!
1'
1/
#561390000000
0!
0'
0/
#561400000000
1!
1'
1/
#561410000000
0!
0'
0/
#561420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#561430000000
0!
0'
0/
#561440000000
1!
1'
1/
#561450000000
0!
0'
0/
#561460000000
1!
1'
1/
#561470000000
0!
0'
0/
#561480000000
1!
1'
1/
#561490000000
0!
0'
0/
#561500000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#561510000000
0!
0'
0/
#561520000000
1!
1'
1/
#561530000000
0!
0'
0/
#561540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#561550000000
0!
0'
0/
#561560000000
1!
1'
1/
#561570000000
0!
0'
0/
#561580000000
#561590000000
1!
1'
1/
#561600000000
0!
0'
0/
#561610000000
1!
1'
1/
#561620000000
0!
1"
0'
1(
0/
10
#561630000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#561640000000
0!
0'
0/
#561650000000
1!
1'
1/
#561660000000
0!
0'
0/
#561670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#561680000000
0!
0'
0/
#561690000000
1!
1'
1/
#561700000000
0!
1"
0'
1(
0/
10
#561710000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#561720000000
0!
1$
0'
1+
0/
#561730000000
1!
1'
1/
#561740000000
0!
0'
0/
#561750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#561760000000
0!
0'
0/
#561770000000
1!
1'
1/
#561780000000
0!
0'
0/
#561790000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#561800000000
0!
0'
0/
#561810000000
1!
1'
1/
#561820000000
0!
0'
0/
#561830000000
1!
1'
1/
#561840000000
0!
0'
0/
#561850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#561860000000
0!
0'
0/
#561870000000
1!
1'
1/
#561880000000
0!
0'
0/
#561890000000
1!
1'
1/
#561900000000
0!
0'
0/
#561910000000
1!
1'
1/
#561920000000
0!
0'
0/
#561930000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#561940000000
0!
0'
0/
#561950000000
1!
1'
1/
#561960000000
0!
0'
0/
#561970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#561980000000
0!
0'
0/
#561990000000
1!
1'
1/
#562000000000
0!
0'
0/
#562010000000
#562020000000
1!
1'
1/
#562030000000
0!
0'
0/
#562040000000
1!
1'
1/
#562050000000
0!
1"
0'
1(
0/
10
#562060000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#562070000000
0!
0'
0/
#562080000000
1!
1'
1/
#562090000000
0!
0'
0/
#562100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#562110000000
0!
0'
0/
#562120000000
1!
1'
1/
#562130000000
0!
1"
0'
1(
0/
10
#562140000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#562150000000
0!
1$
0'
1+
0/
#562160000000
1!
1'
1/
#562170000000
0!
0'
0/
#562180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#562190000000
0!
0'
0/
#562200000000
1!
1'
1/
#562210000000
0!
0'
0/
#562220000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#562230000000
0!
0'
0/
#562240000000
1!
1'
1/
#562250000000
0!
0'
0/
#562260000000
1!
1'
1/
#562270000000
0!
0'
0/
#562280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#562290000000
0!
0'
0/
#562300000000
1!
1'
1/
#562310000000
0!
0'
0/
#562320000000
1!
1'
1/
#562330000000
0!
0'
0/
#562340000000
1!
1'
1/
#562350000000
0!
0'
0/
#562360000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#562370000000
0!
0'
0/
#562380000000
1!
1'
1/
#562390000000
0!
0'
0/
#562400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#562410000000
0!
0'
0/
#562420000000
1!
1'
1/
#562430000000
0!
0'
0/
#562440000000
#562450000000
1!
1'
1/
#562460000000
0!
0'
0/
#562470000000
1!
1'
1/
#562480000000
0!
1"
0'
1(
0/
10
#562490000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#562500000000
0!
0'
0/
#562510000000
1!
1'
1/
#562520000000
0!
0'
0/
#562530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#562540000000
0!
0'
0/
#562550000000
1!
1'
1/
#562560000000
0!
1"
0'
1(
0/
10
#562570000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#562580000000
0!
1$
0'
1+
0/
#562590000000
1!
1'
1/
#562600000000
0!
0'
0/
#562610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#562620000000
0!
0'
0/
#562630000000
1!
1'
1/
#562640000000
0!
0'
0/
#562650000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#562660000000
0!
0'
0/
#562670000000
1!
1'
1/
#562680000000
0!
0'
0/
#562690000000
1!
1'
1/
#562700000000
0!
0'
0/
#562710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#562720000000
0!
0'
0/
#562730000000
1!
1'
1/
#562740000000
0!
0'
0/
#562750000000
1!
1'
1/
#562760000000
0!
0'
0/
#562770000000
1!
1'
1/
#562780000000
0!
0'
0/
#562790000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#562800000000
0!
0'
0/
#562810000000
1!
1'
1/
#562820000000
0!
0'
0/
#562830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#562840000000
0!
0'
0/
#562850000000
1!
1'
1/
#562860000000
0!
0'
0/
#562870000000
#562880000000
1!
1'
1/
#562890000000
0!
0'
0/
#562900000000
1!
1'
1/
#562910000000
0!
1"
0'
1(
0/
10
#562920000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#562930000000
0!
0'
0/
#562940000000
1!
1'
1/
#562950000000
0!
0'
0/
#562960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#562970000000
0!
0'
0/
#562980000000
1!
1'
1/
#562990000000
0!
1"
0'
1(
0/
10
#563000000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#563010000000
0!
1$
0'
1+
0/
#563020000000
1!
1'
1/
#563030000000
0!
0'
0/
#563040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#563050000000
0!
0'
0/
#563060000000
1!
1'
1/
#563070000000
0!
0'
0/
#563080000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#563090000000
0!
0'
0/
#563100000000
1!
1'
1/
#563110000000
0!
0'
0/
#563120000000
1!
1'
1/
#563130000000
0!
0'
0/
#563140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#563150000000
0!
0'
0/
#563160000000
1!
1'
1/
#563170000000
0!
0'
0/
#563180000000
1!
1'
1/
#563190000000
0!
0'
0/
#563200000000
1!
1'
1/
#563210000000
0!
0'
0/
#563220000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#563230000000
0!
0'
0/
#563240000000
1!
1'
1/
#563250000000
0!
0'
0/
#563260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#563270000000
0!
0'
0/
#563280000000
1!
1'
1/
#563290000000
0!
0'
0/
#563300000000
#563310000000
1!
1'
1/
#563320000000
0!
0'
0/
#563330000000
1!
1'
1/
#563340000000
0!
1"
0'
1(
0/
10
#563350000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#563360000000
0!
0'
0/
#563370000000
1!
1'
1/
#563380000000
0!
0'
0/
#563390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#563400000000
0!
0'
0/
#563410000000
1!
1'
1/
#563420000000
0!
1"
0'
1(
0/
10
#563430000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#563440000000
0!
1$
0'
1+
0/
#563450000000
1!
1'
1/
#563460000000
0!
0'
0/
#563470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#563480000000
0!
0'
0/
#563490000000
1!
1'
1/
#563500000000
0!
0'
0/
#563510000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#563520000000
0!
0'
0/
#563530000000
1!
1'
1/
#563540000000
0!
0'
0/
#563550000000
1!
1'
1/
#563560000000
0!
0'
0/
#563570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#563580000000
0!
0'
0/
#563590000000
1!
1'
1/
#563600000000
0!
0'
0/
#563610000000
1!
1'
1/
#563620000000
0!
0'
0/
#563630000000
1!
1'
1/
#563640000000
0!
0'
0/
#563650000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#563660000000
0!
0'
0/
#563670000000
1!
1'
1/
#563680000000
0!
0'
0/
#563690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#563700000000
0!
0'
0/
#563710000000
1!
1'
1/
#563720000000
0!
0'
0/
#563730000000
#563740000000
1!
1'
1/
#563750000000
0!
0'
0/
#563760000000
1!
1'
1/
#563770000000
0!
1"
0'
1(
0/
10
#563780000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#563790000000
0!
0'
0/
#563800000000
1!
1'
1/
#563810000000
0!
0'
0/
#563820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#563830000000
0!
0'
0/
#563840000000
1!
1'
1/
#563850000000
0!
1"
0'
1(
0/
10
#563860000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#563870000000
0!
1$
0'
1+
0/
#563880000000
1!
1'
1/
#563890000000
0!
0'
0/
#563900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#563910000000
0!
0'
0/
#563920000000
1!
1'
1/
#563930000000
0!
0'
0/
#563940000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#563950000000
0!
0'
0/
#563960000000
1!
1'
1/
#563970000000
0!
0'
0/
#563980000000
1!
1'
1/
#563990000000
0!
0'
0/
#564000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#564010000000
0!
0'
0/
#564020000000
1!
1'
1/
#564030000000
0!
0'
0/
#564040000000
1!
1'
1/
#564050000000
0!
0'
0/
#564060000000
1!
1'
1/
#564070000000
0!
0'
0/
#564080000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#564090000000
0!
0'
0/
#564100000000
1!
1'
1/
#564110000000
0!
0'
0/
#564120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#564130000000
0!
0'
0/
#564140000000
1!
1'
1/
#564150000000
0!
0'
0/
#564160000000
#564170000000
1!
1'
1/
#564180000000
0!
0'
0/
#564190000000
1!
1'
1/
#564200000000
0!
1"
0'
1(
0/
10
#564210000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#564220000000
0!
0'
0/
#564230000000
1!
1'
1/
#564240000000
0!
0'
0/
#564250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#564260000000
0!
0'
0/
#564270000000
1!
1'
1/
#564280000000
0!
1"
0'
1(
0/
10
#564290000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#564300000000
0!
1$
0'
1+
0/
#564310000000
1!
1'
1/
#564320000000
0!
0'
0/
#564330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#564340000000
0!
0'
0/
#564350000000
1!
1'
1/
#564360000000
0!
0'
0/
#564370000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#564380000000
0!
0'
0/
#564390000000
1!
1'
1/
#564400000000
0!
0'
0/
#564410000000
1!
1'
1/
#564420000000
0!
0'
0/
#564430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#564440000000
0!
0'
0/
#564450000000
1!
1'
1/
#564460000000
0!
0'
0/
#564470000000
1!
1'
1/
#564480000000
0!
0'
0/
#564490000000
1!
1'
1/
#564500000000
0!
0'
0/
#564510000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#564520000000
0!
0'
0/
#564530000000
1!
1'
1/
#564540000000
0!
0'
0/
#564550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#564560000000
0!
0'
0/
#564570000000
1!
1'
1/
#564580000000
0!
0'
0/
#564590000000
#564600000000
1!
1'
1/
#564610000000
0!
0'
0/
#564620000000
1!
1'
1/
#564630000000
0!
1"
0'
1(
0/
10
#564640000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#564650000000
0!
0'
0/
#564660000000
1!
1'
1/
#564670000000
0!
0'
0/
#564680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#564690000000
0!
0'
0/
#564700000000
1!
1'
1/
#564710000000
0!
1"
0'
1(
0/
10
#564720000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#564730000000
0!
1$
0'
1+
0/
#564740000000
1!
1'
1/
#564750000000
0!
0'
0/
#564760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#564770000000
0!
0'
0/
#564780000000
1!
1'
1/
#564790000000
0!
0'
0/
#564800000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#564810000000
0!
0'
0/
#564820000000
1!
1'
1/
#564830000000
0!
0'
0/
#564840000000
1!
1'
1/
#564850000000
0!
0'
0/
#564860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#564870000000
0!
0'
0/
#564880000000
1!
1'
1/
#564890000000
0!
0'
0/
#564900000000
1!
1'
1/
#564910000000
0!
0'
0/
#564920000000
1!
1'
1/
#564930000000
0!
0'
0/
#564940000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#564950000000
0!
0'
0/
#564960000000
1!
1'
1/
#564970000000
0!
0'
0/
#564980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#564990000000
0!
0'
0/
#565000000000
1!
1'
1/
#565010000000
0!
0'
0/
#565020000000
#565030000000
1!
1'
1/
#565040000000
0!
0'
0/
#565050000000
1!
1'
1/
#565060000000
0!
1"
0'
1(
0/
10
#565070000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#565080000000
0!
0'
0/
#565090000000
1!
1'
1/
#565100000000
0!
0'
0/
#565110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#565120000000
0!
0'
0/
#565130000000
1!
1'
1/
#565140000000
0!
1"
0'
1(
0/
10
#565150000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#565160000000
0!
1$
0'
1+
0/
#565170000000
1!
1'
1/
#565180000000
0!
0'
0/
#565190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#565200000000
0!
0'
0/
#565210000000
1!
1'
1/
#565220000000
0!
0'
0/
#565230000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#565240000000
0!
0'
0/
#565250000000
1!
1'
1/
#565260000000
0!
0'
0/
#565270000000
1!
1'
1/
#565280000000
0!
0'
0/
#565290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#565300000000
0!
0'
0/
#565310000000
1!
1'
1/
#565320000000
0!
0'
0/
#565330000000
1!
1'
1/
#565340000000
0!
0'
0/
#565350000000
1!
1'
1/
#565360000000
0!
0'
0/
#565370000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#565380000000
0!
0'
0/
#565390000000
1!
1'
1/
#565400000000
0!
0'
0/
#565410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#565420000000
0!
0'
0/
#565430000000
1!
1'
1/
#565440000000
0!
0'
0/
#565450000000
#565460000000
1!
1'
1/
#565470000000
0!
0'
0/
#565480000000
1!
1'
1/
#565490000000
0!
1"
0'
1(
0/
10
#565500000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#565510000000
0!
0'
0/
#565520000000
1!
1'
1/
#565530000000
0!
0'
0/
#565540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#565550000000
0!
0'
0/
#565560000000
1!
1'
1/
#565570000000
0!
1"
0'
1(
0/
10
#565580000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#565590000000
0!
1$
0'
1+
0/
#565600000000
1!
1'
1/
#565610000000
0!
0'
0/
#565620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#565630000000
0!
0'
0/
#565640000000
1!
1'
1/
#565650000000
0!
0'
0/
#565660000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#565670000000
0!
0'
0/
#565680000000
1!
1'
1/
#565690000000
0!
0'
0/
#565700000000
1!
1'
1/
#565710000000
0!
0'
0/
#565720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#565730000000
0!
0'
0/
#565740000000
1!
1'
1/
#565750000000
0!
0'
0/
#565760000000
1!
1'
1/
#565770000000
0!
0'
0/
#565780000000
1!
1'
1/
#565790000000
0!
0'
0/
#565800000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#565810000000
0!
0'
0/
#565820000000
1!
1'
1/
#565830000000
0!
0'
0/
#565840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#565850000000
0!
0'
0/
#565860000000
1!
1'
1/
#565870000000
0!
0'
0/
#565880000000
#565890000000
1!
1'
1/
#565900000000
0!
0'
0/
#565910000000
1!
1'
1/
#565920000000
0!
1"
0'
1(
0/
10
#565930000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#565940000000
0!
0'
0/
#565950000000
1!
1'
1/
#565960000000
0!
0'
0/
#565970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#565980000000
0!
0'
0/
#565990000000
1!
1'
1/
#566000000000
0!
1"
0'
1(
0/
10
#566010000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#566020000000
0!
1$
0'
1+
0/
#566030000000
1!
1'
1/
#566040000000
0!
0'
0/
#566050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#566060000000
0!
0'
0/
#566070000000
1!
1'
1/
#566080000000
0!
0'
0/
#566090000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#566100000000
0!
0'
0/
#566110000000
1!
1'
1/
#566120000000
0!
0'
0/
#566130000000
1!
1'
1/
#566140000000
0!
0'
0/
#566150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#566160000000
0!
0'
0/
#566170000000
1!
1'
1/
#566180000000
0!
0'
0/
#566190000000
1!
1'
1/
#566200000000
0!
0'
0/
#566210000000
1!
1'
1/
#566220000000
0!
0'
0/
#566230000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#566240000000
0!
0'
0/
#566250000000
1!
1'
1/
#566260000000
0!
0'
0/
#566270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#566280000000
0!
0'
0/
#566290000000
1!
1'
1/
#566300000000
0!
0'
0/
#566310000000
#566320000000
1!
1'
1/
#566330000000
0!
0'
0/
#566340000000
1!
1'
1/
#566350000000
0!
1"
0'
1(
0/
10
#566360000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#566370000000
0!
0'
0/
#566380000000
1!
1'
1/
#566390000000
0!
0'
0/
#566400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#566410000000
0!
0'
0/
#566420000000
1!
1'
1/
#566430000000
0!
1"
0'
1(
0/
10
#566440000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#566450000000
0!
1$
0'
1+
0/
#566460000000
1!
1'
1/
#566470000000
0!
0'
0/
#566480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#566490000000
0!
0'
0/
#566500000000
1!
1'
1/
#566510000000
0!
0'
0/
#566520000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#566530000000
0!
0'
0/
#566540000000
1!
1'
1/
#566550000000
0!
0'
0/
#566560000000
1!
1'
1/
#566570000000
0!
0'
0/
#566580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#566590000000
0!
0'
0/
#566600000000
1!
1'
1/
#566610000000
0!
0'
0/
#566620000000
1!
1'
1/
#566630000000
0!
0'
0/
#566640000000
1!
1'
1/
#566650000000
0!
0'
0/
#566660000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#566670000000
0!
0'
0/
#566680000000
1!
1'
1/
#566690000000
0!
0'
0/
#566700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#566710000000
0!
0'
0/
#566720000000
1!
1'
1/
#566730000000
0!
0'
0/
#566740000000
#566750000000
1!
1'
1/
#566760000000
0!
0'
0/
#566770000000
1!
1'
1/
#566780000000
0!
1"
0'
1(
0/
10
#566790000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#566800000000
0!
0'
0/
#566810000000
1!
1'
1/
#566820000000
0!
0'
0/
#566830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#566840000000
0!
0'
0/
#566850000000
1!
1'
1/
#566860000000
0!
1"
0'
1(
0/
10
#566870000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#566880000000
0!
1$
0'
1+
0/
#566890000000
1!
1'
1/
#566900000000
0!
0'
0/
#566910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#566920000000
0!
0'
0/
#566930000000
1!
1'
1/
#566940000000
0!
0'
0/
#566950000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#566960000000
0!
0'
0/
#566970000000
1!
1'
1/
#566980000000
0!
0'
0/
#566990000000
1!
1'
1/
#567000000000
0!
0'
0/
#567010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#567020000000
0!
0'
0/
#567030000000
1!
1'
1/
#567040000000
0!
0'
0/
#567050000000
1!
1'
1/
#567060000000
0!
0'
0/
#567070000000
1!
1'
1/
#567080000000
0!
0'
0/
#567090000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#567100000000
0!
0'
0/
#567110000000
1!
1'
1/
#567120000000
0!
0'
0/
#567130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#567140000000
0!
0'
0/
#567150000000
1!
1'
1/
#567160000000
0!
0'
0/
#567170000000
#567180000000
1!
1'
1/
#567190000000
0!
0'
0/
#567200000000
1!
1'
1/
#567210000000
0!
1"
0'
1(
0/
10
#567220000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#567230000000
0!
0'
0/
#567240000000
1!
1'
1/
#567250000000
0!
0'
0/
#567260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#567270000000
0!
0'
0/
#567280000000
1!
1'
1/
#567290000000
0!
1"
0'
1(
0/
10
#567300000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#567310000000
0!
1$
0'
1+
0/
#567320000000
1!
1'
1/
#567330000000
0!
0'
0/
#567340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#567350000000
0!
0'
0/
#567360000000
1!
1'
1/
#567370000000
0!
0'
0/
#567380000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#567390000000
0!
0'
0/
#567400000000
1!
1'
1/
#567410000000
0!
0'
0/
#567420000000
1!
1'
1/
#567430000000
0!
0'
0/
#567440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#567450000000
0!
0'
0/
#567460000000
1!
1'
1/
#567470000000
0!
0'
0/
#567480000000
1!
1'
1/
#567490000000
0!
0'
0/
#567500000000
1!
1'
1/
#567510000000
0!
0'
0/
#567520000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#567530000000
0!
0'
0/
#567540000000
1!
1'
1/
#567550000000
0!
0'
0/
#567560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#567570000000
0!
0'
0/
#567580000000
1!
1'
1/
#567590000000
0!
0'
0/
#567600000000
#567610000000
1!
1'
1/
#567620000000
0!
0'
0/
#567630000000
1!
1'
1/
#567640000000
0!
1"
0'
1(
0/
10
#567650000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#567660000000
0!
0'
0/
#567670000000
1!
1'
1/
#567680000000
0!
0'
0/
#567690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#567700000000
0!
0'
0/
#567710000000
1!
1'
1/
#567720000000
0!
1"
0'
1(
0/
10
#567730000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#567740000000
0!
1$
0'
1+
0/
#567750000000
1!
1'
1/
#567760000000
0!
0'
0/
#567770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#567780000000
0!
0'
0/
#567790000000
1!
1'
1/
#567800000000
0!
0'
0/
#567810000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#567820000000
0!
0'
0/
#567830000000
1!
1'
1/
#567840000000
0!
0'
0/
#567850000000
1!
1'
1/
#567860000000
0!
0'
0/
#567870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#567880000000
0!
0'
0/
#567890000000
1!
1'
1/
#567900000000
0!
0'
0/
#567910000000
1!
1'
1/
#567920000000
0!
0'
0/
#567930000000
1!
1'
1/
#567940000000
0!
0'
0/
#567950000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#567960000000
0!
0'
0/
#567970000000
1!
1'
1/
#567980000000
0!
0'
0/
#567990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#568000000000
0!
0'
0/
#568010000000
1!
1'
1/
#568020000000
0!
0'
0/
#568030000000
#568040000000
1!
1'
1/
#568050000000
0!
0'
0/
#568060000000
1!
1'
1/
#568070000000
0!
1"
0'
1(
0/
10
#568080000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#568090000000
0!
0'
0/
#568100000000
1!
1'
1/
#568110000000
0!
0'
0/
#568120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#568130000000
0!
0'
0/
#568140000000
1!
1'
1/
#568150000000
0!
1"
0'
1(
0/
10
#568160000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#568170000000
0!
1$
0'
1+
0/
#568180000000
1!
1'
1/
#568190000000
0!
0'
0/
#568200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#568210000000
0!
0'
0/
#568220000000
1!
1'
1/
#568230000000
0!
0'
0/
#568240000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#568250000000
0!
0'
0/
#568260000000
1!
1'
1/
#568270000000
0!
0'
0/
#568280000000
1!
1'
1/
#568290000000
0!
0'
0/
#568300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#568310000000
0!
0'
0/
#568320000000
1!
1'
1/
#568330000000
0!
0'
0/
#568340000000
1!
1'
1/
#568350000000
0!
0'
0/
#568360000000
1!
1'
1/
#568370000000
0!
0'
0/
#568380000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#568390000000
0!
0'
0/
#568400000000
1!
1'
1/
#568410000000
0!
0'
0/
#568420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#568430000000
0!
0'
0/
#568440000000
1!
1'
1/
#568450000000
0!
0'
0/
#568460000000
#568470000000
1!
1'
1/
#568480000000
0!
0'
0/
#568490000000
1!
1'
1/
#568500000000
0!
1"
0'
1(
0/
10
#568510000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#568520000000
0!
0'
0/
#568530000000
1!
1'
1/
#568540000000
0!
0'
0/
#568550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#568560000000
0!
0'
0/
#568570000000
1!
1'
1/
#568580000000
0!
1"
0'
1(
0/
10
#568590000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#568600000000
0!
1$
0'
1+
0/
#568610000000
1!
1'
1/
#568620000000
0!
0'
0/
#568630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#568640000000
0!
0'
0/
#568650000000
1!
1'
1/
#568660000000
0!
0'
0/
#568670000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#568680000000
0!
0'
0/
#568690000000
1!
1'
1/
#568700000000
0!
0'
0/
#568710000000
1!
1'
1/
#568720000000
0!
0'
0/
#568730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#568740000000
0!
0'
0/
#568750000000
1!
1'
1/
#568760000000
0!
0'
0/
#568770000000
1!
1'
1/
#568780000000
0!
0'
0/
#568790000000
1!
1'
1/
#568800000000
0!
0'
0/
#568810000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#568820000000
0!
0'
0/
#568830000000
1!
1'
1/
#568840000000
0!
0'
0/
#568850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#568860000000
0!
0'
0/
#568870000000
1!
1'
1/
#568880000000
0!
0'
0/
#568890000000
#568900000000
1!
1'
1/
#568910000000
0!
0'
0/
#568920000000
1!
1'
1/
#568930000000
0!
1"
0'
1(
0/
10
#568940000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#568950000000
0!
0'
0/
#568960000000
1!
1'
1/
#568970000000
0!
0'
0/
#568980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#568990000000
0!
0'
0/
#569000000000
1!
1'
1/
#569010000000
0!
1"
0'
1(
0/
10
#569020000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#569030000000
0!
1$
0'
1+
0/
#569040000000
1!
1'
1/
#569050000000
0!
0'
0/
#569060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#569070000000
0!
0'
0/
#569080000000
1!
1'
1/
#569090000000
0!
0'
0/
#569100000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#569110000000
0!
0'
0/
#569120000000
1!
1'
1/
#569130000000
0!
0'
0/
#569140000000
1!
1'
1/
#569150000000
0!
0'
0/
#569160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#569170000000
0!
0'
0/
#569180000000
1!
1'
1/
#569190000000
0!
0'
0/
#569200000000
1!
1'
1/
#569210000000
0!
0'
0/
#569220000000
1!
1'
1/
#569230000000
0!
0'
0/
#569240000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#569250000000
0!
0'
0/
#569260000000
1!
1'
1/
#569270000000
0!
0'
0/
#569280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#569290000000
0!
0'
0/
#569300000000
1!
1'
1/
#569310000000
0!
0'
0/
#569320000000
#569330000000
1!
1'
1/
#569340000000
0!
0'
0/
#569350000000
1!
1'
1/
#569360000000
0!
1"
0'
1(
0/
10
#569370000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#569380000000
0!
0'
0/
#569390000000
1!
1'
1/
#569400000000
0!
0'
0/
#569410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#569420000000
0!
0'
0/
#569430000000
1!
1'
1/
#569440000000
0!
1"
0'
1(
0/
10
#569450000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#569460000000
0!
1$
0'
1+
0/
#569470000000
1!
1'
1/
#569480000000
0!
0'
0/
#569490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#569500000000
0!
0'
0/
#569510000000
1!
1'
1/
#569520000000
0!
0'
0/
#569530000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#569540000000
0!
0'
0/
#569550000000
1!
1'
1/
#569560000000
0!
0'
0/
#569570000000
1!
1'
1/
#569580000000
0!
0'
0/
#569590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#569600000000
0!
0'
0/
#569610000000
1!
1'
1/
#569620000000
0!
0'
0/
#569630000000
1!
1'
1/
#569640000000
0!
0'
0/
#569650000000
1!
1'
1/
#569660000000
0!
0'
0/
#569670000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#569680000000
0!
0'
0/
#569690000000
1!
1'
1/
#569700000000
0!
0'
0/
#569710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#569720000000
0!
0'
0/
#569730000000
1!
1'
1/
#569740000000
0!
0'
0/
#569750000000
#569760000000
1!
1'
1/
#569770000000
0!
0'
0/
#569780000000
1!
1'
1/
#569790000000
0!
1"
0'
1(
0/
10
#569800000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#569810000000
0!
0'
0/
#569820000000
1!
1'
1/
#569830000000
0!
0'
0/
#569840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#569850000000
0!
0'
0/
#569860000000
1!
1'
1/
#569870000000
0!
1"
0'
1(
0/
10
#569880000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#569890000000
0!
1$
0'
1+
0/
#569900000000
1!
1'
1/
#569910000000
0!
0'
0/
#569920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#569930000000
0!
0'
0/
#569940000000
1!
1'
1/
#569950000000
0!
0'
0/
#569960000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#569970000000
0!
0'
0/
#569980000000
1!
1'
1/
#569990000000
0!
0'
0/
#570000000000
1!
1'
1/
#570010000000
0!
0'
0/
#570020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#570030000000
0!
0'
0/
#570040000000
1!
1'
1/
#570050000000
0!
0'
0/
#570060000000
1!
1'
1/
#570070000000
0!
0'
0/
#570080000000
1!
1'
1/
#570090000000
0!
0'
0/
#570100000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#570110000000
0!
0'
0/
#570120000000
1!
1'
1/
#570130000000
0!
0'
0/
#570140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#570150000000
0!
0'
0/
#570160000000
1!
1'
1/
#570170000000
0!
0'
0/
#570180000000
#570190000000
1!
1'
1/
#570200000000
0!
0'
0/
#570210000000
1!
1'
1/
#570220000000
0!
1"
0'
1(
0/
10
#570230000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#570240000000
0!
0'
0/
#570250000000
1!
1'
1/
#570260000000
0!
0'
0/
#570270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#570280000000
0!
0'
0/
#570290000000
1!
1'
1/
#570300000000
0!
1"
0'
1(
0/
10
#570310000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#570320000000
0!
1$
0'
1+
0/
#570330000000
1!
1'
1/
#570340000000
0!
0'
0/
#570350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#570360000000
0!
0'
0/
#570370000000
1!
1'
1/
#570380000000
0!
0'
0/
#570390000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#570400000000
0!
0'
0/
#570410000000
1!
1'
1/
#570420000000
0!
0'
0/
#570430000000
1!
1'
1/
#570440000000
0!
0'
0/
#570450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#570460000000
0!
0'
0/
#570470000000
1!
1'
1/
#570480000000
0!
0'
0/
#570490000000
1!
1'
1/
#570500000000
0!
0'
0/
#570510000000
1!
1'
1/
#570520000000
0!
0'
0/
#570530000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#570540000000
0!
0'
0/
#570550000000
1!
1'
1/
#570560000000
0!
0'
0/
#570570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#570580000000
0!
0'
0/
#570590000000
1!
1'
1/
#570600000000
0!
0'
0/
#570610000000
#570620000000
1!
1'
1/
#570630000000
0!
0'
0/
#570640000000
1!
1'
1/
#570650000000
0!
1"
0'
1(
0/
10
#570660000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#570670000000
0!
0'
0/
#570680000000
1!
1'
1/
#570690000000
0!
0'
0/
#570700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#570710000000
0!
0'
0/
#570720000000
1!
1'
1/
#570730000000
0!
1"
0'
1(
0/
10
#570740000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#570750000000
0!
1$
0'
1+
0/
#570760000000
1!
1'
1/
#570770000000
0!
0'
0/
#570780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#570790000000
0!
0'
0/
#570800000000
1!
1'
1/
#570810000000
0!
0'
0/
#570820000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#570830000000
0!
0'
0/
#570840000000
1!
1'
1/
#570850000000
0!
0'
0/
#570860000000
1!
1'
1/
#570870000000
0!
0'
0/
#570880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#570890000000
0!
0'
0/
#570900000000
1!
1'
1/
#570910000000
0!
0'
0/
#570920000000
1!
1'
1/
#570930000000
0!
0'
0/
#570940000000
1!
1'
1/
#570950000000
0!
0'
0/
#570960000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#570970000000
0!
0'
0/
#570980000000
1!
1'
1/
#570990000000
0!
0'
0/
#571000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#571010000000
0!
0'
0/
#571020000000
1!
1'
1/
#571030000000
0!
0'
0/
#571040000000
#571050000000
1!
1'
1/
#571060000000
0!
0'
0/
#571070000000
1!
1'
1/
#571080000000
0!
1"
0'
1(
0/
10
#571090000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#571100000000
0!
0'
0/
#571110000000
1!
1'
1/
#571120000000
0!
0'
0/
#571130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#571140000000
0!
0'
0/
#571150000000
1!
1'
1/
#571160000000
0!
1"
0'
1(
0/
10
#571170000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#571180000000
0!
1$
0'
1+
0/
#571190000000
1!
1'
1/
#571200000000
0!
0'
0/
#571210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#571220000000
0!
0'
0/
#571230000000
1!
1'
1/
#571240000000
0!
0'
0/
#571250000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#571260000000
0!
0'
0/
#571270000000
1!
1'
1/
#571280000000
0!
0'
0/
#571290000000
1!
1'
1/
#571300000000
0!
0'
0/
#571310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#571320000000
0!
0'
0/
#571330000000
1!
1'
1/
#571340000000
0!
0'
0/
#571350000000
1!
1'
1/
#571360000000
0!
0'
0/
#571370000000
1!
1'
1/
#571380000000
0!
0'
0/
#571390000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#571400000000
0!
0'
0/
#571410000000
1!
1'
1/
#571420000000
0!
0'
0/
#571430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#571440000000
0!
0'
0/
#571450000000
1!
1'
1/
#571460000000
0!
0'
0/
#571470000000
#571480000000
1!
1'
1/
#571490000000
0!
0'
0/
#571500000000
1!
1'
1/
#571510000000
0!
1"
0'
1(
0/
10
#571520000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#571530000000
0!
0'
0/
#571540000000
1!
1'
1/
#571550000000
0!
0'
0/
#571560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#571570000000
0!
0'
0/
#571580000000
1!
1'
1/
#571590000000
0!
1"
0'
1(
0/
10
#571600000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#571610000000
0!
1$
0'
1+
0/
#571620000000
1!
1'
1/
#571630000000
0!
0'
0/
#571640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#571650000000
0!
0'
0/
#571660000000
1!
1'
1/
#571670000000
0!
0'
0/
#571680000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#571690000000
0!
0'
0/
#571700000000
1!
1'
1/
#571710000000
0!
0'
0/
#571720000000
1!
1'
1/
#571730000000
0!
0'
0/
#571740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#571750000000
0!
0'
0/
#571760000000
1!
1'
1/
#571770000000
0!
0'
0/
#571780000000
1!
1'
1/
#571790000000
0!
0'
0/
#571800000000
1!
1'
1/
#571810000000
0!
0'
0/
#571820000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#571830000000
0!
0'
0/
#571840000000
1!
1'
1/
#571850000000
0!
0'
0/
#571860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#571870000000
0!
0'
0/
#571880000000
1!
1'
1/
#571890000000
0!
0'
0/
#571900000000
#571910000000
1!
1'
1/
#571920000000
0!
0'
0/
#571930000000
1!
1'
1/
#571940000000
0!
1"
0'
1(
0/
10
#571950000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#571960000000
0!
0'
0/
#571970000000
1!
1'
1/
#571980000000
0!
0'
0/
#571990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#572000000000
0!
0'
0/
#572010000000
1!
1'
1/
#572020000000
0!
1"
0'
1(
0/
10
#572030000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#572040000000
0!
1$
0'
1+
0/
#572050000000
1!
1'
1/
#572060000000
0!
0'
0/
#572070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#572080000000
0!
0'
0/
#572090000000
1!
1'
1/
#572100000000
0!
0'
0/
#572110000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#572120000000
0!
0'
0/
#572130000000
1!
1'
1/
#572140000000
0!
0'
0/
#572150000000
1!
1'
1/
#572160000000
0!
0'
0/
#572170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#572180000000
0!
0'
0/
#572190000000
1!
1'
1/
#572200000000
0!
0'
0/
#572210000000
1!
1'
1/
#572220000000
0!
0'
0/
#572230000000
1!
1'
1/
#572240000000
0!
0'
0/
#572250000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#572260000000
0!
0'
0/
#572270000000
1!
1'
1/
#572280000000
0!
0'
0/
#572290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#572300000000
0!
0'
0/
#572310000000
1!
1'
1/
#572320000000
0!
0'
0/
#572330000000
#572340000000
1!
1'
1/
#572350000000
0!
0'
0/
#572360000000
1!
1'
1/
#572370000000
0!
1"
0'
1(
0/
10
#572380000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#572390000000
0!
0'
0/
#572400000000
1!
1'
1/
#572410000000
0!
0'
0/
#572420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#572430000000
0!
0'
0/
#572440000000
1!
1'
1/
#572450000000
0!
1"
0'
1(
0/
10
#572460000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#572470000000
0!
1$
0'
1+
0/
#572480000000
1!
1'
1/
#572490000000
0!
0'
0/
#572500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#572510000000
0!
0'
0/
#572520000000
1!
1'
1/
#572530000000
0!
0'
0/
#572540000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#572550000000
0!
0'
0/
#572560000000
1!
1'
1/
#572570000000
0!
0'
0/
#572580000000
1!
1'
1/
#572590000000
0!
0'
0/
#572600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#572610000000
0!
0'
0/
#572620000000
1!
1'
1/
#572630000000
0!
0'
0/
#572640000000
1!
1'
1/
#572650000000
0!
0'
0/
#572660000000
1!
1'
1/
#572670000000
0!
0'
0/
#572680000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#572690000000
0!
0'
0/
#572700000000
1!
1'
1/
#572710000000
0!
0'
0/
#572720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#572730000000
0!
0'
0/
#572740000000
1!
1'
1/
#572750000000
0!
0'
0/
#572760000000
#572770000000
1!
1'
1/
#572780000000
0!
0'
0/
#572790000000
1!
1'
1/
#572800000000
0!
1"
0'
1(
0/
10
#572810000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#572820000000
0!
0'
0/
#572830000000
1!
1'
1/
#572840000000
0!
0'
0/
#572850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#572860000000
0!
0'
0/
#572870000000
1!
1'
1/
#572880000000
0!
1"
0'
1(
0/
10
#572890000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#572900000000
0!
1$
0'
1+
0/
#572910000000
1!
1'
1/
#572920000000
0!
0'
0/
#572930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#572940000000
0!
0'
0/
#572950000000
1!
1'
1/
#572960000000
0!
0'
0/
#572970000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#572980000000
0!
0'
0/
#572990000000
1!
1'
1/
#573000000000
0!
0'
0/
#573010000000
1!
1'
1/
#573020000000
0!
0'
0/
#573030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#573040000000
0!
0'
0/
#573050000000
1!
1'
1/
#573060000000
0!
0'
0/
#573070000000
1!
1'
1/
#573080000000
0!
0'
0/
#573090000000
1!
1'
1/
#573100000000
0!
0'
0/
#573110000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#573120000000
0!
0'
0/
#573130000000
1!
1'
1/
#573140000000
0!
0'
0/
#573150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#573160000000
0!
0'
0/
#573170000000
1!
1'
1/
#573180000000
0!
0'
0/
#573190000000
#573200000000
1!
1'
1/
#573210000000
0!
0'
0/
#573220000000
1!
1'
1/
#573230000000
0!
1"
0'
1(
0/
10
#573240000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#573250000000
0!
0'
0/
#573260000000
1!
1'
1/
#573270000000
0!
0'
0/
#573280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#573290000000
0!
0'
0/
#573300000000
1!
1'
1/
#573310000000
0!
1"
0'
1(
0/
10
#573320000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#573330000000
0!
1$
0'
1+
0/
#573340000000
1!
1'
1/
#573350000000
0!
0'
0/
#573360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#573370000000
0!
0'
0/
#573380000000
1!
1'
1/
#573390000000
0!
0'
0/
#573400000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#573410000000
0!
0'
0/
#573420000000
1!
1'
1/
#573430000000
0!
0'
0/
#573440000000
1!
1'
1/
#573450000000
0!
0'
0/
#573460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#573470000000
0!
0'
0/
#573480000000
1!
1'
1/
#573490000000
0!
0'
0/
#573500000000
1!
1'
1/
#573510000000
0!
0'
0/
#573520000000
1!
1'
1/
#573530000000
0!
0'
0/
#573540000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#573550000000
0!
0'
0/
#573560000000
1!
1'
1/
#573570000000
0!
0'
0/
#573580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#573590000000
0!
0'
0/
#573600000000
1!
1'
1/
#573610000000
0!
0'
0/
#573620000000
#573630000000
1!
1'
1/
#573640000000
0!
0'
0/
#573650000000
1!
1'
1/
#573660000000
0!
1"
0'
1(
0/
10
#573670000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#573680000000
0!
0'
0/
#573690000000
1!
1'
1/
#573700000000
0!
0'
0/
#573710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#573720000000
0!
0'
0/
#573730000000
1!
1'
1/
#573740000000
0!
1"
0'
1(
0/
10
#573750000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#573760000000
0!
1$
0'
1+
0/
#573770000000
1!
1'
1/
#573780000000
0!
0'
0/
#573790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#573800000000
0!
0'
0/
#573810000000
1!
1'
1/
#573820000000
0!
0'
0/
#573830000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#573840000000
0!
0'
0/
#573850000000
1!
1'
1/
#573860000000
0!
0'
0/
#573870000000
1!
1'
1/
#573880000000
0!
0'
0/
#573890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#573900000000
0!
0'
0/
#573910000000
1!
1'
1/
#573920000000
0!
0'
0/
#573930000000
1!
1'
1/
#573940000000
0!
0'
0/
#573950000000
1!
1'
1/
#573960000000
0!
0'
0/
#573970000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#573980000000
0!
0'
0/
#573990000000
1!
1'
1/
#574000000000
0!
0'
0/
#574010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#574020000000
0!
0'
0/
#574030000000
1!
1'
1/
#574040000000
0!
0'
0/
#574050000000
#574060000000
1!
1'
1/
#574070000000
0!
0'
0/
#574080000000
1!
1'
1/
#574090000000
0!
1"
0'
1(
0/
10
#574100000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#574110000000
0!
0'
0/
#574120000000
1!
1'
1/
#574130000000
0!
0'
0/
#574140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#574150000000
0!
0'
0/
#574160000000
1!
1'
1/
#574170000000
0!
1"
0'
1(
0/
10
#574180000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#574190000000
0!
1$
0'
1+
0/
#574200000000
1!
1'
1/
#574210000000
0!
0'
0/
#574220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#574230000000
0!
0'
0/
#574240000000
1!
1'
1/
#574250000000
0!
0'
0/
#574260000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#574270000000
0!
0'
0/
#574280000000
1!
1'
1/
#574290000000
0!
0'
0/
#574300000000
1!
1'
1/
#574310000000
0!
0'
0/
#574320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#574330000000
0!
0'
0/
#574340000000
1!
1'
1/
#574350000000
0!
0'
0/
#574360000000
1!
1'
1/
#574370000000
0!
0'
0/
#574380000000
1!
1'
1/
#574390000000
0!
0'
0/
#574400000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#574410000000
0!
0'
0/
#574420000000
1!
1'
1/
#574430000000
0!
0'
0/
#574440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#574450000000
0!
0'
0/
#574460000000
1!
1'
1/
#574470000000
0!
0'
0/
#574480000000
#574490000000
1!
1'
1/
#574500000000
0!
0'
0/
#574510000000
1!
1'
1/
#574520000000
0!
1"
0'
1(
0/
10
#574530000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#574540000000
0!
0'
0/
#574550000000
1!
1'
1/
#574560000000
0!
0'
0/
#574570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#574580000000
0!
0'
0/
#574590000000
1!
1'
1/
#574600000000
0!
1"
0'
1(
0/
10
#574610000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#574620000000
0!
1$
0'
1+
0/
#574630000000
1!
1'
1/
#574640000000
0!
0'
0/
#574650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#574660000000
0!
0'
0/
#574670000000
1!
1'
1/
#574680000000
0!
0'
0/
#574690000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#574700000000
0!
0'
0/
#574710000000
1!
1'
1/
#574720000000
0!
0'
0/
#574730000000
1!
1'
1/
#574740000000
0!
0'
0/
#574750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#574760000000
0!
0'
0/
#574770000000
1!
1'
1/
#574780000000
0!
0'
0/
#574790000000
1!
1'
1/
#574800000000
0!
0'
0/
#574810000000
1!
1'
1/
#574820000000
0!
0'
0/
#574830000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#574840000000
0!
0'
0/
#574850000000
1!
1'
1/
#574860000000
0!
0'
0/
#574870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#574880000000
0!
0'
0/
#574890000000
1!
1'
1/
#574900000000
0!
0'
0/
#574910000000
#574920000000
1!
1'
1/
#574930000000
0!
0'
0/
#574940000000
1!
1'
1/
#574950000000
0!
1"
0'
1(
0/
10
#574960000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#574970000000
0!
0'
0/
#574980000000
1!
1'
1/
#574990000000
0!
0'
0/
#575000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#575010000000
0!
0'
0/
#575020000000
1!
1'
1/
#575030000000
0!
1"
0'
1(
0/
10
#575040000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#575050000000
0!
1$
0'
1+
0/
#575060000000
1!
1'
1/
#575070000000
0!
0'
0/
#575080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#575090000000
0!
0'
0/
#575100000000
1!
1'
1/
#575110000000
0!
0'
0/
#575120000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#575130000000
0!
0'
0/
#575140000000
1!
1'
1/
#575150000000
0!
0'
0/
#575160000000
1!
1'
1/
#575170000000
0!
0'
0/
#575180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#575190000000
0!
0'
0/
#575200000000
1!
1'
1/
#575210000000
0!
0'
0/
#575220000000
1!
1'
1/
#575230000000
0!
0'
0/
#575240000000
1!
1'
1/
#575250000000
0!
0'
0/
#575260000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#575270000000
0!
0'
0/
#575280000000
1!
1'
1/
#575290000000
0!
0'
0/
#575300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#575310000000
0!
0'
0/
#575320000000
1!
1'
1/
#575330000000
0!
0'
0/
#575340000000
#575350000000
1!
1'
1/
#575360000000
0!
0'
0/
#575370000000
1!
1'
1/
#575380000000
0!
1"
0'
1(
0/
10
#575390000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#575400000000
0!
0'
0/
#575410000000
1!
1'
1/
#575420000000
0!
0'
0/
#575430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#575440000000
0!
0'
0/
#575450000000
1!
1'
1/
#575460000000
0!
1"
0'
1(
0/
10
#575470000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#575480000000
0!
1$
0'
1+
0/
#575490000000
1!
1'
1/
#575500000000
0!
0'
0/
#575510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#575520000000
0!
0'
0/
#575530000000
1!
1'
1/
#575540000000
0!
0'
0/
#575550000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#575560000000
0!
0'
0/
#575570000000
1!
1'
1/
#575580000000
0!
0'
0/
#575590000000
1!
1'
1/
#575600000000
0!
0'
0/
#575610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#575620000000
0!
0'
0/
#575630000000
1!
1'
1/
#575640000000
0!
0'
0/
#575650000000
1!
1'
1/
#575660000000
0!
0'
0/
#575670000000
1!
1'
1/
#575680000000
0!
0'
0/
#575690000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#575700000000
0!
0'
0/
#575710000000
1!
1'
1/
#575720000000
0!
0'
0/
#575730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#575740000000
0!
0'
0/
#575750000000
1!
1'
1/
#575760000000
0!
0'
0/
#575770000000
#575780000000
1!
1'
1/
#575790000000
0!
0'
0/
#575800000000
1!
1'
1/
#575810000000
0!
1"
0'
1(
0/
10
#575820000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#575830000000
0!
0'
0/
#575840000000
1!
1'
1/
#575850000000
0!
0'
0/
#575860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#575870000000
0!
0'
0/
#575880000000
1!
1'
1/
#575890000000
0!
1"
0'
1(
0/
10
#575900000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#575910000000
0!
1$
0'
1+
0/
#575920000000
1!
1'
1/
#575930000000
0!
0'
0/
#575940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#575950000000
0!
0'
0/
#575960000000
1!
1'
1/
#575970000000
0!
0'
0/
#575980000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#575990000000
0!
0'
0/
#576000000000
1!
1'
1/
#576010000000
0!
0'
0/
#576020000000
1!
1'
1/
#576030000000
0!
0'
0/
#576040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#576050000000
0!
0'
0/
#576060000000
1!
1'
1/
#576070000000
0!
0'
0/
#576080000000
1!
1'
1/
#576090000000
0!
0'
0/
#576100000000
1!
1'
1/
#576110000000
0!
0'
0/
#576120000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#576130000000
0!
0'
0/
#576140000000
1!
1'
1/
#576150000000
0!
0'
0/
#576160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#576170000000
0!
0'
0/
#576180000000
1!
1'
1/
#576190000000
0!
0'
0/
#576200000000
#576210000000
1!
1'
1/
#576220000000
0!
0'
0/
#576230000000
1!
1'
1/
#576240000000
0!
1"
0'
1(
0/
10
#576250000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#576260000000
0!
0'
0/
#576270000000
1!
1'
1/
#576280000000
0!
0'
0/
#576290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#576300000000
0!
0'
0/
#576310000000
1!
1'
1/
#576320000000
0!
1"
0'
1(
0/
10
#576330000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#576340000000
0!
1$
0'
1+
0/
#576350000000
1!
1'
1/
#576360000000
0!
0'
0/
#576370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#576380000000
0!
0'
0/
#576390000000
1!
1'
1/
#576400000000
0!
0'
0/
#576410000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#576420000000
0!
0'
0/
#576430000000
1!
1'
1/
#576440000000
0!
0'
0/
#576450000000
1!
1'
1/
#576460000000
0!
0'
0/
#576470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#576480000000
0!
0'
0/
#576490000000
1!
1'
1/
#576500000000
0!
0'
0/
#576510000000
1!
1'
1/
#576520000000
0!
0'
0/
#576530000000
1!
1'
1/
#576540000000
0!
0'
0/
#576550000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#576560000000
0!
0'
0/
#576570000000
1!
1'
1/
#576580000000
0!
0'
0/
#576590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#576600000000
0!
0'
0/
#576610000000
1!
1'
1/
#576620000000
0!
0'
0/
#576630000000
#576640000000
1!
1'
1/
#576650000000
0!
0'
0/
#576660000000
1!
1'
1/
#576670000000
0!
1"
0'
1(
0/
10
#576680000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#576690000000
0!
0'
0/
#576700000000
1!
1'
1/
#576710000000
0!
0'
0/
#576720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#576730000000
0!
0'
0/
#576740000000
1!
1'
1/
#576750000000
0!
1"
0'
1(
0/
10
#576760000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#576770000000
0!
1$
0'
1+
0/
#576780000000
1!
1'
1/
#576790000000
0!
0'
0/
#576800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#576810000000
0!
0'
0/
#576820000000
1!
1'
1/
#576830000000
0!
0'
0/
#576840000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#576850000000
0!
0'
0/
#576860000000
1!
1'
1/
#576870000000
0!
0'
0/
#576880000000
1!
1'
1/
#576890000000
0!
0'
0/
#576900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#576910000000
0!
0'
0/
#576920000000
1!
1'
1/
#576930000000
0!
0'
0/
#576940000000
1!
1'
1/
#576950000000
0!
0'
0/
#576960000000
1!
1'
1/
#576970000000
0!
0'
0/
#576980000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#576990000000
0!
0'
0/
#577000000000
1!
1'
1/
#577010000000
0!
0'
0/
#577020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#577030000000
0!
0'
0/
#577040000000
1!
1'
1/
#577050000000
0!
0'
0/
#577060000000
#577070000000
1!
1'
1/
#577080000000
0!
0'
0/
#577090000000
1!
1'
1/
#577100000000
0!
1"
0'
1(
0/
10
#577110000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#577120000000
0!
0'
0/
#577130000000
1!
1'
1/
#577140000000
0!
0'
0/
#577150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#577160000000
0!
0'
0/
#577170000000
1!
1'
1/
#577180000000
0!
1"
0'
1(
0/
10
#577190000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#577200000000
0!
1$
0'
1+
0/
#577210000000
1!
1'
1/
#577220000000
0!
0'
0/
#577230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#577240000000
0!
0'
0/
#577250000000
1!
1'
1/
#577260000000
0!
0'
0/
#577270000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#577280000000
0!
0'
0/
#577290000000
1!
1'
1/
#577300000000
0!
0'
0/
#577310000000
1!
1'
1/
#577320000000
0!
0'
0/
#577330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#577340000000
0!
0'
0/
#577350000000
1!
1'
1/
#577360000000
0!
0'
0/
#577370000000
1!
1'
1/
#577380000000
0!
0'
0/
#577390000000
1!
1'
1/
#577400000000
0!
0'
0/
#577410000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#577420000000
0!
0'
0/
#577430000000
1!
1'
1/
#577440000000
0!
0'
0/
#577450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#577460000000
0!
0'
0/
#577470000000
1!
1'
1/
#577480000000
0!
0'
0/
#577490000000
#577500000000
1!
1'
1/
#577510000000
0!
0'
0/
#577520000000
1!
1'
1/
#577530000000
0!
1"
0'
1(
0/
10
#577540000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#577550000000
0!
0'
0/
#577560000000
1!
1'
1/
#577570000000
0!
0'
0/
#577580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#577590000000
0!
0'
0/
#577600000000
1!
1'
1/
#577610000000
0!
1"
0'
1(
0/
10
#577620000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#577630000000
0!
1$
0'
1+
0/
#577640000000
1!
1'
1/
#577650000000
0!
0'
0/
#577660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#577670000000
0!
0'
0/
#577680000000
1!
1'
1/
#577690000000
0!
0'
0/
#577700000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#577710000000
0!
0'
0/
#577720000000
1!
1'
1/
#577730000000
0!
0'
0/
#577740000000
1!
1'
1/
#577750000000
0!
0'
0/
#577760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#577770000000
0!
0'
0/
#577780000000
1!
1'
1/
#577790000000
0!
0'
0/
#577800000000
1!
1'
1/
#577810000000
0!
0'
0/
#577820000000
1!
1'
1/
#577830000000
0!
0'
0/
#577840000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#577850000000
0!
0'
0/
#577860000000
1!
1'
1/
#577870000000
0!
0'
0/
#577880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#577890000000
0!
0'
0/
#577900000000
1!
1'
1/
#577910000000
0!
0'
0/
#577920000000
#577930000000
1!
1'
1/
#577940000000
0!
0'
0/
#577950000000
1!
1'
1/
#577960000000
0!
1"
0'
1(
0/
10
#577970000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#577980000000
0!
0'
0/
#577990000000
1!
1'
1/
#578000000000
0!
0'
0/
#578010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#578020000000
0!
0'
0/
#578030000000
1!
1'
1/
#578040000000
0!
1"
0'
1(
0/
10
#578050000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#578060000000
0!
1$
0'
1+
0/
#578070000000
1!
1'
1/
#578080000000
0!
0'
0/
#578090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#578100000000
0!
0'
0/
#578110000000
1!
1'
1/
#578120000000
0!
0'
0/
#578130000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#578140000000
0!
0'
0/
#578150000000
1!
1'
1/
#578160000000
0!
0'
0/
#578170000000
1!
1'
1/
#578180000000
0!
0'
0/
#578190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#578200000000
0!
0'
0/
#578210000000
1!
1'
1/
#578220000000
0!
0'
0/
#578230000000
1!
1'
1/
#578240000000
0!
0'
0/
#578250000000
1!
1'
1/
#578260000000
0!
0'
0/
#578270000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#578280000000
0!
0'
0/
#578290000000
1!
1'
1/
#578300000000
0!
0'
0/
#578310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#578320000000
0!
0'
0/
#578330000000
1!
1'
1/
#578340000000
0!
0'
0/
#578350000000
#578360000000
1!
1'
1/
#578370000000
0!
0'
0/
#578380000000
1!
1'
1/
#578390000000
0!
1"
0'
1(
0/
10
#578400000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#578410000000
0!
0'
0/
#578420000000
1!
1'
1/
#578430000000
0!
0'
0/
#578440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#578450000000
0!
0'
0/
#578460000000
1!
1'
1/
#578470000000
0!
1"
0'
1(
0/
10
#578480000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#578490000000
0!
1$
0'
1+
0/
#578500000000
1!
1'
1/
#578510000000
0!
0'
0/
#578520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#578530000000
0!
0'
0/
#578540000000
1!
1'
1/
#578550000000
0!
0'
0/
#578560000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#578570000000
0!
0'
0/
#578580000000
1!
1'
1/
#578590000000
0!
0'
0/
#578600000000
1!
1'
1/
#578610000000
0!
0'
0/
#578620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#578630000000
0!
0'
0/
#578640000000
1!
1'
1/
#578650000000
0!
0'
0/
#578660000000
1!
1'
1/
#578670000000
0!
0'
0/
#578680000000
1!
1'
1/
#578690000000
0!
0'
0/
#578700000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#578710000000
0!
0'
0/
#578720000000
1!
1'
1/
#578730000000
0!
0'
0/
#578740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#578750000000
0!
0'
0/
#578760000000
1!
1'
1/
#578770000000
0!
0'
0/
#578780000000
#578790000000
1!
1'
1/
#578800000000
0!
0'
0/
#578810000000
1!
1'
1/
#578820000000
0!
1"
0'
1(
0/
10
#578830000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#578840000000
0!
0'
0/
#578850000000
1!
1'
1/
#578860000000
0!
0'
0/
#578870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#578880000000
0!
0'
0/
#578890000000
1!
1'
1/
#578900000000
0!
1"
0'
1(
0/
10
#578910000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#578920000000
0!
1$
0'
1+
0/
#578930000000
1!
1'
1/
#578940000000
0!
0'
0/
#578950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#578960000000
0!
0'
0/
#578970000000
1!
1'
1/
#578980000000
0!
0'
0/
#578990000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#579000000000
0!
0'
0/
#579010000000
1!
1'
1/
#579020000000
0!
0'
0/
#579030000000
1!
1'
1/
#579040000000
0!
0'
0/
#579050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#579060000000
0!
0'
0/
#579070000000
1!
1'
1/
#579080000000
0!
0'
0/
#579090000000
1!
1'
1/
#579100000000
0!
0'
0/
#579110000000
1!
1'
1/
#579120000000
0!
0'
0/
#579130000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#579140000000
0!
0'
0/
#579150000000
1!
1'
1/
#579160000000
0!
0'
0/
#579170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#579180000000
0!
0'
0/
#579190000000
1!
1'
1/
#579200000000
0!
0'
0/
#579210000000
#579220000000
1!
1'
1/
#579230000000
0!
0'
0/
#579240000000
1!
1'
1/
#579250000000
0!
1"
0'
1(
0/
10
#579260000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#579270000000
0!
0'
0/
#579280000000
1!
1'
1/
#579290000000
0!
0'
0/
#579300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#579310000000
0!
0'
0/
#579320000000
1!
1'
1/
#579330000000
0!
1"
0'
1(
0/
10
#579340000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#579350000000
0!
1$
0'
1+
0/
#579360000000
1!
1'
1/
#579370000000
0!
0'
0/
#579380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#579390000000
0!
0'
0/
#579400000000
1!
1'
1/
#579410000000
0!
0'
0/
#579420000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#579430000000
0!
0'
0/
#579440000000
1!
1'
1/
#579450000000
0!
0'
0/
#579460000000
1!
1'
1/
#579470000000
0!
0'
0/
#579480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#579490000000
0!
0'
0/
#579500000000
1!
1'
1/
#579510000000
0!
0'
0/
#579520000000
1!
1'
1/
#579530000000
0!
0'
0/
#579540000000
1!
1'
1/
#579550000000
0!
0'
0/
#579560000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#579570000000
0!
0'
0/
#579580000000
1!
1'
1/
#579590000000
0!
0'
0/
#579600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#579610000000
0!
0'
0/
#579620000000
1!
1'
1/
#579630000000
0!
0'
0/
#579640000000
#579650000000
1!
1'
1/
#579660000000
0!
0'
0/
#579670000000
1!
1'
1/
#579680000000
0!
1"
0'
1(
0/
10
#579690000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#579700000000
0!
0'
0/
#579710000000
1!
1'
1/
#579720000000
0!
0'
0/
#579730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#579740000000
0!
0'
0/
#579750000000
1!
1'
1/
#579760000000
0!
1"
0'
1(
0/
10
#579770000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#579780000000
0!
1$
0'
1+
0/
#579790000000
1!
1'
1/
#579800000000
0!
0'
0/
#579810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#579820000000
0!
0'
0/
#579830000000
1!
1'
1/
#579840000000
0!
0'
0/
#579850000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#579860000000
0!
0'
0/
#579870000000
1!
1'
1/
#579880000000
0!
0'
0/
#579890000000
1!
1'
1/
#579900000000
0!
0'
0/
#579910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#579920000000
0!
0'
0/
#579930000000
1!
1'
1/
#579940000000
0!
0'
0/
#579950000000
1!
1'
1/
#579960000000
0!
0'
0/
#579970000000
1!
1'
1/
#579980000000
0!
0'
0/
#579990000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#580000000000
0!
0'
0/
#580010000000
1!
1'
1/
#580020000000
0!
0'
0/
#580030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#580040000000
0!
0'
0/
#580050000000
1!
1'
1/
#580060000000
0!
0'
0/
#580070000000
#580080000000
1!
1'
1/
#580090000000
0!
0'
0/
#580100000000
1!
1'
1/
#580110000000
0!
1"
0'
1(
0/
10
#580120000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#580130000000
0!
0'
0/
#580140000000
1!
1'
1/
#580150000000
0!
0'
0/
#580160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#580170000000
0!
0'
0/
#580180000000
1!
1'
1/
#580190000000
0!
1"
0'
1(
0/
10
#580200000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#580210000000
0!
1$
0'
1+
0/
#580220000000
1!
1'
1/
#580230000000
0!
0'
0/
#580240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#580250000000
0!
0'
0/
#580260000000
1!
1'
1/
#580270000000
0!
0'
0/
#580280000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#580290000000
0!
0'
0/
#580300000000
1!
1'
1/
#580310000000
0!
0'
0/
#580320000000
1!
1'
1/
#580330000000
0!
0'
0/
#580340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#580350000000
0!
0'
0/
#580360000000
1!
1'
1/
#580370000000
0!
0'
0/
#580380000000
1!
1'
1/
#580390000000
0!
0'
0/
#580400000000
1!
1'
1/
#580410000000
0!
0'
0/
#580420000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#580430000000
0!
0'
0/
#580440000000
1!
1'
1/
#580450000000
0!
0'
0/
#580460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#580470000000
0!
0'
0/
#580480000000
1!
1'
1/
#580490000000
0!
0'
0/
#580500000000
#580510000000
1!
1'
1/
#580520000000
0!
0'
0/
#580530000000
1!
1'
1/
#580540000000
0!
1"
0'
1(
0/
10
#580550000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#580560000000
0!
0'
0/
#580570000000
1!
1'
1/
#580580000000
0!
0'
0/
#580590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#580600000000
0!
0'
0/
#580610000000
1!
1'
1/
#580620000000
0!
1"
0'
1(
0/
10
#580630000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#580640000000
0!
1$
0'
1+
0/
#580650000000
1!
1'
1/
#580660000000
0!
0'
0/
#580670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#580680000000
0!
0'
0/
#580690000000
1!
1'
1/
#580700000000
0!
0'
0/
#580710000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#580720000000
0!
0'
0/
#580730000000
1!
1'
1/
#580740000000
0!
0'
0/
#580750000000
1!
1'
1/
#580760000000
0!
0'
0/
#580770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#580780000000
0!
0'
0/
#580790000000
1!
1'
1/
#580800000000
0!
0'
0/
#580810000000
1!
1'
1/
#580820000000
0!
0'
0/
#580830000000
1!
1'
1/
#580840000000
0!
0'
0/
#580850000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#580860000000
0!
0'
0/
#580870000000
1!
1'
1/
#580880000000
0!
0'
0/
#580890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#580900000000
0!
0'
0/
#580910000000
1!
1'
1/
#580920000000
0!
0'
0/
#580930000000
#580940000000
1!
1'
1/
#580950000000
0!
0'
0/
#580960000000
1!
1'
1/
#580970000000
0!
1"
0'
1(
0/
10
#580980000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#580990000000
0!
0'
0/
#581000000000
1!
1'
1/
#581010000000
0!
0'
0/
#581020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#581030000000
0!
0'
0/
#581040000000
1!
1'
1/
#581050000000
0!
1"
0'
1(
0/
10
#581060000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#581070000000
0!
1$
0'
1+
0/
#581080000000
1!
1'
1/
#581090000000
0!
0'
0/
#581100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#581110000000
0!
0'
0/
#581120000000
1!
1'
1/
#581130000000
0!
0'
0/
#581140000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#581150000000
0!
0'
0/
#581160000000
1!
1'
1/
#581170000000
0!
0'
0/
#581180000000
1!
1'
1/
#581190000000
0!
0'
0/
#581200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#581210000000
0!
0'
0/
#581220000000
1!
1'
1/
#581230000000
0!
0'
0/
#581240000000
1!
1'
1/
#581250000000
0!
0'
0/
#581260000000
1!
1'
1/
#581270000000
0!
0'
0/
#581280000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#581290000000
0!
0'
0/
#581300000000
1!
1'
1/
#581310000000
0!
0'
0/
#581320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#581330000000
0!
0'
0/
#581340000000
1!
1'
1/
#581350000000
0!
0'
0/
#581360000000
#581370000000
1!
1'
1/
#581380000000
0!
0'
0/
#581390000000
1!
1'
1/
#581400000000
0!
1"
0'
1(
0/
10
#581410000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#581420000000
0!
0'
0/
#581430000000
1!
1'
1/
#581440000000
0!
0'
0/
#581450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#581460000000
0!
0'
0/
#581470000000
1!
1'
1/
#581480000000
0!
1"
0'
1(
0/
10
#581490000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#581500000000
0!
1$
0'
1+
0/
#581510000000
1!
1'
1/
#581520000000
0!
0'
0/
#581530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#581540000000
0!
0'
0/
#581550000000
1!
1'
1/
#581560000000
0!
0'
0/
#581570000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#581580000000
0!
0'
0/
#581590000000
1!
1'
1/
#581600000000
0!
0'
0/
#581610000000
1!
1'
1/
#581620000000
0!
0'
0/
#581630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#581640000000
0!
0'
0/
#581650000000
1!
1'
1/
#581660000000
0!
0'
0/
#581670000000
1!
1'
1/
#581680000000
0!
0'
0/
#581690000000
1!
1'
1/
#581700000000
0!
0'
0/
#581710000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#581720000000
0!
0'
0/
#581730000000
1!
1'
1/
#581740000000
0!
0'
0/
#581750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#581760000000
0!
0'
0/
#581770000000
1!
1'
1/
#581780000000
0!
0'
0/
#581790000000
#581800000000
1!
1'
1/
#581810000000
0!
0'
0/
#581820000000
1!
1'
1/
#581830000000
0!
1"
0'
1(
0/
10
#581840000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#581850000000
0!
0'
0/
#581860000000
1!
1'
1/
#581870000000
0!
0'
0/
#581880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#581890000000
0!
0'
0/
#581900000000
1!
1'
1/
#581910000000
0!
1"
0'
1(
0/
10
#581920000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#581930000000
0!
1$
0'
1+
0/
#581940000000
1!
1'
1/
#581950000000
0!
0'
0/
#581960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#581970000000
0!
0'
0/
#581980000000
1!
1'
1/
#581990000000
0!
0'
0/
#582000000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#582010000000
0!
0'
0/
#582020000000
1!
1'
1/
#582030000000
0!
0'
0/
#582040000000
1!
1'
1/
#582050000000
0!
0'
0/
#582060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#582070000000
0!
0'
0/
#582080000000
1!
1'
1/
#582090000000
0!
0'
0/
#582100000000
1!
1'
1/
#582110000000
0!
0'
0/
#582120000000
1!
1'
1/
#582130000000
0!
0'
0/
#582140000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#582150000000
0!
0'
0/
#582160000000
1!
1'
1/
#582170000000
0!
0'
0/
#582180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#582190000000
0!
0'
0/
#582200000000
1!
1'
1/
#582210000000
0!
0'
0/
#582220000000
#582230000000
1!
1'
1/
#582240000000
0!
0'
0/
#582250000000
1!
1'
1/
#582260000000
0!
1"
0'
1(
0/
10
#582270000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#582280000000
0!
0'
0/
#582290000000
1!
1'
1/
#582300000000
0!
0'
0/
#582310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#582320000000
0!
0'
0/
#582330000000
1!
1'
1/
#582340000000
0!
1"
0'
1(
0/
10
#582350000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#582360000000
0!
1$
0'
1+
0/
#582370000000
1!
1'
1/
#582380000000
0!
0'
0/
#582390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#582400000000
0!
0'
0/
#582410000000
1!
1'
1/
#582420000000
0!
0'
0/
#582430000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#582440000000
0!
0'
0/
#582450000000
1!
1'
1/
#582460000000
0!
0'
0/
#582470000000
1!
1'
1/
#582480000000
0!
0'
0/
#582490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#582500000000
0!
0'
0/
#582510000000
1!
1'
1/
#582520000000
0!
0'
0/
#582530000000
1!
1'
1/
#582540000000
0!
0'
0/
#582550000000
1!
1'
1/
#582560000000
0!
0'
0/
#582570000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#582580000000
0!
0'
0/
#582590000000
1!
1'
1/
#582600000000
0!
0'
0/
#582610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#582620000000
0!
0'
0/
#582630000000
1!
1'
1/
#582640000000
0!
0'
0/
#582650000000
#582660000000
1!
1'
1/
#582670000000
0!
0'
0/
#582680000000
1!
1'
1/
#582690000000
0!
1"
0'
1(
0/
10
#582700000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#582710000000
0!
0'
0/
#582720000000
1!
1'
1/
#582730000000
0!
0'
0/
#582740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#582750000000
0!
0'
0/
#582760000000
1!
1'
1/
#582770000000
0!
1"
0'
1(
0/
10
#582780000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#582790000000
0!
1$
0'
1+
0/
#582800000000
1!
1'
1/
#582810000000
0!
0'
0/
#582820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#582830000000
0!
0'
0/
#582840000000
1!
1'
1/
#582850000000
0!
0'
0/
#582860000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#582870000000
0!
0'
0/
#582880000000
1!
1'
1/
#582890000000
0!
0'
0/
#582900000000
1!
1'
1/
#582910000000
0!
0'
0/
#582920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#582930000000
0!
0'
0/
#582940000000
1!
1'
1/
#582950000000
0!
0'
0/
#582960000000
1!
1'
1/
#582970000000
0!
0'
0/
#582980000000
1!
1'
1/
#582990000000
0!
0'
0/
#583000000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#583010000000
0!
0'
0/
#583020000000
1!
1'
1/
#583030000000
0!
0'
0/
#583040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#583050000000
0!
0'
0/
#583060000000
1!
1'
1/
#583070000000
0!
0'
0/
#583080000000
#583090000000
1!
1'
1/
#583100000000
0!
0'
0/
#583110000000
1!
1'
1/
#583120000000
0!
1"
0'
1(
0/
10
#583130000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#583140000000
0!
0'
0/
#583150000000
1!
1'
1/
#583160000000
0!
0'
0/
#583170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#583180000000
0!
0'
0/
#583190000000
1!
1'
1/
#583200000000
0!
1"
0'
1(
0/
10
#583210000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#583220000000
0!
1$
0'
1+
0/
#583230000000
1!
1'
1/
#583240000000
0!
0'
0/
#583250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#583260000000
0!
0'
0/
#583270000000
1!
1'
1/
#583280000000
0!
0'
0/
#583290000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#583300000000
0!
0'
0/
#583310000000
1!
1'
1/
#583320000000
0!
0'
0/
#583330000000
1!
1'
1/
#583340000000
0!
0'
0/
#583350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#583360000000
0!
0'
0/
#583370000000
1!
1'
1/
#583380000000
0!
0'
0/
#583390000000
1!
1'
1/
#583400000000
0!
0'
0/
#583410000000
1!
1'
1/
#583420000000
0!
0'
0/
#583430000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#583440000000
0!
0'
0/
#583450000000
1!
1'
1/
#583460000000
0!
0'
0/
#583470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#583480000000
0!
0'
0/
#583490000000
1!
1'
1/
#583500000000
0!
0'
0/
#583510000000
#583520000000
1!
1'
1/
#583530000000
0!
0'
0/
#583540000000
1!
1'
1/
#583550000000
0!
1"
0'
1(
0/
10
#583560000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#583570000000
0!
0'
0/
#583580000000
1!
1'
1/
#583590000000
0!
0'
0/
#583600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#583610000000
0!
0'
0/
#583620000000
1!
1'
1/
#583630000000
0!
1"
0'
1(
0/
10
#583640000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#583650000000
0!
1$
0'
1+
0/
#583660000000
1!
1'
1/
#583670000000
0!
0'
0/
#583680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#583690000000
0!
0'
0/
#583700000000
1!
1'
1/
#583710000000
0!
0'
0/
#583720000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#583730000000
0!
0'
0/
#583740000000
1!
1'
1/
#583750000000
0!
0'
0/
#583760000000
1!
1'
1/
#583770000000
0!
0'
0/
#583780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#583790000000
0!
0'
0/
#583800000000
1!
1'
1/
#583810000000
0!
0'
0/
#583820000000
1!
1'
1/
#583830000000
0!
0'
0/
#583840000000
1!
1'
1/
#583850000000
0!
0'
0/
#583860000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#583870000000
0!
0'
0/
#583880000000
1!
1'
1/
#583890000000
0!
0'
0/
#583900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#583910000000
0!
0'
0/
#583920000000
1!
1'
1/
#583930000000
0!
0'
0/
#583940000000
#583950000000
1!
1'
1/
#583960000000
0!
0'
0/
#583970000000
1!
1'
1/
#583980000000
0!
1"
0'
1(
0/
10
#583990000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#584000000000
0!
0'
0/
#584010000000
1!
1'
1/
#584020000000
0!
0'
0/
#584030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#584040000000
0!
0'
0/
#584050000000
1!
1'
1/
#584060000000
0!
1"
0'
1(
0/
10
#584070000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#584080000000
0!
1$
0'
1+
0/
#584090000000
1!
1'
1/
#584100000000
0!
0'
0/
#584110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#584120000000
0!
0'
0/
#584130000000
1!
1'
1/
#584140000000
0!
0'
0/
#584150000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#584160000000
0!
0'
0/
#584170000000
1!
1'
1/
#584180000000
0!
0'
0/
#584190000000
1!
1'
1/
#584200000000
0!
0'
0/
#584210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#584220000000
0!
0'
0/
#584230000000
1!
1'
1/
#584240000000
0!
0'
0/
#584250000000
1!
1'
1/
#584260000000
0!
0'
0/
#584270000000
1!
1'
1/
#584280000000
0!
0'
0/
#584290000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#584300000000
0!
0'
0/
#584310000000
1!
1'
1/
#584320000000
0!
0'
0/
#584330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#584340000000
0!
0'
0/
#584350000000
1!
1'
1/
#584360000000
0!
0'
0/
#584370000000
#584380000000
1!
1'
1/
#584390000000
0!
0'
0/
#584400000000
1!
1'
1/
#584410000000
0!
1"
0'
1(
0/
10
#584420000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#584430000000
0!
0'
0/
#584440000000
1!
1'
1/
#584450000000
0!
0'
0/
#584460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#584470000000
0!
0'
0/
#584480000000
1!
1'
1/
#584490000000
0!
1"
0'
1(
0/
10
#584500000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#584510000000
0!
1$
0'
1+
0/
#584520000000
1!
1'
1/
#584530000000
0!
0'
0/
#584540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#584550000000
0!
0'
0/
#584560000000
1!
1'
1/
#584570000000
0!
0'
0/
#584580000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#584590000000
0!
0'
0/
#584600000000
1!
1'
1/
#584610000000
0!
0'
0/
#584620000000
1!
1'
1/
#584630000000
0!
0'
0/
#584640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#584650000000
0!
0'
0/
#584660000000
1!
1'
1/
#584670000000
0!
0'
0/
#584680000000
1!
1'
1/
#584690000000
0!
0'
0/
#584700000000
1!
1'
1/
#584710000000
0!
0'
0/
#584720000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#584730000000
0!
0'
0/
#584740000000
1!
1'
1/
#584750000000
0!
0'
0/
#584760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#584770000000
0!
0'
0/
#584780000000
1!
1'
1/
#584790000000
0!
0'
0/
#584800000000
#584810000000
1!
1'
1/
#584820000000
0!
0'
0/
#584830000000
1!
1'
1/
#584840000000
0!
1"
0'
1(
0/
10
#584850000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#584860000000
0!
0'
0/
#584870000000
1!
1'
1/
#584880000000
0!
0'
0/
#584890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#584900000000
0!
0'
0/
#584910000000
1!
1'
1/
#584920000000
0!
1"
0'
1(
0/
10
#584930000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#584940000000
0!
1$
0'
1+
0/
#584950000000
1!
1'
1/
#584960000000
0!
0'
0/
#584970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#584980000000
0!
0'
0/
#584990000000
1!
1'
1/
#585000000000
0!
0'
0/
#585010000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#585020000000
0!
0'
0/
#585030000000
1!
1'
1/
#585040000000
0!
0'
0/
#585050000000
1!
1'
1/
#585060000000
0!
0'
0/
#585070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#585080000000
0!
0'
0/
#585090000000
1!
1'
1/
#585100000000
0!
0'
0/
#585110000000
1!
1'
1/
#585120000000
0!
0'
0/
#585130000000
1!
1'
1/
#585140000000
0!
0'
0/
#585150000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#585160000000
0!
0'
0/
#585170000000
1!
1'
1/
#585180000000
0!
0'
0/
#585190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#585200000000
0!
0'
0/
#585210000000
1!
1'
1/
#585220000000
0!
0'
0/
#585230000000
#585240000000
1!
1'
1/
#585250000000
0!
0'
0/
#585260000000
1!
1'
1/
#585270000000
0!
1"
0'
1(
0/
10
#585280000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#585290000000
0!
0'
0/
#585300000000
1!
1'
1/
#585310000000
0!
0'
0/
#585320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#585330000000
0!
0'
0/
#585340000000
1!
1'
1/
#585350000000
0!
1"
0'
1(
0/
10
#585360000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#585370000000
0!
1$
0'
1+
0/
#585380000000
1!
1'
1/
#585390000000
0!
0'
0/
#585400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#585410000000
0!
0'
0/
#585420000000
1!
1'
1/
#585430000000
0!
0'
0/
#585440000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#585450000000
0!
0'
0/
#585460000000
1!
1'
1/
#585470000000
0!
0'
0/
#585480000000
1!
1'
1/
#585490000000
0!
0'
0/
#585500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#585510000000
0!
0'
0/
#585520000000
1!
1'
1/
#585530000000
0!
0'
0/
#585540000000
1!
1'
1/
#585550000000
0!
0'
0/
#585560000000
1!
1'
1/
#585570000000
0!
0'
0/
#585580000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#585590000000
0!
0'
0/
#585600000000
1!
1'
1/
#585610000000
0!
0'
0/
#585620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#585630000000
0!
0'
0/
#585640000000
1!
1'
1/
#585650000000
0!
0'
0/
#585660000000
#585670000000
1!
1'
1/
#585680000000
0!
0'
0/
#585690000000
1!
1'
1/
#585700000000
0!
1"
0'
1(
0/
10
#585710000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#585720000000
0!
0'
0/
#585730000000
1!
1'
1/
#585740000000
0!
0'
0/
#585750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#585760000000
0!
0'
0/
#585770000000
1!
1'
1/
#585780000000
0!
1"
0'
1(
0/
10
#585790000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#585800000000
0!
1$
0'
1+
0/
#585810000000
1!
1'
1/
#585820000000
0!
0'
0/
#585830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#585840000000
0!
0'
0/
#585850000000
1!
1'
1/
#585860000000
0!
0'
0/
#585870000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#585880000000
0!
0'
0/
#585890000000
1!
1'
1/
#585900000000
0!
0'
0/
#585910000000
1!
1'
1/
#585920000000
0!
0'
0/
#585930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#585940000000
0!
0'
0/
#585950000000
1!
1'
1/
#585960000000
0!
0'
0/
#585970000000
1!
1'
1/
#585980000000
0!
0'
0/
#585990000000
1!
1'
1/
#586000000000
0!
0'
0/
#586010000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#586020000000
0!
0'
0/
#586030000000
1!
1'
1/
#586040000000
0!
0'
0/
#586050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#586060000000
0!
0'
0/
#586070000000
1!
1'
1/
#586080000000
0!
0'
0/
#586090000000
#586100000000
1!
1'
1/
#586110000000
0!
0'
0/
#586120000000
1!
1'
1/
#586130000000
0!
1"
0'
1(
0/
10
#586140000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#586150000000
0!
0'
0/
#586160000000
1!
1'
1/
#586170000000
0!
0'
0/
#586180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#586190000000
0!
0'
0/
#586200000000
1!
1'
1/
#586210000000
0!
1"
0'
1(
0/
10
#586220000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#586230000000
0!
1$
0'
1+
0/
#586240000000
1!
1'
1/
#586250000000
0!
0'
0/
#586260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#586270000000
0!
0'
0/
#586280000000
1!
1'
1/
#586290000000
0!
0'
0/
#586300000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#586310000000
0!
0'
0/
#586320000000
1!
1'
1/
#586330000000
0!
0'
0/
#586340000000
1!
1'
1/
#586350000000
0!
0'
0/
#586360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#586370000000
0!
0'
0/
#586380000000
1!
1'
1/
#586390000000
0!
0'
0/
#586400000000
1!
1'
1/
#586410000000
0!
0'
0/
#586420000000
1!
1'
1/
#586430000000
0!
0'
0/
#586440000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#586450000000
0!
0'
0/
#586460000000
1!
1'
1/
#586470000000
0!
0'
0/
#586480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#586490000000
0!
0'
0/
#586500000000
1!
1'
1/
#586510000000
0!
0'
0/
#586520000000
#586530000000
1!
1'
1/
#586540000000
0!
0'
0/
#586550000000
1!
1'
1/
#586560000000
0!
1"
0'
1(
0/
10
#586570000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#586580000000
0!
0'
0/
#586590000000
1!
1'
1/
#586600000000
0!
0'
0/
#586610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#586620000000
0!
0'
0/
#586630000000
1!
1'
1/
#586640000000
0!
1"
0'
1(
0/
10
#586650000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#586660000000
0!
1$
0'
1+
0/
#586670000000
1!
1'
1/
#586680000000
0!
0'
0/
#586690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#586700000000
0!
0'
0/
#586710000000
1!
1'
1/
#586720000000
0!
0'
0/
#586730000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#586740000000
0!
0'
0/
#586750000000
1!
1'
1/
#586760000000
0!
0'
0/
#586770000000
1!
1'
1/
#586780000000
0!
0'
0/
#586790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#586800000000
0!
0'
0/
#586810000000
1!
1'
1/
#586820000000
0!
0'
0/
#586830000000
1!
1'
1/
#586840000000
0!
0'
0/
#586850000000
1!
1'
1/
#586860000000
0!
0'
0/
#586870000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#586880000000
0!
0'
0/
#586890000000
1!
1'
1/
#586900000000
0!
0'
0/
#586910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#586920000000
0!
0'
0/
#586930000000
1!
1'
1/
#586940000000
0!
0'
0/
#586950000000
#586960000000
1!
1'
1/
#586970000000
0!
0'
0/
#586980000000
1!
1'
1/
#586990000000
0!
1"
0'
1(
0/
10
#587000000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#587010000000
0!
0'
0/
#587020000000
1!
1'
1/
#587030000000
0!
0'
0/
#587040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#587050000000
0!
0'
0/
#587060000000
1!
1'
1/
#587070000000
0!
1"
0'
1(
0/
10
#587080000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#587090000000
0!
1$
0'
1+
0/
#587100000000
1!
1'
1/
#587110000000
0!
0'
0/
#587120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#587130000000
0!
0'
0/
#587140000000
1!
1'
1/
#587150000000
0!
0'
0/
#587160000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#587170000000
0!
0'
0/
#587180000000
1!
1'
1/
#587190000000
0!
0'
0/
#587200000000
1!
1'
1/
#587210000000
0!
0'
0/
#587220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#587230000000
0!
0'
0/
#587240000000
1!
1'
1/
#587250000000
0!
0'
0/
#587260000000
1!
1'
1/
#587270000000
0!
0'
0/
#587280000000
1!
1'
1/
#587290000000
0!
0'
0/
#587300000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#587310000000
0!
0'
0/
#587320000000
1!
1'
1/
#587330000000
0!
0'
0/
#587340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#587350000000
0!
0'
0/
#587360000000
1!
1'
1/
#587370000000
0!
0'
0/
#587380000000
#587390000000
1!
1'
1/
#587400000000
0!
0'
0/
#587410000000
1!
1'
1/
#587420000000
0!
1"
0'
1(
0/
10
#587430000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#587440000000
0!
0'
0/
#587450000000
1!
1'
1/
#587460000000
0!
0'
0/
#587470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#587480000000
0!
0'
0/
#587490000000
1!
1'
1/
#587500000000
0!
1"
0'
1(
0/
10
#587510000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#587520000000
0!
1$
0'
1+
0/
#587530000000
1!
1'
1/
#587540000000
0!
0'
0/
#587550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#587560000000
0!
0'
0/
#587570000000
1!
1'
1/
#587580000000
0!
0'
0/
#587590000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#587600000000
0!
0'
0/
#587610000000
1!
1'
1/
#587620000000
0!
0'
0/
#587630000000
1!
1'
1/
#587640000000
0!
0'
0/
#587650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#587660000000
0!
0'
0/
#587670000000
1!
1'
1/
#587680000000
0!
0'
0/
#587690000000
1!
1'
1/
#587700000000
0!
0'
0/
#587710000000
1!
1'
1/
#587720000000
0!
0'
0/
#587730000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#587740000000
0!
0'
0/
#587750000000
1!
1'
1/
#587760000000
0!
0'
0/
#587770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#587780000000
0!
0'
0/
#587790000000
1!
1'
1/
#587800000000
0!
0'
0/
#587810000000
#587820000000
1!
1'
1/
#587830000000
0!
0'
0/
#587840000000
1!
1'
1/
#587850000000
0!
1"
0'
1(
0/
10
#587860000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#587870000000
0!
0'
0/
#587880000000
1!
1'
1/
#587890000000
0!
0'
0/
#587900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#587910000000
0!
0'
0/
#587920000000
1!
1'
1/
#587930000000
0!
1"
0'
1(
0/
10
#587940000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#587950000000
0!
1$
0'
1+
0/
#587960000000
1!
1'
1/
#587970000000
0!
0'
0/
#587980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#587990000000
0!
0'
0/
#588000000000
1!
1'
1/
#588010000000
0!
0'
0/
#588020000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#588030000000
0!
0'
0/
#588040000000
1!
1'
1/
#588050000000
0!
0'
0/
#588060000000
1!
1'
1/
#588070000000
0!
0'
0/
#588080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#588090000000
0!
0'
0/
#588100000000
1!
1'
1/
#588110000000
0!
0'
0/
#588120000000
1!
1'
1/
#588130000000
0!
0'
0/
#588140000000
1!
1'
1/
#588150000000
0!
0'
0/
#588160000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#588170000000
0!
0'
0/
#588180000000
1!
1'
1/
#588190000000
0!
0'
0/
#588200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#588210000000
0!
0'
0/
#588220000000
1!
1'
1/
#588230000000
0!
0'
0/
#588240000000
#588250000000
1!
1'
1/
#588260000000
0!
0'
0/
#588270000000
1!
1'
1/
#588280000000
0!
1"
0'
1(
0/
10
#588290000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#588300000000
0!
0'
0/
#588310000000
1!
1'
1/
#588320000000
0!
0'
0/
#588330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#588340000000
0!
0'
0/
#588350000000
1!
1'
1/
#588360000000
0!
1"
0'
1(
0/
10
#588370000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#588380000000
0!
1$
0'
1+
0/
#588390000000
1!
1'
1/
#588400000000
0!
0'
0/
#588410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#588420000000
0!
0'
0/
#588430000000
1!
1'
1/
#588440000000
0!
0'
0/
#588450000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#588460000000
0!
0'
0/
#588470000000
1!
1'
1/
#588480000000
0!
0'
0/
#588490000000
1!
1'
1/
#588500000000
0!
0'
0/
#588510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#588520000000
0!
0'
0/
#588530000000
1!
1'
1/
#588540000000
0!
0'
0/
#588550000000
1!
1'
1/
#588560000000
0!
0'
0/
#588570000000
1!
1'
1/
#588580000000
0!
0'
0/
#588590000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#588600000000
0!
0'
0/
#588610000000
1!
1'
1/
#588620000000
0!
0'
0/
#588630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#588640000000
0!
0'
0/
#588650000000
1!
1'
1/
#588660000000
0!
0'
0/
#588670000000
#588680000000
1!
1'
1/
#588690000000
0!
0'
0/
#588700000000
1!
1'
1/
#588710000000
0!
1"
0'
1(
0/
10
#588720000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#588730000000
0!
0'
0/
#588740000000
1!
1'
1/
#588750000000
0!
0'
0/
#588760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#588770000000
0!
0'
0/
#588780000000
1!
1'
1/
#588790000000
0!
1"
0'
1(
0/
10
#588800000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#588810000000
0!
1$
0'
1+
0/
#588820000000
1!
1'
1/
#588830000000
0!
0'
0/
#588840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#588850000000
0!
0'
0/
#588860000000
1!
1'
1/
#588870000000
0!
0'
0/
#588880000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#588890000000
0!
0'
0/
#588900000000
1!
1'
1/
#588910000000
0!
0'
0/
#588920000000
1!
1'
1/
#588930000000
0!
0'
0/
#588940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#588950000000
0!
0'
0/
#588960000000
1!
1'
1/
#588970000000
0!
0'
0/
#588980000000
1!
1'
1/
#588990000000
0!
0'
0/
#589000000000
1!
1'
1/
#589010000000
0!
0'
0/
#589020000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#589030000000
0!
0'
0/
#589040000000
1!
1'
1/
#589050000000
0!
0'
0/
#589060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#589070000000
0!
0'
0/
#589080000000
1!
1'
1/
#589090000000
0!
0'
0/
#589100000000
#589110000000
1!
1'
1/
#589120000000
0!
0'
0/
#589130000000
1!
1'
1/
#589140000000
0!
1"
0'
1(
0/
10
#589150000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#589160000000
0!
0'
0/
#589170000000
1!
1'
1/
#589180000000
0!
0'
0/
#589190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#589200000000
0!
0'
0/
#589210000000
1!
1'
1/
#589220000000
0!
1"
0'
1(
0/
10
#589230000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#589240000000
0!
1$
0'
1+
0/
#589250000000
1!
1'
1/
#589260000000
0!
0'
0/
#589270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#589280000000
0!
0'
0/
#589290000000
1!
1'
1/
#589300000000
0!
0'
0/
#589310000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#589320000000
0!
0'
0/
#589330000000
1!
1'
1/
#589340000000
0!
0'
0/
#589350000000
1!
1'
1/
#589360000000
0!
0'
0/
#589370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#589380000000
0!
0'
0/
#589390000000
1!
1'
1/
#589400000000
0!
0'
0/
#589410000000
1!
1'
1/
#589420000000
0!
0'
0/
#589430000000
1!
1'
1/
#589440000000
0!
0'
0/
#589450000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#589460000000
0!
0'
0/
#589470000000
1!
1'
1/
#589480000000
0!
0'
0/
#589490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#589500000000
0!
0'
0/
#589510000000
1!
1'
1/
#589520000000
0!
0'
0/
#589530000000
#589540000000
1!
1'
1/
#589550000000
0!
0'
0/
#589560000000
1!
1'
1/
#589570000000
0!
1"
0'
1(
0/
10
#589580000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#589590000000
0!
0'
0/
#589600000000
1!
1'
1/
#589610000000
0!
0'
0/
#589620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#589630000000
0!
0'
0/
#589640000000
1!
1'
1/
#589650000000
0!
1"
0'
1(
0/
10
#589660000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#589670000000
0!
1$
0'
1+
0/
#589680000000
1!
1'
1/
#589690000000
0!
0'
0/
#589700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#589710000000
0!
0'
0/
#589720000000
1!
1'
1/
#589730000000
0!
0'
0/
#589740000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#589750000000
0!
0'
0/
#589760000000
1!
1'
1/
#589770000000
0!
0'
0/
#589780000000
1!
1'
1/
#589790000000
0!
0'
0/
#589800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#589810000000
0!
0'
0/
#589820000000
1!
1'
1/
#589830000000
0!
0'
0/
#589840000000
1!
1'
1/
#589850000000
0!
0'
0/
#589860000000
1!
1'
1/
#589870000000
0!
0'
0/
#589880000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#589890000000
0!
0'
0/
#589900000000
1!
1'
1/
#589910000000
0!
0'
0/
#589920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#589930000000
0!
0'
0/
#589940000000
1!
1'
1/
#589950000000
0!
0'
0/
#589960000000
#589970000000
1!
1'
1/
#589980000000
0!
0'
0/
#589990000000
1!
1'
1/
#590000000000
0!
1"
0'
1(
0/
10
#590010000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#590020000000
0!
0'
0/
#590030000000
1!
1'
1/
#590040000000
0!
0'
0/
#590050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#590060000000
0!
0'
0/
#590070000000
1!
1'
1/
#590080000000
0!
1"
0'
1(
0/
10
#590090000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#590100000000
0!
1$
0'
1+
0/
#590110000000
1!
1'
1/
#590120000000
0!
0'
0/
#590130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#590140000000
0!
0'
0/
#590150000000
1!
1'
1/
#590160000000
0!
0'
0/
#590170000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#590180000000
0!
0'
0/
#590190000000
1!
1'
1/
#590200000000
0!
0'
0/
#590210000000
1!
1'
1/
#590220000000
0!
0'
0/
#590230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#590240000000
0!
0'
0/
#590250000000
1!
1'
1/
#590260000000
0!
0'
0/
#590270000000
1!
1'
1/
#590280000000
0!
0'
0/
#590290000000
1!
1'
1/
#590300000000
0!
0'
0/
#590310000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#590320000000
0!
0'
0/
#590330000000
1!
1'
1/
#590340000000
0!
0'
0/
#590350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#590360000000
0!
0'
0/
#590370000000
1!
1'
1/
#590380000000
0!
0'
0/
#590390000000
#590400000000
1!
1'
1/
#590410000000
0!
0'
0/
#590420000000
1!
1'
1/
#590430000000
0!
1"
0'
1(
0/
10
#590440000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#590450000000
0!
0'
0/
#590460000000
1!
1'
1/
#590470000000
0!
0'
0/
#590480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#590490000000
0!
0'
0/
#590500000000
1!
1'
1/
#590510000000
0!
1"
0'
1(
0/
10
#590520000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#590530000000
0!
1$
0'
1+
0/
#590540000000
1!
1'
1/
#590550000000
0!
0'
0/
#590560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#590570000000
0!
0'
0/
#590580000000
1!
1'
1/
#590590000000
0!
0'
0/
#590600000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#590610000000
0!
0'
0/
#590620000000
1!
1'
1/
#590630000000
0!
0'
0/
#590640000000
1!
1'
1/
#590650000000
0!
0'
0/
#590660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#590670000000
0!
0'
0/
#590680000000
1!
1'
1/
#590690000000
0!
0'
0/
#590700000000
1!
1'
1/
#590710000000
0!
0'
0/
#590720000000
1!
1'
1/
#590730000000
0!
0'
0/
#590740000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#590750000000
0!
0'
0/
#590760000000
1!
1'
1/
#590770000000
0!
0'
0/
#590780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#590790000000
0!
0'
0/
#590800000000
1!
1'
1/
#590810000000
0!
0'
0/
#590820000000
#590830000000
1!
1'
1/
#590840000000
0!
0'
0/
#590850000000
1!
1'
1/
#590860000000
0!
1"
0'
1(
0/
10
#590870000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#590880000000
0!
0'
0/
#590890000000
1!
1'
1/
#590900000000
0!
0'
0/
#590910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#590920000000
0!
0'
0/
#590930000000
1!
1'
1/
#590940000000
0!
1"
0'
1(
0/
10
#590950000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#590960000000
0!
1$
0'
1+
0/
#590970000000
1!
1'
1/
#590980000000
0!
0'
0/
#590990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#591000000000
0!
0'
0/
#591010000000
1!
1'
1/
#591020000000
0!
0'
0/
#591030000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#591040000000
0!
0'
0/
#591050000000
1!
1'
1/
#591060000000
0!
0'
0/
#591070000000
1!
1'
1/
#591080000000
0!
0'
0/
#591090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#591100000000
0!
0'
0/
#591110000000
1!
1'
1/
#591120000000
0!
0'
0/
#591130000000
1!
1'
1/
#591140000000
0!
0'
0/
#591150000000
1!
1'
1/
#591160000000
0!
0'
0/
#591170000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#591180000000
0!
0'
0/
#591190000000
1!
1'
1/
#591200000000
0!
0'
0/
#591210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#591220000000
0!
0'
0/
#591230000000
1!
1'
1/
#591240000000
0!
0'
0/
#591250000000
#591260000000
1!
1'
1/
#591270000000
0!
0'
0/
#591280000000
1!
1'
1/
#591290000000
0!
1"
0'
1(
0/
10
#591300000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#591310000000
0!
0'
0/
#591320000000
1!
1'
1/
#591330000000
0!
0'
0/
#591340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#591350000000
0!
0'
0/
#591360000000
1!
1'
1/
#591370000000
0!
1"
0'
1(
0/
10
#591380000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#591390000000
0!
1$
0'
1+
0/
#591400000000
1!
1'
1/
#591410000000
0!
0'
0/
#591420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#591430000000
0!
0'
0/
#591440000000
1!
1'
1/
#591450000000
0!
0'
0/
#591460000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#591470000000
0!
0'
0/
#591480000000
1!
1'
1/
#591490000000
0!
0'
0/
#591500000000
1!
1'
1/
#591510000000
0!
0'
0/
#591520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#591530000000
0!
0'
0/
#591540000000
1!
1'
1/
#591550000000
0!
0'
0/
#591560000000
1!
1'
1/
#591570000000
0!
0'
0/
#591580000000
1!
1'
1/
#591590000000
0!
0'
0/
#591600000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#591610000000
0!
0'
0/
#591620000000
1!
1'
1/
#591630000000
0!
0'
0/
#591640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#591650000000
0!
0'
0/
#591660000000
1!
1'
1/
#591670000000
0!
0'
0/
#591680000000
#591690000000
1!
1'
1/
#591700000000
0!
0'
0/
#591710000000
1!
1'
1/
#591720000000
0!
1"
0'
1(
0/
10
#591730000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#591740000000
0!
0'
0/
#591750000000
1!
1'
1/
#591760000000
0!
0'
0/
#591770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#591780000000
0!
0'
0/
#591790000000
1!
1'
1/
#591800000000
0!
1"
0'
1(
0/
10
#591810000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#591820000000
0!
1$
0'
1+
0/
#591830000000
1!
1'
1/
#591840000000
0!
0'
0/
#591850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#591860000000
0!
0'
0/
#591870000000
1!
1'
1/
#591880000000
0!
0'
0/
#591890000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#591900000000
0!
0'
0/
#591910000000
1!
1'
1/
#591920000000
0!
0'
0/
#591930000000
1!
1'
1/
#591940000000
0!
0'
0/
#591950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#591960000000
0!
0'
0/
#591970000000
1!
1'
1/
#591980000000
0!
0'
0/
#591990000000
1!
1'
1/
#592000000000
0!
0'
0/
#592010000000
1!
1'
1/
#592020000000
0!
0'
0/
#592030000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#592040000000
0!
0'
0/
#592050000000
1!
1'
1/
#592060000000
0!
0'
0/
#592070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#592080000000
0!
0'
0/
#592090000000
1!
1'
1/
#592100000000
0!
0'
0/
#592110000000
#592120000000
1!
1'
1/
#592130000000
0!
0'
0/
#592140000000
1!
1'
1/
#592150000000
0!
1"
0'
1(
0/
10
#592160000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#592170000000
0!
0'
0/
#592180000000
1!
1'
1/
#592190000000
0!
0'
0/
#592200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#592210000000
0!
0'
0/
#592220000000
1!
1'
1/
#592230000000
0!
1"
0'
1(
0/
10
#592240000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#592250000000
0!
1$
0'
1+
0/
#592260000000
1!
1'
1/
#592270000000
0!
0'
0/
#592280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#592290000000
0!
0'
0/
#592300000000
1!
1'
1/
#592310000000
0!
0'
0/
#592320000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#592330000000
0!
0'
0/
#592340000000
1!
1'
1/
#592350000000
0!
0'
0/
#592360000000
1!
1'
1/
#592370000000
0!
0'
0/
#592380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#592390000000
0!
0'
0/
#592400000000
1!
1'
1/
#592410000000
0!
0'
0/
#592420000000
1!
1'
1/
#592430000000
0!
0'
0/
#592440000000
1!
1'
1/
#592450000000
0!
0'
0/
#592460000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#592470000000
0!
0'
0/
#592480000000
1!
1'
1/
#592490000000
0!
0'
0/
#592500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#592510000000
0!
0'
0/
#592520000000
1!
1'
1/
#592530000000
0!
0'
0/
#592540000000
#592550000000
1!
1'
1/
#592560000000
0!
0'
0/
#592570000000
1!
1'
1/
#592580000000
0!
1"
0'
1(
0/
10
#592590000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#592600000000
0!
0'
0/
#592610000000
1!
1'
1/
#592620000000
0!
0'
0/
#592630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#592640000000
0!
0'
0/
#592650000000
1!
1'
1/
#592660000000
0!
1"
0'
1(
0/
10
#592670000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#592680000000
0!
1$
0'
1+
0/
#592690000000
1!
1'
1/
#592700000000
0!
0'
0/
#592710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#592720000000
0!
0'
0/
#592730000000
1!
1'
1/
#592740000000
0!
0'
0/
#592750000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#592760000000
0!
0'
0/
#592770000000
1!
1'
1/
#592780000000
0!
0'
0/
#592790000000
1!
1'
1/
#592800000000
0!
0'
0/
#592810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#592820000000
0!
0'
0/
#592830000000
1!
1'
1/
#592840000000
0!
0'
0/
#592850000000
1!
1'
1/
#592860000000
0!
0'
0/
#592870000000
1!
1'
1/
#592880000000
0!
0'
0/
#592890000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#592900000000
0!
0'
0/
#592910000000
1!
1'
1/
#592920000000
0!
0'
0/
#592930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#592940000000
0!
0'
0/
#592950000000
1!
1'
1/
#592960000000
0!
0'
0/
#592970000000
#592980000000
1!
1'
1/
#592990000000
0!
0'
0/
#593000000000
1!
1'
1/
#593010000000
0!
1"
0'
1(
0/
10
#593020000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#593030000000
0!
0'
0/
#593040000000
1!
1'
1/
#593050000000
0!
0'
0/
#593060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#593070000000
0!
0'
0/
#593080000000
1!
1'
1/
#593090000000
0!
1"
0'
1(
0/
10
#593100000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#593110000000
0!
1$
0'
1+
0/
#593120000000
1!
1'
1/
#593130000000
0!
0'
0/
#593140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#593150000000
0!
0'
0/
#593160000000
1!
1'
1/
#593170000000
0!
0'
0/
#593180000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#593190000000
0!
0'
0/
#593200000000
1!
1'
1/
#593210000000
0!
0'
0/
#593220000000
1!
1'
1/
#593230000000
0!
0'
0/
#593240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#593250000000
0!
0'
0/
#593260000000
1!
1'
1/
#593270000000
0!
0'
0/
#593280000000
1!
1'
1/
#593290000000
0!
0'
0/
#593300000000
1!
1'
1/
#593310000000
0!
0'
0/
#593320000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#593330000000
0!
0'
0/
#593340000000
1!
1'
1/
#593350000000
0!
0'
0/
#593360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#593370000000
0!
0'
0/
#593380000000
1!
1'
1/
#593390000000
0!
0'
0/
#593400000000
#593410000000
1!
1'
1/
#593420000000
0!
0'
0/
#593430000000
1!
1'
1/
#593440000000
0!
1"
0'
1(
0/
10
#593450000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#593460000000
0!
0'
0/
#593470000000
1!
1'
1/
#593480000000
0!
0'
0/
#593490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#593500000000
0!
0'
0/
#593510000000
1!
1'
1/
#593520000000
0!
1"
0'
1(
0/
10
#593530000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#593540000000
0!
1$
0'
1+
0/
#593550000000
1!
1'
1/
#593560000000
0!
0'
0/
#593570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#593580000000
0!
0'
0/
#593590000000
1!
1'
1/
#593600000000
0!
0'
0/
#593610000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#593620000000
0!
0'
0/
#593630000000
1!
1'
1/
#593640000000
0!
0'
0/
#593650000000
1!
1'
1/
#593660000000
0!
0'
0/
#593670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#593680000000
0!
0'
0/
#593690000000
1!
1'
1/
#593700000000
0!
0'
0/
#593710000000
1!
1'
1/
#593720000000
0!
0'
0/
#593730000000
1!
1'
1/
#593740000000
0!
0'
0/
#593750000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#593760000000
0!
0'
0/
#593770000000
1!
1'
1/
#593780000000
0!
0'
0/
#593790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#593800000000
0!
0'
0/
#593810000000
1!
1'
1/
#593820000000
0!
0'
0/
#593830000000
#593840000000
1!
1'
1/
#593850000000
0!
0'
0/
#593860000000
1!
1'
1/
#593870000000
0!
1"
0'
1(
0/
10
#593880000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#593890000000
0!
0'
0/
#593900000000
1!
1'
1/
#593910000000
0!
0'
0/
#593920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#593930000000
0!
0'
0/
#593940000000
1!
1'
1/
#593950000000
0!
1"
0'
1(
0/
10
#593960000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#593970000000
0!
1$
0'
1+
0/
#593980000000
1!
1'
1/
#593990000000
0!
0'
0/
#594000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#594010000000
0!
0'
0/
#594020000000
1!
1'
1/
#594030000000
0!
0'
0/
#594040000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#594050000000
0!
0'
0/
#594060000000
1!
1'
1/
#594070000000
0!
0'
0/
#594080000000
1!
1'
1/
#594090000000
0!
0'
0/
#594100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#594110000000
0!
0'
0/
#594120000000
1!
1'
1/
#594130000000
0!
0'
0/
#594140000000
1!
1'
1/
#594150000000
0!
0'
0/
#594160000000
1!
1'
1/
#594170000000
0!
0'
0/
#594180000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#594190000000
0!
0'
0/
#594200000000
1!
1'
1/
#594210000000
0!
0'
0/
#594220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#594230000000
0!
0'
0/
#594240000000
1!
1'
1/
#594250000000
0!
0'
0/
#594260000000
#594270000000
1!
1'
1/
#594280000000
0!
0'
0/
#594290000000
1!
1'
1/
#594300000000
0!
1"
0'
1(
0/
10
#594310000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#594320000000
0!
0'
0/
#594330000000
1!
1'
1/
#594340000000
0!
0'
0/
#594350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#594360000000
0!
0'
0/
#594370000000
1!
1'
1/
#594380000000
0!
1"
0'
1(
0/
10
#594390000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#594400000000
0!
1$
0'
1+
0/
#594410000000
1!
1'
1/
#594420000000
0!
0'
0/
#594430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#594440000000
0!
0'
0/
#594450000000
1!
1'
1/
#594460000000
0!
0'
0/
#594470000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#594480000000
0!
0'
0/
#594490000000
1!
1'
1/
#594500000000
0!
0'
0/
#594510000000
1!
1'
1/
#594520000000
0!
0'
0/
#594530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#594540000000
0!
0'
0/
#594550000000
1!
1'
1/
#594560000000
0!
0'
0/
#594570000000
1!
1'
1/
#594580000000
0!
0'
0/
#594590000000
1!
1'
1/
#594600000000
0!
0'
0/
#594610000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#594620000000
0!
0'
0/
#594630000000
1!
1'
1/
#594640000000
0!
0'
0/
#594650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#594660000000
0!
0'
0/
#594670000000
1!
1'
1/
#594680000000
0!
0'
0/
#594690000000
#594700000000
1!
1'
1/
#594710000000
0!
0'
0/
#594720000000
1!
1'
1/
#594730000000
0!
1"
0'
1(
0/
10
#594740000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#594750000000
0!
0'
0/
#594760000000
1!
1'
1/
#594770000000
0!
0'
0/
#594780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#594790000000
0!
0'
0/
#594800000000
1!
1'
1/
#594810000000
0!
1"
0'
1(
0/
10
#594820000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#594830000000
0!
1$
0'
1+
0/
#594840000000
1!
1'
1/
#594850000000
0!
0'
0/
#594860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#594870000000
0!
0'
0/
#594880000000
1!
1'
1/
#594890000000
0!
0'
0/
#594900000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#594910000000
0!
0'
0/
#594920000000
1!
1'
1/
#594930000000
0!
0'
0/
#594940000000
1!
1'
1/
#594950000000
0!
0'
0/
#594960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#594970000000
0!
0'
0/
#594980000000
1!
1'
1/
#594990000000
0!
0'
0/
#595000000000
1!
1'
1/
#595010000000
0!
0'
0/
#595020000000
1!
1'
1/
#595030000000
0!
0'
0/
#595040000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#595050000000
0!
0'
0/
#595060000000
1!
1'
1/
#595070000000
0!
0'
0/
#595080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#595090000000
0!
0'
0/
#595100000000
1!
1'
1/
#595110000000
0!
0'
0/
#595120000000
#595130000000
1!
1'
1/
#595140000000
0!
0'
0/
#595150000000
1!
1'
1/
#595160000000
0!
1"
0'
1(
0/
10
#595170000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#595180000000
0!
0'
0/
#595190000000
1!
1'
1/
#595200000000
0!
0'
0/
#595210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#595220000000
0!
0'
0/
#595230000000
1!
1'
1/
#595240000000
0!
1"
0'
1(
0/
10
#595250000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#595260000000
0!
1$
0'
1+
0/
#595270000000
1!
1'
1/
#595280000000
0!
0'
0/
#595290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#595300000000
0!
0'
0/
#595310000000
1!
1'
1/
#595320000000
0!
0'
0/
#595330000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#595340000000
0!
0'
0/
#595350000000
1!
1'
1/
#595360000000
0!
0'
0/
#595370000000
1!
1'
1/
#595380000000
0!
0'
0/
#595390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#595400000000
0!
0'
0/
#595410000000
1!
1'
1/
#595420000000
0!
0'
0/
#595430000000
1!
1'
1/
#595440000000
0!
0'
0/
#595450000000
1!
1'
1/
#595460000000
0!
0'
0/
#595470000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#595480000000
0!
0'
0/
#595490000000
1!
1'
1/
#595500000000
0!
0'
0/
#595510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#595520000000
0!
0'
0/
#595530000000
1!
1'
1/
#595540000000
0!
0'
0/
#595550000000
#595560000000
1!
1'
1/
#595570000000
0!
0'
0/
#595580000000
1!
1'
1/
#595590000000
0!
1"
0'
1(
0/
10
#595600000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#595610000000
0!
0'
0/
#595620000000
1!
1'
1/
#595630000000
0!
0'
0/
#595640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#595650000000
0!
0'
0/
#595660000000
1!
1'
1/
#595670000000
0!
1"
0'
1(
0/
10
#595680000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#595690000000
0!
1$
0'
1+
0/
#595700000000
1!
1'
1/
#595710000000
0!
0'
0/
#595720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#595730000000
0!
0'
0/
#595740000000
1!
1'
1/
#595750000000
0!
0'
0/
#595760000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#595770000000
0!
0'
0/
#595780000000
1!
1'
1/
#595790000000
0!
0'
0/
#595800000000
1!
1'
1/
#595810000000
0!
0'
0/
#595820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#595830000000
0!
0'
0/
#595840000000
1!
1'
1/
#595850000000
0!
0'
0/
#595860000000
1!
1'
1/
#595870000000
0!
0'
0/
#595880000000
1!
1'
1/
#595890000000
0!
0'
0/
#595900000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#595910000000
0!
0'
0/
#595920000000
1!
1'
1/
#595930000000
0!
0'
0/
#595940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#595950000000
0!
0'
0/
#595960000000
1!
1'
1/
#595970000000
0!
0'
0/
#595980000000
#595990000000
1!
1'
1/
#596000000000
0!
0'
0/
#596010000000
1!
1'
1/
#596020000000
0!
1"
0'
1(
0/
10
#596030000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#596040000000
0!
0'
0/
#596050000000
1!
1'
1/
#596060000000
0!
0'
0/
#596070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#596080000000
0!
0'
0/
#596090000000
1!
1'
1/
#596100000000
0!
1"
0'
1(
0/
10
#596110000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#596120000000
0!
1$
0'
1+
0/
#596130000000
1!
1'
1/
#596140000000
0!
0'
0/
#596150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#596160000000
0!
0'
0/
#596170000000
1!
1'
1/
#596180000000
0!
0'
0/
#596190000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#596200000000
0!
0'
0/
#596210000000
1!
1'
1/
#596220000000
0!
0'
0/
#596230000000
1!
1'
1/
#596240000000
0!
0'
0/
#596250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#596260000000
0!
0'
0/
#596270000000
1!
1'
1/
#596280000000
0!
0'
0/
#596290000000
1!
1'
1/
#596300000000
0!
0'
0/
#596310000000
1!
1'
1/
#596320000000
0!
0'
0/
#596330000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#596340000000
0!
0'
0/
#596350000000
1!
1'
1/
#596360000000
0!
0'
0/
#596370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#596380000000
0!
0'
0/
#596390000000
1!
1'
1/
#596400000000
0!
0'
0/
#596410000000
#596420000000
1!
1'
1/
#596430000000
0!
0'
0/
#596440000000
1!
1'
1/
#596450000000
0!
1"
0'
1(
0/
10
#596460000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#596470000000
0!
0'
0/
#596480000000
1!
1'
1/
#596490000000
0!
0'
0/
#596500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#596510000000
0!
0'
0/
#596520000000
1!
1'
1/
#596530000000
0!
1"
0'
1(
0/
10
#596540000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#596550000000
0!
1$
0'
1+
0/
#596560000000
1!
1'
1/
#596570000000
0!
0'
0/
#596580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#596590000000
0!
0'
0/
#596600000000
1!
1'
1/
#596610000000
0!
0'
0/
#596620000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#596630000000
0!
0'
0/
#596640000000
1!
1'
1/
#596650000000
0!
0'
0/
#596660000000
1!
1'
1/
#596670000000
0!
0'
0/
#596680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#596690000000
0!
0'
0/
#596700000000
1!
1'
1/
#596710000000
0!
0'
0/
#596720000000
1!
1'
1/
#596730000000
0!
0'
0/
#596740000000
1!
1'
1/
#596750000000
0!
0'
0/
#596760000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#596770000000
0!
0'
0/
#596780000000
1!
1'
1/
#596790000000
0!
0'
0/
#596800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#596810000000
0!
0'
0/
#596820000000
1!
1'
1/
#596830000000
0!
0'
0/
#596840000000
#596850000000
1!
1'
1/
#596860000000
0!
0'
0/
#596870000000
1!
1'
1/
#596880000000
0!
1"
0'
1(
0/
10
#596890000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#596900000000
0!
0'
0/
#596910000000
1!
1'
1/
#596920000000
0!
0'
0/
#596930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#596940000000
0!
0'
0/
#596950000000
1!
1'
1/
#596960000000
0!
1"
0'
1(
0/
10
#596970000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#596980000000
0!
1$
0'
1+
0/
#596990000000
1!
1'
1/
#597000000000
0!
0'
0/
#597010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#597020000000
0!
0'
0/
#597030000000
1!
1'
1/
#597040000000
0!
0'
0/
#597050000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#597060000000
0!
0'
0/
#597070000000
1!
1'
1/
#597080000000
0!
0'
0/
#597090000000
1!
1'
1/
#597100000000
0!
0'
0/
#597110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#597120000000
0!
0'
0/
#597130000000
1!
1'
1/
#597140000000
0!
0'
0/
#597150000000
1!
1'
1/
#597160000000
0!
0'
0/
#597170000000
1!
1'
1/
#597180000000
0!
0'
0/
#597190000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#597200000000
0!
0'
0/
#597210000000
1!
1'
1/
#597220000000
0!
0'
0/
#597230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#597240000000
0!
0'
0/
#597250000000
1!
1'
1/
#597260000000
0!
0'
0/
#597270000000
#597280000000
1!
1'
1/
#597290000000
0!
0'
0/
#597300000000
1!
1'
1/
#597310000000
0!
1"
0'
1(
0/
10
#597320000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#597330000000
0!
0'
0/
#597340000000
1!
1'
1/
#597350000000
0!
0'
0/
#597360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#597370000000
0!
0'
0/
#597380000000
1!
1'
1/
#597390000000
0!
1"
0'
1(
0/
10
#597400000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#597410000000
0!
1$
0'
1+
0/
#597420000000
1!
1'
1/
#597430000000
0!
0'
0/
#597440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#597450000000
0!
0'
0/
#597460000000
1!
1'
1/
#597470000000
0!
0'
0/
#597480000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#597490000000
0!
0'
0/
#597500000000
1!
1'
1/
#597510000000
0!
0'
0/
#597520000000
1!
1'
1/
#597530000000
0!
0'
0/
#597540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#597550000000
0!
0'
0/
#597560000000
1!
1'
1/
#597570000000
0!
0'
0/
#597580000000
1!
1'
1/
#597590000000
0!
0'
0/
#597600000000
1!
1'
1/
#597610000000
0!
0'
0/
#597620000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#597630000000
0!
0'
0/
#597640000000
1!
1'
1/
#597650000000
0!
0'
0/
#597660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#597670000000
0!
0'
0/
#597680000000
1!
1'
1/
#597690000000
0!
0'
0/
#597700000000
#597710000000
1!
1'
1/
#597720000000
0!
0'
0/
#597730000000
1!
1'
1/
#597740000000
0!
1"
0'
1(
0/
10
#597750000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#597760000000
0!
0'
0/
#597770000000
1!
1'
1/
#597780000000
0!
0'
0/
#597790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#597800000000
0!
0'
0/
#597810000000
1!
1'
1/
#597820000000
0!
1"
0'
1(
0/
10
#597830000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#597840000000
0!
1$
0'
1+
0/
#597850000000
1!
1'
1/
#597860000000
0!
0'
0/
#597870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#597880000000
0!
0'
0/
#597890000000
1!
1'
1/
#597900000000
0!
0'
0/
#597910000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#597920000000
0!
0'
0/
#597930000000
1!
1'
1/
#597940000000
0!
0'
0/
#597950000000
1!
1'
1/
#597960000000
0!
0'
0/
#597970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#597980000000
0!
0'
0/
#597990000000
1!
1'
1/
#598000000000
0!
0'
0/
#598010000000
1!
1'
1/
#598020000000
0!
0'
0/
#598030000000
1!
1'
1/
#598040000000
0!
0'
0/
#598050000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#598060000000
0!
0'
0/
#598070000000
1!
1'
1/
#598080000000
0!
0'
0/
#598090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#598100000000
0!
0'
0/
#598110000000
1!
1'
1/
#598120000000
0!
0'
0/
#598130000000
#598140000000
1!
1'
1/
#598150000000
0!
0'
0/
#598160000000
1!
1'
1/
#598170000000
0!
1"
0'
1(
0/
10
#598180000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#598190000000
0!
0'
0/
#598200000000
1!
1'
1/
#598210000000
0!
0'
0/
#598220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#598230000000
0!
0'
0/
#598240000000
1!
1'
1/
#598250000000
0!
1"
0'
1(
0/
10
#598260000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#598270000000
0!
1$
0'
1+
0/
#598280000000
1!
1'
1/
#598290000000
0!
0'
0/
#598300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#598310000000
0!
0'
0/
#598320000000
1!
1'
1/
#598330000000
0!
0'
0/
#598340000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#598350000000
0!
0'
0/
#598360000000
1!
1'
1/
#598370000000
0!
0'
0/
#598380000000
1!
1'
1/
#598390000000
0!
0'
0/
#598400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#598410000000
0!
0'
0/
#598420000000
1!
1'
1/
#598430000000
0!
0'
0/
#598440000000
1!
1'
1/
#598450000000
0!
0'
0/
#598460000000
1!
1'
1/
#598470000000
0!
0'
0/
#598480000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#598490000000
0!
0'
0/
#598500000000
1!
1'
1/
#598510000000
0!
0'
0/
#598520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#598530000000
0!
0'
0/
#598540000000
1!
1'
1/
#598550000000
0!
0'
0/
#598560000000
#598570000000
1!
1'
1/
#598580000000
0!
0'
0/
#598590000000
1!
1'
1/
#598600000000
0!
1"
0'
1(
0/
10
#598610000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#598620000000
0!
0'
0/
#598630000000
1!
1'
1/
#598640000000
0!
0'
0/
#598650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#598660000000
0!
0'
0/
#598670000000
1!
1'
1/
#598680000000
0!
1"
0'
1(
0/
10
#598690000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#598700000000
0!
1$
0'
1+
0/
#598710000000
1!
1'
1/
#598720000000
0!
0'
0/
#598730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#598740000000
0!
0'
0/
#598750000000
1!
1'
1/
#598760000000
0!
0'
0/
#598770000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#598780000000
0!
0'
0/
#598790000000
1!
1'
1/
#598800000000
0!
0'
0/
#598810000000
1!
1'
1/
#598820000000
0!
0'
0/
#598830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#598840000000
0!
0'
0/
#598850000000
1!
1'
1/
#598860000000
0!
0'
0/
#598870000000
1!
1'
1/
#598880000000
0!
0'
0/
#598890000000
1!
1'
1/
#598900000000
0!
0'
0/
#598910000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#598920000000
0!
0'
0/
#598930000000
1!
1'
1/
#598940000000
0!
0'
0/
#598950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#598960000000
0!
0'
0/
#598970000000
1!
1'
1/
#598980000000
0!
0'
0/
#598990000000
#599000000000
1!
1'
1/
#599010000000
0!
0'
0/
#599020000000
1!
1'
1/
#599030000000
0!
1"
0'
1(
0/
10
#599040000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#599050000000
0!
0'
0/
#599060000000
1!
1'
1/
#599070000000
0!
0'
0/
#599080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#599090000000
0!
0'
0/
#599100000000
1!
1'
1/
#599110000000
0!
1"
0'
1(
0/
10
#599120000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#599130000000
0!
1$
0'
1+
0/
#599140000000
1!
1'
1/
#599150000000
0!
0'
0/
#599160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#599170000000
0!
0'
0/
#599180000000
1!
1'
1/
#599190000000
0!
0'
0/
#599200000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#599210000000
0!
0'
0/
#599220000000
1!
1'
1/
#599230000000
0!
0'
0/
#599240000000
1!
1'
1/
#599250000000
0!
0'
0/
#599260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#599270000000
0!
0'
0/
#599280000000
1!
1'
1/
#599290000000
0!
0'
0/
#599300000000
1!
1'
1/
#599310000000
0!
0'
0/
#599320000000
1!
1'
1/
#599330000000
0!
0'
0/
#599340000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#599350000000
0!
0'
0/
#599360000000
1!
1'
1/
#599370000000
0!
0'
0/
#599380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#599390000000
0!
0'
0/
#599400000000
1!
1'
1/
#599410000000
0!
0'
0/
#599420000000
#599430000000
1!
1'
1/
#599440000000
0!
0'
0/
#599450000000
1!
1'
1/
#599460000000
0!
1"
0'
1(
0/
10
#599470000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#599480000000
0!
0'
0/
#599490000000
1!
1'
1/
#599500000000
0!
0'
0/
#599510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#599520000000
0!
0'
0/
#599530000000
1!
1'
1/
#599540000000
0!
1"
0'
1(
0/
10
#599550000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#599560000000
0!
1$
0'
1+
0/
#599570000000
1!
1'
1/
#599580000000
0!
0'
0/
#599590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#599600000000
0!
0'
0/
#599610000000
1!
1'
1/
#599620000000
0!
0'
0/
#599630000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#599640000000
0!
0'
0/
#599650000000
1!
1'
1/
#599660000000
0!
0'
0/
#599670000000
1!
1'
1/
#599680000000
0!
0'
0/
#599690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#599700000000
0!
0'
0/
#599710000000
1!
1'
1/
#599720000000
0!
0'
0/
#599730000000
1!
1'
1/
#599740000000
0!
0'
0/
#599750000000
1!
1'
1/
#599760000000
0!
0'
0/
#599770000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#599780000000
0!
0'
0/
#599790000000
1!
1'
1/
#599800000000
0!
0'
0/
#599810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#599820000000
0!
0'
0/
#599830000000
1!
1'
1/
#599840000000
0!
0'
0/
#599850000000
#599860000000
1!
1'
1/
#599870000000
0!
0'
0/
#599880000000
1!
1'
1/
#599890000000
0!
1"
0'
1(
0/
10
#599900000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#599910000000
0!
0'
0/
#599920000000
1!
1'
1/
#599930000000
0!
0'
0/
#599940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#599950000000
0!
0'
0/
#599960000000
1!
1'
1/
#599970000000
0!
1"
0'
1(
0/
10
#599980000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#599990000000
0!
1$
0'
1+
0/
#600000000000
1!
1'
1/
#600010000000
0!
0'
0/
#600020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#600030000000
0!
0'
0/
#600040000000
1!
1'
1/
#600050000000
0!
0'
0/
#600060000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#600070000000
0!
0'
0/
#600080000000
1!
1'
1/
#600090000000
0!
0'
0/
#600100000000
1!
1'
1/
#600110000000
0!
0'
0/
#600120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#600130000000
0!
0'
0/
#600140000000
1!
1'
1/
#600150000000
0!
0'
0/
#600160000000
1!
1'
1/
#600170000000
0!
0'
0/
#600180000000
1!
1'
1/
#600190000000
0!
0'
0/
#600200000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#600210000000
0!
0'
0/
#600220000000
1!
1'
1/
#600230000000
0!
0'
0/
#600240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#600250000000
0!
0'
0/
#600260000000
1!
1'
1/
#600270000000
0!
0'
0/
#600280000000
#600290000000
1!
1'
1/
#600300000000
0!
0'
0/
#600310000000
1!
1'
1/
#600320000000
0!
1"
0'
1(
0/
10
#600330000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#600340000000
0!
0'
0/
#600350000000
1!
1'
1/
#600360000000
0!
0'
0/
#600370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#600380000000
0!
0'
0/
#600390000000
1!
1'
1/
#600400000000
0!
1"
0'
1(
0/
10
#600410000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#600420000000
0!
1$
0'
1+
0/
#600430000000
1!
1'
1/
#600440000000
0!
0'
0/
#600450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#600460000000
0!
0'
0/
#600470000000
1!
1'
1/
#600480000000
0!
0'
0/
#600490000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#600500000000
0!
0'
0/
#600510000000
1!
1'
1/
#600520000000
0!
0'
0/
#600530000000
1!
1'
1/
#600540000000
0!
0'
0/
#600550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#600560000000
0!
0'
0/
#600570000000
1!
1'
1/
#600580000000
0!
0'
0/
#600590000000
1!
1'
1/
#600600000000
0!
0'
0/
#600610000000
1!
1'
1/
#600620000000
0!
0'
0/
#600630000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#600640000000
0!
0'
0/
#600650000000
1!
1'
1/
#600660000000
0!
0'
0/
#600670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#600680000000
0!
0'
0/
#600690000000
1!
1'
1/
#600700000000
0!
0'
0/
#600710000000
#600720000000
1!
1'
1/
#600730000000
0!
0'
0/
#600740000000
1!
1'
1/
#600750000000
0!
1"
0'
1(
0/
10
#600760000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#600770000000
0!
0'
0/
#600780000000
1!
1'
1/
#600790000000
0!
0'
0/
#600800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#600810000000
0!
0'
0/
#600820000000
1!
1'
1/
#600830000000
0!
1"
0'
1(
0/
10
#600840000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#600850000000
0!
1$
0'
1+
0/
#600860000000
1!
1'
1/
#600870000000
0!
0'
0/
#600880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#600890000000
0!
0'
0/
#600900000000
1!
1'
1/
#600910000000
0!
0'
0/
#600920000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#600930000000
0!
0'
0/
#600940000000
1!
1'
1/
#600950000000
0!
0'
0/
#600960000000
1!
1'
1/
#600970000000
0!
0'
0/
#600980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#600990000000
0!
0'
0/
#601000000000
1!
1'
1/
#601010000000
0!
0'
0/
#601020000000
1!
1'
1/
#601030000000
0!
0'
0/
#601040000000
1!
1'
1/
#601050000000
0!
0'
0/
#601060000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#601070000000
0!
0'
0/
#601080000000
1!
1'
1/
#601090000000
0!
0'
0/
#601100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#601110000000
0!
0'
0/
#601120000000
1!
1'
1/
#601130000000
0!
0'
0/
#601140000000
#601150000000
1!
1'
1/
#601160000000
0!
0'
0/
#601170000000
1!
1'
1/
#601180000000
0!
1"
0'
1(
0/
10
#601190000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#601200000000
0!
0'
0/
#601210000000
1!
1'
1/
#601220000000
0!
0'
0/
#601230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#601240000000
0!
0'
0/
#601250000000
1!
1'
1/
#601260000000
0!
1"
0'
1(
0/
10
#601270000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#601280000000
0!
1$
0'
1+
0/
#601290000000
1!
1'
1/
#601300000000
0!
0'
0/
#601310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#601320000000
0!
0'
0/
#601330000000
1!
1'
1/
#601340000000
0!
0'
0/
#601350000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#601360000000
0!
0'
0/
#601370000000
1!
1'
1/
#601380000000
0!
0'
0/
#601390000000
1!
1'
1/
#601400000000
0!
0'
0/
#601410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#601420000000
0!
0'
0/
#601430000000
1!
1'
1/
#601440000000
0!
0'
0/
#601450000000
1!
1'
1/
#601460000000
0!
0'
0/
#601470000000
1!
1'
1/
#601480000000
0!
0'
0/
#601490000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#601500000000
0!
0'
0/
#601510000000
1!
1'
1/
#601520000000
0!
0'
0/
#601530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#601540000000
0!
0'
0/
#601550000000
1!
1'
1/
#601560000000
0!
0'
0/
#601570000000
#601580000000
1!
1'
1/
#601590000000
0!
0'
0/
#601600000000
1!
1'
1/
#601610000000
0!
1"
0'
1(
0/
10
#601620000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#601630000000
0!
0'
0/
#601640000000
1!
1'
1/
#601650000000
0!
0'
0/
#601660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#601670000000
0!
0'
0/
#601680000000
1!
1'
1/
#601690000000
0!
1"
0'
1(
0/
10
#601700000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#601710000000
0!
1$
0'
1+
0/
#601720000000
1!
1'
1/
#601730000000
0!
0'
0/
#601740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#601750000000
0!
0'
0/
#601760000000
1!
1'
1/
#601770000000
0!
0'
0/
#601780000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#601790000000
0!
0'
0/
#601800000000
1!
1'
1/
#601810000000
0!
0'
0/
#601820000000
1!
1'
1/
#601830000000
0!
0'
0/
#601840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#601850000000
0!
0'
0/
#601860000000
1!
1'
1/
#601870000000
0!
0'
0/
#601880000000
1!
1'
1/
#601890000000
0!
0'
0/
#601900000000
1!
1'
1/
#601910000000
0!
0'
0/
#601920000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#601930000000
0!
0'
0/
#601940000000
1!
1'
1/
#601950000000
0!
0'
0/
#601960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#601970000000
0!
0'
0/
#601980000000
1!
1'
1/
#601990000000
0!
0'
0/
#602000000000
#602010000000
1!
1'
1/
#602020000000
0!
0'
0/
#602030000000
1!
1'
1/
#602040000000
0!
1"
0'
1(
0/
10
#602050000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#602060000000
0!
0'
0/
#602070000000
1!
1'
1/
#602080000000
0!
0'
0/
#602090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#602100000000
0!
0'
0/
#602110000000
1!
1'
1/
#602120000000
0!
1"
0'
1(
0/
10
#602130000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#602140000000
0!
1$
0'
1+
0/
#602150000000
1!
1'
1/
#602160000000
0!
0'
0/
#602170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#602180000000
0!
0'
0/
#602190000000
1!
1'
1/
#602200000000
0!
0'
0/
#602210000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#602220000000
0!
0'
0/
#602230000000
1!
1'
1/
#602240000000
0!
0'
0/
#602250000000
1!
1'
1/
#602260000000
0!
0'
0/
#602270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#602280000000
0!
0'
0/
#602290000000
1!
1'
1/
#602300000000
0!
0'
0/
#602310000000
1!
1'
1/
#602320000000
0!
0'
0/
#602330000000
1!
1'
1/
#602340000000
0!
0'
0/
#602350000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#602360000000
0!
0'
0/
#602370000000
1!
1'
1/
#602380000000
0!
0'
0/
#602390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#602400000000
0!
0'
0/
#602410000000
1!
1'
1/
#602420000000
0!
0'
0/
#602430000000
#602440000000
1!
1'
1/
#602450000000
0!
0'
0/
#602460000000
1!
1'
1/
#602470000000
0!
1"
0'
1(
0/
10
#602480000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#602490000000
0!
0'
0/
#602500000000
1!
1'
1/
#602510000000
0!
0'
0/
#602520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#602530000000
0!
0'
0/
#602540000000
1!
1'
1/
#602550000000
0!
1"
0'
1(
0/
10
#602560000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#602570000000
0!
1$
0'
1+
0/
#602580000000
1!
1'
1/
#602590000000
0!
0'
0/
#602600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#602610000000
0!
0'
0/
#602620000000
1!
1'
1/
#602630000000
0!
0'
0/
#602640000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#602650000000
0!
0'
0/
#602660000000
1!
1'
1/
#602670000000
0!
0'
0/
#602680000000
1!
1'
1/
#602690000000
0!
0'
0/
#602700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#602710000000
0!
0'
0/
#602720000000
1!
1'
1/
#602730000000
0!
0'
0/
#602740000000
1!
1'
1/
#602750000000
0!
0'
0/
#602760000000
1!
1'
1/
#602770000000
0!
0'
0/
#602780000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#602790000000
0!
0'
0/
#602800000000
1!
1'
1/
#602810000000
0!
0'
0/
#602820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#602830000000
0!
0'
0/
#602840000000
1!
1'
1/
#602850000000
0!
0'
0/
#602860000000
#602870000000
1!
1'
1/
#602880000000
0!
0'
0/
#602890000000
1!
1'
1/
#602900000000
0!
1"
0'
1(
0/
10
#602910000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#602920000000
0!
0'
0/
#602930000000
1!
1'
1/
#602940000000
0!
0'
0/
#602950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#602960000000
0!
0'
0/
#602970000000
1!
1'
1/
#602980000000
0!
1"
0'
1(
0/
10
#602990000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#603000000000
0!
1$
0'
1+
0/
#603010000000
1!
1'
1/
#603020000000
0!
0'
0/
#603030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#603040000000
0!
0'
0/
#603050000000
1!
1'
1/
#603060000000
0!
0'
0/
#603070000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#603080000000
0!
0'
0/
#603090000000
1!
1'
1/
#603100000000
0!
0'
0/
#603110000000
1!
1'
1/
#603120000000
0!
0'
0/
#603130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#603140000000
0!
0'
0/
#603150000000
1!
1'
1/
#603160000000
0!
0'
0/
#603170000000
1!
1'
1/
#603180000000
0!
0'
0/
#603190000000
1!
1'
1/
#603200000000
0!
0'
0/
#603210000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#603220000000
0!
0'
0/
#603230000000
1!
1'
1/
#603240000000
0!
0'
0/
#603250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#603260000000
0!
0'
0/
#603270000000
1!
1'
1/
#603280000000
0!
0'
0/
#603290000000
#603300000000
1!
1'
1/
#603310000000
0!
0'
0/
#603320000000
1!
1'
1/
#603330000000
0!
1"
0'
1(
0/
10
#603340000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#603350000000
0!
0'
0/
#603360000000
1!
1'
1/
#603370000000
0!
0'
0/
#603380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#603390000000
0!
0'
0/
#603400000000
1!
1'
1/
#603410000000
0!
1"
0'
1(
0/
10
#603420000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#603430000000
0!
1$
0'
1+
0/
#603440000000
1!
1'
1/
#603450000000
0!
0'
0/
#603460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#603470000000
0!
0'
0/
#603480000000
1!
1'
1/
#603490000000
0!
0'
0/
#603500000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#603510000000
0!
0'
0/
#603520000000
1!
1'
1/
#603530000000
0!
0'
0/
#603540000000
1!
1'
1/
#603550000000
0!
0'
0/
#603560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#603570000000
0!
0'
0/
#603580000000
1!
1'
1/
#603590000000
0!
0'
0/
#603600000000
1!
1'
1/
#603610000000
0!
0'
0/
#603620000000
1!
1'
1/
#603630000000
0!
0'
0/
#603640000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#603650000000
0!
0'
0/
#603660000000
1!
1'
1/
#603670000000
0!
0'
0/
#603680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#603690000000
0!
0'
0/
#603700000000
1!
1'
1/
#603710000000
0!
0'
0/
#603720000000
#603730000000
1!
1'
1/
#603740000000
0!
0'
0/
#603750000000
1!
1'
1/
#603760000000
0!
1"
0'
1(
0/
10
#603770000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#603780000000
0!
0'
0/
#603790000000
1!
1'
1/
#603800000000
0!
0'
0/
#603810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#603820000000
0!
0'
0/
#603830000000
1!
1'
1/
#603840000000
0!
1"
0'
1(
0/
10
#603850000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#603860000000
0!
1$
0'
1+
0/
#603870000000
1!
1'
1/
#603880000000
0!
0'
0/
#603890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#603900000000
0!
0'
0/
#603910000000
1!
1'
1/
#603920000000
0!
0'
0/
#603930000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#603940000000
0!
0'
0/
#603950000000
1!
1'
1/
#603960000000
0!
0'
0/
#603970000000
1!
1'
1/
#603980000000
0!
0'
0/
#603990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#604000000000
0!
0'
0/
#604010000000
1!
1'
1/
#604020000000
0!
0'
0/
#604030000000
1!
1'
1/
#604040000000
0!
0'
0/
#604050000000
1!
1'
1/
#604060000000
0!
0'
0/
#604070000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#604080000000
0!
0'
0/
#604090000000
1!
1'
1/
#604100000000
0!
0'
0/
#604110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#604120000000
0!
0'
0/
#604130000000
1!
1'
1/
#604140000000
0!
0'
0/
#604150000000
#604160000000
1!
1'
1/
#604170000000
0!
0'
0/
#604180000000
1!
1'
1/
#604190000000
0!
1"
0'
1(
0/
10
#604200000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#604210000000
0!
0'
0/
#604220000000
1!
1'
1/
#604230000000
0!
0'
0/
#604240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#604250000000
0!
0'
0/
#604260000000
1!
1'
1/
#604270000000
0!
1"
0'
1(
0/
10
#604280000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#604290000000
0!
1$
0'
1+
0/
#604300000000
1!
1'
1/
#604310000000
0!
0'
0/
#604320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#604330000000
0!
0'
0/
#604340000000
1!
1'
1/
#604350000000
0!
0'
0/
#604360000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#604370000000
0!
0'
0/
#604380000000
1!
1'
1/
#604390000000
0!
0'
0/
#604400000000
1!
1'
1/
#604410000000
0!
0'
0/
#604420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#604430000000
0!
0'
0/
#604440000000
1!
1'
1/
#604450000000
0!
0'
0/
#604460000000
1!
1'
1/
#604470000000
0!
0'
0/
#604480000000
1!
1'
1/
#604490000000
0!
0'
0/
#604500000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#604510000000
0!
0'
0/
#604520000000
1!
1'
1/
#604530000000
0!
0'
0/
#604540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#604550000000
0!
0'
0/
#604560000000
1!
1'
1/
#604570000000
0!
0'
0/
#604580000000
#604590000000
1!
1'
1/
#604600000000
0!
0'
0/
#604610000000
1!
1'
1/
#604620000000
0!
1"
0'
1(
0/
10
#604630000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#604640000000
0!
0'
0/
#604650000000
1!
1'
1/
#604660000000
0!
0'
0/
#604670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#604680000000
0!
0'
0/
#604690000000
1!
1'
1/
#604700000000
0!
1"
0'
1(
0/
10
#604710000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#604720000000
0!
1$
0'
1+
0/
#604730000000
1!
1'
1/
#604740000000
0!
0'
0/
#604750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#604760000000
0!
0'
0/
#604770000000
1!
1'
1/
#604780000000
0!
0'
0/
#604790000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#604800000000
0!
0'
0/
#604810000000
1!
1'
1/
#604820000000
0!
0'
0/
#604830000000
1!
1'
1/
#604840000000
0!
0'
0/
#604850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#604860000000
0!
0'
0/
#604870000000
1!
1'
1/
#604880000000
0!
0'
0/
#604890000000
1!
1'
1/
#604900000000
0!
0'
0/
#604910000000
1!
1'
1/
#604920000000
0!
0'
0/
#604930000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#604940000000
0!
0'
0/
#604950000000
1!
1'
1/
#604960000000
0!
0'
0/
#604970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#604980000000
0!
0'
0/
#604990000000
1!
1'
1/
#605000000000
0!
0'
0/
#605010000000
#605020000000
1!
1'
1/
#605030000000
0!
0'
0/
#605040000000
1!
1'
1/
#605050000000
0!
1"
0'
1(
0/
10
#605060000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#605070000000
0!
0'
0/
#605080000000
1!
1'
1/
#605090000000
0!
0'
0/
#605100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#605110000000
0!
0'
0/
#605120000000
1!
1'
1/
#605130000000
0!
1"
0'
1(
0/
10
#605140000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#605150000000
0!
1$
0'
1+
0/
#605160000000
1!
1'
1/
#605170000000
0!
0'
0/
#605180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#605190000000
0!
0'
0/
#605200000000
1!
1'
1/
#605210000000
0!
0'
0/
#605220000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#605230000000
0!
0'
0/
#605240000000
1!
1'
1/
#605250000000
0!
0'
0/
#605260000000
1!
1'
1/
#605270000000
0!
0'
0/
#605280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#605290000000
0!
0'
0/
#605300000000
1!
1'
1/
#605310000000
0!
0'
0/
#605320000000
1!
1'
1/
#605330000000
0!
0'
0/
#605340000000
1!
1'
1/
#605350000000
0!
0'
0/
#605360000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#605370000000
0!
0'
0/
#605380000000
1!
1'
1/
#605390000000
0!
0'
0/
#605400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#605410000000
0!
0'
0/
#605420000000
1!
1'
1/
#605430000000
0!
0'
0/
#605440000000
#605450000000
1!
1'
1/
#605460000000
0!
0'
0/
#605470000000
1!
1'
1/
#605480000000
0!
1"
0'
1(
0/
10
#605490000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#605500000000
0!
0'
0/
#605510000000
1!
1'
1/
#605520000000
0!
0'
0/
#605530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#605540000000
0!
0'
0/
#605550000000
1!
1'
1/
#605560000000
0!
1"
0'
1(
0/
10
#605570000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#605580000000
0!
1$
0'
1+
0/
#605590000000
1!
1'
1/
#605600000000
0!
0'
0/
#605610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#605620000000
0!
0'
0/
#605630000000
1!
1'
1/
#605640000000
0!
0'
0/
#605650000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#605660000000
0!
0'
0/
#605670000000
1!
1'
1/
#605680000000
0!
0'
0/
#605690000000
1!
1'
1/
#605700000000
0!
0'
0/
#605710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#605720000000
0!
0'
0/
#605730000000
1!
1'
1/
#605740000000
0!
0'
0/
#605750000000
1!
1'
1/
#605760000000
0!
0'
0/
#605770000000
1!
1'
1/
#605780000000
0!
0'
0/
#605790000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#605800000000
0!
0'
0/
#605810000000
1!
1'
1/
#605820000000
0!
0'
0/
#605830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#605840000000
0!
0'
0/
#605850000000
1!
1'
1/
#605860000000
0!
0'
0/
#605870000000
#605880000000
1!
1'
1/
#605890000000
0!
0'
0/
#605900000000
1!
1'
1/
#605910000000
0!
1"
0'
1(
0/
10
#605920000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#605930000000
0!
0'
0/
#605940000000
1!
1'
1/
#605950000000
0!
0'
0/
#605960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#605970000000
0!
0'
0/
#605980000000
1!
1'
1/
#605990000000
0!
1"
0'
1(
0/
10
#606000000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#606010000000
0!
1$
0'
1+
0/
#606020000000
1!
1'
1/
#606030000000
0!
0'
0/
#606040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#606050000000
0!
0'
0/
#606060000000
1!
1'
1/
#606070000000
0!
0'
0/
#606080000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#606090000000
0!
0'
0/
#606100000000
1!
1'
1/
#606110000000
0!
0'
0/
#606120000000
1!
1'
1/
#606130000000
0!
0'
0/
#606140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#606150000000
0!
0'
0/
#606160000000
1!
1'
1/
#606170000000
0!
0'
0/
#606180000000
1!
1'
1/
#606190000000
0!
0'
0/
#606200000000
1!
1'
1/
#606210000000
0!
0'
0/
#606220000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#606230000000
0!
0'
0/
#606240000000
1!
1'
1/
#606250000000
0!
0'
0/
#606260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#606270000000
0!
0'
0/
#606280000000
1!
1'
1/
#606290000000
0!
0'
0/
#606300000000
#606310000000
1!
1'
1/
#606320000000
0!
0'
0/
#606330000000
1!
1'
1/
#606340000000
0!
1"
0'
1(
0/
10
#606350000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#606360000000
0!
0'
0/
#606370000000
1!
1'
1/
#606380000000
0!
0'
0/
#606390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#606400000000
0!
0'
0/
#606410000000
1!
1'
1/
#606420000000
0!
1"
0'
1(
0/
10
#606430000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#606440000000
0!
1$
0'
1+
0/
#606450000000
1!
1'
1/
#606460000000
0!
0'
0/
#606470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#606480000000
0!
0'
0/
#606490000000
1!
1'
1/
#606500000000
0!
0'
0/
#606510000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#606520000000
0!
0'
0/
#606530000000
1!
1'
1/
#606540000000
0!
0'
0/
#606550000000
1!
1'
1/
#606560000000
0!
0'
0/
#606570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#606580000000
0!
0'
0/
#606590000000
1!
1'
1/
#606600000000
0!
0'
0/
#606610000000
1!
1'
1/
#606620000000
0!
0'
0/
#606630000000
1!
1'
1/
#606640000000
0!
0'
0/
#606650000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#606660000000
0!
0'
0/
#606670000000
1!
1'
1/
#606680000000
0!
0'
0/
#606690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#606700000000
0!
0'
0/
#606710000000
1!
1'
1/
#606720000000
0!
0'
0/
#606730000000
#606740000000
1!
1'
1/
#606750000000
0!
0'
0/
#606760000000
1!
1'
1/
#606770000000
0!
1"
0'
1(
0/
10
#606780000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#606790000000
0!
0'
0/
#606800000000
1!
1'
1/
#606810000000
0!
0'
0/
#606820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#606830000000
0!
0'
0/
#606840000000
1!
1'
1/
#606850000000
0!
1"
0'
1(
0/
10
#606860000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#606870000000
0!
1$
0'
1+
0/
#606880000000
1!
1'
1/
#606890000000
0!
0'
0/
#606900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#606910000000
0!
0'
0/
#606920000000
1!
1'
1/
#606930000000
0!
0'
0/
#606940000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#606950000000
0!
0'
0/
#606960000000
1!
1'
1/
#606970000000
0!
0'
0/
#606980000000
1!
1'
1/
#606990000000
0!
0'
0/
#607000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#607010000000
0!
0'
0/
#607020000000
1!
1'
1/
#607030000000
0!
0'
0/
#607040000000
1!
1'
1/
#607050000000
0!
0'
0/
#607060000000
1!
1'
1/
#607070000000
0!
0'
0/
#607080000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#607090000000
0!
0'
0/
#607100000000
1!
1'
1/
#607110000000
0!
0'
0/
#607120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#607130000000
0!
0'
0/
#607140000000
1!
1'
1/
#607150000000
0!
0'
0/
#607160000000
#607170000000
1!
1'
1/
#607180000000
0!
0'
0/
#607190000000
1!
1'
1/
#607200000000
0!
1"
0'
1(
0/
10
#607210000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#607220000000
0!
0'
0/
#607230000000
1!
1'
1/
#607240000000
0!
0'
0/
#607250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#607260000000
0!
0'
0/
#607270000000
1!
1'
1/
#607280000000
0!
1"
0'
1(
0/
10
#607290000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#607300000000
0!
1$
0'
1+
0/
#607310000000
1!
1'
1/
#607320000000
0!
0'
0/
#607330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#607340000000
0!
0'
0/
#607350000000
1!
1'
1/
#607360000000
0!
0'
0/
#607370000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#607380000000
0!
0'
0/
#607390000000
1!
1'
1/
#607400000000
0!
0'
0/
#607410000000
1!
1'
1/
#607420000000
0!
0'
0/
#607430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#607440000000
0!
0'
0/
#607450000000
1!
1'
1/
#607460000000
0!
0'
0/
#607470000000
1!
1'
1/
#607480000000
0!
0'
0/
#607490000000
1!
1'
1/
#607500000000
0!
0'
0/
#607510000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#607520000000
0!
0'
0/
#607530000000
1!
1'
1/
#607540000000
0!
0'
0/
#607550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#607560000000
0!
0'
0/
#607570000000
1!
1'
1/
#607580000000
0!
0'
0/
#607590000000
#607600000000
1!
1'
1/
#607610000000
0!
0'
0/
#607620000000
1!
1'
1/
#607630000000
0!
1"
0'
1(
0/
10
#607640000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#607650000000
0!
0'
0/
#607660000000
1!
1'
1/
#607670000000
0!
0'
0/
#607680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#607690000000
0!
0'
0/
#607700000000
1!
1'
1/
#607710000000
0!
1"
0'
1(
0/
10
#607720000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#607730000000
0!
1$
0'
1+
0/
#607740000000
1!
1'
1/
#607750000000
0!
0'
0/
#607760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#607770000000
0!
0'
0/
#607780000000
1!
1'
1/
#607790000000
0!
0'
0/
#607800000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#607810000000
0!
0'
0/
#607820000000
1!
1'
1/
#607830000000
0!
0'
0/
#607840000000
1!
1'
1/
#607850000000
0!
0'
0/
#607860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#607870000000
0!
0'
0/
#607880000000
1!
1'
1/
#607890000000
0!
0'
0/
#607900000000
1!
1'
1/
#607910000000
0!
0'
0/
#607920000000
1!
1'
1/
#607930000000
0!
0'
0/
#607940000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#607950000000
0!
0'
0/
#607960000000
1!
1'
1/
#607970000000
0!
0'
0/
#607980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#607990000000
0!
0'
0/
#608000000000
1!
1'
1/
#608010000000
0!
0'
0/
#608020000000
#608030000000
1!
1'
1/
#608040000000
0!
0'
0/
#608050000000
1!
1'
1/
#608060000000
0!
1"
0'
1(
0/
10
#608070000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#608080000000
0!
0'
0/
#608090000000
1!
1'
1/
#608100000000
0!
0'
0/
#608110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#608120000000
0!
0'
0/
#608130000000
1!
1'
1/
#608140000000
0!
1"
0'
1(
0/
10
#608150000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#608160000000
0!
1$
0'
1+
0/
#608170000000
1!
1'
1/
#608180000000
0!
0'
0/
#608190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#608200000000
0!
0'
0/
#608210000000
1!
1'
1/
#608220000000
0!
0'
0/
#608230000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#608240000000
0!
0'
0/
#608250000000
1!
1'
1/
#608260000000
0!
0'
0/
#608270000000
1!
1'
1/
#608280000000
0!
0'
0/
#608290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#608300000000
0!
0'
0/
#608310000000
1!
1'
1/
#608320000000
0!
0'
0/
#608330000000
1!
1'
1/
#608340000000
0!
0'
0/
#608350000000
1!
1'
1/
#608360000000
0!
0'
0/
#608370000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#608380000000
0!
0'
0/
#608390000000
1!
1'
1/
#608400000000
0!
0'
0/
#608410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#608420000000
0!
0'
0/
#608430000000
1!
1'
1/
#608440000000
0!
0'
0/
#608450000000
#608460000000
1!
1'
1/
#608470000000
0!
0'
0/
#608480000000
1!
1'
1/
#608490000000
0!
1"
0'
1(
0/
10
#608500000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#608510000000
0!
0'
0/
#608520000000
1!
1'
1/
#608530000000
0!
0'
0/
#608540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#608550000000
0!
0'
0/
#608560000000
1!
1'
1/
#608570000000
0!
1"
0'
1(
0/
10
#608580000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#608590000000
0!
1$
0'
1+
0/
#608600000000
1!
1'
1/
#608610000000
0!
0'
0/
#608620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#608630000000
0!
0'
0/
#608640000000
1!
1'
1/
#608650000000
0!
0'
0/
#608660000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#608670000000
0!
0'
0/
#608680000000
1!
1'
1/
#608690000000
0!
0'
0/
#608700000000
1!
1'
1/
#608710000000
0!
0'
0/
#608720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#608730000000
0!
0'
0/
#608740000000
1!
1'
1/
#608750000000
0!
0'
0/
#608760000000
1!
1'
1/
#608770000000
0!
0'
0/
#608780000000
1!
1'
1/
#608790000000
0!
0'
0/
#608800000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#608810000000
0!
0'
0/
#608820000000
1!
1'
1/
#608830000000
0!
0'
0/
#608840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#608850000000
0!
0'
0/
#608860000000
1!
1'
1/
#608870000000
0!
0'
0/
#608880000000
#608890000000
1!
1'
1/
#608900000000
0!
0'
0/
#608910000000
1!
1'
1/
#608920000000
0!
1"
0'
1(
0/
10
#608930000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#608940000000
0!
0'
0/
#608950000000
1!
1'
1/
#608960000000
0!
0'
0/
#608970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#608980000000
0!
0'
0/
#608990000000
1!
1'
1/
#609000000000
0!
1"
0'
1(
0/
10
#609010000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#609020000000
0!
1$
0'
1+
0/
#609030000000
1!
1'
1/
#609040000000
0!
0'
0/
#609050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#609060000000
0!
0'
0/
#609070000000
1!
1'
1/
#609080000000
0!
0'
0/
#609090000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#609100000000
0!
0'
0/
#609110000000
1!
1'
1/
#609120000000
0!
0'
0/
#609130000000
1!
1'
1/
#609140000000
0!
0'
0/
#609150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#609160000000
0!
0'
0/
#609170000000
1!
1'
1/
#609180000000
0!
0'
0/
#609190000000
1!
1'
1/
#609200000000
0!
0'
0/
#609210000000
1!
1'
1/
#609220000000
0!
0'
0/
#609230000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#609240000000
0!
0'
0/
#609250000000
1!
1'
1/
#609260000000
0!
0'
0/
#609270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#609280000000
0!
0'
0/
#609290000000
1!
1'
1/
#609300000000
0!
0'
0/
#609310000000
#609320000000
1!
1'
1/
#609330000000
0!
0'
0/
#609340000000
1!
1'
1/
#609350000000
0!
1"
0'
1(
0/
10
#609360000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#609370000000
0!
0'
0/
#609380000000
1!
1'
1/
#609390000000
0!
0'
0/
#609400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#609410000000
0!
0'
0/
#609420000000
1!
1'
1/
#609430000000
0!
1"
0'
1(
0/
10
#609440000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#609450000000
0!
1$
0'
1+
0/
#609460000000
1!
1'
1/
#609470000000
0!
0'
0/
#609480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#609490000000
0!
0'
0/
#609500000000
1!
1'
1/
#609510000000
0!
0'
0/
#609520000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#609530000000
0!
0'
0/
#609540000000
1!
1'
1/
#609550000000
0!
0'
0/
#609560000000
1!
1'
1/
#609570000000
0!
0'
0/
#609580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#609590000000
0!
0'
0/
#609600000000
1!
1'
1/
#609610000000
0!
0'
0/
#609620000000
1!
1'
1/
#609630000000
0!
0'
0/
#609640000000
1!
1'
1/
#609650000000
0!
0'
0/
#609660000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#609670000000
0!
0'
0/
#609680000000
1!
1'
1/
#609690000000
0!
0'
0/
#609700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#609710000000
0!
0'
0/
#609720000000
1!
1'
1/
#609730000000
0!
0'
0/
#609740000000
#609750000000
1!
1'
1/
#609760000000
0!
0'
0/
#609770000000
1!
1'
1/
#609780000000
0!
1"
0'
1(
0/
10
#609790000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#609800000000
0!
0'
0/
#609810000000
1!
1'
1/
#609820000000
0!
0'
0/
#609830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#609840000000
0!
0'
0/
#609850000000
1!
1'
1/
#609860000000
0!
1"
0'
1(
0/
10
#609870000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#609880000000
0!
1$
0'
1+
0/
#609890000000
1!
1'
1/
#609900000000
0!
0'
0/
#609910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#609920000000
0!
0'
0/
#609930000000
1!
1'
1/
#609940000000
0!
0'
0/
#609950000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#609960000000
0!
0'
0/
#609970000000
1!
1'
1/
#609980000000
0!
0'
0/
#609990000000
1!
1'
1/
#610000000000
0!
0'
0/
#610010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#610020000000
0!
0'
0/
#610030000000
1!
1'
1/
#610040000000
0!
0'
0/
#610050000000
1!
1'
1/
#610060000000
0!
0'
0/
#610070000000
1!
1'
1/
#610080000000
0!
0'
0/
#610090000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#610100000000
0!
0'
0/
#610110000000
1!
1'
1/
#610120000000
0!
0'
0/
#610130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#610140000000
0!
0'
0/
#610150000000
1!
1'
1/
#610160000000
0!
0'
0/
#610170000000
#610180000000
1!
1'
1/
#610190000000
0!
0'
0/
#610200000000
1!
1'
1/
#610210000000
0!
1"
0'
1(
0/
10
#610220000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#610230000000
0!
0'
0/
#610240000000
1!
1'
1/
#610250000000
0!
0'
0/
#610260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#610270000000
0!
0'
0/
#610280000000
1!
1'
1/
#610290000000
0!
1"
0'
1(
0/
10
#610300000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#610310000000
0!
1$
0'
1+
0/
#610320000000
1!
1'
1/
#610330000000
0!
0'
0/
#610340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#610350000000
0!
0'
0/
#610360000000
1!
1'
1/
#610370000000
0!
0'
0/
#610380000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#610390000000
0!
0'
0/
#610400000000
1!
1'
1/
#610410000000
0!
0'
0/
#610420000000
1!
1'
1/
#610430000000
0!
0'
0/
#610440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#610450000000
0!
0'
0/
#610460000000
1!
1'
1/
#610470000000
0!
0'
0/
#610480000000
1!
1'
1/
#610490000000
0!
0'
0/
#610500000000
1!
1'
1/
#610510000000
0!
0'
0/
#610520000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#610530000000
0!
0'
0/
#610540000000
1!
1'
1/
#610550000000
0!
0'
0/
#610560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#610570000000
0!
0'
0/
#610580000000
1!
1'
1/
#610590000000
0!
0'
0/
#610600000000
#610610000000
1!
1'
1/
#610620000000
0!
0'
0/
#610630000000
1!
1'
1/
#610640000000
0!
1"
0'
1(
0/
10
#610650000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#610660000000
0!
0'
0/
#610670000000
1!
1'
1/
#610680000000
0!
0'
0/
#610690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#610700000000
0!
0'
0/
#610710000000
1!
1'
1/
#610720000000
0!
1"
0'
1(
0/
10
#610730000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#610740000000
0!
1$
0'
1+
0/
#610750000000
1!
1'
1/
#610760000000
0!
0'
0/
#610770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#610780000000
0!
0'
0/
#610790000000
1!
1'
1/
#610800000000
0!
0'
0/
#610810000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#610820000000
0!
0'
0/
#610830000000
1!
1'
1/
#610840000000
0!
0'
0/
#610850000000
1!
1'
1/
#610860000000
0!
0'
0/
#610870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#610880000000
0!
0'
0/
#610890000000
1!
1'
1/
#610900000000
0!
0'
0/
#610910000000
1!
1'
1/
#610920000000
0!
0'
0/
#610930000000
1!
1'
1/
#610940000000
0!
0'
0/
#610950000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#610960000000
0!
0'
0/
#610970000000
1!
1'
1/
#610980000000
0!
0'
0/
#610990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#611000000000
0!
0'
0/
#611010000000
1!
1'
1/
#611020000000
0!
0'
0/
#611030000000
#611040000000
1!
1'
1/
#611050000000
0!
0'
0/
#611060000000
1!
1'
1/
#611070000000
0!
1"
0'
1(
0/
10
#611080000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#611090000000
0!
0'
0/
#611100000000
1!
1'
1/
#611110000000
0!
0'
0/
#611120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#611130000000
0!
0'
0/
#611140000000
1!
1'
1/
#611150000000
0!
1"
0'
1(
0/
10
#611160000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#611170000000
0!
1$
0'
1+
0/
#611180000000
1!
1'
1/
#611190000000
0!
0'
0/
#611200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#611210000000
0!
0'
0/
#611220000000
1!
1'
1/
#611230000000
0!
0'
0/
#611240000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#611250000000
0!
0'
0/
#611260000000
1!
1'
1/
#611270000000
0!
0'
0/
#611280000000
1!
1'
1/
#611290000000
0!
0'
0/
#611300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#611310000000
0!
0'
0/
#611320000000
1!
1'
1/
#611330000000
0!
0'
0/
#611340000000
1!
1'
1/
#611350000000
0!
0'
0/
#611360000000
1!
1'
1/
#611370000000
0!
0'
0/
#611380000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#611390000000
0!
0'
0/
#611400000000
1!
1'
1/
#611410000000
0!
0'
0/
#611420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#611430000000
0!
0'
0/
#611440000000
1!
1'
1/
#611450000000
0!
0'
0/
#611460000000
#611470000000
1!
1'
1/
#611480000000
0!
0'
0/
#611490000000
1!
1'
1/
#611500000000
0!
1"
0'
1(
0/
10
#611510000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#611520000000
0!
0'
0/
#611530000000
1!
1'
1/
#611540000000
0!
0'
0/
#611550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#611560000000
0!
0'
0/
#611570000000
1!
1'
1/
#611580000000
0!
1"
0'
1(
0/
10
#611590000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#611600000000
0!
1$
0'
1+
0/
#611610000000
1!
1'
1/
#611620000000
0!
0'
0/
#611630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#611640000000
0!
0'
0/
#611650000000
1!
1'
1/
#611660000000
0!
0'
0/
#611670000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#611680000000
0!
0'
0/
#611690000000
1!
1'
1/
#611700000000
0!
0'
0/
#611710000000
1!
1'
1/
#611720000000
0!
0'
0/
#611730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#611740000000
0!
0'
0/
#611750000000
1!
1'
1/
#611760000000
0!
0'
0/
#611770000000
1!
1'
1/
#611780000000
0!
0'
0/
#611790000000
1!
1'
1/
#611800000000
0!
0'
0/
#611810000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#611820000000
0!
0'
0/
#611830000000
1!
1'
1/
#611840000000
0!
0'
0/
#611850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#611860000000
0!
0'
0/
#611870000000
1!
1'
1/
#611880000000
0!
0'
0/
#611890000000
#611900000000
1!
1'
1/
#611910000000
0!
0'
0/
#611920000000
1!
1'
1/
#611930000000
0!
1"
0'
1(
0/
10
#611940000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#611950000000
0!
0'
0/
#611960000000
1!
1'
1/
#611970000000
0!
0'
0/
#611980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#611990000000
0!
0'
0/
#612000000000
1!
1'
1/
#612010000000
0!
1"
0'
1(
0/
10
#612020000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#612030000000
0!
1$
0'
1+
0/
#612040000000
1!
1'
1/
#612050000000
0!
0'
0/
#612060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#612070000000
0!
0'
0/
#612080000000
1!
1'
1/
#612090000000
0!
0'
0/
#612100000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#612110000000
0!
0'
0/
#612120000000
1!
1'
1/
#612130000000
0!
0'
0/
#612140000000
1!
1'
1/
#612150000000
0!
0'
0/
#612160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#612170000000
0!
0'
0/
#612180000000
1!
1'
1/
#612190000000
0!
0'
0/
#612200000000
1!
1'
1/
#612210000000
0!
0'
0/
#612220000000
1!
1'
1/
#612230000000
0!
0'
0/
#612240000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#612250000000
0!
0'
0/
#612260000000
1!
1'
1/
#612270000000
0!
0'
0/
#612280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#612290000000
0!
0'
0/
#612300000000
1!
1'
1/
#612310000000
0!
0'
0/
#612320000000
#612330000000
1!
1'
1/
#612340000000
0!
0'
0/
#612350000000
1!
1'
1/
#612360000000
0!
1"
0'
1(
0/
10
#612370000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#612380000000
0!
0'
0/
#612390000000
1!
1'
1/
#612400000000
0!
0'
0/
#612410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#612420000000
0!
0'
0/
#612430000000
1!
1'
1/
#612440000000
0!
1"
0'
1(
0/
10
#612450000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#612460000000
0!
1$
0'
1+
0/
#612470000000
1!
1'
1/
#612480000000
0!
0'
0/
#612490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#612500000000
0!
0'
0/
#612510000000
1!
1'
1/
#612520000000
0!
0'
0/
#612530000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#612540000000
0!
0'
0/
#612550000000
1!
1'
1/
#612560000000
0!
0'
0/
#612570000000
1!
1'
1/
#612580000000
0!
0'
0/
#612590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#612600000000
0!
0'
0/
#612610000000
1!
1'
1/
#612620000000
0!
0'
0/
#612630000000
1!
1'
1/
#612640000000
0!
0'
0/
#612650000000
1!
1'
1/
#612660000000
0!
0'
0/
#612670000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#612680000000
0!
0'
0/
#612690000000
1!
1'
1/
#612700000000
0!
0'
0/
#612710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#612720000000
0!
0'
0/
#612730000000
1!
1'
1/
#612740000000
0!
0'
0/
#612750000000
#612760000000
1!
1'
1/
#612770000000
0!
0'
0/
#612780000000
1!
1'
1/
#612790000000
0!
1"
0'
1(
0/
10
#612800000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#612810000000
0!
0'
0/
#612820000000
1!
1'
1/
#612830000000
0!
0'
0/
#612840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#612850000000
0!
0'
0/
#612860000000
1!
1'
1/
#612870000000
0!
1"
0'
1(
0/
10
#612880000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#612890000000
0!
1$
0'
1+
0/
#612900000000
1!
1'
1/
#612910000000
0!
0'
0/
#612920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#612930000000
0!
0'
0/
#612940000000
1!
1'
1/
#612950000000
0!
0'
0/
#612960000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#612970000000
0!
0'
0/
#612980000000
1!
1'
1/
#612990000000
0!
0'
0/
#613000000000
1!
1'
1/
#613010000000
0!
0'
0/
#613020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#613030000000
0!
0'
0/
#613040000000
1!
1'
1/
#613050000000
0!
0'
0/
#613060000000
1!
1'
1/
#613070000000
0!
0'
0/
#613080000000
1!
1'
1/
#613090000000
0!
0'
0/
#613100000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#613110000000
0!
0'
0/
#613120000000
1!
1'
1/
#613130000000
0!
0'
0/
#613140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#613150000000
0!
0'
0/
#613160000000
1!
1'
1/
#613170000000
0!
0'
0/
#613180000000
#613190000000
1!
1'
1/
#613200000000
0!
0'
0/
#613210000000
1!
1'
1/
#613220000000
0!
1"
0'
1(
0/
10
#613230000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#613240000000
0!
0'
0/
#613250000000
1!
1'
1/
#613260000000
0!
0'
0/
#613270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#613280000000
0!
0'
0/
#613290000000
1!
1'
1/
#613300000000
0!
1"
0'
1(
0/
10
#613310000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#613320000000
0!
1$
0'
1+
0/
#613330000000
1!
1'
1/
#613340000000
0!
0'
0/
#613350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#613360000000
0!
0'
0/
#613370000000
1!
1'
1/
#613380000000
0!
0'
0/
#613390000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#613400000000
0!
0'
0/
#613410000000
1!
1'
1/
#613420000000
0!
0'
0/
#613430000000
1!
1'
1/
#613440000000
0!
0'
0/
#613450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#613460000000
0!
0'
0/
#613470000000
1!
1'
1/
#613480000000
0!
0'
0/
#613490000000
1!
1'
1/
#613500000000
0!
0'
0/
#613510000000
1!
1'
1/
#613520000000
0!
0'
0/
#613530000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#613540000000
0!
0'
0/
#613550000000
1!
1'
1/
#613560000000
0!
0'
0/
#613570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#613580000000
0!
0'
0/
#613590000000
1!
1'
1/
#613600000000
0!
0'
0/
#613610000000
#613620000000
1!
1'
1/
#613630000000
0!
0'
0/
#613640000000
1!
1'
1/
#613650000000
0!
1"
0'
1(
0/
10
#613660000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#613670000000
0!
0'
0/
#613680000000
1!
1'
1/
#613690000000
0!
0'
0/
#613700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#613710000000
0!
0'
0/
#613720000000
1!
1'
1/
#613730000000
0!
1"
0'
1(
0/
10
#613740000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#613750000000
0!
1$
0'
1+
0/
#613760000000
1!
1'
1/
#613770000000
0!
0'
0/
#613780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#613790000000
0!
0'
0/
#613800000000
1!
1'
1/
#613810000000
0!
0'
0/
#613820000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#613830000000
0!
0'
0/
#613840000000
1!
1'
1/
#613850000000
0!
0'
0/
#613860000000
1!
1'
1/
#613870000000
0!
0'
0/
#613880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#613890000000
0!
0'
0/
#613900000000
1!
1'
1/
#613910000000
0!
0'
0/
#613920000000
1!
1'
1/
#613930000000
0!
0'
0/
#613940000000
1!
1'
1/
#613950000000
0!
0'
0/
#613960000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#613970000000
0!
0'
0/
#613980000000
1!
1'
1/
#613990000000
0!
0'
0/
#614000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#614010000000
0!
0'
0/
#614020000000
1!
1'
1/
#614030000000
0!
0'
0/
#614040000000
#614050000000
1!
1'
1/
#614060000000
0!
0'
0/
#614070000000
1!
1'
1/
#614080000000
0!
1"
0'
1(
0/
10
#614090000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#614100000000
0!
0'
0/
#614110000000
1!
1'
1/
#614120000000
0!
0'
0/
#614130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#614140000000
0!
0'
0/
#614150000000
1!
1'
1/
#614160000000
0!
1"
0'
1(
0/
10
#614170000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#614180000000
0!
1$
0'
1+
0/
#614190000000
1!
1'
1/
#614200000000
0!
0'
0/
#614210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#614220000000
0!
0'
0/
#614230000000
1!
1'
1/
#614240000000
0!
0'
0/
#614250000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#614260000000
0!
0'
0/
#614270000000
1!
1'
1/
#614280000000
0!
0'
0/
#614290000000
1!
1'
1/
#614300000000
0!
0'
0/
#614310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#614320000000
0!
0'
0/
#614330000000
1!
1'
1/
#614340000000
0!
0'
0/
#614350000000
1!
1'
1/
#614360000000
0!
0'
0/
#614370000000
1!
1'
1/
#614380000000
0!
0'
0/
#614390000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#614400000000
0!
0'
0/
#614410000000
1!
1'
1/
#614420000000
0!
0'
0/
#614430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#614440000000
0!
0'
0/
#614450000000
1!
1'
1/
#614460000000
0!
0'
0/
#614470000000
#614480000000
1!
1'
1/
#614490000000
0!
0'
0/
#614500000000
1!
1'
1/
#614510000000
0!
1"
0'
1(
0/
10
#614520000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#614530000000
0!
0'
0/
#614540000000
1!
1'
1/
#614550000000
0!
0'
0/
#614560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#614570000000
0!
0'
0/
#614580000000
1!
1'
1/
#614590000000
0!
1"
0'
1(
0/
10
#614600000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#614610000000
0!
1$
0'
1+
0/
#614620000000
1!
1'
1/
#614630000000
0!
0'
0/
#614640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#614650000000
0!
0'
0/
#614660000000
1!
1'
1/
#614670000000
0!
0'
0/
#614680000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#614690000000
0!
0'
0/
#614700000000
1!
1'
1/
#614710000000
0!
0'
0/
#614720000000
1!
1'
1/
#614730000000
0!
0'
0/
#614740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#614750000000
0!
0'
0/
#614760000000
1!
1'
1/
#614770000000
0!
0'
0/
#614780000000
1!
1'
1/
#614790000000
0!
0'
0/
#614800000000
1!
1'
1/
#614810000000
0!
0'
0/
#614820000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#614830000000
0!
0'
0/
#614840000000
1!
1'
1/
#614850000000
0!
0'
0/
#614860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#614870000000
0!
0'
0/
#614880000000
1!
1'
1/
#614890000000
0!
0'
0/
#614900000000
#614910000000
1!
1'
1/
#614920000000
0!
0'
0/
#614930000000
1!
1'
1/
#614940000000
0!
1"
0'
1(
0/
10
#614950000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#614960000000
0!
0'
0/
#614970000000
1!
1'
1/
#614980000000
0!
0'
0/
#614990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#615000000000
0!
0'
0/
#615010000000
1!
1'
1/
#615020000000
0!
1"
0'
1(
0/
10
#615030000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#615040000000
0!
1$
0'
1+
0/
#615050000000
1!
1'
1/
#615060000000
0!
0'
0/
#615070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#615080000000
0!
0'
0/
#615090000000
1!
1'
1/
#615100000000
0!
0'
0/
#615110000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#615120000000
0!
0'
0/
#615130000000
1!
1'
1/
#615140000000
0!
0'
0/
#615150000000
1!
1'
1/
#615160000000
0!
0'
0/
#615170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#615180000000
0!
0'
0/
#615190000000
1!
1'
1/
#615200000000
0!
0'
0/
#615210000000
1!
1'
1/
#615220000000
0!
0'
0/
#615230000000
1!
1'
1/
#615240000000
0!
0'
0/
#615250000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#615260000000
0!
0'
0/
#615270000000
1!
1'
1/
#615280000000
0!
0'
0/
#615290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#615300000000
0!
0'
0/
#615310000000
1!
1'
1/
#615320000000
0!
0'
0/
#615330000000
#615340000000
1!
1'
1/
#615350000000
0!
0'
0/
#615360000000
1!
1'
1/
#615370000000
0!
1"
0'
1(
0/
10
#615380000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#615390000000
0!
0'
0/
#615400000000
1!
1'
1/
#615410000000
0!
0'
0/
#615420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#615430000000
0!
0'
0/
#615440000000
1!
1'
1/
#615450000000
0!
1"
0'
1(
0/
10
#615460000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#615470000000
0!
1$
0'
1+
0/
#615480000000
1!
1'
1/
#615490000000
0!
0'
0/
#615500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#615510000000
0!
0'
0/
#615520000000
1!
1'
1/
#615530000000
0!
0'
0/
#615540000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#615550000000
0!
0'
0/
#615560000000
1!
1'
1/
#615570000000
0!
0'
0/
#615580000000
1!
1'
1/
#615590000000
0!
0'
0/
#615600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#615610000000
0!
0'
0/
#615620000000
1!
1'
1/
#615630000000
0!
0'
0/
#615640000000
1!
1'
1/
#615650000000
0!
0'
0/
#615660000000
1!
1'
1/
#615670000000
0!
0'
0/
#615680000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#615690000000
0!
0'
0/
#615700000000
1!
1'
1/
#615710000000
0!
0'
0/
#615720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#615730000000
0!
0'
0/
#615740000000
1!
1'
1/
#615750000000
0!
0'
0/
#615760000000
#615770000000
1!
1'
1/
#615780000000
0!
0'
0/
#615790000000
1!
1'
1/
#615800000000
0!
1"
0'
1(
0/
10
#615810000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#615820000000
0!
0'
0/
#615830000000
1!
1'
1/
#615840000000
0!
0'
0/
#615850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#615860000000
0!
0'
0/
#615870000000
1!
1'
1/
#615880000000
0!
1"
0'
1(
0/
10
#615890000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#615900000000
0!
1$
0'
1+
0/
#615910000000
1!
1'
1/
#615920000000
0!
0'
0/
#615930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#615940000000
0!
0'
0/
#615950000000
1!
1'
1/
#615960000000
0!
0'
0/
#615970000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#615980000000
0!
0'
0/
#615990000000
1!
1'
1/
#616000000000
0!
0'
0/
#616010000000
1!
1'
1/
#616020000000
0!
0'
0/
#616030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#616040000000
0!
0'
0/
#616050000000
1!
1'
1/
#616060000000
0!
0'
0/
#616070000000
1!
1'
1/
#616080000000
0!
0'
0/
#616090000000
1!
1'
1/
#616100000000
0!
0'
0/
#616110000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#616120000000
0!
0'
0/
#616130000000
1!
1'
1/
#616140000000
0!
0'
0/
#616150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#616160000000
0!
0'
0/
#616170000000
1!
1'
1/
#616180000000
0!
0'
0/
#616190000000
#616200000000
1!
1'
1/
#616210000000
0!
0'
0/
#616220000000
1!
1'
1/
#616230000000
0!
1"
0'
1(
0/
10
#616240000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#616250000000
0!
0'
0/
#616260000000
1!
1'
1/
#616270000000
0!
0'
0/
#616280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#616290000000
0!
0'
0/
#616300000000
1!
1'
1/
#616310000000
0!
1"
0'
1(
0/
10
#616320000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#616330000000
0!
1$
0'
1+
0/
#616340000000
1!
1'
1/
#616350000000
0!
0'
0/
#616360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#616370000000
0!
0'
0/
#616380000000
1!
1'
1/
#616390000000
0!
0'
0/
#616400000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#616410000000
0!
0'
0/
#616420000000
1!
1'
1/
#616430000000
0!
0'
0/
#616440000000
1!
1'
1/
#616450000000
0!
0'
0/
#616460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#616470000000
0!
0'
0/
#616480000000
1!
1'
1/
#616490000000
0!
0'
0/
#616500000000
1!
1'
1/
#616510000000
0!
0'
0/
#616520000000
1!
1'
1/
#616530000000
0!
0'
0/
#616540000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#616550000000
0!
0'
0/
#616560000000
1!
1'
1/
#616570000000
0!
0'
0/
#616580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#616590000000
0!
0'
0/
#616600000000
1!
1'
1/
#616610000000
0!
0'
0/
#616620000000
#616630000000
1!
1'
1/
#616640000000
0!
0'
0/
#616650000000
1!
1'
1/
#616660000000
0!
1"
0'
1(
0/
10
#616670000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#616680000000
0!
0'
0/
#616690000000
1!
1'
1/
#616700000000
0!
0'
0/
#616710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#616720000000
0!
0'
0/
#616730000000
1!
1'
1/
#616740000000
0!
1"
0'
1(
0/
10
#616750000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#616760000000
0!
1$
0'
1+
0/
#616770000000
1!
1'
1/
#616780000000
0!
0'
0/
#616790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#616800000000
0!
0'
0/
#616810000000
1!
1'
1/
#616820000000
0!
0'
0/
#616830000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#616840000000
0!
0'
0/
#616850000000
1!
1'
1/
#616860000000
0!
0'
0/
#616870000000
1!
1'
1/
#616880000000
0!
0'
0/
#616890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#616900000000
0!
0'
0/
#616910000000
1!
1'
1/
#616920000000
0!
0'
0/
#616930000000
1!
1'
1/
#616940000000
0!
0'
0/
#616950000000
1!
1'
1/
#616960000000
0!
0'
0/
#616970000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#616980000000
0!
0'
0/
#616990000000
1!
1'
1/
#617000000000
0!
0'
0/
#617010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#617020000000
0!
0'
0/
#617030000000
1!
1'
1/
#617040000000
0!
0'
0/
#617050000000
#617060000000
1!
1'
1/
#617070000000
0!
0'
0/
#617080000000
1!
1'
1/
#617090000000
0!
1"
0'
1(
0/
10
#617100000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#617110000000
0!
0'
0/
#617120000000
1!
1'
1/
#617130000000
0!
0'
0/
#617140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#617150000000
0!
0'
0/
#617160000000
1!
1'
1/
#617170000000
0!
1"
0'
1(
0/
10
#617180000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#617190000000
0!
1$
0'
1+
0/
#617200000000
1!
1'
1/
#617210000000
0!
0'
0/
#617220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#617230000000
0!
0'
0/
#617240000000
1!
1'
1/
#617250000000
0!
0'
0/
#617260000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#617270000000
0!
0'
0/
#617280000000
1!
1'
1/
#617290000000
0!
0'
0/
#617300000000
1!
1'
1/
#617310000000
0!
0'
0/
#617320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#617330000000
0!
0'
0/
#617340000000
1!
1'
1/
#617350000000
0!
0'
0/
#617360000000
1!
1'
1/
#617370000000
0!
0'
0/
#617380000000
1!
1'
1/
#617390000000
0!
0'
0/
#617400000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#617410000000
0!
0'
0/
#617420000000
1!
1'
1/
#617430000000
0!
0'
0/
#617440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#617450000000
0!
0'
0/
#617460000000
1!
1'
1/
#617470000000
0!
0'
0/
#617480000000
#617490000000
1!
1'
1/
#617500000000
0!
0'
0/
#617510000000
1!
1'
1/
#617520000000
0!
1"
0'
1(
0/
10
#617530000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#617540000000
0!
0'
0/
#617550000000
1!
1'
1/
#617560000000
0!
0'
0/
#617570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#617580000000
0!
0'
0/
#617590000000
1!
1'
1/
#617600000000
0!
1"
0'
1(
0/
10
#617610000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#617620000000
0!
1$
0'
1+
0/
#617630000000
1!
1'
1/
#617640000000
0!
0'
0/
#617650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#617660000000
0!
0'
0/
#617670000000
1!
1'
1/
#617680000000
0!
0'
0/
#617690000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#617700000000
0!
0'
0/
#617710000000
1!
1'
1/
#617720000000
0!
0'
0/
#617730000000
1!
1'
1/
#617740000000
0!
0'
0/
#617750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#617760000000
0!
0'
0/
#617770000000
1!
1'
1/
#617780000000
0!
0'
0/
#617790000000
1!
1'
1/
#617800000000
0!
0'
0/
#617810000000
1!
1'
1/
#617820000000
0!
0'
0/
#617830000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#617840000000
0!
0'
0/
#617850000000
1!
1'
1/
#617860000000
0!
0'
0/
#617870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#617880000000
0!
0'
0/
#617890000000
1!
1'
1/
#617900000000
0!
0'
0/
#617910000000
#617920000000
1!
1'
1/
#617930000000
0!
0'
0/
#617940000000
1!
1'
1/
#617950000000
0!
1"
0'
1(
0/
10
#617960000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#617970000000
0!
0'
0/
#617980000000
1!
1'
1/
#617990000000
0!
0'
0/
#618000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#618010000000
0!
0'
0/
#618020000000
1!
1'
1/
#618030000000
0!
1"
0'
1(
0/
10
#618040000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#618050000000
0!
1$
0'
1+
0/
#618060000000
1!
1'
1/
#618070000000
0!
0'
0/
#618080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#618090000000
0!
0'
0/
#618100000000
1!
1'
1/
#618110000000
0!
0'
0/
#618120000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#618130000000
0!
0'
0/
#618140000000
1!
1'
1/
#618150000000
0!
0'
0/
#618160000000
1!
1'
1/
#618170000000
0!
0'
0/
#618180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#618190000000
0!
0'
0/
#618200000000
1!
1'
1/
#618210000000
0!
0'
0/
#618220000000
1!
1'
1/
#618230000000
0!
0'
0/
#618240000000
1!
1'
1/
#618250000000
0!
0'
0/
#618260000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#618270000000
0!
0'
0/
#618280000000
1!
1'
1/
#618290000000
0!
0'
0/
#618300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#618310000000
0!
0'
0/
#618320000000
1!
1'
1/
#618330000000
0!
0'
0/
#618340000000
#618350000000
1!
1'
1/
#618360000000
0!
0'
0/
#618370000000
1!
1'
1/
#618380000000
0!
1"
0'
1(
0/
10
#618390000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#618400000000
0!
0'
0/
#618410000000
1!
1'
1/
#618420000000
0!
0'
0/
#618430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#618440000000
0!
0'
0/
#618450000000
1!
1'
1/
#618460000000
0!
1"
0'
1(
0/
10
#618470000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#618480000000
0!
1$
0'
1+
0/
#618490000000
1!
1'
1/
#618500000000
0!
0'
0/
#618510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#618520000000
0!
0'
0/
#618530000000
1!
1'
1/
#618540000000
0!
0'
0/
#618550000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#618560000000
0!
0'
0/
#618570000000
1!
1'
1/
#618580000000
0!
0'
0/
#618590000000
1!
1'
1/
#618600000000
0!
0'
0/
#618610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#618620000000
0!
0'
0/
#618630000000
1!
1'
1/
#618640000000
0!
0'
0/
#618650000000
1!
1'
1/
#618660000000
0!
0'
0/
#618670000000
1!
1'
1/
#618680000000
0!
0'
0/
#618690000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#618700000000
0!
0'
0/
#618710000000
1!
1'
1/
#618720000000
0!
0'
0/
#618730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#618740000000
0!
0'
0/
#618750000000
1!
1'
1/
#618760000000
0!
0'
0/
#618770000000
#618780000000
1!
1'
1/
#618790000000
0!
0'
0/
#618800000000
1!
1'
1/
#618810000000
0!
1"
0'
1(
0/
10
#618820000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#618830000000
0!
0'
0/
#618840000000
1!
1'
1/
#618850000000
0!
0'
0/
#618860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#618870000000
0!
0'
0/
#618880000000
1!
1'
1/
#618890000000
0!
1"
0'
1(
0/
10
#618900000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#618910000000
0!
1$
0'
1+
0/
#618920000000
1!
1'
1/
#618930000000
0!
0'
0/
#618940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#618950000000
0!
0'
0/
#618960000000
1!
1'
1/
#618970000000
0!
0'
0/
#618980000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#618990000000
0!
0'
0/
#619000000000
1!
1'
1/
#619010000000
0!
0'
0/
#619020000000
1!
1'
1/
#619030000000
0!
0'
0/
#619040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#619050000000
0!
0'
0/
#619060000000
1!
1'
1/
#619070000000
0!
0'
0/
#619080000000
1!
1'
1/
#619090000000
0!
0'
0/
#619100000000
1!
1'
1/
#619110000000
0!
0'
0/
#619120000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#619130000000
0!
0'
0/
#619140000000
1!
1'
1/
#619150000000
0!
0'
0/
#619160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#619170000000
0!
0'
0/
#619180000000
1!
1'
1/
#619190000000
0!
0'
0/
#619200000000
#619210000000
1!
1'
1/
#619220000000
0!
0'
0/
#619230000000
1!
1'
1/
#619240000000
0!
1"
0'
1(
0/
10
#619250000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#619260000000
0!
0'
0/
#619270000000
1!
1'
1/
#619280000000
0!
0'
0/
#619290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#619300000000
0!
0'
0/
#619310000000
1!
1'
1/
#619320000000
0!
1"
0'
1(
0/
10
#619330000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#619340000000
0!
1$
0'
1+
0/
#619350000000
1!
1'
1/
#619360000000
0!
0'
0/
#619370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#619380000000
0!
0'
0/
#619390000000
1!
1'
1/
#619400000000
0!
0'
0/
#619410000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#619420000000
0!
0'
0/
#619430000000
1!
1'
1/
#619440000000
0!
0'
0/
#619450000000
1!
1'
1/
#619460000000
0!
0'
0/
#619470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#619480000000
0!
0'
0/
#619490000000
1!
1'
1/
#619500000000
0!
0'
0/
#619510000000
1!
1'
1/
#619520000000
0!
0'
0/
#619530000000
1!
1'
1/
#619540000000
0!
0'
0/
#619550000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#619560000000
0!
0'
0/
#619570000000
1!
1'
1/
#619580000000
0!
0'
0/
#619590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#619600000000
0!
0'
0/
#619610000000
1!
1'
1/
#619620000000
0!
0'
0/
#619630000000
#619640000000
1!
1'
1/
#619650000000
0!
0'
0/
#619660000000
1!
1'
1/
#619670000000
0!
1"
0'
1(
0/
10
#619680000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#619690000000
0!
0'
0/
#619700000000
1!
1'
1/
#619710000000
0!
0'
0/
#619720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#619730000000
0!
0'
0/
#619740000000
1!
1'
1/
#619750000000
0!
1"
0'
1(
0/
10
#619760000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#619770000000
0!
1$
0'
1+
0/
#619780000000
1!
1'
1/
#619790000000
0!
0'
0/
#619800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#619810000000
0!
0'
0/
#619820000000
1!
1'
1/
#619830000000
0!
0'
0/
#619840000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#619850000000
0!
0'
0/
#619860000000
1!
1'
1/
#619870000000
0!
0'
0/
#619880000000
1!
1'
1/
#619890000000
0!
0'
0/
#619900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#619910000000
0!
0'
0/
#619920000000
1!
1'
1/
#619930000000
0!
0'
0/
#619940000000
1!
1'
1/
#619950000000
0!
0'
0/
#619960000000
1!
1'
1/
#619970000000
0!
0'
0/
#619980000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#619990000000
0!
0'
0/
#620000000000
1!
1'
1/
#620010000000
0!
0'
0/
#620020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#620030000000
0!
0'
0/
#620040000000
1!
1'
1/
#620050000000
0!
0'
0/
#620060000000
#620070000000
1!
1'
1/
#620080000000
0!
0'
0/
#620090000000
1!
1'
1/
#620100000000
0!
1"
0'
1(
0/
10
#620110000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#620120000000
0!
0'
0/
#620130000000
1!
1'
1/
#620140000000
0!
0'
0/
#620150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#620160000000
0!
0'
0/
#620170000000
1!
1'
1/
#620180000000
0!
1"
0'
1(
0/
10
#620190000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#620200000000
0!
1$
0'
1+
0/
#620210000000
1!
1'
1/
#620220000000
0!
0'
0/
#620230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#620240000000
0!
0'
0/
#620250000000
1!
1'
1/
#620260000000
0!
0'
0/
#620270000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#620280000000
0!
0'
0/
#620290000000
1!
1'
1/
#620300000000
0!
0'
0/
#620310000000
1!
1'
1/
#620320000000
0!
0'
0/
#620330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#620340000000
0!
0'
0/
#620350000000
1!
1'
1/
#620360000000
0!
0'
0/
#620370000000
1!
1'
1/
#620380000000
0!
0'
0/
#620390000000
1!
1'
1/
#620400000000
0!
0'
0/
#620410000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#620420000000
0!
0'
0/
#620430000000
1!
1'
1/
#620440000000
0!
0'
0/
#620450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#620460000000
0!
0'
0/
#620470000000
1!
1'
1/
#620480000000
0!
0'
0/
#620490000000
#620500000000
1!
1'
1/
#620510000000
0!
0'
0/
#620520000000
1!
1'
1/
#620530000000
0!
1"
0'
1(
0/
10
#620540000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#620550000000
0!
0'
0/
#620560000000
1!
1'
1/
#620570000000
0!
0'
0/
#620580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#620590000000
0!
0'
0/
#620600000000
1!
1'
1/
#620610000000
0!
1"
0'
1(
0/
10
#620620000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#620630000000
0!
1$
0'
1+
0/
#620640000000
1!
1'
1/
#620650000000
0!
0'
0/
#620660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#620670000000
0!
0'
0/
#620680000000
1!
1'
1/
#620690000000
0!
0'
0/
#620700000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#620710000000
0!
0'
0/
#620720000000
1!
1'
1/
#620730000000
0!
0'
0/
#620740000000
1!
1'
1/
#620750000000
0!
0'
0/
#620760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#620770000000
0!
0'
0/
#620780000000
1!
1'
1/
#620790000000
0!
0'
0/
#620800000000
1!
1'
1/
#620810000000
0!
0'
0/
#620820000000
1!
1'
1/
#620830000000
0!
0'
0/
#620840000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#620850000000
0!
0'
0/
#620860000000
1!
1'
1/
#620870000000
0!
0'
0/
#620880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#620890000000
0!
0'
0/
#620900000000
1!
1'
1/
#620910000000
0!
0'
0/
#620920000000
#620930000000
1!
1'
1/
#620940000000
0!
0'
0/
#620950000000
1!
1'
1/
#620960000000
0!
1"
0'
1(
0/
10
#620970000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#620980000000
0!
0'
0/
#620990000000
1!
1'
1/
#621000000000
0!
0'
0/
#621010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#621020000000
0!
0'
0/
#621030000000
1!
1'
1/
#621040000000
0!
1"
0'
1(
0/
10
#621050000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#621060000000
0!
1$
0'
1+
0/
#621070000000
1!
1'
1/
#621080000000
0!
0'
0/
#621090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#621100000000
0!
0'
0/
#621110000000
1!
1'
1/
#621120000000
0!
0'
0/
#621130000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#621140000000
0!
0'
0/
#621150000000
1!
1'
1/
#621160000000
0!
0'
0/
#621170000000
1!
1'
1/
#621180000000
0!
0'
0/
#621190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#621200000000
0!
0'
0/
#621210000000
1!
1'
1/
#621220000000
0!
0'
0/
#621230000000
1!
1'
1/
#621240000000
0!
0'
0/
#621250000000
1!
1'
1/
#621260000000
0!
0'
0/
#621270000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#621280000000
0!
0'
0/
#621290000000
1!
1'
1/
#621300000000
0!
0'
0/
#621310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#621320000000
0!
0'
0/
#621330000000
1!
1'
1/
#621340000000
0!
0'
0/
#621350000000
#621360000000
1!
1'
1/
#621370000000
0!
0'
0/
#621380000000
1!
1'
1/
#621390000000
0!
1"
0'
1(
0/
10
#621400000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#621410000000
0!
0'
0/
#621420000000
1!
1'
1/
#621430000000
0!
0'
0/
#621440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#621450000000
0!
0'
0/
#621460000000
1!
1'
1/
#621470000000
0!
1"
0'
1(
0/
10
#621480000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#621490000000
0!
1$
0'
1+
0/
#621500000000
1!
1'
1/
#621510000000
0!
0'
0/
#621520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#621530000000
0!
0'
0/
#621540000000
1!
1'
1/
#621550000000
0!
0'
0/
#621560000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#621570000000
0!
0'
0/
#621580000000
1!
1'
1/
#621590000000
0!
0'
0/
#621600000000
1!
1'
1/
#621610000000
0!
0'
0/
#621620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#621630000000
0!
0'
0/
#621640000000
1!
1'
1/
#621650000000
0!
0'
0/
#621660000000
1!
1'
1/
#621670000000
0!
0'
0/
#621680000000
1!
1'
1/
#621690000000
0!
0'
0/
#621700000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#621710000000
0!
0'
0/
#621720000000
1!
1'
1/
#621730000000
0!
0'
0/
#621740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#621750000000
0!
0'
0/
#621760000000
1!
1'
1/
#621770000000
0!
0'
0/
#621780000000
#621790000000
1!
1'
1/
#621800000000
0!
0'
0/
#621810000000
1!
1'
1/
#621820000000
0!
1"
0'
1(
0/
10
#621830000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#621840000000
0!
0'
0/
#621850000000
1!
1'
1/
#621860000000
0!
0'
0/
#621870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#621880000000
0!
0'
0/
#621890000000
1!
1'
1/
#621900000000
0!
1"
0'
1(
0/
10
#621910000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#621920000000
0!
1$
0'
1+
0/
#621930000000
1!
1'
1/
#621940000000
0!
0'
0/
#621950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#621960000000
0!
0'
0/
#621970000000
1!
1'
1/
#621980000000
0!
0'
0/
#621990000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#622000000000
0!
0'
0/
#622010000000
1!
1'
1/
#622020000000
0!
0'
0/
#622030000000
1!
1'
1/
#622040000000
0!
0'
0/
#622050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#622060000000
0!
0'
0/
#622070000000
1!
1'
1/
#622080000000
0!
0'
0/
#622090000000
1!
1'
1/
#622100000000
0!
0'
0/
#622110000000
1!
1'
1/
#622120000000
0!
0'
0/
#622130000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#622140000000
0!
0'
0/
#622150000000
1!
1'
1/
#622160000000
0!
0'
0/
#622170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#622180000000
0!
0'
0/
#622190000000
1!
1'
1/
#622200000000
0!
0'
0/
#622210000000
#622220000000
1!
1'
1/
#622230000000
0!
0'
0/
#622240000000
1!
1'
1/
#622250000000
0!
1"
0'
1(
0/
10
#622260000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#622270000000
0!
0'
0/
#622280000000
1!
1'
1/
#622290000000
0!
0'
0/
#622300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#622310000000
0!
0'
0/
#622320000000
1!
1'
1/
#622330000000
0!
1"
0'
1(
0/
10
#622340000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#622350000000
0!
1$
0'
1+
0/
#622360000000
1!
1'
1/
#622370000000
0!
0'
0/
#622380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#622390000000
0!
0'
0/
#622400000000
1!
1'
1/
#622410000000
0!
0'
0/
#622420000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#622430000000
0!
0'
0/
#622440000000
1!
1'
1/
#622450000000
0!
0'
0/
#622460000000
1!
1'
1/
#622470000000
0!
0'
0/
#622480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#622490000000
0!
0'
0/
#622500000000
1!
1'
1/
#622510000000
0!
0'
0/
#622520000000
1!
1'
1/
#622530000000
0!
0'
0/
#622540000000
1!
1'
1/
#622550000000
0!
0'
0/
#622560000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#622570000000
0!
0'
0/
#622580000000
1!
1'
1/
#622590000000
0!
0'
0/
#622600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#622610000000
0!
0'
0/
#622620000000
1!
1'
1/
#622630000000
0!
0'
0/
#622640000000
#622650000000
1!
1'
1/
#622660000000
0!
0'
0/
#622670000000
1!
1'
1/
#622680000000
0!
1"
0'
1(
0/
10
#622690000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#622700000000
0!
0'
0/
#622710000000
1!
1'
1/
#622720000000
0!
0'
0/
#622730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#622740000000
0!
0'
0/
#622750000000
1!
1'
1/
#622760000000
0!
1"
0'
1(
0/
10
#622770000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#622780000000
0!
1$
0'
1+
0/
#622790000000
1!
1'
1/
#622800000000
0!
0'
0/
#622810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#622820000000
0!
0'
0/
#622830000000
1!
1'
1/
#622840000000
0!
0'
0/
#622850000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#622860000000
0!
0'
0/
#622870000000
1!
1'
1/
#622880000000
0!
0'
0/
#622890000000
1!
1'
1/
#622900000000
0!
0'
0/
#622910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#622920000000
0!
0'
0/
#622930000000
1!
1'
1/
#622940000000
0!
0'
0/
#622950000000
1!
1'
1/
#622960000000
0!
0'
0/
#622970000000
1!
1'
1/
#622980000000
0!
0'
0/
#622990000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#623000000000
0!
0'
0/
#623010000000
1!
1'
1/
#623020000000
0!
0'
0/
#623030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#623040000000
0!
0'
0/
#623050000000
1!
1'
1/
#623060000000
0!
0'
0/
#623070000000
#623080000000
1!
1'
1/
#623090000000
0!
0'
0/
#623100000000
1!
1'
1/
#623110000000
0!
1"
0'
1(
0/
10
#623120000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#623130000000
0!
0'
0/
#623140000000
1!
1'
1/
#623150000000
0!
0'
0/
#623160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#623170000000
0!
0'
0/
#623180000000
1!
1'
1/
#623190000000
0!
1"
0'
1(
0/
10
#623200000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#623210000000
0!
1$
0'
1+
0/
#623220000000
1!
1'
1/
#623230000000
0!
0'
0/
#623240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#623250000000
0!
0'
0/
#623260000000
1!
1'
1/
#623270000000
0!
0'
0/
#623280000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#623290000000
0!
0'
0/
#623300000000
1!
1'
1/
#623310000000
0!
0'
0/
#623320000000
1!
1'
1/
#623330000000
0!
0'
0/
#623340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#623350000000
0!
0'
0/
#623360000000
1!
1'
1/
#623370000000
0!
0'
0/
#623380000000
1!
1'
1/
#623390000000
0!
0'
0/
#623400000000
1!
1'
1/
#623410000000
0!
0'
0/
#623420000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#623430000000
0!
0'
0/
#623440000000
1!
1'
1/
#623450000000
0!
0'
0/
#623460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#623470000000
0!
0'
0/
#623480000000
1!
1'
1/
#623490000000
0!
0'
0/
#623500000000
#623510000000
1!
1'
1/
#623520000000
0!
0'
0/
#623530000000
1!
1'
1/
#623540000000
0!
1"
0'
1(
0/
10
#623550000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#623560000000
0!
0'
0/
#623570000000
1!
1'
1/
#623580000000
0!
0'
0/
#623590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#623600000000
0!
0'
0/
#623610000000
1!
1'
1/
#623620000000
0!
1"
0'
1(
0/
10
#623630000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#623640000000
0!
1$
0'
1+
0/
#623650000000
1!
1'
1/
#623660000000
0!
0'
0/
#623670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#623680000000
0!
0'
0/
#623690000000
1!
1'
1/
#623700000000
0!
0'
0/
#623710000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#623720000000
0!
0'
0/
#623730000000
1!
1'
1/
#623740000000
0!
0'
0/
#623750000000
1!
1'
1/
#623760000000
0!
0'
0/
#623770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#623780000000
0!
0'
0/
#623790000000
1!
1'
1/
#623800000000
0!
0'
0/
#623810000000
1!
1'
1/
#623820000000
0!
0'
0/
#623830000000
1!
1'
1/
#623840000000
0!
0'
0/
#623850000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#623860000000
0!
0'
0/
#623870000000
1!
1'
1/
#623880000000
0!
0'
0/
#623890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#623900000000
0!
0'
0/
#623910000000
1!
1'
1/
#623920000000
0!
0'
0/
#623930000000
#623940000000
1!
1'
1/
#623950000000
0!
0'
0/
#623960000000
1!
1'
1/
#623970000000
0!
1"
0'
1(
0/
10
#623980000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#623990000000
0!
0'
0/
#624000000000
1!
1'
1/
#624010000000
0!
0'
0/
#624020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#624030000000
0!
0'
0/
#624040000000
1!
1'
1/
#624050000000
0!
1"
0'
1(
0/
10
#624060000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#624070000000
0!
1$
0'
1+
0/
#624080000000
1!
1'
1/
#624090000000
0!
0'
0/
#624100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#624110000000
0!
0'
0/
#624120000000
1!
1'
1/
#624130000000
0!
0'
0/
#624140000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#624150000000
0!
0'
0/
#624160000000
1!
1'
1/
#624170000000
0!
0'
0/
#624180000000
1!
1'
1/
#624190000000
0!
0'
0/
#624200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#624210000000
0!
0'
0/
#624220000000
1!
1'
1/
#624230000000
0!
0'
0/
#624240000000
1!
1'
1/
#624250000000
0!
0'
0/
#624260000000
1!
1'
1/
#624270000000
0!
0'
0/
#624280000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#624290000000
0!
0'
0/
#624300000000
1!
1'
1/
#624310000000
0!
0'
0/
#624320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#624330000000
0!
0'
0/
#624340000000
1!
1'
1/
#624350000000
0!
0'
0/
#624360000000
#624370000000
1!
1'
1/
#624380000000
0!
0'
0/
#624390000000
1!
1'
1/
#624400000000
0!
1"
0'
1(
0/
10
#624410000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#624420000000
0!
0'
0/
#624430000000
1!
1'
1/
#624440000000
0!
0'
0/
#624450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#624460000000
0!
0'
0/
#624470000000
1!
1'
1/
#624480000000
0!
1"
0'
1(
0/
10
#624490000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#624500000000
0!
1$
0'
1+
0/
#624510000000
1!
1'
1/
#624520000000
0!
0'
0/
#624530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#624540000000
0!
0'
0/
#624550000000
1!
1'
1/
#624560000000
0!
0'
0/
#624570000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#624580000000
0!
0'
0/
#624590000000
1!
1'
1/
#624600000000
0!
0'
0/
#624610000000
1!
1'
1/
#624620000000
0!
0'
0/
#624630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#624640000000
0!
0'
0/
#624650000000
1!
1'
1/
#624660000000
0!
0'
0/
#624670000000
1!
1'
1/
#624680000000
0!
0'
0/
#624690000000
1!
1'
1/
#624700000000
0!
0'
0/
#624710000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#624720000000
0!
0'
0/
#624730000000
1!
1'
1/
#624740000000
0!
0'
0/
#624750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#624760000000
0!
0'
0/
#624770000000
1!
1'
1/
#624780000000
0!
0'
0/
#624790000000
#624800000000
1!
1'
1/
#624810000000
0!
0'
0/
#624820000000
1!
1'
1/
#624830000000
0!
1"
0'
1(
0/
10
#624840000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#624850000000
0!
0'
0/
#624860000000
1!
1'
1/
#624870000000
0!
0'
0/
#624880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#624890000000
0!
0'
0/
#624900000000
1!
1'
1/
#624910000000
0!
1"
0'
1(
0/
10
#624920000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#624930000000
0!
1$
0'
1+
0/
#624940000000
1!
1'
1/
#624950000000
0!
0'
0/
#624960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#624970000000
0!
0'
0/
#624980000000
1!
1'
1/
#624990000000
0!
0'
0/
#625000000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#625010000000
0!
0'
0/
#625020000000
1!
1'
1/
#625030000000
0!
0'
0/
#625040000000
1!
1'
1/
#625050000000
0!
0'
0/
#625060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#625070000000
0!
0'
0/
#625080000000
1!
1'
1/
#625090000000
0!
0'
0/
#625100000000
1!
1'
1/
#625110000000
0!
0'
0/
#625120000000
1!
1'
1/
#625130000000
0!
0'
0/
#625140000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#625150000000
0!
0'
0/
#625160000000
1!
1'
1/
#625170000000
0!
0'
0/
#625180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#625190000000
0!
0'
0/
#625200000000
1!
1'
1/
#625210000000
0!
0'
0/
#625220000000
#625230000000
1!
1'
1/
#625240000000
0!
0'
0/
#625250000000
1!
1'
1/
#625260000000
0!
1"
0'
1(
0/
10
#625270000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#625280000000
0!
0'
0/
#625290000000
1!
1'
1/
#625300000000
0!
0'
0/
#625310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#625320000000
0!
0'
0/
#625330000000
1!
1'
1/
#625340000000
0!
1"
0'
1(
0/
10
#625350000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#625360000000
0!
1$
0'
1+
0/
#625370000000
1!
1'
1/
#625380000000
0!
0'
0/
#625390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#625400000000
0!
0'
0/
#625410000000
1!
1'
1/
#625420000000
0!
0'
0/
#625430000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#625440000000
0!
0'
0/
#625450000000
1!
1'
1/
#625460000000
0!
0'
0/
#625470000000
1!
1'
1/
#625480000000
0!
0'
0/
#625490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#625500000000
0!
0'
0/
#625510000000
1!
1'
1/
#625520000000
0!
0'
0/
#625530000000
1!
1'
1/
#625540000000
0!
0'
0/
#625550000000
1!
1'
1/
#625560000000
0!
0'
0/
#625570000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#625580000000
0!
0'
0/
#625590000000
1!
1'
1/
#625600000000
0!
0'
0/
#625610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#625620000000
0!
0'
0/
#625630000000
1!
1'
1/
#625640000000
0!
0'
0/
#625650000000
#625660000000
1!
1'
1/
#625670000000
0!
0'
0/
#625680000000
1!
1'
1/
#625690000000
0!
1"
0'
1(
0/
10
#625700000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#625710000000
0!
0'
0/
#625720000000
1!
1'
1/
#625730000000
0!
0'
0/
#625740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#625750000000
0!
0'
0/
#625760000000
1!
1'
1/
#625770000000
0!
1"
0'
1(
0/
10
#625780000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#625790000000
0!
1$
0'
1+
0/
#625800000000
1!
1'
1/
#625810000000
0!
0'
0/
#625820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#625830000000
0!
0'
0/
#625840000000
1!
1'
1/
#625850000000
0!
0'
0/
#625860000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#625870000000
0!
0'
0/
#625880000000
1!
1'
1/
#625890000000
0!
0'
0/
#625900000000
1!
1'
1/
#625910000000
0!
0'
0/
#625920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#625930000000
0!
0'
0/
#625940000000
1!
1'
1/
#625950000000
0!
0'
0/
#625960000000
1!
1'
1/
#625970000000
0!
0'
0/
#625980000000
1!
1'
1/
#625990000000
0!
0'
0/
#626000000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#626010000000
0!
0'
0/
#626020000000
1!
1'
1/
#626030000000
0!
0'
0/
#626040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#626050000000
0!
0'
0/
#626060000000
1!
1'
1/
#626070000000
0!
0'
0/
#626080000000
#626090000000
1!
1'
1/
#626100000000
0!
0'
0/
#626110000000
1!
1'
1/
#626120000000
0!
1"
0'
1(
0/
10
#626130000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#626140000000
0!
0'
0/
#626150000000
1!
1'
1/
#626160000000
0!
0'
0/
#626170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#626180000000
0!
0'
0/
#626190000000
1!
1'
1/
#626200000000
0!
1"
0'
1(
0/
10
#626210000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#626220000000
0!
1$
0'
1+
0/
#626230000000
1!
1'
1/
#626240000000
0!
0'
0/
#626250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#626260000000
0!
0'
0/
#626270000000
1!
1'
1/
#626280000000
0!
0'
0/
#626290000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#626300000000
0!
0'
0/
#626310000000
1!
1'
1/
#626320000000
0!
0'
0/
#626330000000
1!
1'
1/
#626340000000
0!
0'
0/
#626350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#626360000000
0!
0'
0/
#626370000000
1!
1'
1/
#626380000000
0!
0'
0/
#626390000000
1!
1'
1/
#626400000000
0!
0'
0/
#626410000000
1!
1'
1/
#626420000000
0!
0'
0/
#626430000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#626440000000
0!
0'
0/
#626450000000
1!
1'
1/
#626460000000
0!
0'
0/
#626470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#626480000000
0!
0'
0/
#626490000000
1!
1'
1/
#626500000000
0!
0'
0/
#626510000000
#626520000000
1!
1'
1/
#626530000000
0!
0'
0/
#626540000000
1!
1'
1/
#626550000000
0!
1"
0'
1(
0/
10
#626560000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#626570000000
0!
0'
0/
#626580000000
1!
1'
1/
#626590000000
0!
0'
0/
#626600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#626610000000
0!
0'
0/
#626620000000
1!
1'
1/
#626630000000
0!
1"
0'
1(
0/
10
#626640000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#626650000000
0!
1$
0'
1+
0/
#626660000000
1!
1'
1/
#626670000000
0!
0'
0/
#626680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#626690000000
0!
0'
0/
#626700000000
1!
1'
1/
#626710000000
0!
0'
0/
#626720000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#626730000000
0!
0'
0/
#626740000000
1!
1'
1/
#626750000000
0!
0'
0/
#626760000000
1!
1'
1/
#626770000000
0!
0'
0/
#626780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#626790000000
0!
0'
0/
#626800000000
1!
1'
1/
#626810000000
0!
0'
0/
#626820000000
1!
1'
1/
#626830000000
0!
0'
0/
#626840000000
1!
1'
1/
#626850000000
0!
0'
0/
#626860000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#626870000000
0!
0'
0/
#626880000000
1!
1'
1/
#626890000000
0!
0'
0/
#626900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#626910000000
0!
0'
0/
#626920000000
1!
1'
1/
#626930000000
0!
0'
0/
#626940000000
#626950000000
1!
1'
1/
#626960000000
0!
0'
0/
#626970000000
1!
1'
1/
#626980000000
0!
1"
0'
1(
0/
10
#626990000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#627000000000
0!
0'
0/
#627010000000
1!
1'
1/
#627020000000
0!
0'
0/
#627030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#627040000000
0!
0'
0/
#627050000000
1!
1'
1/
#627060000000
0!
1"
0'
1(
0/
10
#627070000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#627080000000
0!
1$
0'
1+
0/
#627090000000
1!
1'
1/
#627100000000
0!
0'
0/
#627110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#627120000000
0!
0'
0/
#627130000000
1!
1'
1/
#627140000000
0!
0'
0/
#627150000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#627160000000
0!
0'
0/
#627170000000
1!
1'
1/
#627180000000
0!
0'
0/
#627190000000
1!
1'
1/
#627200000000
0!
0'
0/
#627210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#627220000000
0!
0'
0/
#627230000000
1!
1'
1/
#627240000000
0!
0'
0/
#627250000000
1!
1'
1/
#627260000000
0!
0'
0/
#627270000000
1!
1'
1/
#627280000000
0!
0'
0/
#627290000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#627300000000
0!
0'
0/
#627310000000
1!
1'
1/
#627320000000
0!
0'
0/
#627330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#627340000000
0!
0'
0/
#627350000000
1!
1'
1/
#627360000000
0!
0'
0/
#627370000000
#627380000000
1!
1'
1/
#627390000000
0!
0'
0/
#627400000000
1!
1'
1/
#627410000000
0!
1"
0'
1(
0/
10
#627420000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#627430000000
0!
0'
0/
#627440000000
1!
1'
1/
#627450000000
0!
0'
0/
#627460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#627470000000
0!
0'
0/
#627480000000
1!
1'
1/
#627490000000
0!
1"
0'
1(
0/
10
#627500000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#627510000000
0!
1$
0'
1+
0/
#627520000000
1!
1'
1/
#627530000000
0!
0'
0/
#627540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#627550000000
0!
0'
0/
#627560000000
1!
1'
1/
#627570000000
0!
0'
0/
#627580000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#627590000000
0!
0'
0/
#627600000000
1!
1'
1/
#627610000000
0!
0'
0/
#627620000000
1!
1'
1/
#627630000000
0!
0'
0/
#627640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#627650000000
0!
0'
0/
#627660000000
1!
1'
1/
#627670000000
0!
0'
0/
#627680000000
1!
1'
1/
#627690000000
0!
0'
0/
#627700000000
1!
1'
1/
#627710000000
0!
0'
0/
#627720000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#627730000000
0!
0'
0/
#627740000000
1!
1'
1/
#627750000000
0!
0'
0/
#627760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#627770000000
0!
0'
0/
#627780000000
1!
1'
1/
#627790000000
0!
0'
0/
#627800000000
#627810000000
1!
1'
1/
#627820000000
0!
0'
0/
#627830000000
1!
1'
1/
#627840000000
0!
1"
0'
1(
0/
10
#627850000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#627860000000
0!
0'
0/
#627870000000
1!
1'
1/
#627880000000
0!
0'
0/
#627890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#627900000000
0!
0'
0/
#627910000000
1!
1'
1/
#627920000000
0!
1"
0'
1(
0/
10
#627930000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#627940000000
0!
1$
0'
1+
0/
#627950000000
1!
1'
1/
#627960000000
0!
0'
0/
#627970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#627980000000
0!
0'
0/
#627990000000
1!
1'
1/
#628000000000
0!
0'
0/
#628010000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#628020000000
0!
0'
0/
#628030000000
1!
1'
1/
#628040000000
0!
0'
0/
#628050000000
1!
1'
1/
#628060000000
0!
0'
0/
#628070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#628080000000
0!
0'
0/
#628090000000
1!
1'
1/
#628100000000
0!
0'
0/
#628110000000
1!
1'
1/
#628120000000
0!
0'
0/
#628130000000
1!
1'
1/
#628140000000
0!
0'
0/
#628150000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#628160000000
0!
0'
0/
#628170000000
1!
1'
1/
#628180000000
0!
0'
0/
#628190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#628200000000
0!
0'
0/
#628210000000
1!
1'
1/
#628220000000
0!
0'
0/
#628230000000
#628240000000
1!
1'
1/
#628250000000
0!
0'
0/
#628260000000
1!
1'
1/
#628270000000
0!
1"
0'
1(
0/
10
#628280000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#628290000000
0!
0'
0/
#628300000000
1!
1'
1/
#628310000000
0!
0'
0/
#628320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#628330000000
0!
0'
0/
#628340000000
1!
1'
1/
#628350000000
0!
1"
0'
1(
0/
10
#628360000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#628370000000
0!
1$
0'
1+
0/
#628380000000
1!
1'
1/
#628390000000
0!
0'
0/
#628400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#628410000000
0!
0'
0/
#628420000000
1!
1'
1/
#628430000000
0!
0'
0/
#628440000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#628450000000
0!
0'
0/
#628460000000
1!
1'
1/
#628470000000
0!
0'
0/
#628480000000
1!
1'
1/
#628490000000
0!
0'
0/
#628500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#628510000000
0!
0'
0/
#628520000000
1!
1'
1/
#628530000000
0!
0'
0/
#628540000000
1!
1'
1/
#628550000000
0!
0'
0/
#628560000000
1!
1'
1/
#628570000000
0!
0'
0/
#628580000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#628590000000
0!
0'
0/
#628600000000
1!
1'
1/
#628610000000
0!
0'
0/
#628620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#628630000000
0!
0'
0/
#628640000000
1!
1'
1/
#628650000000
0!
0'
0/
#628660000000
#628670000000
1!
1'
1/
#628680000000
0!
0'
0/
#628690000000
1!
1'
1/
#628700000000
0!
1"
0'
1(
0/
10
#628710000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#628720000000
0!
0'
0/
#628730000000
1!
1'
1/
#628740000000
0!
0'
0/
#628750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#628760000000
0!
0'
0/
#628770000000
1!
1'
1/
#628780000000
0!
1"
0'
1(
0/
10
#628790000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#628800000000
0!
1$
0'
1+
0/
#628810000000
1!
1'
1/
#628820000000
0!
0'
0/
#628830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#628840000000
0!
0'
0/
#628850000000
1!
1'
1/
#628860000000
0!
0'
0/
#628870000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#628880000000
0!
0'
0/
#628890000000
1!
1'
1/
#628900000000
0!
0'
0/
#628910000000
1!
1'
1/
#628920000000
0!
0'
0/
#628930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#628940000000
0!
0'
0/
#628950000000
1!
1'
1/
#628960000000
0!
0'
0/
#628970000000
1!
1'
1/
#628980000000
0!
0'
0/
#628990000000
1!
1'
1/
#629000000000
0!
0'
0/
#629010000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#629020000000
0!
0'
0/
#629030000000
1!
1'
1/
#629040000000
0!
0'
0/
#629050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#629060000000
0!
0'
0/
#629070000000
1!
1'
1/
#629080000000
0!
0'
0/
#629090000000
#629100000000
1!
1'
1/
#629110000000
0!
0'
0/
#629120000000
1!
1'
1/
#629130000000
0!
1"
0'
1(
0/
10
#629140000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#629150000000
0!
0'
0/
#629160000000
1!
1'
1/
#629170000000
0!
0'
0/
#629180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#629190000000
0!
0'
0/
#629200000000
1!
1'
1/
#629210000000
0!
1"
0'
1(
0/
10
#629220000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#629230000000
0!
1$
0'
1+
0/
#629240000000
1!
1'
1/
#629250000000
0!
0'
0/
#629260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#629270000000
0!
0'
0/
#629280000000
1!
1'
1/
#629290000000
0!
0'
0/
#629300000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#629310000000
0!
0'
0/
#629320000000
1!
1'
1/
#629330000000
0!
0'
0/
#629340000000
1!
1'
1/
#629350000000
0!
0'
0/
#629360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#629370000000
0!
0'
0/
#629380000000
1!
1'
1/
#629390000000
0!
0'
0/
#629400000000
1!
1'
1/
#629410000000
0!
0'
0/
#629420000000
1!
1'
1/
#629430000000
0!
0'
0/
#629440000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#629450000000
0!
0'
0/
#629460000000
1!
1'
1/
#629470000000
0!
0'
0/
#629480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#629490000000
0!
0'
0/
#629500000000
1!
1'
1/
#629510000000
0!
0'
0/
#629520000000
#629530000000
1!
1'
1/
#629540000000
0!
0'
0/
#629550000000
1!
1'
1/
#629560000000
0!
1"
0'
1(
0/
10
#629570000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#629580000000
0!
0'
0/
#629590000000
1!
1'
1/
#629600000000
0!
0'
0/
#629610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#629620000000
0!
0'
0/
#629630000000
1!
1'
1/
#629640000000
0!
1"
0'
1(
0/
10
#629650000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#629660000000
0!
1$
0'
1+
0/
#629670000000
1!
1'
1/
#629680000000
0!
0'
0/
#629690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#629700000000
0!
0'
0/
#629710000000
1!
1'
1/
#629720000000
0!
0'
0/
#629730000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#629740000000
0!
0'
0/
#629750000000
1!
1'
1/
#629760000000
0!
0'
0/
#629770000000
1!
1'
1/
#629780000000
0!
0'
0/
#629790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#629800000000
0!
0'
0/
#629810000000
1!
1'
1/
#629820000000
0!
0'
0/
#629830000000
1!
1'
1/
#629840000000
0!
0'
0/
#629850000000
1!
1'
1/
#629860000000
0!
0'
0/
#629870000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#629880000000
0!
0'
0/
#629890000000
1!
1'
1/
#629900000000
0!
0'
0/
#629910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#629920000000
0!
0'
0/
#629930000000
1!
1'
1/
#629940000000
0!
0'
0/
#629950000000
#629960000000
1!
1'
1/
#629970000000
0!
0'
0/
#629980000000
1!
1'
1/
#629990000000
0!
1"
0'
1(
0/
10
#630000000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#630010000000
0!
0'
0/
#630020000000
1!
1'
1/
#630030000000
0!
0'
0/
#630040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#630050000000
0!
0'
0/
#630060000000
1!
1'
1/
#630070000000
0!
1"
0'
1(
0/
10
#630080000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#630090000000
0!
1$
0'
1+
0/
#630100000000
1!
1'
1/
#630110000000
0!
0'
0/
#630120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#630130000000
0!
0'
0/
#630140000000
1!
1'
1/
#630150000000
0!
0'
0/
#630160000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#630170000000
0!
0'
0/
#630180000000
1!
1'
1/
#630190000000
0!
0'
0/
#630200000000
1!
1'
1/
#630210000000
0!
0'
0/
#630220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#630230000000
0!
0'
0/
#630240000000
1!
1'
1/
#630250000000
0!
0'
0/
#630260000000
1!
1'
1/
#630270000000
0!
0'
0/
#630280000000
1!
1'
1/
#630290000000
0!
0'
0/
#630300000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#630310000000
0!
0'
0/
#630320000000
1!
1'
1/
#630330000000
0!
0'
0/
#630340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#630350000000
0!
0'
0/
#630360000000
1!
1'
1/
#630370000000
0!
0'
0/
#630380000000
#630390000000
1!
1'
1/
#630400000000
0!
0'
0/
#630410000000
1!
1'
1/
#630420000000
0!
1"
0'
1(
0/
10
#630430000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#630440000000
0!
0'
0/
#630450000000
1!
1'
1/
#630460000000
0!
0'
0/
#630470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#630480000000
0!
0'
0/
#630490000000
1!
1'
1/
#630500000000
0!
1"
0'
1(
0/
10
#630510000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#630520000000
0!
1$
0'
1+
0/
#630530000000
1!
1'
1/
#630540000000
0!
0'
0/
#630550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#630560000000
0!
0'
0/
#630570000000
1!
1'
1/
#630580000000
0!
0'
0/
#630590000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#630600000000
0!
0'
0/
#630610000000
1!
1'
1/
#630620000000
0!
0'
0/
#630630000000
1!
1'
1/
#630640000000
0!
0'
0/
#630650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#630660000000
0!
0'
0/
#630670000000
1!
1'
1/
#630680000000
0!
0'
0/
#630690000000
1!
1'
1/
#630700000000
0!
0'
0/
#630710000000
1!
1'
1/
#630720000000
0!
0'
0/
#630730000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#630740000000
0!
0'
0/
#630750000000
1!
1'
1/
#630760000000
0!
0'
0/
#630770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#630780000000
0!
0'
0/
#630790000000
1!
1'
1/
#630800000000
0!
0'
0/
#630810000000
#630820000000
1!
1'
1/
#630830000000
0!
0'
0/
#630840000000
1!
1'
1/
#630850000000
0!
1"
0'
1(
0/
10
#630860000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#630870000000
0!
0'
0/
#630880000000
1!
1'
1/
#630890000000
0!
0'
0/
#630900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#630910000000
0!
0'
0/
#630920000000
1!
1'
1/
#630930000000
0!
1"
0'
1(
0/
10
#630940000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#630950000000
0!
1$
0'
1+
0/
#630960000000
1!
1'
1/
#630970000000
0!
0'
0/
#630980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#630990000000
0!
0'
0/
#631000000000
1!
1'
1/
#631010000000
0!
0'
0/
#631020000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#631030000000
0!
0'
0/
#631040000000
1!
1'
1/
#631050000000
0!
0'
0/
#631060000000
1!
1'
1/
#631070000000
0!
0'
0/
#631080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#631090000000
0!
0'
0/
#631100000000
1!
1'
1/
#631110000000
0!
0'
0/
#631120000000
1!
1'
1/
#631130000000
0!
0'
0/
#631140000000
1!
1'
1/
#631150000000
0!
0'
0/
#631160000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#631170000000
0!
0'
0/
#631180000000
1!
1'
1/
#631190000000
0!
0'
0/
#631200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#631210000000
0!
0'
0/
#631220000000
1!
1'
1/
#631230000000
0!
0'
0/
#631240000000
#631250000000
1!
1'
1/
#631260000000
0!
0'
0/
#631270000000
1!
1'
1/
#631280000000
0!
1"
0'
1(
0/
10
#631290000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#631300000000
0!
0'
0/
#631310000000
1!
1'
1/
#631320000000
0!
0'
0/
#631330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#631340000000
0!
0'
0/
#631350000000
1!
1'
1/
#631360000000
0!
1"
0'
1(
0/
10
#631370000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#631380000000
0!
1$
0'
1+
0/
#631390000000
1!
1'
1/
#631400000000
0!
0'
0/
#631410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#631420000000
0!
0'
0/
#631430000000
1!
1'
1/
#631440000000
0!
0'
0/
#631450000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#631460000000
0!
0'
0/
#631470000000
1!
1'
1/
#631480000000
0!
0'
0/
#631490000000
1!
1'
1/
#631500000000
0!
0'
0/
#631510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#631520000000
0!
0'
0/
#631530000000
1!
1'
1/
#631540000000
0!
0'
0/
#631550000000
1!
1'
1/
#631560000000
0!
0'
0/
#631570000000
1!
1'
1/
#631580000000
0!
0'
0/
#631590000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#631600000000
0!
0'
0/
#631610000000
1!
1'
1/
#631620000000
0!
0'
0/
#631630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#631640000000
0!
0'
0/
#631650000000
1!
1'
1/
#631660000000
0!
0'
0/
#631670000000
#631680000000
1!
1'
1/
#631690000000
0!
0'
0/
#631700000000
1!
1'
1/
#631710000000
0!
1"
0'
1(
0/
10
#631720000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#631730000000
0!
0'
0/
#631740000000
1!
1'
1/
#631750000000
0!
0'
0/
#631760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#631770000000
0!
0'
0/
#631780000000
1!
1'
1/
#631790000000
0!
1"
0'
1(
0/
10
#631800000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#631810000000
0!
1$
0'
1+
0/
#631820000000
1!
1'
1/
#631830000000
0!
0'
0/
#631840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#631850000000
0!
0'
0/
#631860000000
1!
1'
1/
#631870000000
0!
0'
0/
#631880000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#631890000000
0!
0'
0/
#631900000000
1!
1'
1/
#631910000000
0!
0'
0/
#631920000000
1!
1'
1/
#631930000000
0!
0'
0/
#631940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#631950000000
0!
0'
0/
#631960000000
1!
1'
1/
#631970000000
0!
0'
0/
#631980000000
1!
1'
1/
#631990000000
0!
0'
0/
#632000000000
1!
1'
1/
#632010000000
0!
0'
0/
#632020000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#632030000000
0!
0'
0/
#632040000000
1!
1'
1/
#632050000000
0!
0'
0/
#632060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#632070000000
0!
0'
0/
#632080000000
1!
1'
1/
#632090000000
0!
0'
0/
#632100000000
#632110000000
1!
1'
1/
#632120000000
0!
0'
0/
#632130000000
1!
1'
1/
#632140000000
0!
1"
0'
1(
0/
10
#632150000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#632160000000
0!
0'
0/
#632170000000
1!
1'
1/
#632180000000
0!
0'
0/
#632190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#632200000000
0!
0'
0/
#632210000000
1!
1'
1/
#632220000000
0!
1"
0'
1(
0/
10
#632230000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#632240000000
0!
1$
0'
1+
0/
#632250000000
1!
1'
1/
#632260000000
0!
0'
0/
#632270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#632280000000
0!
0'
0/
#632290000000
1!
1'
1/
#632300000000
0!
0'
0/
#632310000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#632320000000
0!
0'
0/
#632330000000
1!
1'
1/
#632340000000
0!
0'
0/
#632350000000
1!
1'
1/
#632360000000
0!
0'
0/
#632370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#632380000000
0!
0'
0/
#632390000000
1!
1'
1/
#632400000000
0!
0'
0/
#632410000000
1!
1'
1/
#632420000000
0!
0'
0/
#632430000000
1!
1'
1/
#632440000000
0!
0'
0/
#632450000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#632460000000
0!
0'
0/
#632470000000
1!
1'
1/
#632480000000
0!
0'
0/
#632490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#632500000000
0!
0'
0/
#632510000000
1!
1'
1/
#632520000000
0!
0'
0/
#632530000000
#632540000000
1!
1'
1/
#632550000000
0!
0'
0/
#632560000000
1!
1'
1/
#632570000000
0!
1"
0'
1(
0/
10
#632580000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#632590000000
0!
0'
0/
#632600000000
1!
1'
1/
#632610000000
0!
0'
0/
#632620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#632630000000
0!
0'
0/
#632640000000
1!
1'
1/
#632650000000
0!
1"
0'
1(
0/
10
#632660000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#632670000000
0!
1$
0'
1+
0/
#632680000000
1!
1'
1/
#632690000000
0!
0'
0/
#632700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#632710000000
0!
0'
0/
#632720000000
1!
1'
1/
#632730000000
0!
0'
0/
#632740000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#632750000000
0!
0'
0/
#632760000000
1!
1'
1/
#632770000000
0!
0'
0/
#632780000000
1!
1'
1/
#632790000000
0!
0'
0/
#632800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#632810000000
0!
0'
0/
#632820000000
1!
1'
1/
#632830000000
0!
0'
0/
#632840000000
1!
1'
1/
#632850000000
0!
0'
0/
#632860000000
1!
1'
1/
#632870000000
0!
0'
0/
#632880000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#632890000000
0!
0'
0/
#632900000000
1!
1'
1/
#632910000000
0!
0'
0/
#632920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#632930000000
0!
0'
0/
#632940000000
1!
1'
1/
#632950000000
0!
0'
0/
#632960000000
#632970000000
1!
1'
1/
#632980000000
0!
0'
0/
#632990000000
1!
1'
1/
#633000000000
0!
1"
0'
1(
0/
10
#633010000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#633020000000
0!
0'
0/
#633030000000
1!
1'
1/
#633040000000
0!
0'
0/
#633050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#633060000000
0!
0'
0/
#633070000000
1!
1'
1/
#633080000000
0!
1"
0'
1(
0/
10
#633090000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#633100000000
0!
1$
0'
1+
0/
#633110000000
1!
1'
1/
#633120000000
0!
0'
0/
#633130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#633140000000
0!
0'
0/
#633150000000
1!
1'
1/
#633160000000
0!
0'
0/
#633170000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#633180000000
0!
0'
0/
#633190000000
1!
1'
1/
#633200000000
0!
0'
0/
#633210000000
1!
1'
1/
#633220000000
0!
0'
0/
#633230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#633240000000
0!
0'
0/
#633250000000
1!
1'
1/
#633260000000
0!
0'
0/
#633270000000
1!
1'
1/
#633280000000
0!
0'
0/
#633290000000
1!
1'
1/
#633300000000
0!
0'
0/
#633310000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#633320000000
0!
0'
0/
#633330000000
1!
1'
1/
#633340000000
0!
0'
0/
#633350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#633360000000
0!
0'
0/
#633370000000
1!
1'
1/
#633380000000
0!
0'
0/
#633390000000
#633400000000
1!
1'
1/
#633410000000
0!
0'
0/
#633420000000
1!
1'
1/
#633430000000
0!
1"
0'
1(
0/
10
#633440000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#633450000000
0!
0'
0/
#633460000000
1!
1'
1/
#633470000000
0!
0'
0/
#633480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#633490000000
0!
0'
0/
#633500000000
1!
1'
1/
#633510000000
0!
1"
0'
1(
0/
10
#633520000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#633530000000
0!
1$
0'
1+
0/
#633540000000
1!
1'
1/
#633550000000
0!
0'
0/
#633560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#633570000000
0!
0'
0/
#633580000000
1!
1'
1/
#633590000000
0!
0'
0/
#633600000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#633610000000
0!
0'
0/
#633620000000
1!
1'
1/
#633630000000
0!
0'
0/
#633640000000
1!
1'
1/
#633650000000
0!
0'
0/
#633660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#633670000000
0!
0'
0/
#633680000000
1!
1'
1/
#633690000000
0!
0'
0/
#633700000000
1!
1'
1/
#633710000000
0!
0'
0/
#633720000000
1!
1'
1/
#633730000000
0!
0'
0/
#633740000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#633750000000
0!
0'
0/
#633760000000
1!
1'
1/
#633770000000
0!
0'
0/
#633780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#633790000000
0!
0'
0/
#633800000000
1!
1'
1/
#633810000000
0!
0'
0/
#633820000000
#633830000000
1!
1'
1/
#633840000000
0!
0'
0/
#633850000000
1!
1'
1/
#633860000000
0!
1"
0'
1(
0/
10
#633870000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#633880000000
0!
0'
0/
#633890000000
1!
1'
1/
#633900000000
0!
0'
0/
#633910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#633920000000
0!
0'
0/
#633930000000
1!
1'
1/
#633940000000
0!
1"
0'
1(
0/
10
#633950000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#633960000000
0!
1$
0'
1+
0/
#633970000000
1!
1'
1/
#633980000000
0!
0'
0/
#633990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#634000000000
0!
0'
0/
#634010000000
1!
1'
1/
#634020000000
0!
0'
0/
#634030000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#634040000000
0!
0'
0/
#634050000000
1!
1'
1/
#634060000000
0!
0'
0/
#634070000000
1!
1'
1/
#634080000000
0!
0'
0/
#634090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#634100000000
0!
0'
0/
#634110000000
1!
1'
1/
#634120000000
0!
0'
0/
#634130000000
1!
1'
1/
#634140000000
0!
0'
0/
#634150000000
1!
1'
1/
#634160000000
0!
0'
0/
#634170000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#634180000000
0!
0'
0/
#634190000000
1!
1'
1/
#634200000000
0!
0'
0/
#634210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#634220000000
0!
0'
0/
#634230000000
1!
1'
1/
#634240000000
0!
0'
0/
#634250000000
#634260000000
1!
1'
1/
#634270000000
0!
0'
0/
#634280000000
1!
1'
1/
#634290000000
0!
1"
0'
1(
0/
10
#634300000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#634310000000
0!
0'
0/
#634320000000
1!
1'
1/
#634330000000
0!
0'
0/
#634340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#634350000000
0!
0'
0/
#634360000000
1!
1'
1/
#634370000000
0!
1"
0'
1(
0/
10
#634380000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#634390000000
0!
1$
0'
1+
0/
#634400000000
1!
1'
1/
#634410000000
0!
0'
0/
#634420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#634430000000
0!
0'
0/
#634440000000
1!
1'
1/
#634450000000
0!
0'
0/
#634460000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#634470000000
0!
0'
0/
#634480000000
1!
1'
1/
#634490000000
0!
0'
0/
#634500000000
1!
1'
1/
#634510000000
0!
0'
0/
#634520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#634530000000
0!
0'
0/
#634540000000
1!
1'
1/
#634550000000
0!
0'
0/
#634560000000
1!
1'
1/
#634570000000
0!
0'
0/
#634580000000
1!
1'
1/
#634590000000
0!
0'
0/
#634600000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#634610000000
0!
0'
0/
#634620000000
1!
1'
1/
#634630000000
0!
0'
0/
#634640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#634650000000
0!
0'
0/
#634660000000
1!
1'
1/
#634670000000
0!
0'
0/
#634680000000
#634690000000
1!
1'
1/
#634700000000
0!
0'
0/
#634710000000
1!
1'
1/
#634720000000
0!
1"
0'
1(
0/
10
#634730000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#634740000000
0!
0'
0/
#634750000000
1!
1'
1/
#634760000000
0!
0'
0/
#634770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#634780000000
0!
0'
0/
#634790000000
1!
1'
1/
#634800000000
0!
1"
0'
1(
0/
10
#634810000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#634820000000
0!
1$
0'
1+
0/
#634830000000
1!
1'
1/
#634840000000
0!
0'
0/
#634850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#634860000000
0!
0'
0/
#634870000000
1!
1'
1/
#634880000000
0!
0'
0/
#634890000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#634900000000
0!
0'
0/
#634910000000
1!
1'
1/
#634920000000
0!
0'
0/
#634930000000
1!
1'
1/
#634940000000
0!
0'
0/
#634950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#634960000000
0!
0'
0/
#634970000000
1!
1'
1/
#634980000000
0!
0'
0/
#634990000000
1!
1'
1/
#635000000000
0!
0'
0/
#635010000000
1!
1'
1/
#635020000000
0!
0'
0/
#635030000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#635040000000
0!
0'
0/
#635050000000
1!
1'
1/
#635060000000
0!
0'
0/
#635070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#635080000000
0!
0'
0/
#635090000000
1!
1'
1/
#635100000000
0!
0'
0/
#635110000000
#635120000000
1!
1'
1/
#635130000000
0!
0'
0/
#635140000000
1!
1'
1/
#635150000000
0!
1"
0'
1(
0/
10
#635160000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#635170000000
0!
0'
0/
#635180000000
1!
1'
1/
#635190000000
0!
0'
0/
#635200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#635210000000
0!
0'
0/
#635220000000
1!
1'
1/
#635230000000
0!
1"
0'
1(
0/
10
#635240000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#635250000000
0!
1$
0'
1+
0/
#635260000000
1!
1'
1/
#635270000000
0!
0'
0/
#635280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#635290000000
0!
0'
0/
#635300000000
1!
1'
1/
#635310000000
0!
0'
0/
#635320000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#635330000000
0!
0'
0/
#635340000000
1!
1'
1/
#635350000000
0!
0'
0/
#635360000000
1!
1'
1/
#635370000000
0!
0'
0/
#635380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#635390000000
0!
0'
0/
#635400000000
1!
1'
1/
#635410000000
0!
0'
0/
#635420000000
1!
1'
1/
#635430000000
0!
0'
0/
#635440000000
1!
1'
1/
#635450000000
0!
0'
0/
#635460000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#635470000000
0!
0'
0/
#635480000000
1!
1'
1/
#635490000000
0!
0'
0/
#635500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#635510000000
0!
0'
0/
#635520000000
1!
1'
1/
#635530000000
0!
0'
0/
#635540000000
#635550000000
1!
1'
1/
#635560000000
0!
0'
0/
#635570000000
1!
1'
1/
#635580000000
0!
1"
0'
1(
0/
10
#635590000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#635600000000
0!
0'
0/
#635610000000
1!
1'
1/
#635620000000
0!
0'
0/
#635630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#635640000000
0!
0'
0/
#635650000000
1!
1'
1/
#635660000000
0!
1"
0'
1(
0/
10
#635670000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#635680000000
0!
1$
0'
1+
0/
#635690000000
1!
1'
1/
#635700000000
0!
0'
0/
#635710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#635720000000
0!
0'
0/
#635730000000
1!
1'
1/
#635740000000
0!
0'
0/
#635750000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#635760000000
0!
0'
0/
#635770000000
1!
1'
1/
#635780000000
0!
0'
0/
#635790000000
1!
1'
1/
#635800000000
0!
0'
0/
#635810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#635820000000
0!
0'
0/
#635830000000
1!
1'
1/
#635840000000
0!
0'
0/
#635850000000
1!
1'
1/
#635860000000
0!
0'
0/
#635870000000
1!
1'
1/
#635880000000
0!
0'
0/
#635890000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#635900000000
0!
0'
0/
#635910000000
1!
1'
1/
#635920000000
0!
0'
0/
#635930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#635940000000
0!
0'
0/
#635950000000
1!
1'
1/
#635960000000
0!
0'
0/
#635970000000
#635980000000
1!
1'
1/
#635990000000
0!
0'
0/
#636000000000
1!
1'
1/
#636010000000
0!
1"
0'
1(
0/
10
#636020000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#636030000000
0!
0'
0/
#636040000000
1!
1'
1/
#636050000000
0!
0'
0/
#636060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#636070000000
0!
0'
0/
#636080000000
1!
1'
1/
#636090000000
0!
1"
0'
1(
0/
10
#636100000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#636110000000
0!
1$
0'
1+
0/
#636120000000
1!
1'
1/
#636130000000
0!
0'
0/
#636140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#636150000000
0!
0'
0/
#636160000000
1!
1'
1/
#636170000000
0!
0'
0/
#636180000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#636190000000
0!
0'
0/
#636200000000
1!
1'
1/
#636210000000
0!
0'
0/
#636220000000
1!
1'
1/
#636230000000
0!
0'
0/
#636240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#636250000000
0!
0'
0/
#636260000000
1!
1'
1/
#636270000000
0!
0'
0/
#636280000000
1!
1'
1/
#636290000000
0!
0'
0/
#636300000000
1!
1'
1/
#636310000000
0!
0'
0/
#636320000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#636330000000
0!
0'
0/
#636340000000
1!
1'
1/
#636350000000
0!
0'
0/
#636360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#636370000000
0!
0'
0/
#636380000000
1!
1'
1/
#636390000000
0!
0'
0/
#636400000000
#636410000000
1!
1'
1/
#636420000000
0!
0'
0/
#636430000000
1!
1'
1/
#636440000000
0!
1"
0'
1(
0/
10
#636450000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#636460000000
0!
0'
0/
#636470000000
1!
1'
1/
#636480000000
0!
0'
0/
#636490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#636500000000
0!
0'
0/
#636510000000
1!
1'
1/
#636520000000
0!
1"
0'
1(
0/
10
#636530000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#636540000000
0!
1$
0'
1+
0/
#636550000000
1!
1'
1/
#636560000000
0!
0'
0/
#636570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#636580000000
0!
0'
0/
#636590000000
1!
1'
1/
#636600000000
0!
0'
0/
#636610000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#636620000000
0!
0'
0/
#636630000000
1!
1'
1/
#636640000000
0!
0'
0/
#636650000000
1!
1'
1/
#636660000000
0!
0'
0/
#636670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#636680000000
0!
0'
0/
#636690000000
1!
1'
1/
#636700000000
0!
0'
0/
#636710000000
1!
1'
1/
#636720000000
0!
0'
0/
#636730000000
1!
1'
1/
#636740000000
0!
0'
0/
#636750000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#636760000000
0!
0'
0/
#636770000000
1!
1'
1/
#636780000000
0!
0'
0/
#636790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#636800000000
0!
0'
0/
#636810000000
1!
1'
1/
#636820000000
0!
0'
0/
#636830000000
#636840000000
1!
1'
1/
#636850000000
0!
0'
0/
#636860000000
1!
1'
1/
#636870000000
0!
1"
0'
1(
0/
10
#636880000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#636890000000
0!
0'
0/
#636900000000
1!
1'
1/
#636910000000
0!
0'
0/
#636920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#636930000000
0!
0'
0/
#636940000000
1!
1'
1/
#636950000000
0!
1"
0'
1(
0/
10
#636960000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#636970000000
0!
1$
0'
1+
0/
#636980000000
1!
1'
1/
#636990000000
0!
0'
0/
#637000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#637010000000
0!
0'
0/
#637020000000
1!
1'
1/
#637030000000
0!
0'
0/
#637040000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#637050000000
0!
0'
0/
#637060000000
1!
1'
1/
#637070000000
0!
0'
0/
#637080000000
1!
1'
1/
#637090000000
0!
0'
0/
#637100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#637110000000
0!
0'
0/
#637120000000
1!
1'
1/
#637130000000
0!
0'
0/
#637140000000
1!
1'
1/
#637150000000
0!
0'
0/
#637160000000
1!
1'
1/
#637170000000
0!
0'
0/
#637180000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#637190000000
0!
0'
0/
#637200000000
1!
1'
1/
#637210000000
0!
0'
0/
#637220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#637230000000
0!
0'
0/
#637240000000
1!
1'
1/
#637250000000
0!
0'
0/
#637260000000
#637270000000
1!
1'
1/
#637280000000
0!
0'
0/
#637290000000
1!
1'
1/
#637300000000
0!
1"
0'
1(
0/
10
#637310000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#637320000000
0!
0'
0/
#637330000000
1!
1'
1/
#637340000000
0!
0'
0/
#637350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#637360000000
0!
0'
0/
#637370000000
1!
1'
1/
#637380000000
0!
1"
0'
1(
0/
10
#637390000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#637400000000
0!
1$
0'
1+
0/
#637410000000
1!
1'
1/
#637420000000
0!
0'
0/
#637430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#637440000000
0!
0'
0/
#637450000000
1!
1'
1/
#637460000000
0!
0'
0/
#637470000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#637480000000
0!
0'
0/
#637490000000
1!
1'
1/
#637500000000
0!
0'
0/
#637510000000
1!
1'
1/
#637520000000
0!
0'
0/
#637530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#637540000000
0!
0'
0/
#637550000000
1!
1'
1/
#637560000000
0!
0'
0/
#637570000000
1!
1'
1/
#637580000000
0!
0'
0/
#637590000000
1!
1'
1/
#637600000000
0!
0'
0/
#637610000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#637620000000
0!
0'
0/
#637630000000
1!
1'
1/
#637640000000
0!
0'
0/
#637650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#637660000000
0!
0'
0/
#637670000000
1!
1'
1/
#637680000000
0!
0'
0/
#637690000000
#637700000000
1!
1'
1/
#637710000000
0!
0'
0/
#637720000000
1!
1'
1/
#637730000000
0!
1"
0'
1(
0/
10
#637740000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#637750000000
0!
0'
0/
#637760000000
1!
1'
1/
#637770000000
0!
0'
0/
#637780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#637790000000
0!
0'
0/
#637800000000
1!
1'
1/
#637810000000
0!
1"
0'
1(
0/
10
#637820000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#637830000000
0!
1$
0'
1+
0/
#637840000000
1!
1'
1/
#637850000000
0!
0'
0/
#637860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#637870000000
0!
0'
0/
#637880000000
1!
1'
1/
#637890000000
0!
0'
0/
#637900000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#637910000000
0!
0'
0/
#637920000000
1!
1'
1/
#637930000000
0!
0'
0/
#637940000000
1!
1'
1/
#637950000000
0!
0'
0/
#637960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#637970000000
0!
0'
0/
#637980000000
1!
1'
1/
#637990000000
0!
0'
0/
#638000000000
1!
1'
1/
#638010000000
0!
0'
0/
#638020000000
1!
1'
1/
#638030000000
0!
0'
0/
#638040000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#638050000000
0!
0'
0/
#638060000000
1!
1'
1/
#638070000000
0!
0'
0/
#638080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#638090000000
0!
0'
0/
#638100000000
1!
1'
1/
#638110000000
0!
0'
0/
#638120000000
#638130000000
1!
1'
1/
#638140000000
0!
0'
0/
#638150000000
1!
1'
1/
#638160000000
0!
1"
0'
1(
0/
10
#638170000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#638180000000
0!
0'
0/
#638190000000
1!
1'
1/
#638200000000
0!
0'
0/
#638210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#638220000000
0!
0'
0/
#638230000000
1!
1'
1/
#638240000000
0!
1"
0'
1(
0/
10
#638250000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#638260000000
0!
1$
0'
1+
0/
#638270000000
1!
1'
1/
#638280000000
0!
0'
0/
#638290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#638300000000
0!
0'
0/
#638310000000
1!
1'
1/
#638320000000
0!
0'
0/
#638330000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#638340000000
0!
0'
0/
#638350000000
1!
1'
1/
#638360000000
0!
0'
0/
#638370000000
1!
1'
1/
#638380000000
0!
0'
0/
#638390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#638400000000
0!
0'
0/
#638410000000
1!
1'
1/
#638420000000
0!
0'
0/
#638430000000
1!
1'
1/
#638440000000
0!
0'
0/
#638450000000
1!
1'
1/
#638460000000
0!
0'
0/
#638470000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#638480000000
0!
0'
0/
#638490000000
1!
1'
1/
#638500000000
0!
0'
0/
#638510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#638520000000
0!
0'
0/
#638530000000
1!
1'
1/
#638540000000
0!
0'
0/
#638550000000
#638560000000
1!
1'
1/
#638570000000
0!
0'
0/
#638580000000
1!
1'
1/
#638590000000
0!
1"
0'
1(
0/
10
#638600000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#638610000000
0!
0'
0/
#638620000000
1!
1'
1/
#638630000000
0!
0'
0/
#638640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#638650000000
0!
0'
0/
#638660000000
1!
1'
1/
#638670000000
0!
1"
0'
1(
0/
10
#638680000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#638690000000
0!
1$
0'
1+
0/
#638700000000
1!
1'
1/
#638710000000
0!
0'
0/
#638720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#638730000000
0!
0'
0/
#638740000000
1!
1'
1/
#638750000000
0!
0'
0/
#638760000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#638770000000
0!
0'
0/
#638780000000
1!
1'
1/
#638790000000
0!
0'
0/
#638800000000
1!
1'
1/
#638810000000
0!
0'
0/
#638820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#638830000000
0!
0'
0/
#638840000000
1!
1'
1/
#638850000000
0!
0'
0/
#638860000000
1!
1'
1/
#638870000000
0!
0'
0/
#638880000000
1!
1'
1/
#638890000000
0!
0'
0/
#638900000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#638910000000
0!
0'
0/
#638920000000
1!
1'
1/
#638930000000
0!
0'
0/
#638940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#638950000000
0!
0'
0/
#638960000000
1!
1'
1/
#638970000000
0!
0'
0/
#638980000000
#638990000000
1!
1'
1/
#639000000000
0!
0'
0/
#639010000000
1!
1'
1/
#639020000000
0!
1"
0'
1(
0/
10
#639030000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#639040000000
0!
0'
0/
#639050000000
1!
1'
1/
#639060000000
0!
0'
0/
#639070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#639080000000
0!
0'
0/
#639090000000
1!
1'
1/
#639100000000
0!
1"
0'
1(
0/
10
#639110000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#639120000000
0!
1$
0'
1+
0/
#639130000000
1!
1'
1/
#639140000000
0!
0'
0/
#639150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#639160000000
0!
0'
0/
#639170000000
1!
1'
1/
#639180000000
0!
0'
0/
#639190000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#639200000000
0!
0'
0/
#639210000000
1!
1'
1/
#639220000000
0!
0'
0/
#639230000000
1!
1'
1/
#639240000000
0!
0'
0/
#639250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#639260000000
0!
0'
0/
#639270000000
1!
1'
1/
#639280000000
0!
0'
0/
#639290000000
1!
1'
1/
#639300000000
0!
0'
0/
#639310000000
1!
1'
1/
#639320000000
0!
0'
0/
#639330000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#639340000000
0!
0'
0/
#639350000000
1!
1'
1/
#639360000000
0!
0'
0/
#639370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#639380000000
0!
0'
0/
#639390000000
1!
1'
1/
#639400000000
0!
0'
0/
#639410000000
#639420000000
1!
1'
1/
#639430000000
0!
0'
0/
#639440000000
1!
1'
1/
#639450000000
0!
1"
0'
1(
0/
10
#639460000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#639470000000
0!
0'
0/
#639480000000
1!
1'
1/
#639490000000
0!
0'
0/
#639500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#639510000000
0!
0'
0/
#639520000000
1!
1'
1/
#639530000000
0!
1"
0'
1(
0/
10
#639540000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#639550000000
0!
1$
0'
1+
0/
#639560000000
1!
1'
1/
#639570000000
0!
0'
0/
#639580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#639590000000
0!
0'
0/
#639600000000
1!
1'
1/
#639610000000
0!
0'
0/
#639620000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#639630000000
0!
0'
0/
#639640000000
1!
1'
1/
#639650000000
0!
0'
0/
#639660000000
1!
1'
1/
#639670000000
0!
0'
0/
#639680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#639690000000
0!
0'
0/
#639700000000
1!
1'
1/
#639710000000
0!
0'
0/
#639720000000
1!
1'
1/
#639730000000
0!
0'
0/
#639740000000
1!
1'
1/
#639750000000
0!
0'
0/
#639760000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#639770000000
0!
0'
0/
#639780000000
1!
1'
1/
#639790000000
0!
0'
0/
#639800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#639810000000
0!
0'
0/
#639820000000
1!
1'
1/
#639830000000
0!
0'
0/
#639840000000
#639850000000
1!
1'
1/
#639860000000
0!
0'
0/
#639870000000
1!
1'
1/
#639880000000
0!
1"
0'
1(
0/
10
#639890000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#639900000000
0!
0'
0/
#639910000000
1!
1'
1/
#639920000000
0!
0'
0/
#639930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#639940000000
0!
0'
0/
#639950000000
1!
1'
1/
#639960000000
0!
1"
0'
1(
0/
10
#639970000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#639980000000
0!
1$
0'
1+
0/
#639990000000
1!
1'
1/
#640000000000
0!
0'
0/
#640010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#640020000000
0!
0'
0/
#640030000000
1!
1'
1/
#640040000000
0!
0'
0/
#640050000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#640060000000
0!
0'
0/
#640070000000
1!
1'
1/
#640080000000
0!
0'
0/
#640090000000
1!
1'
1/
#640100000000
0!
0'
0/
#640110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#640120000000
0!
0'
0/
#640130000000
1!
1'
1/
#640140000000
0!
0'
0/
#640150000000
1!
1'
1/
#640160000000
0!
0'
0/
#640170000000
1!
1'
1/
#640180000000
0!
0'
0/
#640190000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#640200000000
0!
0'
0/
#640210000000
1!
1'
1/
#640220000000
0!
0'
0/
#640230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#640240000000
0!
0'
0/
#640250000000
1!
1'
1/
#640260000000
0!
0'
0/
#640270000000
#640280000000
1!
1'
1/
#640290000000
0!
0'
0/
#640300000000
1!
1'
1/
#640310000000
0!
1"
0'
1(
0/
10
#640320000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#640330000000
0!
0'
0/
#640340000000
1!
1'
1/
#640350000000
0!
0'
0/
#640360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#640370000000
0!
0'
0/
#640380000000
1!
1'
1/
#640390000000
0!
1"
0'
1(
0/
10
#640400000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#640410000000
0!
1$
0'
1+
0/
#640420000000
1!
1'
1/
#640430000000
0!
0'
0/
#640440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#640450000000
0!
0'
0/
#640460000000
1!
1'
1/
#640470000000
0!
0'
0/
#640480000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#640490000000
0!
0'
0/
#640500000000
1!
1'
1/
#640510000000
0!
0'
0/
#640520000000
1!
1'
1/
#640530000000
0!
0'
0/
#640540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#640550000000
0!
0'
0/
#640560000000
1!
1'
1/
#640570000000
0!
0'
0/
#640580000000
1!
1'
1/
#640590000000
0!
0'
0/
#640600000000
1!
1'
1/
#640610000000
0!
0'
0/
#640620000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#640630000000
0!
0'
0/
#640640000000
1!
1'
1/
#640650000000
0!
0'
0/
#640660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#640670000000
0!
0'
0/
#640680000000
1!
1'
1/
#640690000000
0!
0'
0/
#640700000000
#640710000000
1!
1'
1/
#640720000000
0!
0'
0/
#640730000000
1!
1'
1/
#640740000000
0!
1"
0'
1(
0/
10
#640750000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#640760000000
0!
0'
0/
#640770000000
1!
1'
1/
#640780000000
0!
0'
0/
#640790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#640800000000
0!
0'
0/
#640810000000
1!
1'
1/
#640820000000
0!
1"
0'
1(
0/
10
#640830000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#640840000000
0!
1$
0'
1+
0/
#640850000000
1!
1'
1/
#640860000000
0!
0'
0/
#640870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#640880000000
0!
0'
0/
#640890000000
1!
1'
1/
#640900000000
0!
0'
0/
#640910000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#640920000000
0!
0'
0/
#640930000000
1!
1'
1/
#640940000000
0!
0'
0/
#640950000000
1!
1'
1/
#640960000000
0!
0'
0/
#640970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#640980000000
0!
0'
0/
#640990000000
1!
1'
1/
#641000000000
0!
0'
0/
#641010000000
1!
1'
1/
#641020000000
0!
0'
0/
#641030000000
1!
1'
1/
#641040000000
0!
0'
0/
#641050000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#641060000000
0!
0'
0/
#641070000000
1!
1'
1/
#641080000000
0!
0'
0/
#641090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#641100000000
0!
0'
0/
#641110000000
1!
1'
1/
#641120000000
0!
0'
0/
#641130000000
#641140000000
1!
1'
1/
#641150000000
0!
0'
0/
#641160000000
1!
1'
1/
#641170000000
0!
1"
0'
1(
0/
10
#641180000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#641190000000
0!
0'
0/
#641200000000
1!
1'
1/
#641210000000
0!
0'
0/
#641220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#641230000000
0!
0'
0/
#641240000000
1!
1'
1/
#641250000000
0!
1"
0'
1(
0/
10
#641260000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#641270000000
0!
1$
0'
1+
0/
#641280000000
1!
1'
1/
#641290000000
0!
0'
0/
#641300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#641310000000
0!
0'
0/
#641320000000
1!
1'
1/
#641330000000
0!
0'
0/
#641340000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#641350000000
0!
0'
0/
#641360000000
1!
1'
1/
#641370000000
0!
0'
0/
#641380000000
1!
1'
1/
#641390000000
0!
0'
0/
#641400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#641410000000
0!
0'
0/
#641420000000
1!
1'
1/
#641430000000
0!
0'
0/
#641440000000
1!
1'
1/
#641450000000
0!
0'
0/
#641460000000
1!
1'
1/
#641470000000
0!
0'
0/
#641480000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#641490000000
0!
0'
0/
#641500000000
1!
1'
1/
#641510000000
0!
0'
0/
#641520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#641530000000
0!
0'
0/
#641540000000
1!
1'
1/
#641550000000
0!
0'
0/
#641560000000
#641570000000
1!
1'
1/
#641580000000
0!
0'
0/
#641590000000
1!
1'
1/
#641600000000
0!
1"
0'
1(
0/
10
#641610000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#641620000000
0!
0'
0/
#641630000000
1!
1'
1/
#641640000000
0!
0'
0/
#641650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#641660000000
0!
0'
0/
#641670000000
1!
1'
1/
#641680000000
0!
1"
0'
1(
0/
10
#641690000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#641700000000
0!
1$
0'
1+
0/
#641710000000
1!
1'
1/
#641720000000
0!
0'
0/
#641730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#641740000000
0!
0'
0/
#641750000000
1!
1'
1/
#641760000000
0!
0'
0/
#641770000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#641780000000
0!
0'
0/
#641790000000
1!
1'
1/
#641800000000
0!
0'
0/
#641810000000
1!
1'
1/
#641820000000
0!
0'
0/
#641830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#641840000000
0!
0'
0/
#641850000000
1!
1'
1/
#641860000000
0!
0'
0/
#641870000000
1!
1'
1/
#641880000000
0!
0'
0/
#641890000000
1!
1'
1/
#641900000000
0!
0'
0/
#641910000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#641920000000
0!
0'
0/
#641930000000
1!
1'
1/
#641940000000
0!
0'
0/
#641950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#641960000000
0!
0'
0/
#641970000000
1!
1'
1/
#641980000000
0!
0'
0/
#641990000000
#642000000000
1!
1'
1/
#642010000000
0!
0'
0/
#642020000000
1!
1'
1/
#642030000000
0!
1"
0'
1(
0/
10
#642040000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#642050000000
0!
0'
0/
#642060000000
1!
1'
1/
#642070000000
0!
0'
0/
#642080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#642090000000
0!
0'
0/
#642100000000
1!
1'
1/
#642110000000
0!
1"
0'
1(
0/
10
#642120000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#642130000000
0!
1$
0'
1+
0/
#642140000000
1!
1'
1/
#642150000000
0!
0'
0/
#642160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#642170000000
0!
0'
0/
#642180000000
1!
1'
1/
#642190000000
0!
0'
0/
#642200000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#642210000000
0!
0'
0/
#642220000000
1!
1'
1/
#642230000000
0!
0'
0/
#642240000000
1!
1'
1/
#642250000000
0!
0'
0/
#642260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#642270000000
0!
0'
0/
#642280000000
1!
1'
1/
#642290000000
0!
0'
0/
#642300000000
1!
1'
1/
#642310000000
0!
0'
0/
#642320000000
1!
1'
1/
#642330000000
0!
0'
0/
#642340000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#642350000000
0!
0'
0/
#642360000000
1!
1'
1/
#642370000000
0!
0'
0/
#642380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#642390000000
0!
0'
0/
#642400000000
1!
1'
1/
#642410000000
0!
0'
0/
#642420000000
#642430000000
1!
1'
1/
#642440000000
0!
0'
0/
#642450000000
1!
1'
1/
#642460000000
0!
1"
0'
1(
0/
10
#642470000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#642480000000
0!
0'
0/
#642490000000
1!
1'
1/
#642500000000
0!
0'
0/
#642510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#642520000000
0!
0'
0/
#642530000000
1!
1'
1/
#642540000000
0!
1"
0'
1(
0/
10
#642550000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#642560000000
0!
1$
0'
1+
0/
#642570000000
1!
1'
1/
#642580000000
0!
0'
0/
#642590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#642600000000
0!
0'
0/
#642610000000
1!
1'
1/
#642620000000
0!
0'
0/
#642630000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#642640000000
0!
0'
0/
#642650000000
1!
1'
1/
#642660000000
0!
0'
0/
#642670000000
1!
1'
1/
#642680000000
0!
0'
0/
#642690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#642700000000
0!
0'
0/
#642710000000
1!
1'
1/
#642720000000
0!
0'
0/
#642730000000
1!
1'
1/
#642740000000
0!
0'
0/
#642750000000
1!
1'
1/
#642760000000
0!
0'
0/
#642770000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#642780000000
0!
0'
0/
#642790000000
1!
1'
1/
#642800000000
0!
0'
0/
#642810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#642820000000
0!
0'
0/
#642830000000
1!
1'
1/
#642840000000
0!
0'
0/
#642850000000
#642860000000
1!
1'
1/
#642870000000
0!
0'
0/
#642880000000
1!
1'
1/
#642890000000
0!
1"
0'
1(
0/
10
#642900000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#642910000000
0!
0'
0/
#642920000000
1!
1'
1/
#642930000000
0!
0'
0/
#642940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#642950000000
0!
0'
0/
#642960000000
1!
1'
1/
#642970000000
0!
1"
0'
1(
0/
10
#642980000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#642990000000
0!
1$
0'
1+
0/
#643000000000
1!
1'
1/
#643010000000
0!
0'
0/
#643020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#643030000000
0!
0'
0/
#643040000000
1!
1'
1/
#643050000000
0!
0'
0/
#643060000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#643070000000
0!
0'
0/
#643080000000
1!
1'
1/
#643090000000
0!
0'
0/
#643100000000
1!
1'
1/
#643110000000
0!
0'
0/
#643120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#643130000000
0!
0'
0/
#643140000000
1!
1'
1/
#643150000000
0!
0'
0/
#643160000000
1!
1'
1/
#643170000000
0!
0'
0/
#643180000000
1!
1'
1/
#643190000000
0!
0'
0/
#643200000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#643210000000
0!
0'
0/
#643220000000
1!
1'
1/
#643230000000
0!
0'
0/
#643240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#643250000000
0!
0'
0/
#643260000000
1!
1'
1/
#643270000000
0!
0'
0/
#643280000000
#643290000000
1!
1'
1/
#643300000000
0!
0'
0/
#643310000000
1!
1'
1/
#643320000000
0!
1"
0'
1(
0/
10
#643330000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#643340000000
0!
0'
0/
#643350000000
1!
1'
1/
#643360000000
0!
0'
0/
#643370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#643380000000
0!
0'
0/
#643390000000
1!
1'
1/
#643400000000
0!
1"
0'
1(
0/
10
#643410000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#643420000000
0!
1$
0'
1+
0/
#643430000000
1!
1'
1/
#643440000000
0!
0'
0/
#643450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#643460000000
0!
0'
0/
#643470000000
1!
1'
1/
#643480000000
0!
0'
0/
#643490000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#643500000000
0!
0'
0/
#643510000000
1!
1'
1/
#643520000000
0!
0'
0/
#643530000000
1!
1'
1/
#643540000000
0!
0'
0/
#643550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#643560000000
0!
0'
0/
#643570000000
1!
1'
1/
#643580000000
0!
0'
0/
#643590000000
1!
1'
1/
#643600000000
0!
0'
0/
#643610000000
1!
1'
1/
#643620000000
0!
0'
0/
#643630000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#643640000000
0!
0'
0/
#643650000000
1!
1'
1/
#643660000000
0!
0'
0/
#643670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#643680000000
0!
0'
0/
#643690000000
1!
1'
1/
#643700000000
0!
0'
0/
#643710000000
#643720000000
1!
1'
1/
#643730000000
0!
0'
0/
#643740000000
1!
1'
1/
#643750000000
0!
1"
0'
1(
0/
10
#643760000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#643770000000
0!
0'
0/
#643780000000
1!
1'
1/
#643790000000
0!
0'
0/
#643800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#643810000000
0!
0'
0/
#643820000000
1!
1'
1/
#643830000000
0!
1"
0'
1(
0/
10
#643840000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#643850000000
0!
1$
0'
1+
0/
#643860000000
1!
1'
1/
#643870000000
0!
0'
0/
#643880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#643890000000
0!
0'
0/
#643900000000
1!
1'
1/
#643910000000
0!
0'
0/
#643920000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#643930000000
0!
0'
0/
#643940000000
1!
1'
1/
#643950000000
0!
0'
0/
#643960000000
1!
1'
1/
#643970000000
0!
0'
0/
#643980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#643990000000
0!
0'
0/
#644000000000
1!
1'
1/
#644010000000
0!
0'
0/
#644020000000
1!
1'
1/
#644030000000
0!
0'
0/
#644040000000
1!
1'
1/
#644050000000
0!
0'
0/
#644060000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#644070000000
0!
0'
0/
#644080000000
1!
1'
1/
#644090000000
0!
0'
0/
#644100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#644110000000
0!
0'
0/
#644120000000
1!
1'
1/
#644130000000
0!
0'
0/
#644140000000
#644150000000
1!
1'
1/
#644160000000
0!
0'
0/
#644170000000
1!
1'
1/
#644180000000
0!
1"
0'
1(
0/
10
#644190000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#644200000000
0!
0'
0/
#644210000000
1!
1'
1/
#644220000000
0!
0'
0/
#644230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#644240000000
0!
0'
0/
#644250000000
1!
1'
1/
#644260000000
0!
1"
0'
1(
0/
10
#644270000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#644280000000
0!
1$
0'
1+
0/
#644290000000
1!
1'
1/
#644300000000
0!
0'
0/
#644310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#644320000000
0!
0'
0/
#644330000000
1!
1'
1/
#644340000000
0!
0'
0/
#644350000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#644360000000
0!
0'
0/
#644370000000
1!
1'
1/
#644380000000
0!
0'
0/
#644390000000
1!
1'
1/
#644400000000
0!
0'
0/
#644410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#644420000000
0!
0'
0/
#644430000000
1!
1'
1/
#644440000000
0!
0'
0/
#644450000000
1!
1'
1/
#644460000000
0!
0'
0/
#644470000000
1!
1'
1/
#644480000000
0!
0'
0/
#644490000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#644500000000
0!
0'
0/
#644510000000
1!
1'
1/
#644520000000
0!
0'
0/
#644530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#644540000000
0!
0'
0/
#644550000000
1!
1'
1/
#644560000000
0!
0'
0/
#644570000000
#644580000000
1!
1'
1/
#644590000000
0!
0'
0/
#644600000000
1!
1'
1/
#644610000000
0!
1"
0'
1(
0/
10
#644620000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#644630000000
0!
0'
0/
#644640000000
1!
1'
1/
#644650000000
0!
0'
0/
#644660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#644670000000
0!
0'
0/
#644680000000
1!
1'
1/
#644690000000
0!
1"
0'
1(
0/
10
#644700000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#644710000000
0!
1$
0'
1+
0/
#644720000000
1!
1'
1/
#644730000000
0!
0'
0/
#644740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#644750000000
0!
0'
0/
#644760000000
1!
1'
1/
#644770000000
0!
0'
0/
#644780000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#644790000000
0!
0'
0/
#644800000000
1!
1'
1/
#644810000000
0!
0'
0/
#644820000000
1!
1'
1/
#644830000000
0!
0'
0/
#644840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#644850000000
0!
0'
0/
#644860000000
1!
1'
1/
#644870000000
0!
0'
0/
#644880000000
1!
1'
1/
#644890000000
0!
0'
0/
#644900000000
1!
1'
1/
#644910000000
0!
0'
0/
#644920000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#644930000000
0!
0'
0/
#644940000000
1!
1'
1/
#644950000000
0!
0'
0/
#644960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#644970000000
0!
0'
0/
#644980000000
1!
1'
1/
#644990000000
0!
0'
0/
#645000000000
#645010000000
1!
1'
1/
#645020000000
0!
0'
0/
#645030000000
1!
1'
1/
#645040000000
0!
1"
0'
1(
0/
10
#645050000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#645060000000
0!
0'
0/
#645070000000
1!
1'
1/
#645080000000
0!
0'
0/
#645090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#645100000000
0!
0'
0/
#645110000000
1!
1'
1/
#645120000000
0!
1"
0'
1(
0/
10
#645130000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#645140000000
0!
1$
0'
1+
0/
#645150000000
1!
1'
1/
#645160000000
0!
0'
0/
#645170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#645180000000
0!
0'
0/
#645190000000
1!
1'
1/
#645200000000
0!
0'
0/
#645210000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#645220000000
0!
0'
0/
#645230000000
1!
1'
1/
#645240000000
0!
0'
0/
#645250000000
1!
1'
1/
#645260000000
0!
0'
0/
#645270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#645280000000
0!
0'
0/
#645290000000
1!
1'
1/
#645300000000
0!
0'
0/
#645310000000
1!
1'
1/
#645320000000
0!
0'
0/
#645330000000
1!
1'
1/
#645340000000
0!
0'
0/
#645350000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#645360000000
0!
0'
0/
#645370000000
1!
1'
1/
#645380000000
0!
0'
0/
#645390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#645400000000
0!
0'
0/
#645410000000
1!
1'
1/
#645420000000
0!
0'
0/
#645430000000
#645440000000
1!
1'
1/
#645450000000
0!
0'
0/
#645460000000
1!
1'
1/
#645470000000
0!
1"
0'
1(
0/
10
#645480000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#645490000000
0!
0'
0/
#645500000000
1!
1'
1/
#645510000000
0!
0'
0/
#645520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#645530000000
0!
0'
0/
#645540000000
1!
1'
1/
#645550000000
0!
1"
0'
1(
0/
10
#645560000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#645570000000
0!
1$
0'
1+
0/
#645580000000
1!
1'
1/
#645590000000
0!
0'
0/
#645600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#645610000000
0!
0'
0/
#645620000000
1!
1'
1/
#645630000000
0!
0'
0/
#645640000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#645650000000
0!
0'
0/
#645660000000
1!
1'
1/
#645670000000
0!
0'
0/
#645680000000
1!
1'
1/
#645690000000
0!
0'
0/
#645700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#645710000000
0!
0'
0/
#645720000000
1!
1'
1/
#645730000000
0!
0'
0/
#645740000000
1!
1'
1/
#645750000000
0!
0'
0/
#645760000000
1!
1'
1/
#645770000000
0!
0'
0/
#645780000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#645790000000
0!
0'
0/
#645800000000
1!
1'
1/
#645810000000
0!
0'
0/
#645820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#645830000000
0!
0'
0/
#645840000000
1!
1'
1/
#645850000000
0!
0'
0/
#645860000000
#645870000000
1!
1'
1/
#645880000000
0!
0'
0/
#645890000000
1!
1'
1/
#645900000000
0!
1"
0'
1(
0/
10
#645910000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#645920000000
0!
0'
0/
#645930000000
1!
1'
1/
#645940000000
0!
0'
0/
#645950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#645960000000
0!
0'
0/
#645970000000
1!
1'
1/
#645980000000
0!
1"
0'
1(
0/
10
#645990000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#646000000000
0!
1$
0'
1+
0/
#646010000000
1!
1'
1/
#646020000000
0!
0'
0/
#646030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#646040000000
0!
0'
0/
#646050000000
1!
1'
1/
#646060000000
0!
0'
0/
#646070000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#646080000000
0!
0'
0/
#646090000000
1!
1'
1/
#646100000000
0!
0'
0/
#646110000000
1!
1'
1/
#646120000000
0!
0'
0/
#646130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#646140000000
0!
0'
0/
#646150000000
1!
1'
1/
#646160000000
0!
0'
0/
#646170000000
1!
1'
1/
#646180000000
0!
0'
0/
#646190000000
1!
1'
1/
#646200000000
0!
0'
0/
#646210000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#646220000000
0!
0'
0/
#646230000000
1!
1'
1/
#646240000000
0!
0'
0/
#646250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#646260000000
0!
0'
0/
#646270000000
1!
1'
1/
#646280000000
0!
0'
0/
#646290000000
#646300000000
1!
1'
1/
#646310000000
0!
0'
0/
#646320000000
1!
1'
1/
#646330000000
0!
1"
0'
1(
0/
10
#646340000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#646350000000
0!
0'
0/
#646360000000
1!
1'
1/
#646370000000
0!
0'
0/
#646380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#646390000000
0!
0'
0/
#646400000000
1!
1'
1/
#646410000000
0!
1"
0'
1(
0/
10
#646420000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#646430000000
0!
1$
0'
1+
0/
#646440000000
1!
1'
1/
#646450000000
0!
0'
0/
#646460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#646470000000
0!
0'
0/
#646480000000
1!
1'
1/
#646490000000
0!
0'
0/
#646500000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#646510000000
0!
0'
0/
#646520000000
1!
1'
1/
#646530000000
0!
0'
0/
#646540000000
1!
1'
1/
#646550000000
0!
0'
0/
#646560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#646570000000
0!
0'
0/
#646580000000
1!
1'
1/
#646590000000
0!
0'
0/
#646600000000
1!
1'
1/
#646610000000
0!
0'
0/
#646620000000
1!
1'
1/
#646630000000
0!
0'
0/
#646640000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#646650000000
0!
0'
0/
#646660000000
1!
1'
1/
#646670000000
0!
0'
0/
#646680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#646690000000
0!
0'
0/
#646700000000
1!
1'
1/
#646710000000
0!
0'
0/
#646720000000
#646730000000
1!
1'
1/
#646740000000
0!
0'
0/
#646750000000
1!
1'
1/
#646760000000
0!
1"
0'
1(
0/
10
#646770000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#646780000000
0!
0'
0/
#646790000000
1!
1'
1/
#646800000000
0!
0'
0/
#646810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#646820000000
0!
0'
0/
#646830000000
1!
1'
1/
#646840000000
0!
1"
0'
1(
0/
10
#646850000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#646860000000
0!
1$
0'
1+
0/
#646870000000
1!
1'
1/
#646880000000
0!
0'
0/
#646890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#646900000000
0!
0'
0/
#646910000000
1!
1'
1/
#646920000000
0!
0'
0/
#646930000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#646940000000
0!
0'
0/
#646950000000
1!
1'
1/
#646960000000
0!
0'
0/
#646970000000
1!
1'
1/
#646980000000
0!
0'
0/
#646990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#647000000000
0!
0'
0/
#647010000000
1!
1'
1/
#647020000000
0!
0'
0/
#647030000000
1!
1'
1/
#647040000000
0!
0'
0/
#647050000000
1!
1'
1/
#647060000000
0!
0'
0/
#647070000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#647080000000
0!
0'
0/
#647090000000
1!
1'
1/
#647100000000
0!
0'
0/
#647110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#647120000000
0!
0'
0/
#647130000000
1!
1'
1/
#647140000000
0!
0'
0/
#647150000000
#647160000000
1!
1'
1/
#647170000000
0!
0'
0/
#647180000000
1!
1'
1/
#647190000000
0!
1"
0'
1(
0/
10
#647200000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#647210000000
0!
0'
0/
#647220000000
1!
1'
1/
#647230000000
0!
0'
0/
#647240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#647250000000
0!
0'
0/
#647260000000
1!
1'
1/
#647270000000
0!
1"
0'
1(
0/
10
#647280000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#647290000000
0!
1$
0'
1+
0/
#647300000000
1!
1'
1/
#647310000000
0!
0'
0/
#647320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#647330000000
0!
0'
0/
#647340000000
1!
1'
1/
#647350000000
0!
0'
0/
#647360000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#647370000000
0!
0'
0/
#647380000000
1!
1'
1/
#647390000000
0!
0'
0/
#647400000000
1!
1'
1/
#647410000000
0!
0'
0/
#647420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#647430000000
0!
0'
0/
#647440000000
1!
1'
1/
#647450000000
0!
0'
0/
#647460000000
1!
1'
1/
#647470000000
0!
0'
0/
#647480000000
1!
1'
1/
#647490000000
0!
0'
0/
#647500000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#647510000000
0!
0'
0/
#647520000000
1!
1'
1/
#647530000000
0!
0'
0/
#647540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#647550000000
0!
0'
0/
#647560000000
1!
1'
1/
#647570000000
0!
0'
0/
#647580000000
#647590000000
1!
1'
1/
#647600000000
0!
0'
0/
#647610000000
1!
1'
1/
#647620000000
0!
1"
0'
1(
0/
10
#647630000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#647640000000
0!
0'
0/
#647650000000
1!
1'
1/
#647660000000
0!
0'
0/
#647670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#647680000000
0!
0'
0/
#647690000000
1!
1'
1/
#647700000000
0!
1"
0'
1(
0/
10
#647710000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#647720000000
0!
1$
0'
1+
0/
#647730000000
1!
1'
1/
#647740000000
0!
0'
0/
#647750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#647760000000
0!
0'
0/
#647770000000
1!
1'
1/
#647780000000
0!
0'
0/
#647790000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#647800000000
0!
0'
0/
#647810000000
1!
1'
1/
#647820000000
0!
0'
0/
#647830000000
1!
1'
1/
#647840000000
0!
0'
0/
#647850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#647860000000
0!
0'
0/
#647870000000
1!
1'
1/
#647880000000
0!
0'
0/
#647890000000
1!
1'
1/
#647900000000
0!
0'
0/
#647910000000
1!
1'
1/
#647920000000
0!
0'
0/
#647930000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#647940000000
0!
0'
0/
#647950000000
1!
1'
1/
#647960000000
0!
0'
0/
#647970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#647980000000
0!
0'
0/
#647990000000
1!
1'
1/
#648000000000
0!
0'
0/
#648010000000
#648020000000
1!
1'
1/
#648030000000
0!
0'
0/
#648040000000
1!
1'
1/
#648050000000
0!
1"
0'
1(
0/
10
#648060000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#648070000000
0!
0'
0/
#648080000000
1!
1'
1/
#648090000000
0!
0'
0/
#648100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#648110000000
0!
0'
0/
#648120000000
1!
1'
1/
#648130000000
0!
1"
0'
1(
0/
10
#648140000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#648150000000
0!
1$
0'
1+
0/
#648160000000
1!
1'
1/
#648170000000
0!
0'
0/
#648180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#648190000000
0!
0'
0/
#648200000000
1!
1'
1/
#648210000000
0!
0'
0/
#648220000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#648230000000
0!
0'
0/
#648240000000
1!
1'
1/
#648250000000
0!
0'
0/
#648260000000
1!
1'
1/
#648270000000
0!
0'
0/
#648280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#648290000000
0!
0'
0/
#648300000000
1!
1'
1/
#648310000000
0!
0'
0/
#648320000000
1!
1'
1/
#648330000000
0!
0'
0/
#648340000000
1!
1'
1/
#648350000000
0!
0'
0/
#648360000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#648370000000
0!
0'
0/
#648380000000
1!
1'
1/
#648390000000
0!
0'
0/
#648400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#648410000000
0!
0'
0/
#648420000000
1!
1'
1/
#648430000000
0!
0'
0/
#648440000000
#648450000000
1!
1'
1/
#648460000000
0!
0'
0/
#648470000000
1!
1'
1/
#648480000000
0!
1"
0'
1(
0/
10
#648490000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#648500000000
0!
0'
0/
#648510000000
1!
1'
1/
#648520000000
0!
0'
0/
#648530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#648540000000
0!
0'
0/
#648550000000
1!
1'
1/
#648560000000
0!
1"
0'
1(
0/
10
#648570000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#648580000000
0!
1$
0'
1+
0/
#648590000000
1!
1'
1/
#648600000000
0!
0'
0/
#648610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#648620000000
0!
0'
0/
#648630000000
1!
1'
1/
#648640000000
0!
0'
0/
#648650000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#648660000000
0!
0'
0/
#648670000000
1!
1'
1/
#648680000000
0!
0'
0/
#648690000000
1!
1'
1/
#648700000000
0!
0'
0/
#648710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#648720000000
0!
0'
0/
#648730000000
1!
1'
1/
#648740000000
0!
0'
0/
#648750000000
1!
1'
1/
#648760000000
0!
0'
0/
#648770000000
1!
1'
1/
#648780000000
0!
0'
0/
#648790000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#648800000000
0!
0'
0/
#648810000000
1!
1'
1/
#648820000000
0!
0'
0/
#648830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#648840000000
0!
0'
0/
#648850000000
1!
1'
1/
#648860000000
0!
0'
0/
#648870000000
#648880000000
1!
1'
1/
#648890000000
0!
0'
0/
#648900000000
1!
1'
1/
#648910000000
0!
1"
0'
1(
0/
10
#648920000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#648930000000
0!
0'
0/
#648940000000
1!
1'
1/
#648950000000
0!
0'
0/
#648960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#648970000000
0!
0'
0/
#648980000000
1!
1'
1/
#648990000000
0!
1"
0'
1(
0/
10
#649000000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#649010000000
0!
1$
0'
1+
0/
#649020000000
1!
1'
1/
#649030000000
0!
0'
0/
#649040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#649050000000
0!
0'
0/
#649060000000
1!
1'
1/
#649070000000
0!
0'
0/
#649080000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#649090000000
0!
0'
0/
#649100000000
1!
1'
1/
#649110000000
0!
0'
0/
#649120000000
1!
1'
1/
#649130000000
0!
0'
0/
#649140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#649150000000
0!
0'
0/
#649160000000
1!
1'
1/
#649170000000
0!
0'
0/
#649180000000
1!
1'
1/
#649190000000
0!
0'
0/
#649200000000
1!
1'
1/
#649210000000
0!
0'
0/
#649220000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#649230000000
0!
0'
0/
#649240000000
1!
1'
1/
#649250000000
0!
0'
0/
#649260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#649270000000
0!
0'
0/
#649280000000
1!
1'
1/
#649290000000
0!
0'
0/
#649300000000
#649310000000
1!
1'
1/
#649320000000
0!
0'
0/
#649330000000
1!
1'
1/
#649340000000
0!
1"
0'
1(
0/
10
#649350000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#649360000000
0!
0'
0/
#649370000000
1!
1'
1/
#649380000000
0!
0'
0/
#649390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#649400000000
0!
0'
0/
#649410000000
1!
1'
1/
#649420000000
0!
1"
0'
1(
0/
10
#649430000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#649440000000
0!
1$
0'
1+
0/
#649450000000
1!
1'
1/
#649460000000
0!
0'
0/
#649470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#649480000000
0!
0'
0/
#649490000000
1!
1'
1/
#649500000000
0!
0'
0/
#649510000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#649520000000
0!
0'
0/
#649530000000
1!
1'
1/
#649540000000
0!
0'
0/
#649550000000
1!
1'
1/
#649560000000
0!
0'
0/
#649570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#649580000000
0!
0'
0/
#649590000000
1!
1'
1/
#649600000000
0!
0'
0/
#649610000000
1!
1'
1/
#649620000000
0!
0'
0/
#649630000000
1!
1'
1/
#649640000000
0!
0'
0/
#649650000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#649660000000
0!
0'
0/
#649670000000
1!
1'
1/
#649680000000
0!
0'
0/
#649690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#649700000000
0!
0'
0/
#649710000000
1!
1'
1/
#649720000000
0!
0'
0/
#649730000000
#649740000000
1!
1'
1/
#649750000000
0!
0'
0/
#649760000000
1!
1'
1/
#649770000000
0!
1"
0'
1(
0/
10
#649780000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#649790000000
0!
0'
0/
#649800000000
1!
1'
1/
#649810000000
0!
0'
0/
#649820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#649830000000
0!
0'
0/
#649840000000
1!
1'
1/
#649850000000
0!
1"
0'
1(
0/
10
#649860000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#649870000000
0!
1$
0'
1+
0/
#649880000000
1!
1'
1/
#649890000000
0!
0'
0/
#649900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#649910000000
0!
0'
0/
#649920000000
1!
1'
1/
#649930000000
0!
0'
0/
#649940000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#649950000000
0!
0'
0/
#649960000000
1!
1'
1/
#649970000000
0!
0'
0/
#649980000000
1!
1'
1/
#649990000000
0!
0'
0/
#650000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#650010000000
0!
0'
0/
#650020000000
1!
1'
1/
#650030000000
0!
0'
0/
#650040000000
1!
1'
1/
#650050000000
0!
0'
0/
#650060000000
1!
1'
1/
#650070000000
0!
0'
0/
#650080000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#650090000000
0!
0'
0/
#650100000000
1!
1'
1/
#650110000000
0!
0'
0/
#650120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#650130000000
0!
0'
0/
#650140000000
1!
1'
1/
#650150000000
0!
0'
0/
#650160000000
#650170000000
1!
1'
1/
#650180000000
0!
0'
0/
#650190000000
1!
1'
1/
#650200000000
0!
1"
0'
1(
0/
10
#650210000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#650220000000
0!
0'
0/
#650230000000
1!
1'
1/
#650240000000
0!
0'
0/
#650250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#650260000000
0!
0'
0/
#650270000000
1!
1'
1/
#650280000000
0!
1"
0'
1(
0/
10
#650290000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#650300000000
0!
1$
0'
1+
0/
#650310000000
1!
1'
1/
#650320000000
0!
0'
0/
#650330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#650340000000
0!
0'
0/
#650350000000
1!
1'
1/
#650360000000
0!
0'
0/
#650370000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#650380000000
0!
0'
0/
#650390000000
1!
1'
1/
#650400000000
0!
0'
0/
#650410000000
1!
1'
1/
#650420000000
0!
0'
0/
#650430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#650440000000
0!
0'
0/
#650450000000
1!
1'
1/
#650460000000
0!
0'
0/
#650470000000
1!
1'
1/
#650480000000
0!
0'
0/
#650490000000
1!
1'
1/
#650500000000
0!
0'
0/
#650510000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#650520000000
0!
0'
0/
#650530000000
1!
1'
1/
#650540000000
0!
0'
0/
#650550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#650560000000
0!
0'
0/
#650570000000
1!
1'
1/
#650580000000
0!
0'
0/
#650590000000
#650600000000
1!
1'
1/
#650610000000
0!
0'
0/
#650620000000
1!
1'
1/
#650630000000
0!
1"
0'
1(
0/
10
#650640000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#650650000000
0!
0'
0/
#650660000000
1!
1'
1/
#650670000000
0!
0'
0/
#650680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#650690000000
0!
0'
0/
#650700000000
1!
1'
1/
#650710000000
0!
1"
0'
1(
0/
10
#650720000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#650730000000
0!
1$
0'
1+
0/
#650740000000
1!
1'
1/
#650750000000
0!
0'
0/
#650760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#650770000000
0!
0'
0/
#650780000000
1!
1'
1/
#650790000000
0!
0'
0/
#650800000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#650810000000
0!
0'
0/
#650820000000
1!
1'
1/
#650830000000
0!
0'
0/
#650840000000
1!
1'
1/
#650850000000
0!
0'
0/
#650860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#650870000000
0!
0'
0/
#650880000000
1!
1'
1/
#650890000000
0!
0'
0/
#650900000000
1!
1'
1/
#650910000000
0!
0'
0/
#650920000000
1!
1'
1/
#650930000000
0!
0'
0/
#650940000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#650950000000
0!
0'
0/
#650960000000
1!
1'
1/
#650970000000
0!
0'
0/
#650980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#650990000000
0!
0'
0/
#651000000000
1!
1'
1/
#651010000000
0!
0'
0/
#651020000000
#651030000000
1!
1'
1/
#651040000000
0!
0'
0/
#651050000000
1!
1'
1/
#651060000000
0!
1"
0'
1(
0/
10
#651070000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#651080000000
0!
0'
0/
#651090000000
1!
1'
1/
#651100000000
0!
0'
0/
#651110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#651120000000
0!
0'
0/
#651130000000
1!
1'
1/
#651140000000
0!
1"
0'
1(
0/
10
#651150000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#651160000000
0!
1$
0'
1+
0/
#651170000000
1!
1'
1/
#651180000000
0!
0'
0/
#651190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#651200000000
0!
0'
0/
#651210000000
1!
1'
1/
#651220000000
0!
0'
0/
#651230000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#651240000000
0!
0'
0/
#651250000000
1!
1'
1/
#651260000000
0!
0'
0/
#651270000000
1!
1'
1/
#651280000000
0!
0'
0/
#651290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#651300000000
0!
0'
0/
#651310000000
1!
1'
1/
#651320000000
0!
0'
0/
#651330000000
1!
1'
1/
#651340000000
0!
0'
0/
#651350000000
1!
1'
1/
#651360000000
0!
0'
0/
#651370000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#651380000000
0!
0'
0/
#651390000000
1!
1'
1/
#651400000000
0!
0'
0/
#651410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#651420000000
0!
0'
0/
#651430000000
1!
1'
1/
#651440000000
0!
0'
0/
#651450000000
#651460000000
1!
1'
1/
#651470000000
0!
0'
0/
#651480000000
1!
1'
1/
#651490000000
0!
1"
0'
1(
0/
10
#651500000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#651510000000
0!
0'
0/
#651520000000
1!
1'
1/
#651530000000
0!
0'
0/
#651540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#651550000000
0!
0'
0/
#651560000000
1!
1'
1/
#651570000000
0!
1"
0'
1(
0/
10
#651580000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#651590000000
0!
1$
0'
1+
0/
#651600000000
1!
1'
1/
#651610000000
0!
0'
0/
#651620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#651630000000
0!
0'
0/
#651640000000
1!
1'
1/
#651650000000
0!
0'
0/
#651660000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#651670000000
0!
0'
0/
#651680000000
1!
1'
1/
#651690000000
0!
0'
0/
#651700000000
1!
1'
1/
#651710000000
0!
0'
0/
#651720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#651730000000
0!
0'
0/
#651740000000
1!
1'
1/
#651750000000
0!
0'
0/
#651760000000
1!
1'
1/
#651770000000
0!
0'
0/
#651780000000
1!
1'
1/
#651790000000
0!
0'
0/
#651800000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#651810000000
0!
0'
0/
#651820000000
1!
1'
1/
#651830000000
0!
0'
0/
#651840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#651850000000
0!
0'
0/
#651860000000
1!
1'
1/
#651870000000
0!
0'
0/
#651880000000
#651890000000
1!
1'
1/
#651900000000
0!
0'
0/
#651910000000
1!
1'
1/
#651920000000
0!
1"
0'
1(
0/
10
#651930000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#651940000000
0!
0'
0/
#651950000000
1!
1'
1/
#651960000000
0!
0'
0/
#651970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#651980000000
0!
0'
0/
#651990000000
1!
1'
1/
#652000000000
0!
1"
0'
1(
0/
10
#652010000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#652020000000
0!
1$
0'
1+
0/
#652030000000
1!
1'
1/
#652040000000
0!
0'
0/
#652050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#652060000000
0!
0'
0/
#652070000000
1!
1'
1/
#652080000000
0!
0'
0/
#652090000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#652100000000
0!
0'
0/
#652110000000
1!
1'
1/
#652120000000
0!
0'
0/
#652130000000
1!
1'
1/
#652140000000
0!
0'
0/
#652150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#652160000000
0!
0'
0/
#652170000000
1!
1'
1/
#652180000000
0!
0'
0/
#652190000000
1!
1'
1/
#652200000000
0!
0'
0/
#652210000000
1!
1'
1/
#652220000000
0!
0'
0/
#652230000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#652240000000
0!
0'
0/
#652250000000
1!
1'
1/
#652260000000
0!
0'
0/
#652270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#652280000000
0!
0'
0/
#652290000000
1!
1'
1/
#652300000000
0!
0'
0/
#652310000000
#652320000000
1!
1'
1/
#652330000000
0!
0'
0/
#652340000000
1!
1'
1/
#652350000000
0!
1"
0'
1(
0/
10
#652360000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#652370000000
0!
0'
0/
#652380000000
1!
1'
1/
#652390000000
0!
0'
0/
#652400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#652410000000
0!
0'
0/
#652420000000
1!
1'
1/
#652430000000
0!
1"
0'
1(
0/
10
#652440000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#652450000000
0!
1$
0'
1+
0/
#652460000000
1!
1'
1/
#652470000000
0!
0'
0/
#652480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#652490000000
0!
0'
0/
#652500000000
1!
1'
1/
#652510000000
0!
0'
0/
#652520000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#652530000000
0!
0'
0/
#652540000000
1!
1'
1/
#652550000000
0!
0'
0/
#652560000000
1!
1'
1/
#652570000000
0!
0'
0/
#652580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#652590000000
0!
0'
0/
#652600000000
1!
1'
1/
#652610000000
0!
0'
0/
#652620000000
1!
1'
1/
#652630000000
0!
0'
0/
#652640000000
1!
1'
1/
#652650000000
0!
0'
0/
#652660000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#652670000000
0!
0'
0/
#652680000000
1!
1'
1/
#652690000000
0!
0'
0/
#652700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#652710000000
0!
0'
0/
#652720000000
1!
1'
1/
#652730000000
0!
0'
0/
#652740000000
#652750000000
1!
1'
1/
#652760000000
0!
0'
0/
#652770000000
1!
1'
1/
#652780000000
0!
1"
0'
1(
0/
10
#652790000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#652800000000
0!
0'
0/
#652810000000
1!
1'
1/
#652820000000
0!
0'
0/
#652830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#652840000000
0!
0'
0/
#652850000000
1!
1'
1/
#652860000000
0!
1"
0'
1(
0/
10
#652870000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#652880000000
0!
1$
0'
1+
0/
#652890000000
1!
1'
1/
#652900000000
0!
0'
0/
#652910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#652920000000
0!
0'
0/
#652930000000
1!
1'
1/
#652940000000
0!
0'
0/
#652950000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#652960000000
0!
0'
0/
#652970000000
1!
1'
1/
#652980000000
0!
0'
0/
#652990000000
1!
1'
1/
#653000000000
0!
0'
0/
#653010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#653020000000
0!
0'
0/
#653030000000
1!
1'
1/
#653040000000
0!
0'
0/
#653050000000
1!
1'
1/
#653060000000
0!
0'
0/
#653070000000
1!
1'
1/
#653080000000
0!
0'
0/
#653090000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#653100000000
0!
0'
0/
#653110000000
1!
1'
1/
#653120000000
0!
0'
0/
#653130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#653140000000
0!
0'
0/
#653150000000
1!
1'
1/
#653160000000
0!
0'
0/
#653170000000
#653180000000
1!
1'
1/
#653190000000
0!
0'
0/
#653200000000
1!
1'
1/
#653210000000
0!
1"
0'
1(
0/
10
#653220000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#653230000000
0!
0'
0/
#653240000000
1!
1'
1/
#653250000000
0!
0'
0/
#653260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#653270000000
0!
0'
0/
#653280000000
1!
1'
1/
#653290000000
0!
1"
0'
1(
0/
10
#653300000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#653310000000
0!
1$
0'
1+
0/
#653320000000
1!
1'
1/
#653330000000
0!
0'
0/
#653340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#653350000000
0!
0'
0/
#653360000000
1!
1'
1/
#653370000000
0!
0'
0/
#653380000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#653390000000
0!
0'
0/
#653400000000
1!
1'
1/
#653410000000
0!
0'
0/
#653420000000
1!
1'
1/
#653430000000
0!
0'
0/
#653440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#653450000000
0!
0'
0/
#653460000000
1!
1'
1/
#653470000000
0!
0'
0/
#653480000000
1!
1'
1/
#653490000000
0!
0'
0/
#653500000000
1!
1'
1/
#653510000000
0!
0'
0/
#653520000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#653530000000
0!
0'
0/
#653540000000
1!
1'
1/
#653550000000
0!
0'
0/
#653560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#653570000000
0!
0'
0/
#653580000000
1!
1'
1/
#653590000000
0!
0'
0/
#653600000000
#653610000000
1!
1'
1/
#653620000000
0!
0'
0/
#653630000000
1!
1'
1/
#653640000000
0!
1"
0'
1(
0/
10
#653650000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#653660000000
0!
0'
0/
#653670000000
1!
1'
1/
#653680000000
0!
0'
0/
#653690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#653700000000
0!
0'
0/
#653710000000
1!
1'
1/
#653720000000
0!
1"
0'
1(
0/
10
#653730000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#653740000000
0!
1$
0'
1+
0/
#653750000000
1!
1'
1/
#653760000000
0!
0'
0/
#653770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#653780000000
0!
0'
0/
#653790000000
1!
1'
1/
#653800000000
0!
0'
0/
#653810000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#653820000000
0!
0'
0/
#653830000000
1!
1'
1/
#653840000000
0!
0'
0/
#653850000000
1!
1'
1/
#653860000000
0!
0'
0/
#653870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#653880000000
0!
0'
0/
#653890000000
1!
1'
1/
#653900000000
0!
0'
0/
#653910000000
1!
1'
1/
#653920000000
0!
0'
0/
#653930000000
1!
1'
1/
#653940000000
0!
0'
0/
#653950000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#653960000000
0!
0'
0/
#653970000000
1!
1'
1/
#653980000000
0!
0'
0/
#653990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#654000000000
0!
0'
0/
#654010000000
1!
1'
1/
#654020000000
0!
0'
0/
#654030000000
#654040000000
1!
1'
1/
#654050000000
0!
0'
0/
#654060000000
1!
1'
1/
#654070000000
0!
1"
0'
1(
0/
10
#654080000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#654090000000
0!
0'
0/
#654100000000
1!
1'
1/
#654110000000
0!
0'
0/
#654120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#654130000000
0!
0'
0/
#654140000000
1!
1'
1/
#654150000000
0!
1"
0'
1(
0/
10
#654160000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#654170000000
0!
1$
0'
1+
0/
#654180000000
1!
1'
1/
#654190000000
0!
0'
0/
#654200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#654210000000
0!
0'
0/
#654220000000
1!
1'
1/
#654230000000
0!
0'
0/
#654240000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#654250000000
0!
0'
0/
#654260000000
1!
1'
1/
#654270000000
0!
0'
0/
#654280000000
1!
1'
1/
#654290000000
0!
0'
0/
#654300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#654310000000
0!
0'
0/
#654320000000
1!
1'
1/
#654330000000
0!
0'
0/
#654340000000
1!
1'
1/
#654350000000
0!
0'
0/
#654360000000
1!
1'
1/
#654370000000
0!
0'
0/
#654380000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#654390000000
0!
0'
0/
#654400000000
1!
1'
1/
#654410000000
0!
0'
0/
#654420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#654430000000
0!
0'
0/
#654440000000
1!
1'
1/
#654450000000
0!
0'
0/
#654460000000
#654470000000
1!
1'
1/
#654480000000
0!
0'
0/
#654490000000
1!
1'
1/
#654500000000
0!
1"
0'
1(
0/
10
#654510000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#654520000000
0!
0'
0/
#654530000000
1!
1'
1/
#654540000000
0!
0'
0/
#654550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#654560000000
0!
0'
0/
#654570000000
1!
1'
1/
#654580000000
0!
1"
0'
1(
0/
10
#654590000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#654600000000
0!
1$
0'
1+
0/
#654610000000
1!
1'
1/
#654620000000
0!
0'
0/
#654630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#654640000000
0!
0'
0/
#654650000000
1!
1'
1/
#654660000000
0!
0'
0/
#654670000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#654680000000
0!
0'
0/
#654690000000
1!
1'
1/
#654700000000
0!
0'
0/
#654710000000
1!
1'
1/
#654720000000
0!
0'
0/
#654730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#654740000000
0!
0'
0/
#654750000000
1!
1'
1/
#654760000000
0!
0'
0/
#654770000000
1!
1'
1/
#654780000000
0!
0'
0/
#654790000000
1!
1'
1/
#654800000000
0!
0'
0/
#654810000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#654820000000
0!
0'
0/
#654830000000
1!
1'
1/
#654840000000
0!
0'
0/
#654850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#654860000000
0!
0'
0/
#654870000000
1!
1'
1/
#654880000000
0!
0'
0/
#654890000000
#654900000000
1!
1'
1/
#654910000000
0!
0'
0/
#654920000000
1!
1'
1/
#654930000000
0!
1"
0'
1(
0/
10
#654940000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#654950000000
0!
0'
0/
#654960000000
1!
1'
1/
#654970000000
0!
0'
0/
#654980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#654990000000
0!
0'
0/
#655000000000
1!
1'
1/
#655010000000
0!
1"
0'
1(
0/
10
#655020000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#655030000000
0!
1$
0'
1+
0/
#655040000000
1!
1'
1/
#655050000000
0!
0'
0/
#655060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#655070000000
0!
0'
0/
#655080000000
1!
1'
1/
#655090000000
0!
0'
0/
#655100000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#655110000000
0!
0'
0/
#655120000000
1!
1'
1/
#655130000000
0!
0'
0/
#655140000000
1!
1'
1/
#655150000000
0!
0'
0/
#655160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#655170000000
0!
0'
0/
#655180000000
1!
1'
1/
#655190000000
0!
0'
0/
#655200000000
1!
1'
1/
#655210000000
0!
0'
0/
#655220000000
1!
1'
1/
#655230000000
0!
0'
0/
#655240000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#655250000000
0!
0'
0/
#655260000000
1!
1'
1/
#655270000000
0!
0'
0/
#655280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#655290000000
0!
0'
0/
#655300000000
1!
1'
1/
#655310000000
0!
0'
0/
#655320000000
#655330000000
1!
1'
1/
#655340000000
0!
0'
0/
#655350000000
1!
1'
1/
#655360000000
0!
1"
0'
1(
0/
10
#655370000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#655380000000
0!
0'
0/
#655390000000
1!
1'
1/
#655400000000
0!
0'
0/
#655410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#655420000000
0!
0'
0/
#655430000000
1!
1'
1/
#655440000000
0!
1"
0'
1(
0/
10
#655450000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#655460000000
0!
1$
0'
1+
0/
#655470000000
1!
1'
1/
#655480000000
0!
0'
0/
#655490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#655500000000
0!
0'
0/
#655510000000
1!
1'
1/
#655520000000
0!
0'
0/
#655530000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#655540000000
0!
0'
0/
#655550000000
1!
1'
1/
#655560000000
0!
0'
0/
#655570000000
1!
1'
1/
#655580000000
0!
0'
0/
#655590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#655600000000
0!
0'
0/
#655610000000
1!
1'
1/
#655620000000
0!
0'
0/
#655630000000
1!
1'
1/
#655640000000
0!
0'
0/
#655650000000
1!
1'
1/
#655660000000
0!
0'
0/
#655670000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#655680000000
0!
0'
0/
#655690000000
1!
1'
1/
#655700000000
0!
0'
0/
#655710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#655720000000
0!
0'
0/
#655730000000
1!
1'
1/
#655740000000
0!
0'
0/
#655750000000
#655760000000
1!
1'
1/
#655770000000
0!
0'
0/
#655780000000
1!
1'
1/
#655790000000
0!
1"
0'
1(
0/
10
#655800000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#655810000000
0!
0'
0/
#655820000000
1!
1'
1/
#655830000000
0!
0'
0/
#655840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#655850000000
0!
0'
0/
#655860000000
1!
1'
1/
#655870000000
0!
1"
0'
1(
0/
10
#655880000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#655890000000
0!
1$
0'
1+
0/
#655900000000
1!
1'
1/
#655910000000
0!
0'
0/
#655920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#655930000000
0!
0'
0/
#655940000000
1!
1'
1/
#655950000000
0!
0'
0/
#655960000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#655970000000
0!
0'
0/
#655980000000
1!
1'
1/
#655990000000
0!
0'
0/
#656000000000
1!
1'
1/
#656010000000
0!
0'
0/
#656020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#656030000000
0!
0'
0/
#656040000000
1!
1'
1/
#656050000000
0!
0'
0/
#656060000000
1!
1'
1/
#656070000000
0!
0'
0/
#656080000000
1!
1'
1/
#656090000000
0!
0'
0/
#656100000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#656110000000
0!
0'
0/
#656120000000
1!
1'
1/
#656130000000
0!
0'
0/
#656140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#656150000000
0!
0'
0/
#656160000000
1!
1'
1/
#656170000000
0!
0'
0/
#656180000000
#656190000000
1!
1'
1/
#656200000000
0!
0'
0/
#656210000000
1!
1'
1/
#656220000000
0!
1"
0'
1(
0/
10
#656230000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#656240000000
0!
0'
0/
#656250000000
1!
1'
1/
#656260000000
0!
0'
0/
#656270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#656280000000
0!
0'
0/
#656290000000
1!
1'
1/
#656300000000
0!
1"
0'
1(
0/
10
#656310000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#656320000000
0!
1$
0'
1+
0/
#656330000000
1!
1'
1/
#656340000000
0!
0'
0/
#656350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#656360000000
0!
0'
0/
#656370000000
1!
1'
1/
#656380000000
0!
0'
0/
#656390000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#656400000000
0!
0'
0/
#656410000000
1!
1'
1/
#656420000000
0!
0'
0/
#656430000000
1!
1'
1/
#656440000000
0!
0'
0/
#656450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#656460000000
0!
0'
0/
#656470000000
1!
1'
1/
#656480000000
0!
0'
0/
#656490000000
1!
1'
1/
#656500000000
0!
0'
0/
#656510000000
1!
1'
1/
#656520000000
0!
0'
0/
#656530000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#656540000000
0!
0'
0/
#656550000000
1!
1'
1/
#656560000000
0!
0'
0/
#656570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#656580000000
0!
0'
0/
#656590000000
1!
1'
1/
#656600000000
0!
0'
0/
#656610000000
#656620000000
1!
1'
1/
#656630000000
0!
0'
0/
#656640000000
1!
1'
1/
#656650000000
0!
1"
0'
1(
0/
10
#656660000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#656670000000
0!
0'
0/
#656680000000
1!
1'
1/
#656690000000
0!
0'
0/
#656700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#656710000000
0!
0'
0/
#656720000000
1!
1'
1/
#656730000000
0!
1"
0'
1(
0/
10
#656740000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#656750000000
0!
1$
0'
1+
0/
#656760000000
1!
1'
1/
#656770000000
0!
0'
0/
#656780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#656790000000
0!
0'
0/
#656800000000
1!
1'
1/
#656810000000
0!
0'
0/
#656820000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#656830000000
0!
0'
0/
#656840000000
1!
1'
1/
#656850000000
0!
0'
0/
#656860000000
1!
1'
1/
#656870000000
0!
0'
0/
#656880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#656890000000
0!
0'
0/
#656900000000
1!
1'
1/
#656910000000
0!
0'
0/
#656920000000
1!
1'
1/
#656930000000
0!
0'
0/
#656940000000
1!
1'
1/
#656950000000
0!
0'
0/
#656960000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#656970000000
0!
0'
0/
#656980000000
1!
1'
1/
#656990000000
0!
0'
0/
#657000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#657010000000
0!
0'
0/
#657020000000
1!
1'
1/
#657030000000
0!
0'
0/
#657040000000
#657050000000
1!
1'
1/
#657060000000
0!
0'
0/
#657070000000
1!
1'
1/
#657080000000
0!
1"
0'
1(
0/
10
#657090000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#657100000000
0!
0'
0/
#657110000000
1!
1'
1/
#657120000000
0!
0'
0/
#657130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#657140000000
0!
0'
0/
#657150000000
1!
1'
1/
#657160000000
0!
1"
0'
1(
0/
10
#657170000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#657180000000
0!
1$
0'
1+
0/
#657190000000
1!
1'
1/
#657200000000
0!
0'
0/
#657210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#657220000000
0!
0'
0/
#657230000000
1!
1'
1/
#657240000000
0!
0'
0/
#657250000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#657260000000
0!
0'
0/
#657270000000
1!
1'
1/
#657280000000
0!
0'
0/
#657290000000
1!
1'
1/
#657300000000
0!
0'
0/
#657310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#657320000000
0!
0'
0/
#657330000000
1!
1'
1/
#657340000000
0!
0'
0/
#657350000000
1!
1'
1/
#657360000000
0!
0'
0/
#657370000000
1!
1'
1/
#657380000000
0!
0'
0/
#657390000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#657400000000
0!
0'
0/
#657410000000
1!
1'
1/
#657420000000
0!
0'
0/
#657430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#657440000000
0!
0'
0/
#657450000000
1!
1'
1/
#657460000000
0!
0'
0/
#657470000000
#657480000000
1!
1'
1/
#657490000000
0!
0'
0/
#657500000000
1!
1'
1/
#657510000000
0!
1"
0'
1(
0/
10
#657520000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#657530000000
0!
0'
0/
#657540000000
1!
1'
1/
#657550000000
0!
0'
0/
#657560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#657570000000
0!
0'
0/
#657580000000
1!
1'
1/
#657590000000
0!
1"
0'
1(
0/
10
#657600000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#657610000000
0!
1$
0'
1+
0/
#657620000000
1!
1'
1/
#657630000000
0!
0'
0/
#657640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#657650000000
0!
0'
0/
#657660000000
1!
1'
1/
#657670000000
0!
0'
0/
#657680000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#657690000000
0!
0'
0/
#657700000000
1!
1'
1/
#657710000000
0!
0'
0/
#657720000000
1!
1'
1/
#657730000000
0!
0'
0/
#657740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#657750000000
0!
0'
0/
#657760000000
1!
1'
1/
#657770000000
0!
0'
0/
#657780000000
1!
1'
1/
#657790000000
0!
0'
0/
#657800000000
1!
1'
1/
#657810000000
0!
0'
0/
#657820000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#657830000000
0!
0'
0/
#657840000000
1!
1'
1/
#657850000000
0!
0'
0/
#657860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#657870000000
0!
0'
0/
#657880000000
1!
1'
1/
#657890000000
0!
0'
0/
#657900000000
#657910000000
1!
1'
1/
#657920000000
0!
0'
0/
#657930000000
1!
1'
1/
#657940000000
0!
1"
0'
1(
0/
10
#657950000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#657960000000
0!
0'
0/
#657970000000
1!
1'
1/
#657980000000
0!
0'
0/
#657990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#658000000000
0!
0'
0/
#658010000000
1!
1'
1/
#658020000000
0!
1"
0'
1(
0/
10
#658030000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#658040000000
0!
1$
0'
1+
0/
#658050000000
1!
1'
1/
#658060000000
0!
0'
0/
#658070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#658080000000
0!
0'
0/
#658090000000
1!
1'
1/
#658100000000
0!
0'
0/
#658110000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#658120000000
0!
0'
0/
#658130000000
1!
1'
1/
#658140000000
0!
0'
0/
#658150000000
1!
1'
1/
#658160000000
0!
0'
0/
#658170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#658180000000
0!
0'
0/
#658190000000
1!
1'
1/
#658200000000
0!
0'
0/
#658210000000
1!
1'
1/
#658220000000
0!
0'
0/
#658230000000
1!
1'
1/
#658240000000
0!
0'
0/
#658250000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#658260000000
0!
0'
0/
#658270000000
1!
1'
1/
#658280000000
0!
0'
0/
#658290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#658300000000
0!
0'
0/
#658310000000
1!
1'
1/
#658320000000
0!
0'
0/
#658330000000
#658340000000
1!
1'
1/
#658350000000
0!
0'
0/
#658360000000
1!
1'
1/
#658370000000
0!
1"
0'
1(
0/
10
#658380000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#658390000000
0!
0'
0/
#658400000000
1!
1'
1/
#658410000000
0!
0'
0/
#658420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#658430000000
0!
0'
0/
#658440000000
1!
1'
1/
#658450000000
0!
1"
0'
1(
0/
10
#658460000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#658470000000
0!
1$
0'
1+
0/
#658480000000
1!
1'
1/
#658490000000
0!
0'
0/
#658500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#658510000000
0!
0'
0/
#658520000000
1!
1'
1/
#658530000000
0!
0'
0/
#658540000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#658550000000
0!
0'
0/
#658560000000
1!
1'
1/
#658570000000
0!
0'
0/
#658580000000
1!
1'
1/
#658590000000
0!
0'
0/
#658600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#658610000000
0!
0'
0/
#658620000000
1!
1'
1/
#658630000000
0!
0'
0/
#658640000000
1!
1'
1/
#658650000000
0!
0'
0/
#658660000000
1!
1'
1/
#658670000000
0!
0'
0/
#658680000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#658690000000
0!
0'
0/
#658700000000
1!
1'
1/
#658710000000
0!
0'
0/
#658720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#658730000000
0!
0'
0/
#658740000000
1!
1'
1/
#658750000000
0!
0'
0/
#658760000000
#658770000000
1!
1'
1/
#658780000000
0!
0'
0/
#658790000000
1!
1'
1/
#658800000000
0!
1"
0'
1(
0/
10
#658810000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#658820000000
0!
0'
0/
#658830000000
1!
1'
1/
#658840000000
0!
0'
0/
#658850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#658860000000
0!
0'
0/
#658870000000
1!
1'
1/
#658880000000
0!
1"
0'
1(
0/
10
#658890000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#658900000000
0!
1$
0'
1+
0/
#658910000000
1!
1'
1/
#658920000000
0!
0'
0/
#658930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#658940000000
0!
0'
0/
#658950000000
1!
1'
1/
#658960000000
0!
0'
0/
#658970000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#658980000000
0!
0'
0/
#658990000000
1!
1'
1/
#659000000000
0!
0'
0/
#659010000000
1!
1'
1/
#659020000000
0!
0'
0/
#659030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#659040000000
0!
0'
0/
#659050000000
1!
1'
1/
#659060000000
0!
0'
0/
#659070000000
1!
1'
1/
#659080000000
0!
0'
0/
#659090000000
1!
1'
1/
#659100000000
0!
0'
0/
#659110000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#659120000000
0!
0'
0/
#659130000000
1!
1'
1/
#659140000000
0!
0'
0/
#659150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#659160000000
0!
0'
0/
#659170000000
1!
1'
1/
#659180000000
0!
0'
0/
#659190000000
#659200000000
1!
1'
1/
#659210000000
0!
0'
0/
#659220000000
1!
1'
1/
#659230000000
0!
1"
0'
1(
0/
10
#659240000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#659250000000
0!
0'
0/
#659260000000
1!
1'
1/
#659270000000
0!
0'
0/
#659280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#659290000000
0!
0'
0/
#659300000000
1!
1'
1/
#659310000000
0!
1"
0'
1(
0/
10
#659320000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#659330000000
0!
1$
0'
1+
0/
#659340000000
1!
1'
1/
#659350000000
0!
0'
0/
#659360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#659370000000
0!
0'
0/
#659380000000
1!
1'
1/
#659390000000
0!
0'
0/
#659400000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#659410000000
0!
0'
0/
#659420000000
1!
1'
1/
#659430000000
0!
0'
0/
#659440000000
1!
1'
1/
#659450000000
0!
0'
0/
#659460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#659470000000
0!
0'
0/
#659480000000
1!
1'
1/
#659490000000
0!
0'
0/
#659500000000
1!
1'
1/
#659510000000
0!
0'
0/
#659520000000
1!
1'
1/
#659530000000
0!
0'
0/
#659540000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#659550000000
0!
0'
0/
#659560000000
1!
1'
1/
#659570000000
0!
0'
0/
#659580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#659590000000
0!
0'
0/
#659600000000
1!
1'
1/
#659610000000
0!
0'
0/
#659620000000
#659630000000
1!
1'
1/
#659640000000
0!
0'
0/
#659650000000
1!
1'
1/
#659660000000
0!
1"
0'
1(
0/
10
#659670000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#659680000000
0!
0'
0/
#659690000000
1!
1'
1/
#659700000000
0!
0'
0/
#659710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#659720000000
0!
0'
0/
#659730000000
1!
1'
1/
#659740000000
0!
1"
0'
1(
0/
10
#659750000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#659760000000
0!
1$
0'
1+
0/
#659770000000
1!
1'
1/
#659780000000
0!
0'
0/
#659790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#659800000000
0!
0'
0/
#659810000000
1!
1'
1/
#659820000000
0!
0'
0/
#659830000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#659840000000
0!
0'
0/
#659850000000
1!
1'
1/
#659860000000
0!
0'
0/
#659870000000
1!
1'
1/
#659880000000
0!
0'
0/
#659890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#659900000000
0!
0'
0/
#659910000000
1!
1'
1/
#659920000000
0!
0'
0/
#659930000000
1!
1'
1/
#659940000000
0!
0'
0/
#659950000000
1!
1'
1/
#659960000000
0!
0'
0/
#659970000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#659980000000
0!
0'
0/
#659990000000
1!
1'
1/
#660000000000
0!
0'
0/
#660010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#660020000000
0!
0'
0/
#660030000000
1!
1'
1/
#660040000000
0!
0'
0/
#660050000000
#660060000000
1!
1'
1/
#660070000000
0!
0'
0/
#660080000000
1!
1'
1/
#660090000000
0!
1"
0'
1(
0/
10
#660100000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#660110000000
0!
0'
0/
#660120000000
1!
1'
1/
#660130000000
0!
0'
0/
#660140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#660150000000
0!
0'
0/
#660160000000
1!
1'
1/
#660170000000
0!
1"
0'
1(
0/
10
#660180000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#660190000000
0!
1$
0'
1+
0/
#660200000000
1!
1'
1/
#660210000000
0!
0'
0/
#660220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#660230000000
0!
0'
0/
#660240000000
1!
1'
1/
#660250000000
0!
0'
0/
#660260000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#660270000000
0!
0'
0/
#660280000000
1!
1'
1/
#660290000000
0!
0'
0/
#660300000000
1!
1'
1/
#660310000000
0!
0'
0/
#660320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#660330000000
0!
0'
0/
#660340000000
1!
1'
1/
#660350000000
0!
0'
0/
#660360000000
1!
1'
1/
#660370000000
0!
0'
0/
#660380000000
1!
1'
1/
#660390000000
0!
0'
0/
#660400000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#660410000000
0!
0'
0/
#660420000000
1!
1'
1/
#660430000000
0!
0'
0/
#660440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#660450000000
0!
0'
0/
#660460000000
1!
1'
1/
#660470000000
0!
0'
0/
#660480000000
#660490000000
1!
1'
1/
#660500000000
0!
0'
0/
#660510000000
1!
1'
1/
#660520000000
0!
1"
0'
1(
0/
10
#660530000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#660540000000
0!
0'
0/
#660550000000
1!
1'
1/
#660560000000
0!
0'
0/
#660570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#660580000000
0!
0'
0/
#660590000000
1!
1'
1/
#660600000000
0!
1"
0'
1(
0/
10
#660610000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#660620000000
0!
1$
0'
1+
0/
#660630000000
1!
1'
1/
#660640000000
0!
0'
0/
#660650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#660660000000
0!
0'
0/
#660670000000
1!
1'
1/
#660680000000
0!
0'
0/
#660690000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#660700000000
0!
0'
0/
#660710000000
1!
1'
1/
#660720000000
0!
0'
0/
#660730000000
1!
1'
1/
#660740000000
0!
0'
0/
#660750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#660760000000
0!
0'
0/
#660770000000
1!
1'
1/
#660780000000
0!
0'
0/
#660790000000
1!
1'
1/
#660800000000
0!
0'
0/
#660810000000
1!
1'
1/
#660820000000
0!
0'
0/
#660830000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#660840000000
0!
0'
0/
#660850000000
1!
1'
1/
#660860000000
0!
0'
0/
#660870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#660880000000
0!
0'
0/
#660890000000
1!
1'
1/
#660900000000
0!
0'
0/
#660910000000
#660920000000
1!
1'
1/
#660930000000
0!
0'
0/
#660940000000
1!
1'
1/
#660950000000
0!
1"
0'
1(
0/
10
#660960000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#660970000000
0!
0'
0/
#660980000000
1!
1'
1/
#660990000000
0!
0'
0/
#661000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#661010000000
0!
0'
0/
#661020000000
1!
1'
1/
#661030000000
0!
1"
0'
1(
0/
10
#661040000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#661050000000
0!
1$
0'
1+
0/
#661060000000
1!
1'
1/
#661070000000
0!
0'
0/
#661080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#661090000000
0!
0'
0/
#661100000000
1!
1'
1/
#661110000000
0!
0'
0/
#661120000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#661130000000
0!
0'
0/
#661140000000
1!
1'
1/
#661150000000
0!
0'
0/
#661160000000
1!
1'
1/
#661170000000
0!
0'
0/
#661180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#661190000000
0!
0'
0/
#661200000000
1!
1'
1/
#661210000000
0!
0'
0/
#661220000000
1!
1'
1/
#661230000000
0!
0'
0/
#661240000000
1!
1'
1/
#661250000000
0!
0'
0/
#661260000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#661270000000
0!
0'
0/
#661280000000
1!
1'
1/
#661290000000
0!
0'
0/
#661300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#661310000000
0!
0'
0/
#661320000000
1!
1'
1/
#661330000000
0!
0'
0/
#661340000000
#661350000000
1!
1'
1/
#661360000000
0!
0'
0/
#661370000000
1!
1'
1/
#661380000000
0!
1"
0'
1(
0/
10
#661390000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#661400000000
0!
0'
0/
#661410000000
1!
1'
1/
#661420000000
0!
0'
0/
#661430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#661440000000
0!
0'
0/
#661450000000
1!
1'
1/
#661460000000
0!
1"
0'
1(
0/
10
#661470000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#661480000000
0!
1$
0'
1+
0/
#661490000000
1!
1'
1/
#661500000000
0!
0'
0/
#661510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#661520000000
0!
0'
0/
#661530000000
1!
1'
1/
#661540000000
0!
0'
0/
#661550000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#661560000000
0!
0'
0/
#661570000000
1!
1'
1/
#661580000000
0!
0'
0/
#661590000000
1!
1'
1/
#661600000000
0!
0'
0/
#661610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#661620000000
0!
0'
0/
#661630000000
1!
1'
1/
#661640000000
0!
0'
0/
#661650000000
1!
1'
1/
#661660000000
0!
0'
0/
#661670000000
1!
1'
1/
#661680000000
0!
0'
0/
#661690000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#661700000000
0!
0'
0/
#661710000000
1!
1'
1/
#661720000000
0!
0'
0/
#661730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#661740000000
0!
0'
0/
#661750000000
1!
1'
1/
#661760000000
0!
0'
0/
#661770000000
#661780000000
1!
1'
1/
#661790000000
0!
0'
0/
#661800000000
1!
1'
1/
#661810000000
0!
1"
0'
1(
0/
10
#661820000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#661830000000
0!
0'
0/
#661840000000
1!
1'
1/
#661850000000
0!
0'
0/
#661860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#661870000000
0!
0'
0/
#661880000000
1!
1'
1/
#661890000000
0!
1"
0'
1(
0/
10
#661900000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#661910000000
0!
1$
0'
1+
0/
#661920000000
1!
1'
1/
#661930000000
0!
0'
0/
#661940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#661950000000
0!
0'
0/
#661960000000
1!
1'
1/
#661970000000
0!
0'
0/
#661980000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#661990000000
0!
0'
0/
#662000000000
1!
1'
1/
#662010000000
0!
0'
0/
#662020000000
1!
1'
1/
#662030000000
0!
0'
0/
#662040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#662050000000
0!
0'
0/
#662060000000
1!
1'
1/
#662070000000
0!
0'
0/
#662080000000
1!
1'
1/
#662090000000
0!
0'
0/
#662100000000
1!
1'
1/
#662110000000
0!
0'
0/
#662120000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#662130000000
0!
0'
0/
#662140000000
1!
1'
1/
#662150000000
0!
0'
0/
#662160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#662170000000
0!
0'
0/
#662180000000
1!
1'
1/
#662190000000
0!
0'
0/
#662200000000
#662210000000
1!
1'
1/
#662220000000
0!
0'
0/
#662230000000
1!
1'
1/
#662240000000
0!
1"
0'
1(
0/
10
#662250000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#662260000000
0!
0'
0/
#662270000000
1!
1'
1/
#662280000000
0!
0'
0/
#662290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#662300000000
0!
0'
0/
#662310000000
1!
1'
1/
#662320000000
0!
1"
0'
1(
0/
10
#662330000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#662340000000
0!
1$
0'
1+
0/
#662350000000
1!
1'
1/
#662360000000
0!
0'
0/
#662370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#662380000000
0!
0'
0/
#662390000000
1!
1'
1/
#662400000000
0!
0'
0/
#662410000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#662420000000
0!
0'
0/
#662430000000
1!
1'
1/
#662440000000
0!
0'
0/
#662450000000
1!
1'
1/
#662460000000
0!
0'
0/
#662470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#662480000000
0!
0'
0/
#662490000000
1!
1'
1/
#662500000000
0!
0'
0/
#662510000000
1!
1'
1/
#662520000000
0!
0'
0/
#662530000000
1!
1'
1/
#662540000000
0!
0'
0/
#662550000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#662560000000
0!
0'
0/
#662570000000
1!
1'
1/
#662580000000
0!
0'
0/
#662590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#662600000000
0!
0'
0/
#662610000000
1!
1'
1/
#662620000000
0!
0'
0/
#662630000000
#662640000000
1!
1'
1/
#662650000000
0!
0'
0/
#662660000000
1!
1'
1/
#662670000000
0!
1"
0'
1(
0/
10
#662680000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#662690000000
0!
0'
0/
#662700000000
1!
1'
1/
#662710000000
0!
0'
0/
#662720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#662730000000
0!
0'
0/
#662740000000
1!
1'
1/
#662750000000
0!
1"
0'
1(
0/
10
#662760000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#662770000000
0!
1$
0'
1+
0/
#662780000000
1!
1'
1/
#662790000000
0!
0'
0/
#662800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#662810000000
0!
0'
0/
#662820000000
1!
1'
1/
#662830000000
0!
0'
0/
#662840000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#662850000000
0!
0'
0/
#662860000000
1!
1'
1/
#662870000000
0!
0'
0/
#662880000000
1!
1'
1/
#662890000000
0!
0'
0/
#662900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#662910000000
0!
0'
0/
#662920000000
1!
1'
1/
#662930000000
0!
0'
0/
#662940000000
1!
1'
1/
#662950000000
0!
0'
0/
#662960000000
1!
1'
1/
#662970000000
0!
0'
0/
#662980000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#662990000000
0!
0'
0/
#663000000000
1!
1'
1/
#663010000000
0!
0'
0/
#663020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#663030000000
0!
0'
0/
#663040000000
1!
1'
1/
#663050000000
0!
0'
0/
#663060000000
#663070000000
1!
1'
1/
#663080000000
0!
0'
0/
#663090000000
1!
1'
1/
#663100000000
0!
1"
0'
1(
0/
10
#663110000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#663120000000
0!
0'
0/
#663130000000
1!
1'
1/
#663140000000
0!
0'
0/
#663150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#663160000000
0!
0'
0/
#663170000000
1!
1'
1/
#663180000000
0!
1"
0'
1(
0/
10
#663190000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#663200000000
0!
1$
0'
1+
0/
#663210000000
1!
1'
1/
#663220000000
0!
0'
0/
#663230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#663240000000
0!
0'
0/
#663250000000
1!
1'
1/
#663260000000
0!
0'
0/
#663270000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#663280000000
0!
0'
0/
#663290000000
1!
1'
1/
#663300000000
0!
0'
0/
#663310000000
1!
1'
1/
#663320000000
0!
0'
0/
#663330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#663340000000
0!
0'
0/
#663350000000
1!
1'
1/
#663360000000
0!
0'
0/
#663370000000
1!
1'
1/
#663380000000
0!
0'
0/
#663390000000
1!
1'
1/
#663400000000
0!
0'
0/
#663410000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#663420000000
0!
0'
0/
#663430000000
1!
1'
1/
#663440000000
0!
0'
0/
#663450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#663460000000
0!
0'
0/
#663470000000
1!
1'
1/
#663480000000
0!
0'
0/
#663490000000
#663500000000
1!
1'
1/
#663510000000
0!
0'
0/
#663520000000
1!
1'
1/
#663530000000
0!
1"
0'
1(
0/
10
#663540000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#663550000000
0!
0'
0/
#663560000000
1!
1'
1/
#663570000000
0!
0'
0/
#663580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#663590000000
0!
0'
0/
#663600000000
1!
1'
1/
#663610000000
0!
1"
0'
1(
0/
10
#663620000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#663630000000
0!
1$
0'
1+
0/
#663640000000
1!
1'
1/
#663650000000
0!
0'
0/
#663660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#663670000000
0!
0'
0/
#663680000000
1!
1'
1/
#663690000000
0!
0'
0/
#663700000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#663710000000
0!
0'
0/
#663720000000
1!
1'
1/
#663730000000
0!
0'
0/
#663740000000
1!
1'
1/
#663750000000
0!
0'
0/
#663760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#663770000000
0!
0'
0/
#663780000000
1!
1'
1/
#663790000000
0!
0'
0/
#663800000000
1!
1'
1/
#663810000000
0!
0'
0/
#663820000000
1!
1'
1/
#663830000000
0!
0'
0/
#663840000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#663850000000
0!
0'
0/
#663860000000
1!
1'
1/
#663870000000
0!
0'
0/
#663880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#663890000000
0!
0'
0/
#663900000000
1!
1'
1/
#663910000000
0!
0'
0/
#663920000000
#663930000000
1!
1'
1/
#663940000000
0!
0'
0/
#663950000000
1!
1'
1/
#663960000000
0!
1"
0'
1(
0/
10
#663970000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#663980000000
0!
0'
0/
#663990000000
1!
1'
1/
#664000000000
0!
0'
0/
#664010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#664020000000
0!
0'
0/
#664030000000
1!
1'
1/
#664040000000
0!
1"
0'
1(
0/
10
#664050000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#664060000000
0!
1$
0'
1+
0/
#664070000000
1!
1'
1/
#664080000000
0!
0'
0/
#664090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#664100000000
0!
0'
0/
#664110000000
1!
1'
1/
#664120000000
0!
0'
0/
#664130000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#664140000000
0!
0'
0/
#664150000000
1!
1'
1/
#664160000000
0!
0'
0/
#664170000000
1!
1'
1/
#664180000000
0!
0'
0/
#664190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#664200000000
0!
0'
0/
#664210000000
1!
1'
1/
#664220000000
0!
0'
0/
#664230000000
1!
1'
1/
#664240000000
0!
0'
0/
#664250000000
1!
1'
1/
#664260000000
0!
0'
0/
#664270000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#664280000000
0!
0'
0/
#664290000000
1!
1'
1/
#664300000000
0!
0'
0/
#664310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#664320000000
0!
0'
0/
#664330000000
1!
1'
1/
#664340000000
0!
0'
0/
#664350000000
#664360000000
1!
1'
1/
#664370000000
0!
0'
0/
#664380000000
1!
1'
1/
#664390000000
0!
1"
0'
1(
0/
10
#664400000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#664410000000
0!
0'
0/
#664420000000
1!
1'
1/
#664430000000
0!
0'
0/
#664440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#664450000000
0!
0'
0/
#664460000000
1!
1'
1/
#664470000000
0!
1"
0'
1(
0/
10
#664480000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#664490000000
0!
1$
0'
1+
0/
#664500000000
1!
1'
1/
#664510000000
0!
0'
0/
#664520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#664530000000
0!
0'
0/
#664540000000
1!
1'
1/
#664550000000
0!
0'
0/
#664560000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#664570000000
0!
0'
0/
#664580000000
1!
1'
1/
#664590000000
0!
0'
0/
#664600000000
1!
1'
1/
#664610000000
0!
0'
0/
#664620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#664630000000
0!
0'
0/
#664640000000
1!
1'
1/
#664650000000
0!
0'
0/
#664660000000
1!
1'
1/
#664670000000
0!
0'
0/
#664680000000
1!
1'
1/
#664690000000
0!
0'
0/
#664700000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#664710000000
0!
0'
0/
#664720000000
1!
1'
1/
#664730000000
0!
0'
0/
#664740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#664750000000
0!
0'
0/
#664760000000
1!
1'
1/
#664770000000
0!
0'
0/
#664780000000
#664790000000
1!
1'
1/
#664800000000
0!
0'
0/
#664810000000
1!
1'
1/
#664820000000
0!
1"
0'
1(
0/
10
#664830000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#664840000000
0!
0'
0/
#664850000000
1!
1'
1/
#664860000000
0!
0'
0/
#664870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#664880000000
0!
0'
0/
#664890000000
1!
1'
1/
#664900000000
0!
1"
0'
1(
0/
10
#664910000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#664920000000
0!
1$
0'
1+
0/
#664930000000
1!
1'
1/
#664940000000
0!
0'
0/
#664950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#664960000000
0!
0'
0/
#664970000000
1!
1'
1/
#664980000000
0!
0'
0/
#664990000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#665000000000
0!
0'
0/
#665010000000
1!
1'
1/
#665020000000
0!
0'
0/
#665030000000
1!
1'
1/
#665040000000
0!
0'
0/
#665050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#665060000000
0!
0'
0/
#665070000000
1!
1'
1/
#665080000000
0!
0'
0/
#665090000000
1!
1'
1/
#665100000000
0!
0'
0/
#665110000000
1!
1'
1/
#665120000000
0!
0'
0/
#665130000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#665140000000
0!
0'
0/
#665150000000
1!
1'
1/
#665160000000
0!
0'
0/
#665170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#665180000000
0!
0'
0/
#665190000000
1!
1'
1/
#665200000000
0!
0'
0/
#665210000000
#665220000000
1!
1'
1/
#665230000000
0!
0'
0/
#665240000000
1!
1'
1/
#665250000000
0!
1"
0'
1(
0/
10
#665260000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#665270000000
0!
0'
0/
#665280000000
1!
1'
1/
#665290000000
0!
0'
0/
#665300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#665310000000
0!
0'
0/
#665320000000
1!
1'
1/
#665330000000
0!
1"
0'
1(
0/
10
#665340000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#665350000000
0!
1$
0'
1+
0/
#665360000000
1!
1'
1/
#665370000000
0!
0'
0/
#665380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#665390000000
0!
0'
0/
#665400000000
1!
1'
1/
#665410000000
0!
0'
0/
#665420000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#665430000000
0!
0'
0/
#665440000000
1!
1'
1/
#665450000000
0!
0'
0/
#665460000000
1!
1'
1/
#665470000000
0!
0'
0/
#665480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#665490000000
0!
0'
0/
#665500000000
1!
1'
1/
#665510000000
0!
0'
0/
#665520000000
1!
1'
1/
#665530000000
0!
0'
0/
#665540000000
1!
1'
1/
#665550000000
0!
0'
0/
#665560000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#665570000000
0!
0'
0/
#665580000000
1!
1'
1/
#665590000000
0!
0'
0/
#665600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#665610000000
0!
0'
0/
#665620000000
1!
1'
1/
#665630000000
0!
0'
0/
#665640000000
#665650000000
1!
1'
1/
#665660000000
0!
0'
0/
#665670000000
1!
1'
1/
#665680000000
0!
1"
0'
1(
0/
10
#665690000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#665700000000
0!
0'
0/
#665710000000
1!
1'
1/
#665720000000
0!
0'
0/
#665730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#665740000000
0!
0'
0/
#665750000000
1!
1'
1/
#665760000000
0!
1"
0'
1(
0/
10
#665770000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#665780000000
0!
1$
0'
1+
0/
#665790000000
1!
1'
1/
#665800000000
0!
0'
0/
#665810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#665820000000
0!
0'
0/
#665830000000
1!
1'
1/
#665840000000
0!
0'
0/
#665850000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#665860000000
0!
0'
0/
#665870000000
1!
1'
1/
#665880000000
0!
0'
0/
#665890000000
1!
1'
1/
#665900000000
0!
0'
0/
#665910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#665920000000
0!
0'
0/
#665930000000
1!
1'
1/
#665940000000
0!
0'
0/
#665950000000
1!
1'
1/
#665960000000
0!
0'
0/
#665970000000
1!
1'
1/
#665980000000
0!
0'
0/
#665990000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#666000000000
0!
0'
0/
#666010000000
1!
1'
1/
#666020000000
0!
0'
0/
#666030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#666040000000
0!
0'
0/
#666050000000
1!
1'
1/
#666060000000
0!
0'
0/
#666070000000
#666080000000
1!
1'
1/
#666090000000
0!
0'
0/
#666100000000
1!
1'
1/
#666110000000
0!
1"
0'
1(
0/
10
#666120000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#666130000000
0!
0'
0/
#666140000000
1!
1'
1/
#666150000000
0!
0'
0/
#666160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#666170000000
0!
0'
0/
#666180000000
1!
1'
1/
#666190000000
0!
1"
0'
1(
0/
10
#666200000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#666210000000
0!
1$
0'
1+
0/
#666220000000
1!
1'
1/
#666230000000
0!
0'
0/
#666240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#666250000000
0!
0'
0/
#666260000000
1!
1'
1/
#666270000000
0!
0'
0/
#666280000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#666290000000
0!
0'
0/
#666300000000
1!
1'
1/
#666310000000
0!
0'
0/
#666320000000
1!
1'
1/
#666330000000
0!
0'
0/
#666340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#666350000000
0!
0'
0/
#666360000000
1!
1'
1/
#666370000000
0!
0'
0/
#666380000000
1!
1'
1/
#666390000000
0!
0'
0/
#666400000000
1!
1'
1/
#666410000000
0!
0'
0/
#666420000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#666430000000
0!
0'
0/
#666440000000
1!
1'
1/
#666450000000
0!
0'
0/
#666460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#666470000000
0!
0'
0/
#666480000000
1!
1'
1/
#666490000000
0!
0'
0/
#666500000000
#666510000000
1!
1'
1/
#666520000000
0!
0'
0/
#666530000000
1!
1'
1/
#666540000000
0!
1"
0'
1(
0/
10
#666550000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#666560000000
0!
0'
0/
#666570000000
1!
1'
1/
#666580000000
0!
0'
0/
#666590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#666600000000
0!
0'
0/
#666610000000
1!
1'
1/
#666620000000
0!
1"
0'
1(
0/
10
#666630000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#666640000000
0!
1$
0'
1+
0/
#666650000000
1!
1'
1/
#666660000000
0!
0'
0/
#666670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#666680000000
0!
0'
0/
#666690000000
1!
1'
1/
#666700000000
0!
0'
0/
#666710000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#666720000000
0!
0'
0/
#666730000000
1!
1'
1/
#666740000000
0!
0'
0/
#666750000000
1!
1'
1/
#666760000000
0!
0'
0/
#666770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#666780000000
0!
0'
0/
#666790000000
1!
1'
1/
#666800000000
0!
0'
0/
#666810000000
1!
1'
1/
#666820000000
0!
0'
0/
#666830000000
1!
1'
1/
#666840000000
0!
0'
0/
#666850000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#666860000000
0!
0'
0/
#666870000000
1!
1'
1/
#666880000000
0!
0'
0/
#666890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#666900000000
0!
0'
0/
#666910000000
1!
1'
1/
#666920000000
0!
0'
0/
#666930000000
#666940000000
1!
1'
1/
#666950000000
0!
0'
0/
#666960000000
1!
1'
1/
#666970000000
0!
1"
0'
1(
0/
10
#666980000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#666990000000
0!
0'
0/
#667000000000
1!
1'
1/
#667010000000
0!
0'
0/
#667020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#667030000000
0!
0'
0/
#667040000000
1!
1'
1/
#667050000000
0!
1"
0'
1(
0/
10
#667060000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#667070000000
0!
1$
0'
1+
0/
#667080000000
1!
1'
1/
#667090000000
0!
0'
0/
#667100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#667110000000
0!
0'
0/
#667120000000
1!
1'
1/
#667130000000
0!
0'
0/
#667140000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#667150000000
0!
0'
0/
#667160000000
1!
1'
1/
#667170000000
0!
0'
0/
#667180000000
1!
1'
1/
#667190000000
0!
0'
0/
#667200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#667210000000
0!
0'
0/
#667220000000
1!
1'
1/
#667230000000
0!
0'
0/
#667240000000
1!
1'
1/
#667250000000
0!
0'
0/
#667260000000
1!
1'
1/
#667270000000
0!
0'
0/
#667280000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#667290000000
0!
0'
0/
#667300000000
1!
1'
1/
#667310000000
0!
0'
0/
#667320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#667330000000
0!
0'
0/
#667340000000
1!
1'
1/
#667350000000
0!
0'
0/
#667360000000
#667370000000
1!
1'
1/
#667380000000
0!
0'
0/
#667390000000
1!
1'
1/
#667400000000
0!
1"
0'
1(
0/
10
#667410000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#667420000000
0!
0'
0/
#667430000000
1!
1'
1/
#667440000000
0!
0'
0/
#667450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#667460000000
0!
0'
0/
#667470000000
1!
1'
1/
#667480000000
0!
1"
0'
1(
0/
10
#667490000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#667500000000
0!
1$
0'
1+
0/
#667510000000
1!
1'
1/
#667520000000
0!
0'
0/
#667530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#667540000000
0!
0'
0/
#667550000000
1!
1'
1/
#667560000000
0!
0'
0/
#667570000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#667580000000
0!
0'
0/
#667590000000
1!
1'
1/
#667600000000
0!
0'
0/
#667610000000
1!
1'
1/
#667620000000
0!
0'
0/
#667630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#667640000000
0!
0'
0/
#667650000000
1!
1'
1/
#667660000000
0!
0'
0/
#667670000000
1!
1'
1/
#667680000000
0!
0'
0/
#667690000000
1!
1'
1/
#667700000000
0!
0'
0/
#667710000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#667720000000
0!
0'
0/
#667730000000
1!
1'
1/
#667740000000
0!
0'
0/
#667750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#667760000000
0!
0'
0/
#667770000000
1!
1'
1/
#667780000000
0!
0'
0/
#667790000000
#667800000000
1!
1'
1/
#667810000000
0!
0'
0/
#667820000000
1!
1'
1/
#667830000000
0!
1"
0'
1(
0/
10
#667840000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#667850000000
0!
0'
0/
#667860000000
1!
1'
1/
#667870000000
0!
0'
0/
#667880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#667890000000
0!
0'
0/
#667900000000
1!
1'
1/
#667910000000
0!
1"
0'
1(
0/
10
#667920000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#667930000000
0!
1$
0'
1+
0/
#667940000000
1!
1'
1/
#667950000000
0!
0'
0/
#667960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#667970000000
0!
0'
0/
#667980000000
1!
1'
1/
#667990000000
0!
0'
0/
#668000000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#668010000000
0!
0'
0/
#668020000000
1!
1'
1/
#668030000000
0!
0'
0/
#668040000000
1!
1'
1/
#668050000000
0!
0'
0/
#668060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#668070000000
0!
0'
0/
#668080000000
1!
1'
1/
#668090000000
0!
0'
0/
#668100000000
1!
1'
1/
#668110000000
0!
0'
0/
#668120000000
1!
1'
1/
#668130000000
0!
0'
0/
#668140000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#668150000000
0!
0'
0/
#668160000000
1!
1'
1/
#668170000000
0!
0'
0/
#668180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#668190000000
0!
0'
0/
#668200000000
1!
1'
1/
#668210000000
0!
0'
0/
#668220000000
#668230000000
1!
1'
1/
#668240000000
0!
0'
0/
#668250000000
1!
1'
1/
#668260000000
0!
1"
0'
1(
0/
10
#668270000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#668280000000
0!
0'
0/
#668290000000
1!
1'
1/
#668300000000
0!
0'
0/
#668310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#668320000000
0!
0'
0/
#668330000000
1!
1'
1/
#668340000000
0!
1"
0'
1(
0/
10
#668350000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#668360000000
0!
1$
0'
1+
0/
#668370000000
1!
1'
1/
#668380000000
0!
0'
0/
#668390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#668400000000
0!
0'
0/
#668410000000
1!
1'
1/
#668420000000
0!
0'
0/
#668430000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#668440000000
0!
0'
0/
#668450000000
1!
1'
1/
#668460000000
0!
0'
0/
#668470000000
1!
1'
1/
#668480000000
0!
0'
0/
#668490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#668500000000
0!
0'
0/
#668510000000
1!
1'
1/
#668520000000
0!
0'
0/
#668530000000
1!
1'
1/
#668540000000
0!
0'
0/
#668550000000
1!
1'
1/
#668560000000
0!
0'
0/
#668570000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#668580000000
0!
0'
0/
#668590000000
1!
1'
1/
#668600000000
0!
0'
0/
#668610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#668620000000
0!
0'
0/
#668630000000
1!
1'
1/
#668640000000
0!
0'
0/
#668650000000
#668660000000
1!
1'
1/
#668670000000
0!
0'
0/
#668680000000
1!
1'
1/
#668690000000
0!
1"
0'
1(
0/
10
#668700000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#668710000000
0!
0'
0/
#668720000000
1!
1'
1/
#668730000000
0!
0'
0/
#668740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#668750000000
0!
0'
0/
#668760000000
1!
1'
1/
#668770000000
0!
1"
0'
1(
0/
10
#668780000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#668790000000
0!
1$
0'
1+
0/
#668800000000
1!
1'
1/
#668810000000
0!
0'
0/
#668820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#668830000000
0!
0'
0/
#668840000000
1!
1'
1/
#668850000000
0!
0'
0/
#668860000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#668870000000
0!
0'
0/
#668880000000
1!
1'
1/
#668890000000
0!
0'
0/
#668900000000
1!
1'
1/
#668910000000
0!
0'
0/
#668920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#668930000000
0!
0'
0/
#668940000000
1!
1'
1/
#668950000000
0!
0'
0/
#668960000000
1!
1'
1/
#668970000000
0!
0'
0/
#668980000000
1!
1'
1/
#668990000000
0!
0'
0/
#669000000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#669010000000
0!
0'
0/
#669020000000
1!
1'
1/
#669030000000
0!
0'
0/
#669040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#669050000000
0!
0'
0/
#669060000000
1!
1'
1/
#669070000000
0!
0'
0/
#669080000000
#669090000000
1!
1'
1/
#669100000000
0!
0'
0/
#669110000000
1!
1'
1/
#669120000000
0!
1"
0'
1(
0/
10
#669130000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#669140000000
0!
0'
0/
#669150000000
1!
1'
1/
#669160000000
0!
0'
0/
#669170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#669180000000
0!
0'
0/
#669190000000
1!
1'
1/
#669200000000
0!
1"
0'
1(
0/
10
#669210000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#669220000000
0!
1$
0'
1+
0/
#669230000000
1!
1'
1/
#669240000000
0!
0'
0/
#669250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#669260000000
0!
0'
0/
#669270000000
1!
1'
1/
#669280000000
0!
0'
0/
#669290000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#669300000000
0!
0'
0/
#669310000000
1!
1'
1/
#669320000000
0!
0'
0/
#669330000000
1!
1'
1/
#669340000000
0!
0'
0/
#669350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#669360000000
0!
0'
0/
#669370000000
1!
1'
1/
#669380000000
0!
0'
0/
#669390000000
1!
1'
1/
#669400000000
0!
0'
0/
#669410000000
1!
1'
1/
#669420000000
0!
0'
0/
#669430000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#669440000000
0!
0'
0/
#669450000000
1!
1'
1/
#669460000000
0!
0'
0/
#669470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#669480000000
0!
0'
0/
#669490000000
1!
1'
1/
#669500000000
0!
0'
0/
#669510000000
#669520000000
1!
1'
1/
#669530000000
0!
0'
0/
#669540000000
1!
1'
1/
#669550000000
0!
1"
0'
1(
0/
10
#669560000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#669570000000
0!
0'
0/
#669580000000
1!
1'
1/
#669590000000
0!
0'
0/
#669600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#669610000000
0!
0'
0/
#669620000000
1!
1'
1/
#669630000000
0!
1"
0'
1(
0/
10
#669640000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#669650000000
0!
1$
0'
1+
0/
#669660000000
1!
1'
1/
#669670000000
0!
0'
0/
#669680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#669690000000
0!
0'
0/
#669700000000
1!
1'
1/
#669710000000
0!
0'
0/
#669720000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#669730000000
0!
0'
0/
#669740000000
1!
1'
1/
#669750000000
0!
0'
0/
#669760000000
1!
1'
1/
#669770000000
0!
0'
0/
#669780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#669790000000
0!
0'
0/
#669800000000
1!
1'
1/
#669810000000
0!
0'
0/
#669820000000
1!
1'
1/
#669830000000
0!
0'
0/
#669840000000
1!
1'
1/
#669850000000
0!
0'
0/
#669860000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#669870000000
0!
0'
0/
#669880000000
1!
1'
1/
#669890000000
0!
0'
0/
#669900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#669910000000
0!
0'
0/
#669920000000
1!
1'
1/
#669930000000
0!
0'
0/
#669940000000
#669950000000
1!
1'
1/
#669960000000
0!
0'
0/
#669970000000
1!
1'
1/
#669980000000
0!
1"
0'
1(
0/
10
#669990000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#670000000000
0!
0'
0/
#670010000000
1!
1'
1/
#670020000000
0!
0'
0/
#670030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#670040000000
0!
0'
0/
#670050000000
1!
1'
1/
#670060000000
0!
1"
0'
1(
0/
10
#670070000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#670080000000
0!
1$
0'
1+
0/
#670090000000
1!
1'
1/
#670100000000
0!
0'
0/
#670110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#670120000000
0!
0'
0/
#670130000000
1!
1'
1/
#670140000000
0!
0'
0/
#670150000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#670160000000
0!
0'
0/
#670170000000
1!
1'
1/
#670180000000
0!
0'
0/
#670190000000
1!
1'
1/
#670200000000
0!
0'
0/
#670210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#670220000000
0!
0'
0/
#670230000000
1!
1'
1/
#670240000000
0!
0'
0/
#670250000000
1!
1'
1/
#670260000000
0!
0'
0/
#670270000000
1!
1'
1/
#670280000000
0!
0'
0/
#670290000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#670300000000
0!
0'
0/
#670310000000
1!
1'
1/
#670320000000
0!
0'
0/
#670330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#670340000000
0!
0'
0/
#670350000000
1!
1'
1/
#670360000000
0!
0'
0/
#670370000000
#670380000000
1!
1'
1/
#670390000000
0!
0'
0/
#670400000000
1!
1'
1/
#670410000000
0!
1"
0'
1(
0/
10
#670420000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#670430000000
0!
0'
0/
#670440000000
1!
1'
1/
#670450000000
0!
0'
0/
#670460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#670470000000
0!
0'
0/
#670480000000
1!
1'
1/
#670490000000
0!
1"
0'
1(
0/
10
#670500000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#670510000000
0!
1$
0'
1+
0/
#670520000000
1!
1'
1/
#670530000000
0!
0'
0/
#670540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#670550000000
0!
0'
0/
#670560000000
1!
1'
1/
#670570000000
0!
0'
0/
#670580000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#670590000000
0!
0'
0/
#670600000000
1!
1'
1/
#670610000000
0!
0'
0/
#670620000000
1!
1'
1/
#670630000000
0!
0'
0/
#670640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#670650000000
0!
0'
0/
#670660000000
1!
1'
1/
#670670000000
0!
0'
0/
#670680000000
1!
1'
1/
#670690000000
0!
0'
0/
#670700000000
1!
1'
1/
#670710000000
0!
0'
0/
#670720000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#670730000000
0!
0'
0/
#670740000000
1!
1'
1/
#670750000000
0!
0'
0/
#670760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#670770000000
0!
0'
0/
#670780000000
1!
1'
1/
#670790000000
0!
0'
0/
#670800000000
#670810000000
1!
1'
1/
#670820000000
0!
0'
0/
#670830000000
1!
1'
1/
#670840000000
0!
1"
0'
1(
0/
10
#670850000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#670860000000
0!
0'
0/
#670870000000
1!
1'
1/
#670880000000
0!
0'
0/
#670890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#670900000000
0!
0'
0/
#670910000000
1!
1'
1/
#670920000000
0!
1"
0'
1(
0/
10
#670930000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#670940000000
0!
1$
0'
1+
0/
#670950000000
1!
1'
1/
#670960000000
0!
0'
0/
#670970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#670980000000
0!
0'
0/
#670990000000
1!
1'
1/
#671000000000
0!
0'
0/
#671010000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#671020000000
0!
0'
0/
#671030000000
1!
1'
1/
#671040000000
0!
0'
0/
#671050000000
1!
1'
1/
#671060000000
0!
0'
0/
#671070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#671080000000
0!
0'
0/
#671090000000
1!
1'
1/
#671100000000
0!
0'
0/
#671110000000
1!
1'
1/
#671120000000
0!
0'
0/
#671130000000
1!
1'
1/
#671140000000
0!
0'
0/
#671150000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#671160000000
0!
0'
0/
#671170000000
1!
1'
1/
#671180000000
0!
0'
0/
#671190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#671200000000
0!
0'
0/
#671210000000
1!
1'
1/
#671220000000
0!
0'
0/
#671230000000
#671240000000
1!
1'
1/
#671250000000
0!
0'
0/
#671260000000
1!
1'
1/
#671270000000
0!
1"
0'
1(
0/
10
#671280000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#671290000000
0!
0'
0/
#671300000000
1!
1'
1/
#671310000000
0!
0'
0/
#671320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#671330000000
0!
0'
0/
#671340000000
1!
1'
1/
#671350000000
0!
1"
0'
1(
0/
10
#671360000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#671370000000
0!
1$
0'
1+
0/
#671380000000
1!
1'
1/
#671390000000
0!
0'
0/
#671400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#671410000000
0!
0'
0/
#671420000000
1!
1'
1/
#671430000000
0!
0'
0/
#671440000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#671450000000
0!
0'
0/
#671460000000
1!
1'
1/
#671470000000
0!
0'
0/
#671480000000
1!
1'
1/
#671490000000
0!
0'
0/
#671500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#671510000000
0!
0'
0/
#671520000000
1!
1'
1/
#671530000000
0!
0'
0/
#671540000000
1!
1'
1/
#671550000000
0!
0'
0/
#671560000000
1!
1'
1/
#671570000000
0!
0'
0/
#671580000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#671590000000
0!
0'
0/
#671600000000
1!
1'
1/
#671610000000
0!
0'
0/
#671620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#671630000000
0!
0'
0/
#671640000000
1!
1'
1/
#671650000000
0!
0'
0/
#671660000000
#671670000000
1!
1'
1/
#671680000000
0!
0'
0/
#671690000000
1!
1'
1/
#671700000000
0!
1"
0'
1(
0/
10
#671710000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#671720000000
0!
0'
0/
#671730000000
1!
1'
1/
#671740000000
0!
0'
0/
#671750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#671760000000
0!
0'
0/
#671770000000
1!
1'
1/
#671780000000
0!
1"
0'
1(
0/
10
#671790000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#671800000000
0!
1$
0'
1+
0/
#671810000000
1!
1'
1/
#671820000000
0!
0'
0/
#671830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#671840000000
0!
0'
0/
#671850000000
1!
1'
1/
#671860000000
0!
0'
0/
#671870000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#671880000000
0!
0'
0/
#671890000000
1!
1'
1/
#671900000000
0!
0'
0/
#671910000000
1!
1'
1/
#671920000000
0!
0'
0/
#671930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#671940000000
0!
0'
0/
#671950000000
1!
1'
1/
#671960000000
0!
0'
0/
#671970000000
1!
1'
1/
#671980000000
0!
0'
0/
#671990000000
1!
1'
1/
#672000000000
0!
0'
0/
#672010000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#672020000000
0!
0'
0/
#672030000000
1!
1'
1/
#672040000000
0!
0'
0/
#672050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#672060000000
0!
0'
0/
#672070000000
1!
1'
1/
#672080000000
0!
0'
0/
#672090000000
#672100000000
1!
1'
1/
#672110000000
0!
0'
0/
#672120000000
1!
1'
1/
#672130000000
0!
1"
0'
1(
0/
10
#672140000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#672150000000
0!
0'
0/
#672160000000
1!
1'
1/
#672170000000
0!
0'
0/
#672180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#672190000000
0!
0'
0/
#672200000000
1!
1'
1/
#672210000000
0!
1"
0'
1(
0/
10
#672220000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#672230000000
0!
1$
0'
1+
0/
#672240000000
1!
1'
1/
#672250000000
0!
0'
0/
#672260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#672270000000
0!
0'
0/
#672280000000
1!
1'
1/
#672290000000
0!
0'
0/
#672300000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#672310000000
0!
0'
0/
#672320000000
1!
1'
1/
#672330000000
0!
0'
0/
#672340000000
1!
1'
1/
#672350000000
0!
0'
0/
#672360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#672370000000
0!
0'
0/
#672380000000
1!
1'
1/
#672390000000
0!
0'
0/
#672400000000
1!
1'
1/
#672410000000
0!
0'
0/
#672420000000
1!
1'
1/
#672430000000
0!
0'
0/
#672440000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#672450000000
0!
0'
0/
#672460000000
1!
1'
1/
#672470000000
0!
0'
0/
#672480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#672490000000
0!
0'
0/
#672500000000
1!
1'
1/
#672510000000
0!
0'
0/
#672520000000
#672530000000
1!
1'
1/
#672540000000
0!
0'
0/
#672550000000
1!
1'
1/
#672560000000
0!
1"
0'
1(
0/
10
#672570000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#672580000000
0!
0'
0/
#672590000000
1!
1'
1/
#672600000000
0!
0'
0/
#672610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#672620000000
0!
0'
0/
#672630000000
1!
1'
1/
#672640000000
0!
1"
0'
1(
0/
10
#672650000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#672660000000
0!
1$
0'
1+
0/
#672670000000
1!
1'
1/
#672680000000
0!
0'
0/
#672690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#672700000000
0!
0'
0/
#672710000000
1!
1'
1/
#672720000000
0!
0'
0/
#672730000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#672740000000
0!
0'
0/
#672750000000
1!
1'
1/
#672760000000
0!
0'
0/
#672770000000
1!
1'
1/
#672780000000
0!
0'
0/
#672790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#672800000000
0!
0'
0/
#672810000000
1!
1'
1/
#672820000000
0!
0'
0/
#672830000000
1!
1'
1/
#672840000000
0!
0'
0/
#672850000000
1!
1'
1/
#672860000000
0!
0'
0/
#672870000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#672880000000
0!
0'
0/
#672890000000
1!
1'
1/
#672900000000
0!
0'
0/
#672910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#672920000000
0!
0'
0/
#672930000000
1!
1'
1/
#672940000000
0!
0'
0/
#672950000000
#672960000000
1!
1'
1/
#672970000000
0!
0'
0/
#672980000000
1!
1'
1/
#672990000000
0!
1"
0'
1(
0/
10
#673000000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#673010000000
0!
0'
0/
#673020000000
1!
1'
1/
#673030000000
0!
0'
0/
#673040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#673050000000
0!
0'
0/
#673060000000
1!
1'
1/
#673070000000
0!
1"
0'
1(
0/
10
#673080000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#673090000000
0!
1$
0'
1+
0/
#673100000000
1!
1'
1/
#673110000000
0!
0'
0/
#673120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#673130000000
0!
0'
0/
#673140000000
1!
1'
1/
#673150000000
0!
0'
0/
#673160000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#673170000000
0!
0'
0/
#673180000000
1!
1'
1/
#673190000000
0!
0'
0/
#673200000000
1!
1'
1/
#673210000000
0!
0'
0/
#673220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#673230000000
0!
0'
0/
#673240000000
1!
1'
1/
#673250000000
0!
0'
0/
#673260000000
1!
1'
1/
#673270000000
0!
0'
0/
#673280000000
1!
1'
1/
#673290000000
0!
0'
0/
#673300000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#673310000000
0!
0'
0/
#673320000000
1!
1'
1/
#673330000000
0!
0'
0/
#673340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#673350000000
0!
0'
0/
#673360000000
1!
1'
1/
#673370000000
0!
0'
0/
#673380000000
#673390000000
1!
1'
1/
#673400000000
0!
0'
0/
#673410000000
1!
1'
1/
#673420000000
0!
1"
0'
1(
0/
10
#673430000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#673440000000
0!
0'
0/
#673450000000
1!
1'
1/
#673460000000
0!
0'
0/
#673470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#673480000000
0!
0'
0/
#673490000000
1!
1'
1/
#673500000000
0!
1"
0'
1(
0/
10
#673510000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#673520000000
0!
1$
0'
1+
0/
#673530000000
1!
1'
1/
#673540000000
0!
0'
0/
#673550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#673560000000
0!
0'
0/
#673570000000
1!
1'
1/
#673580000000
0!
0'
0/
#673590000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#673600000000
0!
0'
0/
#673610000000
1!
1'
1/
#673620000000
0!
0'
0/
#673630000000
1!
1'
1/
#673640000000
0!
0'
0/
#673650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#673660000000
0!
0'
0/
#673670000000
1!
1'
1/
#673680000000
0!
0'
0/
#673690000000
1!
1'
1/
#673700000000
0!
0'
0/
#673710000000
1!
1'
1/
#673720000000
0!
0'
0/
#673730000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#673740000000
0!
0'
0/
#673750000000
1!
1'
1/
#673760000000
0!
0'
0/
#673770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#673780000000
0!
0'
0/
#673790000000
1!
1'
1/
#673800000000
0!
0'
0/
#673810000000
#673820000000
1!
1'
1/
#673830000000
0!
0'
0/
#673840000000
1!
1'
1/
#673850000000
0!
1"
0'
1(
0/
10
#673860000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#673870000000
0!
0'
0/
#673880000000
1!
1'
1/
#673890000000
0!
0'
0/
#673900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#673910000000
0!
0'
0/
#673920000000
1!
1'
1/
#673930000000
0!
1"
0'
1(
0/
10
#673940000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#673950000000
0!
1$
0'
1+
0/
#673960000000
1!
1'
1/
#673970000000
0!
0'
0/
#673980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#673990000000
0!
0'
0/
#674000000000
1!
1'
1/
#674010000000
0!
0'
0/
#674020000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#674030000000
0!
0'
0/
#674040000000
1!
1'
1/
#674050000000
0!
0'
0/
#674060000000
1!
1'
1/
#674070000000
0!
0'
0/
#674080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#674090000000
0!
0'
0/
#674100000000
1!
1'
1/
#674110000000
0!
0'
0/
#674120000000
1!
1'
1/
#674130000000
0!
0'
0/
#674140000000
1!
1'
1/
#674150000000
0!
0'
0/
#674160000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#674170000000
0!
0'
0/
#674180000000
1!
1'
1/
#674190000000
0!
0'
0/
#674200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#674210000000
0!
0'
0/
#674220000000
1!
1'
1/
#674230000000
0!
0'
0/
#674240000000
#674250000000
1!
1'
1/
#674260000000
0!
0'
0/
#674270000000
1!
1'
1/
#674280000000
0!
1"
0'
1(
0/
10
#674290000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#674300000000
0!
0'
0/
#674310000000
1!
1'
1/
#674320000000
0!
0'
0/
#674330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#674340000000
0!
0'
0/
#674350000000
1!
1'
1/
#674360000000
0!
1"
0'
1(
0/
10
#674370000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#674380000000
0!
1$
0'
1+
0/
#674390000000
1!
1'
1/
#674400000000
0!
0'
0/
#674410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#674420000000
0!
0'
0/
#674430000000
1!
1'
1/
#674440000000
0!
0'
0/
#674450000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#674460000000
0!
0'
0/
#674470000000
1!
1'
1/
#674480000000
0!
0'
0/
#674490000000
1!
1'
1/
#674500000000
0!
0'
0/
#674510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#674520000000
0!
0'
0/
#674530000000
1!
1'
1/
#674540000000
0!
0'
0/
#674550000000
1!
1'
1/
#674560000000
0!
0'
0/
#674570000000
1!
1'
1/
#674580000000
0!
0'
0/
#674590000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#674600000000
0!
0'
0/
#674610000000
1!
1'
1/
#674620000000
0!
0'
0/
#674630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#674640000000
0!
0'
0/
#674650000000
1!
1'
1/
#674660000000
0!
0'
0/
#674670000000
#674680000000
1!
1'
1/
#674690000000
0!
0'
0/
#674700000000
1!
1'
1/
#674710000000
0!
1"
0'
1(
0/
10
#674720000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#674730000000
0!
0'
0/
#674740000000
1!
1'
1/
#674750000000
0!
0'
0/
#674760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#674770000000
0!
0'
0/
#674780000000
1!
1'
1/
#674790000000
0!
1"
0'
1(
0/
10
#674800000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#674810000000
0!
1$
0'
1+
0/
#674820000000
1!
1'
1/
#674830000000
0!
0'
0/
#674840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#674850000000
0!
0'
0/
#674860000000
1!
1'
1/
#674870000000
0!
0'
0/
#674880000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#674890000000
0!
0'
0/
#674900000000
1!
1'
1/
#674910000000
0!
0'
0/
#674920000000
1!
1'
1/
#674930000000
0!
0'
0/
#674940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#674950000000
0!
0'
0/
#674960000000
1!
1'
1/
#674970000000
0!
0'
0/
#674980000000
1!
1'
1/
#674990000000
0!
0'
0/
#675000000000
1!
1'
1/
#675010000000
0!
0'
0/
#675020000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#675030000000
0!
0'
0/
#675040000000
1!
1'
1/
#675050000000
0!
0'
0/
#675060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#675070000000
0!
0'
0/
#675080000000
1!
1'
1/
#675090000000
0!
0'
0/
#675100000000
#675110000000
1!
1'
1/
#675120000000
0!
0'
0/
#675130000000
1!
1'
1/
#675140000000
0!
1"
0'
1(
0/
10
#675150000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#675160000000
0!
0'
0/
#675170000000
1!
1'
1/
#675180000000
0!
0'
0/
#675190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#675200000000
0!
0'
0/
#675210000000
1!
1'
1/
#675220000000
0!
1"
0'
1(
0/
10
#675230000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#675240000000
0!
1$
0'
1+
0/
#675250000000
1!
1'
1/
#675260000000
0!
0'
0/
#675270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#675280000000
0!
0'
0/
#675290000000
1!
1'
1/
#675300000000
0!
0'
0/
#675310000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#675320000000
0!
0'
0/
#675330000000
1!
1'
1/
#675340000000
0!
0'
0/
#675350000000
1!
1'
1/
#675360000000
0!
0'
0/
#675370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#675380000000
0!
0'
0/
#675390000000
1!
1'
1/
#675400000000
0!
0'
0/
#675410000000
1!
1'
1/
#675420000000
0!
0'
0/
#675430000000
1!
1'
1/
#675440000000
0!
0'
0/
#675450000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#675460000000
0!
0'
0/
#675470000000
1!
1'
1/
#675480000000
0!
0'
0/
#675490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#675500000000
0!
0'
0/
#675510000000
1!
1'
1/
#675520000000
0!
0'
0/
#675530000000
#675540000000
1!
1'
1/
#675550000000
0!
0'
0/
#675560000000
1!
1'
1/
#675570000000
0!
1"
0'
1(
0/
10
#675580000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#675590000000
0!
0'
0/
#675600000000
1!
1'
1/
#675610000000
0!
0'
0/
#675620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#675630000000
0!
0'
0/
#675640000000
1!
1'
1/
#675650000000
0!
1"
0'
1(
0/
10
#675660000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#675670000000
0!
1$
0'
1+
0/
#675680000000
1!
1'
1/
#675690000000
0!
0'
0/
#675700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#675710000000
0!
0'
0/
#675720000000
1!
1'
1/
#675730000000
0!
0'
0/
#675740000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#675750000000
0!
0'
0/
#675760000000
1!
1'
1/
#675770000000
0!
0'
0/
#675780000000
1!
1'
1/
#675790000000
0!
0'
0/
#675800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#675810000000
0!
0'
0/
#675820000000
1!
1'
1/
#675830000000
0!
0'
0/
#675840000000
1!
1'
1/
#675850000000
0!
0'
0/
#675860000000
1!
1'
1/
#675870000000
0!
0'
0/
#675880000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#675890000000
0!
0'
0/
#675900000000
1!
1'
1/
#675910000000
0!
0'
0/
#675920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#675930000000
0!
0'
0/
#675940000000
1!
1'
1/
#675950000000
0!
0'
0/
#675960000000
#675970000000
1!
1'
1/
#675980000000
0!
0'
0/
#675990000000
1!
1'
1/
#676000000000
0!
1"
0'
1(
0/
10
#676010000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#676020000000
0!
0'
0/
#676030000000
1!
1'
1/
#676040000000
0!
0'
0/
#676050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#676060000000
0!
0'
0/
#676070000000
1!
1'
1/
#676080000000
0!
1"
0'
1(
0/
10
#676090000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#676100000000
0!
1$
0'
1+
0/
#676110000000
1!
1'
1/
#676120000000
0!
0'
0/
#676130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#676140000000
0!
0'
0/
#676150000000
1!
1'
1/
#676160000000
0!
0'
0/
#676170000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#676180000000
0!
0'
0/
#676190000000
1!
1'
1/
#676200000000
0!
0'
0/
#676210000000
1!
1'
1/
#676220000000
0!
0'
0/
#676230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#676240000000
0!
0'
0/
#676250000000
1!
1'
1/
#676260000000
0!
0'
0/
#676270000000
1!
1'
1/
#676280000000
0!
0'
0/
#676290000000
1!
1'
1/
#676300000000
0!
0'
0/
#676310000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#676320000000
0!
0'
0/
#676330000000
1!
1'
1/
#676340000000
0!
0'
0/
#676350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#676360000000
0!
0'
0/
#676370000000
1!
1'
1/
#676380000000
0!
0'
0/
#676390000000
#676400000000
1!
1'
1/
#676410000000
0!
0'
0/
#676420000000
1!
1'
1/
#676430000000
0!
1"
0'
1(
0/
10
#676440000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#676450000000
0!
0'
0/
#676460000000
1!
1'
1/
#676470000000
0!
0'
0/
#676480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#676490000000
0!
0'
0/
#676500000000
1!
1'
1/
#676510000000
0!
1"
0'
1(
0/
10
#676520000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#676530000000
0!
1$
0'
1+
0/
#676540000000
1!
1'
1/
#676550000000
0!
0'
0/
#676560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#676570000000
0!
0'
0/
#676580000000
1!
1'
1/
#676590000000
0!
0'
0/
#676600000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#676610000000
0!
0'
0/
#676620000000
1!
1'
1/
#676630000000
0!
0'
0/
#676640000000
1!
1'
1/
#676650000000
0!
0'
0/
#676660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#676670000000
0!
0'
0/
#676680000000
1!
1'
1/
#676690000000
0!
0'
0/
#676700000000
1!
1'
1/
#676710000000
0!
0'
0/
#676720000000
1!
1'
1/
#676730000000
0!
0'
0/
#676740000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#676750000000
0!
0'
0/
#676760000000
1!
1'
1/
#676770000000
0!
0'
0/
#676780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#676790000000
0!
0'
0/
#676800000000
1!
1'
1/
#676810000000
0!
0'
0/
#676820000000
#676830000000
1!
1'
1/
#676840000000
0!
0'
0/
#676850000000
1!
1'
1/
#676860000000
0!
1"
0'
1(
0/
10
#676870000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#676880000000
0!
0'
0/
#676890000000
1!
1'
1/
#676900000000
0!
0'
0/
#676910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#676920000000
0!
0'
0/
#676930000000
1!
1'
1/
#676940000000
0!
1"
0'
1(
0/
10
#676950000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#676960000000
0!
1$
0'
1+
0/
#676970000000
1!
1'
1/
#676980000000
0!
0'
0/
#676990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#677000000000
0!
0'
0/
#677010000000
1!
1'
1/
#677020000000
0!
0'
0/
#677030000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#677040000000
0!
0'
0/
#677050000000
1!
1'
1/
#677060000000
0!
0'
0/
#677070000000
1!
1'
1/
#677080000000
0!
0'
0/
#677090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#677100000000
0!
0'
0/
#677110000000
1!
1'
1/
#677120000000
0!
0'
0/
#677130000000
1!
1'
1/
#677140000000
0!
0'
0/
#677150000000
1!
1'
1/
#677160000000
0!
0'
0/
#677170000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#677180000000
0!
0'
0/
#677190000000
1!
1'
1/
#677200000000
0!
0'
0/
#677210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#677220000000
0!
0'
0/
#677230000000
1!
1'
1/
#677240000000
0!
0'
0/
#677250000000
#677260000000
1!
1'
1/
#677270000000
0!
0'
0/
#677280000000
1!
1'
1/
#677290000000
0!
1"
0'
1(
0/
10
#677300000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#677310000000
0!
0'
0/
#677320000000
1!
1'
1/
#677330000000
0!
0'
0/
#677340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#677350000000
0!
0'
0/
#677360000000
1!
1'
1/
#677370000000
0!
1"
0'
1(
0/
10
#677380000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#677390000000
0!
1$
0'
1+
0/
#677400000000
1!
1'
1/
#677410000000
0!
0'
0/
#677420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#677430000000
0!
0'
0/
#677440000000
1!
1'
1/
#677450000000
0!
0'
0/
#677460000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#677470000000
0!
0'
0/
#677480000000
1!
1'
1/
#677490000000
0!
0'
0/
#677500000000
1!
1'
1/
#677510000000
0!
0'
0/
#677520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#677530000000
0!
0'
0/
#677540000000
1!
1'
1/
#677550000000
0!
0'
0/
#677560000000
1!
1'
1/
#677570000000
0!
0'
0/
#677580000000
1!
1'
1/
#677590000000
0!
0'
0/
#677600000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#677610000000
0!
0'
0/
#677620000000
1!
1'
1/
#677630000000
0!
0'
0/
#677640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#677650000000
0!
0'
0/
#677660000000
1!
1'
1/
#677670000000
0!
0'
0/
#677680000000
#677690000000
1!
1'
1/
#677700000000
0!
0'
0/
#677710000000
1!
1'
1/
#677720000000
0!
1"
0'
1(
0/
10
#677730000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#677740000000
0!
0'
0/
#677750000000
1!
1'
1/
#677760000000
0!
0'
0/
#677770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#677780000000
0!
0'
0/
#677790000000
1!
1'
1/
#677800000000
0!
1"
0'
1(
0/
10
#677810000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#677820000000
0!
1$
0'
1+
0/
#677830000000
1!
1'
1/
#677840000000
0!
0'
0/
#677850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#677860000000
0!
0'
0/
#677870000000
1!
1'
1/
#677880000000
0!
0'
0/
#677890000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#677900000000
0!
0'
0/
#677910000000
1!
1'
1/
#677920000000
0!
0'
0/
#677930000000
1!
1'
1/
#677940000000
0!
0'
0/
#677950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#677960000000
0!
0'
0/
#677970000000
1!
1'
1/
#677980000000
0!
0'
0/
#677990000000
1!
1'
1/
#678000000000
0!
0'
0/
#678010000000
1!
1'
1/
#678020000000
0!
0'
0/
#678030000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#678040000000
0!
0'
0/
#678050000000
1!
1'
1/
#678060000000
0!
0'
0/
#678070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#678080000000
0!
0'
0/
#678090000000
1!
1'
1/
#678100000000
0!
0'
0/
#678110000000
#678120000000
1!
1'
1/
#678130000000
0!
0'
0/
#678140000000
1!
1'
1/
#678150000000
0!
1"
0'
1(
0/
10
#678160000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#678170000000
0!
0'
0/
#678180000000
1!
1'
1/
#678190000000
0!
0'
0/
#678200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#678210000000
0!
0'
0/
#678220000000
1!
1'
1/
#678230000000
0!
1"
0'
1(
0/
10
#678240000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#678250000000
0!
1$
0'
1+
0/
#678260000000
1!
1'
1/
#678270000000
0!
0'
0/
#678280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#678290000000
0!
0'
0/
#678300000000
1!
1'
1/
#678310000000
0!
0'
0/
#678320000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#678330000000
0!
0'
0/
#678340000000
1!
1'
1/
#678350000000
0!
0'
0/
#678360000000
1!
1'
1/
#678370000000
0!
0'
0/
#678380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#678390000000
0!
0'
0/
#678400000000
1!
1'
1/
#678410000000
0!
0'
0/
#678420000000
1!
1'
1/
#678430000000
0!
0'
0/
#678440000000
1!
1'
1/
#678450000000
0!
0'
0/
#678460000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#678470000000
0!
0'
0/
#678480000000
1!
1'
1/
#678490000000
0!
0'
0/
#678500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#678510000000
0!
0'
0/
#678520000000
1!
1'
1/
#678530000000
0!
0'
0/
#678540000000
#678550000000
1!
1'
1/
#678560000000
0!
0'
0/
#678570000000
1!
1'
1/
#678580000000
0!
1"
0'
1(
0/
10
#678590000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#678600000000
0!
0'
0/
#678610000000
1!
1'
1/
#678620000000
0!
0'
0/
#678630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#678640000000
0!
0'
0/
#678650000000
1!
1'
1/
#678660000000
0!
1"
0'
1(
0/
10
#678670000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#678680000000
0!
1$
0'
1+
0/
#678690000000
1!
1'
1/
#678700000000
0!
0'
0/
#678710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#678720000000
0!
0'
0/
#678730000000
1!
1'
1/
#678740000000
0!
0'
0/
#678750000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#678760000000
0!
0'
0/
#678770000000
1!
1'
1/
#678780000000
0!
0'
0/
#678790000000
1!
1'
1/
#678800000000
0!
0'
0/
#678810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#678820000000
0!
0'
0/
#678830000000
1!
1'
1/
#678840000000
0!
0'
0/
#678850000000
1!
1'
1/
#678860000000
0!
0'
0/
#678870000000
1!
1'
1/
#678880000000
0!
0'
0/
#678890000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#678900000000
0!
0'
0/
#678910000000
1!
1'
1/
#678920000000
0!
0'
0/
#678930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#678940000000
0!
0'
0/
#678950000000
1!
1'
1/
#678960000000
0!
0'
0/
#678970000000
#678980000000
1!
1'
1/
#678990000000
0!
0'
0/
#679000000000
1!
1'
1/
#679010000000
0!
1"
0'
1(
0/
10
#679020000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#679030000000
0!
0'
0/
#679040000000
1!
1'
1/
#679050000000
0!
0'
0/
#679060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#679070000000
0!
0'
0/
#679080000000
1!
1'
1/
#679090000000
0!
1"
0'
1(
0/
10
#679100000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#679110000000
0!
1$
0'
1+
0/
#679120000000
1!
1'
1/
#679130000000
0!
0'
0/
#679140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#679150000000
0!
0'
0/
#679160000000
1!
1'
1/
#679170000000
0!
0'
0/
#679180000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#679190000000
0!
0'
0/
#679200000000
1!
1'
1/
#679210000000
0!
0'
0/
#679220000000
1!
1'
1/
#679230000000
0!
0'
0/
#679240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#679250000000
0!
0'
0/
#679260000000
1!
1'
1/
#679270000000
0!
0'
0/
#679280000000
1!
1'
1/
#679290000000
0!
0'
0/
#679300000000
1!
1'
1/
#679310000000
0!
0'
0/
#679320000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#679330000000
0!
0'
0/
#679340000000
1!
1'
1/
#679350000000
0!
0'
0/
#679360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#679370000000
0!
0'
0/
#679380000000
1!
1'
1/
#679390000000
0!
0'
0/
#679400000000
#679410000000
1!
1'
1/
#679420000000
0!
0'
0/
#679430000000
1!
1'
1/
#679440000000
0!
1"
0'
1(
0/
10
#679450000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#679460000000
0!
0'
0/
#679470000000
1!
1'
1/
#679480000000
0!
0'
0/
#679490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#679500000000
0!
0'
0/
#679510000000
1!
1'
1/
#679520000000
0!
1"
0'
1(
0/
10
#679530000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#679540000000
0!
1$
0'
1+
0/
#679550000000
1!
1'
1/
#679560000000
0!
0'
0/
#679570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#679580000000
0!
0'
0/
#679590000000
1!
1'
1/
#679600000000
0!
0'
0/
#679610000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#679620000000
0!
0'
0/
#679630000000
1!
1'
1/
#679640000000
0!
0'
0/
#679650000000
1!
1'
1/
#679660000000
0!
0'
0/
#679670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#679680000000
0!
0'
0/
#679690000000
1!
1'
1/
#679700000000
0!
0'
0/
#679710000000
1!
1'
1/
#679720000000
0!
0'
0/
#679730000000
1!
1'
1/
#679740000000
0!
0'
0/
#679750000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#679760000000
0!
0'
0/
#679770000000
1!
1'
1/
#679780000000
0!
0'
0/
#679790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#679800000000
0!
0'
0/
#679810000000
1!
1'
1/
#679820000000
0!
0'
0/
#679830000000
#679840000000
1!
1'
1/
#679850000000
0!
0'
0/
#679860000000
1!
1'
1/
#679870000000
0!
1"
0'
1(
0/
10
#679880000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#679890000000
0!
0'
0/
#679900000000
1!
1'
1/
#679910000000
0!
0'
0/
#679920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#679930000000
0!
0'
0/
#679940000000
1!
1'
1/
#679950000000
0!
1"
0'
1(
0/
10
#679960000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#679970000000
0!
1$
0'
1+
0/
#679980000000
1!
1'
1/
#679990000000
0!
0'
0/
#680000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#680010000000
0!
0'
0/
#680020000000
1!
1'
1/
#680030000000
0!
0'
0/
#680040000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#680050000000
0!
0'
0/
#680060000000
1!
1'
1/
#680070000000
0!
0'
0/
#680080000000
1!
1'
1/
#680090000000
0!
0'
0/
#680100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#680110000000
0!
0'
0/
#680120000000
1!
1'
1/
#680130000000
0!
0'
0/
#680140000000
1!
1'
1/
#680150000000
0!
0'
0/
#680160000000
1!
1'
1/
#680170000000
0!
0'
0/
#680180000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#680190000000
0!
0'
0/
#680200000000
1!
1'
1/
#680210000000
0!
0'
0/
#680220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#680230000000
0!
0'
0/
#680240000000
1!
1'
1/
#680250000000
0!
0'
0/
#680260000000
#680270000000
1!
1'
1/
#680280000000
0!
0'
0/
#680290000000
1!
1'
1/
#680300000000
0!
1"
0'
1(
0/
10
#680310000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#680320000000
0!
0'
0/
#680330000000
1!
1'
1/
#680340000000
0!
0'
0/
#680350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#680360000000
0!
0'
0/
#680370000000
1!
1'
1/
#680380000000
0!
1"
0'
1(
0/
10
#680390000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#680400000000
0!
1$
0'
1+
0/
#680410000000
1!
1'
1/
#680420000000
0!
0'
0/
#680430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#680440000000
0!
0'
0/
#680450000000
1!
1'
1/
#680460000000
0!
0'
0/
#680470000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#680480000000
0!
0'
0/
#680490000000
1!
1'
1/
#680500000000
0!
0'
0/
#680510000000
1!
1'
1/
#680520000000
0!
0'
0/
#680530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#680540000000
0!
0'
0/
#680550000000
1!
1'
1/
#680560000000
0!
0'
0/
#680570000000
1!
1'
1/
#680580000000
0!
0'
0/
#680590000000
1!
1'
1/
#680600000000
0!
0'
0/
#680610000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#680620000000
0!
0'
0/
#680630000000
1!
1'
1/
#680640000000
0!
0'
0/
#680650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#680660000000
0!
0'
0/
#680670000000
1!
1'
1/
#680680000000
0!
0'
0/
#680690000000
#680700000000
1!
1'
1/
#680710000000
0!
0'
0/
#680720000000
1!
1'
1/
#680730000000
0!
1"
0'
1(
0/
10
#680740000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#680750000000
0!
0'
0/
#680760000000
1!
1'
1/
#680770000000
0!
0'
0/
#680780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#680790000000
0!
0'
0/
#680800000000
1!
1'
1/
#680810000000
0!
1"
0'
1(
0/
10
#680820000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#680830000000
0!
1$
0'
1+
0/
#680840000000
1!
1'
1/
#680850000000
0!
0'
0/
#680860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#680870000000
0!
0'
0/
#680880000000
1!
1'
1/
#680890000000
0!
0'
0/
#680900000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#680910000000
0!
0'
0/
#680920000000
1!
1'
1/
#680930000000
0!
0'
0/
#680940000000
1!
1'
1/
#680950000000
0!
0'
0/
#680960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#680970000000
0!
0'
0/
#680980000000
1!
1'
1/
#680990000000
0!
0'
0/
#681000000000
1!
1'
1/
#681010000000
0!
0'
0/
#681020000000
1!
1'
1/
#681030000000
0!
0'
0/
#681040000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#681050000000
0!
0'
0/
#681060000000
1!
1'
1/
#681070000000
0!
0'
0/
#681080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#681090000000
0!
0'
0/
#681100000000
1!
1'
1/
#681110000000
0!
0'
0/
#681120000000
#681130000000
1!
1'
1/
#681140000000
0!
0'
0/
#681150000000
1!
1'
1/
#681160000000
0!
1"
0'
1(
0/
10
#681170000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#681180000000
0!
0'
0/
#681190000000
1!
1'
1/
#681200000000
0!
0'
0/
#681210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#681220000000
0!
0'
0/
#681230000000
1!
1'
1/
#681240000000
0!
1"
0'
1(
0/
10
#681250000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#681260000000
0!
1$
0'
1+
0/
#681270000000
1!
1'
1/
#681280000000
0!
0'
0/
#681290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#681300000000
0!
0'
0/
#681310000000
1!
1'
1/
#681320000000
0!
0'
0/
#681330000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#681340000000
0!
0'
0/
#681350000000
1!
1'
1/
#681360000000
0!
0'
0/
#681370000000
1!
1'
1/
#681380000000
0!
0'
0/
#681390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#681400000000
0!
0'
0/
#681410000000
1!
1'
1/
#681420000000
0!
0'
0/
#681430000000
1!
1'
1/
#681440000000
0!
0'
0/
#681450000000
1!
1'
1/
#681460000000
0!
0'
0/
#681470000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#681480000000
0!
0'
0/
#681490000000
1!
1'
1/
#681500000000
0!
0'
0/
#681510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#681520000000
0!
0'
0/
#681530000000
1!
1'
1/
#681540000000
0!
0'
0/
#681550000000
#681560000000
1!
1'
1/
#681570000000
0!
0'
0/
#681580000000
1!
1'
1/
#681590000000
0!
1"
0'
1(
0/
10
#681600000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#681610000000
0!
0'
0/
#681620000000
1!
1'
1/
#681630000000
0!
0'
0/
#681640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#681650000000
0!
0'
0/
#681660000000
1!
1'
1/
#681670000000
0!
1"
0'
1(
0/
10
#681680000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#681690000000
0!
1$
0'
1+
0/
#681700000000
1!
1'
1/
#681710000000
0!
0'
0/
#681720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#681730000000
0!
0'
0/
#681740000000
1!
1'
1/
#681750000000
0!
0'
0/
#681760000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#681770000000
0!
0'
0/
#681780000000
1!
1'
1/
#681790000000
0!
0'
0/
#681800000000
1!
1'
1/
#681810000000
0!
0'
0/
#681820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#681830000000
0!
0'
0/
#681840000000
1!
1'
1/
#681850000000
0!
0'
0/
#681860000000
1!
1'
1/
#681870000000
0!
0'
0/
#681880000000
1!
1'
1/
#681890000000
0!
0'
0/
#681900000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#681910000000
0!
0'
0/
#681920000000
1!
1'
1/
#681930000000
0!
0'
0/
#681940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#681950000000
0!
0'
0/
#681960000000
1!
1'
1/
#681970000000
0!
0'
0/
#681980000000
#681990000000
1!
1'
1/
#682000000000
0!
0'
0/
#682010000000
1!
1'
1/
#682020000000
0!
1"
0'
1(
0/
10
#682030000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#682040000000
0!
0'
0/
#682050000000
1!
1'
1/
#682060000000
0!
0'
0/
#682070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#682080000000
0!
0'
0/
#682090000000
1!
1'
1/
#682100000000
0!
1"
0'
1(
0/
10
#682110000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#682120000000
0!
1$
0'
1+
0/
#682130000000
1!
1'
1/
#682140000000
0!
0'
0/
#682150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#682160000000
0!
0'
0/
#682170000000
1!
1'
1/
#682180000000
0!
0'
0/
#682190000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#682200000000
0!
0'
0/
#682210000000
1!
1'
1/
#682220000000
0!
0'
0/
#682230000000
1!
1'
1/
#682240000000
0!
0'
0/
#682250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#682260000000
0!
0'
0/
#682270000000
1!
1'
1/
#682280000000
0!
0'
0/
#682290000000
1!
1'
1/
#682300000000
0!
0'
0/
#682310000000
1!
1'
1/
#682320000000
0!
0'
0/
#682330000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#682340000000
0!
0'
0/
#682350000000
1!
1'
1/
#682360000000
0!
0'
0/
#682370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#682380000000
0!
0'
0/
#682390000000
1!
1'
1/
#682400000000
0!
0'
0/
#682410000000
#682420000000
1!
1'
1/
#682430000000
0!
0'
0/
#682440000000
1!
1'
1/
#682450000000
0!
1"
0'
1(
0/
10
#682460000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#682470000000
0!
0'
0/
#682480000000
1!
1'
1/
#682490000000
0!
0'
0/
#682500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#682510000000
0!
0'
0/
#682520000000
1!
1'
1/
#682530000000
0!
1"
0'
1(
0/
10
#682540000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#682550000000
0!
1$
0'
1+
0/
#682560000000
1!
1'
1/
#682570000000
0!
0'
0/
#682580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#682590000000
0!
0'
0/
#682600000000
1!
1'
1/
#682610000000
0!
0'
0/
#682620000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#682630000000
0!
0'
0/
#682640000000
1!
1'
1/
#682650000000
0!
0'
0/
#682660000000
1!
1'
1/
#682670000000
0!
0'
0/
#682680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#682690000000
0!
0'
0/
#682700000000
1!
1'
1/
#682710000000
0!
0'
0/
#682720000000
1!
1'
1/
#682730000000
0!
0'
0/
#682740000000
1!
1'
1/
#682750000000
0!
0'
0/
#682760000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#682770000000
0!
0'
0/
#682780000000
1!
1'
1/
#682790000000
0!
0'
0/
#682800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#682810000000
0!
0'
0/
#682820000000
1!
1'
1/
#682830000000
0!
0'
0/
#682840000000
#682850000000
1!
1'
1/
#682860000000
0!
0'
0/
#682870000000
1!
1'
1/
#682880000000
0!
1"
0'
1(
0/
10
#682890000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#682900000000
0!
0'
0/
#682910000000
1!
1'
1/
#682920000000
0!
0'
0/
#682930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#682940000000
0!
0'
0/
#682950000000
1!
1'
1/
#682960000000
0!
1"
0'
1(
0/
10
#682970000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#682980000000
0!
1$
0'
1+
0/
#682990000000
1!
1'
1/
#683000000000
0!
0'
0/
#683010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#683020000000
0!
0'
0/
#683030000000
1!
1'
1/
#683040000000
0!
0'
0/
#683050000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#683060000000
0!
0'
0/
#683070000000
1!
1'
1/
#683080000000
0!
0'
0/
#683090000000
1!
1'
1/
#683100000000
0!
0'
0/
#683110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#683120000000
0!
0'
0/
#683130000000
1!
1'
1/
#683140000000
0!
0'
0/
#683150000000
1!
1'
1/
#683160000000
0!
0'
0/
#683170000000
1!
1'
1/
#683180000000
0!
0'
0/
#683190000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#683200000000
0!
0'
0/
#683210000000
1!
1'
1/
#683220000000
0!
0'
0/
#683230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#683240000000
0!
0'
0/
#683250000000
1!
1'
1/
#683260000000
0!
0'
0/
#683270000000
#683280000000
1!
1'
1/
#683290000000
0!
0'
0/
#683300000000
1!
1'
1/
#683310000000
0!
1"
0'
1(
0/
10
#683320000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#683330000000
0!
0'
0/
#683340000000
1!
1'
1/
#683350000000
0!
0'
0/
#683360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#683370000000
0!
0'
0/
#683380000000
1!
1'
1/
#683390000000
0!
1"
0'
1(
0/
10
#683400000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#683410000000
0!
1$
0'
1+
0/
#683420000000
1!
1'
1/
#683430000000
0!
0'
0/
#683440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#683450000000
0!
0'
0/
#683460000000
1!
1'
1/
#683470000000
0!
0'
0/
#683480000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#683490000000
0!
0'
0/
#683500000000
1!
1'
1/
#683510000000
0!
0'
0/
#683520000000
1!
1'
1/
#683530000000
0!
0'
0/
#683540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#683550000000
0!
0'
0/
#683560000000
1!
1'
1/
#683570000000
0!
0'
0/
#683580000000
1!
1'
1/
#683590000000
0!
0'
0/
#683600000000
1!
1'
1/
#683610000000
0!
0'
0/
#683620000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#683630000000
0!
0'
0/
#683640000000
1!
1'
1/
#683650000000
0!
0'
0/
#683660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#683670000000
0!
0'
0/
#683680000000
1!
1'
1/
#683690000000
0!
0'
0/
#683700000000
#683710000000
1!
1'
1/
#683720000000
0!
0'
0/
#683730000000
1!
1'
1/
#683740000000
0!
1"
0'
1(
0/
10
#683750000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#683760000000
0!
0'
0/
#683770000000
1!
1'
1/
#683780000000
0!
0'
0/
#683790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#683800000000
0!
0'
0/
#683810000000
1!
1'
1/
#683820000000
0!
1"
0'
1(
0/
10
#683830000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#683840000000
0!
1$
0'
1+
0/
#683850000000
1!
1'
1/
#683860000000
0!
0'
0/
#683870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#683880000000
0!
0'
0/
#683890000000
1!
1'
1/
#683900000000
0!
0'
0/
#683910000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#683920000000
0!
0'
0/
#683930000000
1!
1'
1/
#683940000000
0!
0'
0/
#683950000000
1!
1'
1/
#683960000000
0!
0'
0/
#683970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#683980000000
0!
0'
0/
#683990000000
1!
1'
1/
#684000000000
0!
0'
0/
#684010000000
1!
1'
1/
#684020000000
0!
0'
0/
#684030000000
1!
1'
1/
#684040000000
0!
0'
0/
#684050000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#684060000000
0!
0'
0/
#684070000000
1!
1'
1/
#684080000000
0!
0'
0/
#684090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#684100000000
0!
0'
0/
#684110000000
1!
1'
1/
#684120000000
0!
0'
0/
#684130000000
#684140000000
1!
1'
1/
#684150000000
0!
0'
0/
#684160000000
1!
1'
1/
#684170000000
0!
1"
0'
1(
0/
10
#684180000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#684190000000
0!
0'
0/
#684200000000
1!
1'
1/
#684210000000
0!
0'
0/
#684220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#684230000000
0!
0'
0/
#684240000000
1!
1'
1/
#684250000000
0!
1"
0'
1(
0/
10
#684260000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#684270000000
0!
1$
0'
1+
0/
#684280000000
1!
1'
1/
#684290000000
0!
0'
0/
#684300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#684310000000
0!
0'
0/
#684320000000
1!
1'
1/
#684330000000
0!
0'
0/
#684340000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#684350000000
0!
0'
0/
#684360000000
1!
1'
1/
#684370000000
0!
0'
0/
#684380000000
1!
1'
1/
#684390000000
0!
0'
0/
#684400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#684410000000
0!
0'
0/
#684420000000
1!
1'
1/
#684430000000
0!
0'
0/
#684440000000
1!
1'
1/
#684450000000
0!
0'
0/
#684460000000
1!
1'
1/
#684470000000
0!
0'
0/
#684480000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#684490000000
0!
0'
0/
#684500000000
1!
1'
1/
#684510000000
0!
0'
0/
#684520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#684530000000
0!
0'
0/
#684540000000
1!
1'
1/
#684550000000
0!
0'
0/
#684560000000
#684570000000
1!
1'
1/
#684580000000
0!
0'
0/
#684590000000
1!
1'
1/
#684600000000
0!
1"
0'
1(
0/
10
#684610000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#684620000000
0!
0'
0/
#684630000000
1!
1'
1/
#684640000000
0!
0'
0/
#684650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#684660000000
0!
0'
0/
#684670000000
1!
1'
1/
#684680000000
0!
1"
0'
1(
0/
10
#684690000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#684700000000
0!
1$
0'
1+
0/
#684710000000
1!
1'
1/
#684720000000
0!
0'
0/
#684730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#684740000000
0!
0'
0/
#684750000000
1!
1'
1/
#684760000000
0!
0'
0/
#684770000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#684780000000
0!
0'
0/
#684790000000
1!
1'
1/
#684800000000
0!
0'
0/
#684810000000
1!
1'
1/
#684820000000
0!
0'
0/
#684830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#684840000000
0!
0'
0/
#684850000000
1!
1'
1/
#684860000000
0!
0'
0/
#684870000000
1!
1'
1/
#684880000000
0!
0'
0/
#684890000000
1!
1'
1/
#684900000000
0!
0'
0/
#684910000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#684920000000
0!
0'
0/
#684930000000
1!
1'
1/
#684940000000
0!
0'
0/
#684950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#684960000000
0!
0'
0/
#684970000000
1!
1'
1/
#684980000000
0!
0'
0/
#684990000000
#685000000000
1!
1'
1/
#685010000000
0!
0'
0/
#685020000000
1!
1'
1/
#685030000000
0!
1"
0'
1(
0/
10
#685040000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#685050000000
0!
0'
0/
#685060000000
1!
1'
1/
#685070000000
0!
0'
0/
#685080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#685090000000
0!
0'
0/
#685100000000
1!
1'
1/
#685110000000
0!
1"
0'
1(
0/
10
#685120000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#685130000000
0!
1$
0'
1+
0/
#685140000000
1!
1'
1/
#685150000000
0!
0'
0/
#685160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#685170000000
0!
0'
0/
#685180000000
1!
1'
1/
#685190000000
0!
0'
0/
#685200000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#685210000000
0!
0'
0/
#685220000000
1!
1'
1/
#685230000000
0!
0'
0/
#685240000000
1!
1'
1/
#685250000000
0!
0'
0/
#685260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#685270000000
0!
0'
0/
#685280000000
1!
1'
1/
#685290000000
0!
0'
0/
#685300000000
1!
1'
1/
#685310000000
0!
0'
0/
#685320000000
1!
1'
1/
#685330000000
0!
0'
0/
#685340000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#685350000000
0!
0'
0/
#685360000000
1!
1'
1/
#685370000000
0!
0'
0/
#685380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#685390000000
0!
0'
0/
#685400000000
1!
1'
1/
#685410000000
0!
0'
0/
#685420000000
#685430000000
1!
1'
1/
#685440000000
0!
0'
0/
#685450000000
1!
1'
1/
#685460000000
0!
1"
0'
1(
0/
10
#685470000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#685480000000
0!
0'
0/
#685490000000
1!
1'
1/
#685500000000
0!
0'
0/
#685510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#685520000000
0!
0'
0/
#685530000000
1!
1'
1/
#685540000000
0!
1"
0'
1(
0/
10
#685550000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#685560000000
0!
1$
0'
1+
0/
#685570000000
1!
1'
1/
#685580000000
0!
0'
0/
#685590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#685600000000
0!
0'
0/
#685610000000
1!
1'
1/
#685620000000
0!
0'
0/
#685630000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#685640000000
0!
0'
0/
#685650000000
1!
1'
1/
#685660000000
0!
0'
0/
#685670000000
1!
1'
1/
#685680000000
0!
0'
0/
#685690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#685700000000
0!
0'
0/
#685710000000
1!
1'
1/
#685720000000
0!
0'
0/
#685730000000
1!
1'
1/
#685740000000
0!
0'
0/
#685750000000
1!
1'
1/
#685760000000
0!
0'
0/
#685770000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#685780000000
0!
0'
0/
#685790000000
1!
1'
1/
#685800000000
0!
0'
0/
#685810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#685820000000
0!
0'
0/
#685830000000
1!
1'
1/
#685840000000
0!
0'
0/
#685850000000
#685860000000
1!
1'
1/
#685870000000
0!
0'
0/
#685880000000
1!
1'
1/
#685890000000
0!
1"
0'
1(
0/
10
#685900000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#685910000000
0!
0'
0/
#685920000000
1!
1'
1/
#685930000000
0!
0'
0/
#685940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#685950000000
0!
0'
0/
#685960000000
1!
1'
1/
#685970000000
0!
1"
0'
1(
0/
10
#685980000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#685990000000
0!
1$
0'
1+
0/
#686000000000
1!
1'
1/
#686010000000
0!
0'
0/
#686020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#686030000000
0!
0'
0/
#686040000000
1!
1'
1/
#686050000000
0!
0'
0/
#686060000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#686070000000
0!
0'
0/
#686080000000
1!
1'
1/
#686090000000
0!
0'
0/
#686100000000
1!
1'
1/
#686110000000
0!
0'
0/
#686120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#686130000000
0!
0'
0/
#686140000000
1!
1'
1/
#686150000000
0!
0'
0/
#686160000000
1!
1'
1/
#686170000000
0!
0'
0/
#686180000000
1!
1'
1/
#686190000000
0!
0'
0/
#686200000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#686210000000
0!
0'
0/
#686220000000
1!
1'
1/
#686230000000
0!
0'
0/
#686240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#686250000000
0!
0'
0/
#686260000000
1!
1'
1/
#686270000000
0!
0'
0/
#686280000000
#686290000000
1!
1'
1/
#686300000000
0!
0'
0/
#686310000000
1!
1'
1/
#686320000000
0!
1"
0'
1(
0/
10
#686330000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#686340000000
0!
0'
0/
#686350000000
1!
1'
1/
#686360000000
0!
0'
0/
#686370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#686380000000
0!
0'
0/
#686390000000
1!
1'
1/
#686400000000
0!
1"
0'
1(
0/
10
#686410000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#686420000000
0!
1$
0'
1+
0/
#686430000000
1!
1'
1/
#686440000000
0!
0'
0/
#686450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#686460000000
0!
0'
0/
#686470000000
1!
1'
1/
#686480000000
0!
0'
0/
#686490000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#686500000000
0!
0'
0/
#686510000000
1!
1'
1/
#686520000000
0!
0'
0/
#686530000000
1!
1'
1/
#686540000000
0!
0'
0/
#686550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#686560000000
0!
0'
0/
#686570000000
1!
1'
1/
#686580000000
0!
0'
0/
#686590000000
1!
1'
1/
#686600000000
0!
0'
0/
#686610000000
1!
1'
1/
#686620000000
0!
0'
0/
#686630000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#686640000000
0!
0'
0/
#686650000000
1!
1'
1/
#686660000000
0!
0'
0/
#686670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#686680000000
0!
0'
0/
#686690000000
1!
1'
1/
#686700000000
0!
0'
0/
#686710000000
#686720000000
1!
1'
1/
#686730000000
0!
0'
0/
#686740000000
1!
1'
1/
#686750000000
0!
1"
0'
1(
0/
10
#686760000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#686770000000
0!
0'
0/
#686780000000
1!
1'
1/
#686790000000
0!
0'
0/
#686800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#686810000000
0!
0'
0/
#686820000000
1!
1'
1/
#686830000000
0!
1"
0'
1(
0/
10
#686840000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#686850000000
0!
1$
0'
1+
0/
#686860000000
1!
1'
1/
#686870000000
0!
0'
0/
#686880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#686890000000
0!
0'
0/
#686900000000
1!
1'
1/
#686910000000
0!
0'
0/
#686920000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#686930000000
0!
0'
0/
#686940000000
1!
1'
1/
#686950000000
0!
0'
0/
#686960000000
1!
1'
1/
#686970000000
0!
0'
0/
#686980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#686990000000
0!
0'
0/
#687000000000
1!
1'
1/
#687010000000
0!
0'
0/
#687020000000
1!
1'
1/
#687030000000
0!
0'
0/
#687040000000
1!
1'
1/
#687050000000
0!
0'
0/
#687060000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#687070000000
0!
0'
0/
#687080000000
1!
1'
1/
#687090000000
0!
0'
0/
#687100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#687110000000
0!
0'
0/
#687120000000
1!
1'
1/
#687130000000
0!
0'
0/
#687140000000
#687150000000
1!
1'
1/
#687160000000
0!
0'
0/
#687170000000
1!
1'
1/
#687180000000
0!
1"
0'
1(
0/
10
#687190000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#687200000000
0!
0'
0/
#687210000000
1!
1'
1/
#687220000000
0!
0'
0/
#687230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#687240000000
0!
0'
0/
#687250000000
1!
1'
1/
#687260000000
0!
1"
0'
1(
0/
10
#687270000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#687280000000
0!
1$
0'
1+
0/
#687290000000
1!
1'
1/
#687300000000
0!
0'
0/
#687310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#687320000000
0!
0'
0/
#687330000000
1!
1'
1/
#687340000000
0!
0'
0/
#687350000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#687360000000
0!
0'
0/
#687370000000
1!
1'
1/
#687380000000
0!
0'
0/
#687390000000
1!
1'
1/
#687400000000
0!
0'
0/
#687410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#687420000000
0!
0'
0/
#687430000000
1!
1'
1/
#687440000000
0!
0'
0/
#687450000000
1!
1'
1/
#687460000000
0!
0'
0/
#687470000000
1!
1'
1/
#687480000000
0!
0'
0/
#687490000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#687500000000
0!
0'
0/
#687510000000
1!
1'
1/
#687520000000
0!
0'
0/
#687530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#687540000000
0!
0'
0/
#687550000000
1!
1'
1/
#687560000000
0!
0'
0/
#687570000000
#687580000000
1!
1'
1/
#687590000000
0!
0'
0/
#687600000000
1!
1'
1/
#687610000000
0!
1"
0'
1(
0/
10
#687620000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#687630000000
0!
0'
0/
#687640000000
1!
1'
1/
#687650000000
0!
0'
0/
#687660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#687670000000
0!
0'
0/
#687680000000
1!
1'
1/
#687690000000
0!
1"
0'
1(
0/
10
#687700000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#687710000000
0!
1$
0'
1+
0/
#687720000000
1!
1'
1/
#687730000000
0!
0'
0/
#687740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#687750000000
0!
0'
0/
#687760000000
1!
1'
1/
#687770000000
0!
0'
0/
#687780000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#687790000000
0!
0'
0/
#687800000000
1!
1'
1/
#687810000000
0!
0'
0/
#687820000000
1!
1'
1/
#687830000000
0!
0'
0/
#687840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#687850000000
0!
0'
0/
#687860000000
1!
1'
1/
#687870000000
0!
0'
0/
#687880000000
1!
1'
1/
#687890000000
0!
0'
0/
#687900000000
1!
1'
1/
#687910000000
0!
0'
0/
#687920000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#687930000000
0!
0'
0/
#687940000000
1!
1'
1/
#687950000000
0!
0'
0/
#687960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#687970000000
0!
0'
0/
#687980000000
1!
1'
1/
#687990000000
0!
0'
0/
#688000000000
#688010000000
1!
1'
1/
#688020000000
0!
0'
0/
#688030000000
1!
1'
1/
#688040000000
0!
1"
0'
1(
0/
10
#688050000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#688060000000
0!
0'
0/
#688070000000
1!
1'
1/
#688080000000
0!
0'
0/
#688090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#688100000000
0!
0'
0/
#688110000000
1!
1'
1/
#688120000000
0!
1"
0'
1(
0/
10
#688130000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#688140000000
0!
1$
0'
1+
0/
#688150000000
1!
1'
1/
#688160000000
0!
0'
0/
#688170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#688180000000
0!
0'
0/
#688190000000
1!
1'
1/
#688200000000
0!
0'
0/
#688210000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#688220000000
0!
0'
0/
#688230000000
1!
1'
1/
#688240000000
0!
0'
0/
#688250000000
1!
1'
1/
#688260000000
0!
0'
0/
#688270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#688280000000
0!
0'
0/
#688290000000
1!
1'
1/
#688300000000
0!
0'
0/
#688310000000
1!
1'
1/
#688320000000
0!
0'
0/
#688330000000
1!
1'
1/
#688340000000
0!
0'
0/
#688350000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#688360000000
0!
0'
0/
#688370000000
1!
1'
1/
#688380000000
0!
0'
0/
#688390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#688400000000
0!
0'
0/
#688410000000
1!
1'
1/
#688420000000
0!
0'
0/
#688430000000
#688440000000
1!
1'
1/
#688450000000
0!
0'
0/
#688460000000
1!
1'
1/
#688470000000
0!
1"
0'
1(
0/
10
#688480000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#688490000000
0!
0'
0/
#688500000000
1!
1'
1/
#688510000000
0!
0'
0/
#688520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#688530000000
0!
0'
0/
#688540000000
1!
1'
1/
#688550000000
0!
1"
0'
1(
0/
10
#688560000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#688570000000
0!
1$
0'
1+
0/
#688580000000
1!
1'
1/
#688590000000
0!
0'
0/
#688600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#688610000000
0!
0'
0/
#688620000000
1!
1'
1/
#688630000000
0!
0'
0/
#688640000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#688650000000
0!
0'
0/
#688660000000
1!
1'
1/
#688670000000
0!
0'
0/
#688680000000
1!
1'
1/
#688690000000
0!
0'
0/
#688700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#688710000000
0!
0'
0/
#688720000000
1!
1'
1/
#688730000000
0!
0'
0/
#688740000000
1!
1'
1/
#688750000000
0!
0'
0/
#688760000000
1!
1'
1/
#688770000000
0!
0'
0/
#688780000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#688790000000
0!
0'
0/
#688800000000
1!
1'
1/
#688810000000
0!
0'
0/
#688820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#688830000000
0!
0'
0/
#688840000000
1!
1'
1/
#688850000000
0!
0'
0/
#688860000000
#688870000000
1!
1'
1/
#688880000000
0!
0'
0/
#688890000000
1!
1'
1/
#688900000000
0!
1"
0'
1(
0/
10
#688910000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#688920000000
0!
0'
0/
#688930000000
1!
1'
1/
#688940000000
0!
0'
0/
#688950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#688960000000
0!
0'
0/
#688970000000
1!
1'
1/
#688980000000
0!
1"
0'
1(
0/
10
#688990000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#689000000000
0!
1$
0'
1+
0/
#689010000000
1!
1'
1/
#689020000000
0!
0'
0/
#689030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#689040000000
0!
0'
0/
#689050000000
1!
1'
1/
#689060000000
0!
0'
0/
#689070000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#689080000000
0!
0'
0/
#689090000000
1!
1'
1/
#689100000000
0!
0'
0/
#689110000000
1!
1'
1/
#689120000000
0!
0'
0/
#689130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#689140000000
0!
0'
0/
#689150000000
1!
1'
1/
#689160000000
0!
0'
0/
#689170000000
1!
1'
1/
#689180000000
0!
0'
0/
#689190000000
1!
1'
1/
#689200000000
0!
0'
0/
#689210000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#689220000000
0!
0'
0/
#689230000000
1!
1'
1/
#689240000000
0!
0'
0/
#689250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#689260000000
0!
0'
0/
#689270000000
1!
1'
1/
#689280000000
0!
0'
0/
#689290000000
#689300000000
1!
1'
1/
#689310000000
0!
0'
0/
#689320000000
1!
1'
1/
#689330000000
0!
1"
0'
1(
0/
10
#689340000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#689350000000
0!
0'
0/
#689360000000
1!
1'
1/
#689370000000
0!
0'
0/
#689380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#689390000000
0!
0'
0/
#689400000000
1!
1'
1/
#689410000000
0!
1"
0'
1(
0/
10
#689420000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#689430000000
0!
1$
0'
1+
0/
#689440000000
1!
1'
1/
#689450000000
0!
0'
0/
#689460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#689470000000
0!
0'
0/
#689480000000
1!
1'
1/
#689490000000
0!
0'
0/
#689500000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#689510000000
0!
0'
0/
#689520000000
1!
1'
1/
#689530000000
0!
0'
0/
#689540000000
1!
1'
1/
#689550000000
0!
0'
0/
#689560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#689570000000
0!
0'
0/
#689580000000
1!
1'
1/
#689590000000
0!
0'
0/
#689600000000
1!
1'
1/
#689610000000
0!
0'
0/
#689620000000
1!
1'
1/
#689630000000
0!
0'
0/
#689640000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#689650000000
0!
0'
0/
#689660000000
1!
1'
1/
#689670000000
0!
0'
0/
#689680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#689690000000
0!
0'
0/
#689700000000
1!
1'
1/
#689710000000
0!
0'
0/
#689720000000
#689730000000
1!
1'
1/
#689740000000
0!
0'
0/
#689750000000
1!
1'
1/
#689760000000
0!
1"
0'
1(
0/
10
#689770000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#689780000000
0!
0'
0/
#689790000000
1!
1'
1/
#689800000000
0!
0'
0/
#689810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#689820000000
0!
0'
0/
#689830000000
1!
1'
1/
#689840000000
0!
1"
0'
1(
0/
10
#689850000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#689860000000
0!
1$
0'
1+
0/
#689870000000
1!
1'
1/
#689880000000
0!
0'
0/
#689890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#689900000000
0!
0'
0/
#689910000000
1!
1'
1/
#689920000000
0!
0'
0/
#689930000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#689940000000
0!
0'
0/
#689950000000
1!
1'
1/
#689960000000
0!
0'
0/
#689970000000
1!
1'
1/
#689980000000
0!
0'
0/
#689990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#690000000000
0!
0'
0/
#690010000000
1!
1'
1/
#690020000000
0!
0'
0/
#690030000000
1!
1'
1/
#690040000000
0!
0'
0/
#690050000000
1!
1'
1/
#690060000000
0!
0'
0/
#690070000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#690080000000
0!
0'
0/
#690090000000
1!
1'
1/
#690100000000
0!
0'
0/
#690110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#690120000000
0!
0'
0/
#690130000000
1!
1'
1/
#690140000000
0!
0'
0/
#690150000000
#690160000000
1!
1'
1/
#690170000000
0!
0'
0/
#690180000000
1!
1'
1/
#690190000000
0!
1"
0'
1(
0/
10
#690200000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#690210000000
0!
0'
0/
#690220000000
1!
1'
1/
#690230000000
0!
0'
0/
#690240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#690250000000
0!
0'
0/
#690260000000
1!
1'
1/
#690270000000
0!
1"
0'
1(
0/
10
#690280000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#690290000000
0!
1$
0'
1+
0/
#690300000000
1!
1'
1/
#690310000000
0!
0'
0/
#690320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#690330000000
0!
0'
0/
#690340000000
1!
1'
1/
#690350000000
0!
0'
0/
#690360000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#690370000000
0!
0'
0/
#690380000000
1!
1'
1/
#690390000000
0!
0'
0/
#690400000000
1!
1'
1/
#690410000000
0!
0'
0/
#690420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#690430000000
0!
0'
0/
#690440000000
1!
1'
1/
#690450000000
0!
0'
0/
#690460000000
1!
1'
1/
#690470000000
0!
0'
0/
#690480000000
1!
1'
1/
#690490000000
0!
0'
0/
#690500000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#690510000000
0!
0'
0/
#690520000000
1!
1'
1/
#690530000000
0!
0'
0/
#690540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#690550000000
0!
0'
0/
#690560000000
1!
1'
1/
#690570000000
0!
0'
0/
#690580000000
#690590000000
1!
1'
1/
#690600000000
0!
0'
0/
#690610000000
1!
1'
1/
#690620000000
0!
1"
0'
1(
0/
10
#690630000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#690640000000
0!
0'
0/
#690650000000
1!
1'
1/
#690660000000
0!
0'
0/
#690670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#690680000000
0!
0'
0/
#690690000000
1!
1'
1/
#690700000000
0!
1"
0'
1(
0/
10
#690710000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#690720000000
0!
1$
0'
1+
0/
#690730000000
1!
1'
1/
#690740000000
0!
0'
0/
#690750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#690760000000
0!
0'
0/
#690770000000
1!
1'
1/
#690780000000
0!
0'
0/
#690790000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#690800000000
0!
0'
0/
#690810000000
1!
1'
1/
#690820000000
0!
0'
0/
#690830000000
1!
1'
1/
#690840000000
0!
0'
0/
#690850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#690860000000
0!
0'
0/
#690870000000
1!
1'
1/
#690880000000
0!
0'
0/
#690890000000
1!
1'
1/
#690900000000
0!
0'
0/
#690910000000
1!
1'
1/
#690920000000
0!
0'
0/
#690930000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#690940000000
0!
0'
0/
#690950000000
1!
1'
1/
#690960000000
0!
0'
0/
#690970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#690980000000
0!
0'
0/
#690990000000
1!
1'
1/
#691000000000
0!
0'
0/
#691010000000
#691020000000
1!
1'
1/
#691030000000
0!
0'
0/
#691040000000
1!
1'
1/
#691050000000
0!
1"
0'
1(
0/
10
#691060000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#691070000000
0!
0'
0/
#691080000000
1!
1'
1/
#691090000000
0!
0'
0/
#691100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#691110000000
0!
0'
0/
#691120000000
1!
1'
1/
#691130000000
0!
1"
0'
1(
0/
10
#691140000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#691150000000
0!
1$
0'
1+
0/
#691160000000
1!
1'
1/
#691170000000
0!
0'
0/
#691180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#691190000000
0!
0'
0/
#691200000000
1!
1'
1/
#691210000000
0!
0'
0/
#691220000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#691230000000
0!
0'
0/
#691240000000
1!
1'
1/
#691250000000
0!
0'
0/
#691260000000
1!
1'
1/
#691270000000
0!
0'
0/
#691280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#691290000000
0!
0'
0/
#691300000000
1!
1'
1/
#691310000000
0!
0'
0/
#691320000000
1!
1'
1/
#691330000000
0!
0'
0/
#691340000000
1!
1'
1/
#691350000000
0!
0'
0/
#691360000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#691370000000
0!
0'
0/
#691380000000
1!
1'
1/
#691390000000
0!
0'
0/
#691400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#691410000000
0!
0'
0/
#691420000000
1!
1'
1/
#691430000000
0!
0'
0/
#691440000000
#691450000000
1!
1'
1/
#691460000000
0!
0'
0/
#691470000000
1!
1'
1/
#691480000000
0!
1"
0'
1(
0/
10
#691490000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#691500000000
0!
0'
0/
#691510000000
1!
1'
1/
#691520000000
0!
0'
0/
#691530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#691540000000
0!
0'
0/
#691550000000
1!
1'
1/
#691560000000
0!
1"
0'
1(
0/
10
#691570000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#691580000000
0!
1$
0'
1+
0/
#691590000000
1!
1'
1/
#691600000000
0!
0'
0/
#691610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#691620000000
0!
0'
0/
#691630000000
1!
1'
1/
#691640000000
0!
0'
0/
#691650000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#691660000000
0!
0'
0/
#691670000000
1!
1'
1/
#691680000000
0!
0'
0/
#691690000000
1!
1'
1/
#691700000000
0!
0'
0/
#691710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#691720000000
0!
0'
0/
#691730000000
1!
1'
1/
#691740000000
0!
0'
0/
#691750000000
1!
1'
1/
#691760000000
0!
0'
0/
#691770000000
1!
1'
1/
#691780000000
0!
0'
0/
#691790000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#691800000000
0!
0'
0/
#691810000000
1!
1'
1/
#691820000000
0!
0'
0/
#691830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#691840000000
0!
0'
0/
#691850000000
1!
1'
1/
#691860000000
0!
0'
0/
#691870000000
#691880000000
1!
1'
1/
#691890000000
0!
0'
0/
#691900000000
1!
1'
1/
#691910000000
0!
1"
0'
1(
0/
10
#691920000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#691930000000
0!
0'
0/
#691940000000
1!
1'
1/
#691950000000
0!
0'
0/
#691960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#691970000000
0!
0'
0/
#691980000000
1!
1'
1/
#691990000000
0!
1"
0'
1(
0/
10
#692000000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#692010000000
0!
1$
0'
1+
0/
#692020000000
1!
1'
1/
#692030000000
0!
0'
0/
#692040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#692050000000
0!
0'
0/
#692060000000
1!
1'
1/
#692070000000
0!
0'
0/
#692080000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#692090000000
0!
0'
0/
#692100000000
1!
1'
1/
#692110000000
0!
0'
0/
#692120000000
1!
1'
1/
#692130000000
0!
0'
0/
#692140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#692150000000
0!
0'
0/
#692160000000
1!
1'
1/
#692170000000
0!
0'
0/
#692180000000
1!
1'
1/
#692190000000
0!
0'
0/
#692200000000
1!
1'
1/
#692210000000
0!
0'
0/
#692220000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#692230000000
0!
0'
0/
#692240000000
1!
1'
1/
#692250000000
0!
0'
0/
#692260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#692270000000
0!
0'
0/
#692280000000
1!
1'
1/
#692290000000
0!
0'
0/
#692300000000
#692310000000
1!
1'
1/
#692320000000
0!
0'
0/
#692330000000
1!
1'
1/
#692340000000
0!
1"
0'
1(
0/
10
#692350000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#692360000000
0!
0'
0/
#692370000000
1!
1'
1/
#692380000000
0!
0'
0/
#692390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#692400000000
0!
0'
0/
#692410000000
1!
1'
1/
#692420000000
0!
1"
0'
1(
0/
10
#692430000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#692440000000
0!
1$
0'
1+
0/
#692450000000
1!
1'
1/
#692460000000
0!
0'
0/
#692470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#692480000000
0!
0'
0/
#692490000000
1!
1'
1/
#692500000000
0!
0'
0/
#692510000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#692520000000
0!
0'
0/
#692530000000
1!
1'
1/
#692540000000
0!
0'
0/
#692550000000
1!
1'
1/
#692560000000
0!
0'
0/
#692570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#692580000000
0!
0'
0/
#692590000000
1!
1'
1/
#692600000000
0!
0'
0/
#692610000000
1!
1'
1/
#692620000000
0!
0'
0/
#692630000000
1!
1'
1/
#692640000000
0!
0'
0/
#692650000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#692660000000
0!
0'
0/
#692670000000
1!
1'
1/
#692680000000
0!
0'
0/
#692690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#692700000000
0!
0'
0/
#692710000000
1!
1'
1/
#692720000000
0!
0'
0/
#692730000000
#692740000000
1!
1'
1/
#692750000000
0!
0'
0/
#692760000000
1!
1'
1/
#692770000000
0!
1"
0'
1(
0/
10
#692780000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#692790000000
0!
0'
0/
#692800000000
1!
1'
1/
#692810000000
0!
0'
0/
#692820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#692830000000
0!
0'
0/
#692840000000
1!
1'
1/
#692850000000
0!
1"
0'
1(
0/
10
#692860000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#692870000000
0!
1$
0'
1+
0/
#692880000000
1!
1'
1/
#692890000000
0!
0'
0/
#692900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#692910000000
0!
0'
0/
#692920000000
1!
1'
1/
#692930000000
0!
0'
0/
#692940000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#692950000000
0!
0'
0/
#692960000000
1!
1'
1/
#692970000000
0!
0'
0/
#692980000000
1!
1'
1/
#692990000000
0!
0'
0/
#693000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#693010000000
0!
0'
0/
#693020000000
1!
1'
1/
#693030000000
0!
0'
0/
#693040000000
1!
1'
1/
#693050000000
0!
0'
0/
#693060000000
1!
1'
1/
#693070000000
0!
0'
0/
#693080000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#693090000000
0!
0'
0/
#693100000000
1!
1'
1/
#693110000000
0!
0'
0/
#693120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#693130000000
0!
0'
0/
#693140000000
1!
1'
1/
#693150000000
0!
0'
0/
#693160000000
#693170000000
1!
1'
1/
#693180000000
0!
0'
0/
#693190000000
1!
1'
1/
#693200000000
0!
1"
0'
1(
0/
10
#693210000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#693220000000
0!
0'
0/
#693230000000
1!
1'
1/
#693240000000
0!
0'
0/
#693250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#693260000000
0!
0'
0/
#693270000000
1!
1'
1/
#693280000000
0!
1"
0'
1(
0/
10
#693290000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#693300000000
0!
1$
0'
1+
0/
#693310000000
1!
1'
1/
#693320000000
0!
0'
0/
#693330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#693340000000
0!
0'
0/
#693350000000
1!
1'
1/
#693360000000
0!
0'
0/
#693370000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#693380000000
0!
0'
0/
#693390000000
1!
1'
1/
#693400000000
0!
0'
0/
#693410000000
1!
1'
1/
#693420000000
0!
0'
0/
#693430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#693440000000
0!
0'
0/
#693450000000
1!
1'
1/
#693460000000
0!
0'
0/
#693470000000
1!
1'
1/
#693480000000
0!
0'
0/
#693490000000
1!
1'
1/
#693500000000
0!
0'
0/
#693510000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#693520000000
0!
0'
0/
#693530000000
1!
1'
1/
#693540000000
0!
0'
0/
#693550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#693560000000
0!
0'
0/
#693570000000
1!
1'
1/
#693580000000
0!
0'
0/
#693590000000
#693600000000
1!
1'
1/
#693610000000
0!
0'
0/
#693620000000
1!
1'
1/
#693630000000
0!
1"
0'
1(
0/
10
#693640000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#693650000000
0!
0'
0/
#693660000000
1!
1'
1/
#693670000000
0!
0'
0/
#693680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#693690000000
0!
0'
0/
#693700000000
1!
1'
1/
#693710000000
0!
1"
0'
1(
0/
10
#693720000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#693730000000
0!
1$
0'
1+
0/
#693740000000
1!
1'
1/
#693750000000
0!
0'
0/
#693760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#693770000000
0!
0'
0/
#693780000000
1!
1'
1/
#693790000000
0!
0'
0/
#693800000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#693810000000
0!
0'
0/
#693820000000
1!
1'
1/
#693830000000
0!
0'
0/
#693840000000
1!
1'
1/
#693850000000
0!
0'
0/
#693860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#693870000000
0!
0'
0/
#693880000000
1!
1'
1/
#693890000000
0!
0'
0/
#693900000000
1!
1'
1/
#693910000000
0!
0'
0/
#693920000000
1!
1'
1/
#693930000000
0!
0'
0/
#693940000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#693950000000
0!
0'
0/
#693960000000
1!
1'
1/
#693970000000
0!
0'
0/
#693980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#693990000000
0!
0'
0/
#694000000000
1!
1'
1/
#694010000000
0!
0'
0/
#694020000000
#694030000000
1!
1'
1/
#694040000000
0!
0'
0/
#694050000000
1!
1'
1/
#694060000000
0!
1"
0'
1(
0/
10
#694070000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#694080000000
0!
0'
0/
#694090000000
1!
1'
1/
#694100000000
0!
0'
0/
#694110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#694120000000
0!
0'
0/
#694130000000
1!
1'
1/
#694140000000
0!
1"
0'
1(
0/
10
#694150000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#694160000000
0!
1$
0'
1+
0/
#694170000000
1!
1'
1/
#694180000000
0!
0'
0/
#694190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#694200000000
0!
0'
0/
#694210000000
1!
1'
1/
#694220000000
0!
0'
0/
#694230000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#694240000000
0!
0'
0/
#694250000000
1!
1'
1/
#694260000000
0!
0'
0/
#694270000000
1!
1'
1/
#694280000000
0!
0'
0/
#694290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#694300000000
0!
0'
0/
#694310000000
1!
1'
1/
#694320000000
0!
0'
0/
#694330000000
1!
1'
1/
#694340000000
0!
0'
0/
#694350000000
1!
1'
1/
#694360000000
0!
0'
0/
#694370000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#694380000000
0!
0'
0/
#694390000000
1!
1'
1/
#694400000000
0!
0'
0/
#694410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#694420000000
0!
0'
0/
#694430000000
1!
1'
1/
#694440000000
0!
0'
0/
#694450000000
#694460000000
1!
1'
1/
#694470000000
0!
0'
0/
#694480000000
1!
1'
1/
#694490000000
0!
1"
0'
1(
0/
10
#694500000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#694510000000
0!
0'
0/
#694520000000
1!
1'
1/
#694530000000
0!
0'
0/
#694540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#694550000000
0!
0'
0/
#694560000000
1!
1'
1/
#694570000000
0!
1"
0'
1(
0/
10
#694580000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#694590000000
0!
1$
0'
1+
0/
#694600000000
1!
1'
1/
#694610000000
0!
0'
0/
#694620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#694630000000
0!
0'
0/
#694640000000
1!
1'
1/
#694650000000
0!
0'
0/
#694660000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#694670000000
0!
0'
0/
#694680000000
1!
1'
1/
#694690000000
0!
0'
0/
#694700000000
1!
1'
1/
#694710000000
0!
0'
0/
#694720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#694730000000
0!
0'
0/
#694740000000
1!
1'
1/
#694750000000
0!
0'
0/
#694760000000
1!
1'
1/
#694770000000
0!
0'
0/
#694780000000
1!
1'
1/
#694790000000
0!
0'
0/
#694800000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#694810000000
0!
0'
0/
#694820000000
1!
1'
1/
#694830000000
0!
0'
0/
#694840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#694850000000
0!
0'
0/
#694860000000
1!
1'
1/
#694870000000
0!
0'
0/
#694880000000
#694890000000
1!
1'
1/
#694900000000
0!
0'
0/
#694910000000
1!
1'
1/
#694920000000
0!
1"
0'
1(
0/
10
#694930000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#694940000000
0!
0'
0/
#694950000000
1!
1'
1/
#694960000000
0!
0'
0/
#694970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#694980000000
0!
0'
0/
#694990000000
1!
1'
1/
#695000000000
0!
1"
0'
1(
0/
10
#695010000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#695020000000
0!
1$
0'
1+
0/
#695030000000
1!
1'
1/
#695040000000
0!
0'
0/
#695050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#695060000000
0!
0'
0/
#695070000000
1!
1'
1/
#695080000000
0!
0'
0/
#695090000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#695100000000
0!
0'
0/
#695110000000
1!
1'
1/
#695120000000
0!
0'
0/
#695130000000
1!
1'
1/
#695140000000
0!
0'
0/
#695150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#695160000000
0!
0'
0/
#695170000000
1!
1'
1/
#695180000000
0!
0'
0/
#695190000000
1!
1'
1/
#695200000000
0!
0'
0/
#695210000000
1!
1'
1/
#695220000000
0!
0'
0/
#695230000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#695240000000
0!
0'
0/
#695250000000
1!
1'
1/
#695260000000
0!
0'
0/
#695270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#695280000000
0!
0'
0/
#695290000000
1!
1'
1/
#695300000000
0!
0'
0/
#695310000000
#695320000000
1!
1'
1/
#695330000000
0!
0'
0/
#695340000000
1!
1'
1/
#695350000000
0!
1"
0'
1(
0/
10
#695360000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#695370000000
0!
0'
0/
#695380000000
1!
1'
1/
#695390000000
0!
0'
0/
#695400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#695410000000
0!
0'
0/
#695420000000
1!
1'
1/
#695430000000
0!
1"
0'
1(
0/
10
#695440000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#695450000000
0!
1$
0'
1+
0/
#695460000000
1!
1'
1/
#695470000000
0!
0'
0/
#695480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#695490000000
0!
0'
0/
#695500000000
1!
1'
1/
#695510000000
0!
0'
0/
#695520000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#695530000000
0!
0'
0/
#695540000000
1!
1'
1/
#695550000000
0!
0'
0/
#695560000000
1!
1'
1/
#695570000000
0!
0'
0/
#695580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#695590000000
0!
0'
0/
#695600000000
1!
1'
1/
#695610000000
0!
0'
0/
#695620000000
1!
1'
1/
#695630000000
0!
0'
0/
#695640000000
1!
1'
1/
#695650000000
0!
0'
0/
#695660000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#695670000000
0!
0'
0/
#695680000000
1!
1'
1/
#695690000000
0!
0'
0/
#695700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#695710000000
0!
0'
0/
#695720000000
1!
1'
1/
#695730000000
0!
0'
0/
#695740000000
#695750000000
1!
1'
1/
#695760000000
0!
0'
0/
#695770000000
1!
1'
1/
#695780000000
0!
1"
0'
1(
0/
10
#695790000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#695800000000
0!
0'
0/
#695810000000
1!
1'
1/
#695820000000
0!
0'
0/
#695830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#695840000000
0!
0'
0/
#695850000000
1!
1'
1/
#695860000000
0!
1"
0'
1(
0/
10
#695870000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#695880000000
0!
1$
0'
1+
0/
#695890000000
1!
1'
1/
#695900000000
0!
0'
0/
#695910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#695920000000
0!
0'
0/
#695930000000
1!
1'
1/
#695940000000
0!
0'
0/
#695950000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#695960000000
0!
0'
0/
#695970000000
1!
1'
1/
#695980000000
0!
0'
0/
#695990000000
1!
1'
1/
#696000000000
0!
0'
0/
#696010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#696020000000
0!
0'
0/
#696030000000
1!
1'
1/
#696040000000
0!
0'
0/
#696050000000
1!
1'
1/
#696060000000
0!
0'
0/
#696070000000
1!
1'
1/
#696080000000
0!
0'
0/
#696090000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#696100000000
0!
0'
0/
#696110000000
1!
1'
1/
#696120000000
0!
0'
0/
#696130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#696140000000
0!
0'
0/
#696150000000
1!
1'
1/
#696160000000
0!
0'
0/
#696170000000
#696180000000
1!
1'
1/
#696190000000
0!
0'
0/
#696200000000
1!
1'
1/
#696210000000
0!
1"
0'
1(
0/
10
#696220000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#696230000000
0!
0'
0/
#696240000000
1!
1'
1/
#696250000000
0!
0'
0/
#696260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#696270000000
0!
0'
0/
#696280000000
1!
1'
1/
#696290000000
0!
1"
0'
1(
0/
10
#696300000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#696310000000
0!
1$
0'
1+
0/
#696320000000
1!
1'
1/
#696330000000
0!
0'
0/
#696340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#696350000000
0!
0'
0/
#696360000000
1!
1'
1/
#696370000000
0!
0'
0/
#696380000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#696390000000
0!
0'
0/
#696400000000
1!
1'
1/
#696410000000
0!
0'
0/
#696420000000
1!
1'
1/
#696430000000
0!
0'
0/
#696440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#696450000000
0!
0'
0/
#696460000000
1!
1'
1/
#696470000000
0!
0'
0/
#696480000000
1!
1'
1/
#696490000000
0!
0'
0/
#696500000000
1!
1'
1/
#696510000000
0!
0'
0/
#696520000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#696530000000
0!
0'
0/
#696540000000
1!
1'
1/
#696550000000
0!
0'
0/
#696560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#696570000000
0!
0'
0/
#696580000000
1!
1'
1/
#696590000000
0!
0'
0/
#696600000000
#696610000000
1!
1'
1/
#696620000000
0!
0'
0/
#696630000000
1!
1'
1/
#696640000000
0!
1"
0'
1(
0/
10
#696650000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#696660000000
0!
0'
0/
#696670000000
1!
1'
1/
#696680000000
0!
0'
0/
#696690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#696700000000
0!
0'
0/
#696710000000
1!
1'
1/
#696720000000
0!
1"
0'
1(
0/
10
#696730000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#696740000000
0!
1$
0'
1+
0/
#696750000000
1!
1'
1/
#696760000000
0!
0'
0/
#696770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#696780000000
0!
0'
0/
#696790000000
1!
1'
1/
#696800000000
0!
0'
0/
#696810000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#696820000000
0!
0'
0/
#696830000000
1!
1'
1/
#696840000000
0!
0'
0/
#696850000000
1!
1'
1/
#696860000000
0!
0'
0/
#696870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#696880000000
0!
0'
0/
#696890000000
1!
1'
1/
#696900000000
0!
0'
0/
#696910000000
1!
1'
1/
#696920000000
0!
0'
0/
#696930000000
1!
1'
1/
#696940000000
0!
0'
0/
#696950000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#696960000000
0!
0'
0/
#696970000000
1!
1'
1/
#696980000000
0!
0'
0/
#696990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#697000000000
0!
0'
0/
#697010000000
1!
1'
1/
#697020000000
0!
0'
0/
#697030000000
#697040000000
1!
1'
1/
#697050000000
0!
0'
0/
#697060000000
1!
1'
1/
#697070000000
0!
1"
0'
1(
0/
10
#697080000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#697090000000
0!
0'
0/
#697100000000
1!
1'
1/
#697110000000
0!
0'
0/
#697120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#697130000000
0!
0'
0/
#697140000000
1!
1'
1/
#697150000000
0!
1"
0'
1(
0/
10
#697160000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#697170000000
0!
1$
0'
1+
0/
#697180000000
1!
1'
1/
#697190000000
0!
0'
0/
#697200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#697210000000
0!
0'
0/
#697220000000
1!
1'
1/
#697230000000
0!
0'
0/
#697240000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#697250000000
0!
0'
0/
#697260000000
1!
1'
1/
#697270000000
0!
0'
0/
#697280000000
1!
1'
1/
#697290000000
0!
0'
0/
#697300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#697310000000
0!
0'
0/
#697320000000
1!
1'
1/
#697330000000
0!
0'
0/
#697340000000
1!
1'
1/
#697350000000
0!
0'
0/
#697360000000
1!
1'
1/
#697370000000
0!
0'
0/
#697380000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#697390000000
0!
0'
0/
#697400000000
1!
1'
1/
#697410000000
0!
0'
0/
#697420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#697430000000
0!
0'
0/
#697440000000
1!
1'
1/
#697450000000
0!
0'
0/
#697460000000
#697470000000
1!
1'
1/
#697480000000
0!
0'
0/
#697490000000
1!
1'
1/
#697500000000
0!
1"
0'
1(
0/
10
#697510000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#697520000000
0!
0'
0/
#697530000000
1!
1'
1/
#697540000000
0!
0'
0/
#697550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#697560000000
0!
0'
0/
#697570000000
1!
1'
1/
#697580000000
0!
1"
0'
1(
0/
10
#697590000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#697600000000
0!
1$
0'
1+
0/
#697610000000
1!
1'
1/
#697620000000
0!
0'
0/
#697630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#697640000000
0!
0'
0/
#697650000000
1!
1'
1/
#697660000000
0!
0'
0/
#697670000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#697680000000
0!
0'
0/
#697690000000
1!
1'
1/
#697700000000
0!
0'
0/
#697710000000
1!
1'
1/
#697720000000
0!
0'
0/
#697730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#697740000000
0!
0'
0/
#697750000000
1!
1'
1/
#697760000000
0!
0'
0/
#697770000000
1!
1'
1/
#697780000000
0!
0'
0/
#697790000000
1!
1'
1/
#697800000000
0!
0'
0/
#697810000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#697820000000
0!
0'
0/
#697830000000
1!
1'
1/
#697840000000
0!
0'
0/
#697850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#697860000000
0!
0'
0/
#697870000000
1!
1'
1/
#697880000000
0!
0'
0/
#697890000000
#697900000000
1!
1'
1/
#697910000000
0!
0'
0/
#697920000000
1!
1'
1/
#697930000000
0!
1"
0'
1(
0/
10
#697940000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#697950000000
0!
0'
0/
#697960000000
1!
1'
1/
#697970000000
0!
0'
0/
#697980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#697990000000
0!
0'
0/
#698000000000
1!
1'
1/
#698010000000
0!
1"
0'
1(
0/
10
#698020000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#698030000000
0!
1$
0'
1+
0/
#698040000000
1!
1'
1/
#698050000000
0!
0'
0/
#698060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#698070000000
0!
0'
0/
#698080000000
1!
1'
1/
#698090000000
0!
0'
0/
#698100000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#698110000000
0!
0'
0/
#698120000000
1!
1'
1/
#698130000000
0!
0'
0/
#698140000000
1!
1'
1/
#698150000000
0!
0'
0/
#698160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#698170000000
0!
0'
0/
#698180000000
1!
1'
1/
#698190000000
0!
0'
0/
#698200000000
1!
1'
1/
#698210000000
0!
0'
0/
#698220000000
1!
1'
1/
#698230000000
0!
0'
0/
#698240000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#698250000000
0!
0'
0/
#698260000000
1!
1'
1/
#698270000000
0!
0'
0/
#698280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#698290000000
0!
0'
0/
#698300000000
1!
1'
1/
#698310000000
0!
0'
0/
#698320000000
#698330000000
1!
1'
1/
#698340000000
0!
0'
0/
#698350000000
1!
1'
1/
#698360000000
0!
1"
0'
1(
0/
10
#698370000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#698380000000
0!
0'
0/
#698390000000
1!
1'
1/
#698400000000
0!
0'
0/
#698410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#698420000000
0!
0'
0/
#698430000000
1!
1'
1/
#698440000000
0!
1"
0'
1(
0/
10
#698450000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#698460000000
0!
1$
0'
1+
0/
#698470000000
1!
1'
1/
#698480000000
0!
0'
0/
#698490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#698500000000
0!
0'
0/
#698510000000
1!
1'
1/
#698520000000
0!
0'
0/
#698530000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#698540000000
0!
0'
0/
#698550000000
1!
1'
1/
#698560000000
0!
0'
0/
#698570000000
1!
1'
1/
#698580000000
0!
0'
0/
#698590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#698600000000
0!
0'
0/
#698610000000
1!
1'
1/
#698620000000
0!
0'
0/
#698630000000
1!
1'
1/
#698640000000
0!
0'
0/
#698650000000
1!
1'
1/
#698660000000
0!
0'
0/
#698670000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#698680000000
0!
0'
0/
#698690000000
1!
1'
1/
#698700000000
0!
0'
0/
#698710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#698720000000
0!
0'
0/
#698730000000
1!
1'
1/
#698740000000
0!
0'
0/
#698750000000
#698760000000
1!
1'
1/
#698770000000
0!
0'
0/
#698780000000
1!
1'
1/
#698790000000
0!
1"
0'
1(
0/
10
#698800000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#698810000000
0!
0'
0/
#698820000000
1!
1'
1/
#698830000000
0!
0'
0/
#698840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#698850000000
0!
0'
0/
#698860000000
1!
1'
1/
#698870000000
0!
1"
0'
1(
0/
10
#698880000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#698890000000
0!
1$
0'
1+
0/
#698900000000
1!
1'
1/
#698910000000
0!
0'
0/
#698920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#698930000000
0!
0'
0/
#698940000000
1!
1'
1/
#698950000000
0!
0'
0/
#698960000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#698970000000
0!
0'
0/
#698980000000
1!
1'
1/
#698990000000
0!
0'
0/
#699000000000
1!
1'
1/
#699010000000
0!
0'
0/
#699020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#699030000000
0!
0'
0/
#699040000000
1!
1'
1/
#699050000000
0!
0'
0/
#699060000000
1!
1'
1/
#699070000000
0!
0'
0/
#699080000000
1!
1'
1/
#699090000000
0!
0'
0/
#699100000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#699110000000
0!
0'
0/
#699120000000
1!
1'
1/
#699130000000
0!
0'
0/
#699140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#699150000000
0!
0'
0/
#699160000000
1!
1'
1/
#699170000000
0!
0'
0/
#699180000000
#699190000000
1!
1'
1/
#699200000000
0!
0'
0/
#699210000000
1!
1'
1/
#699220000000
0!
1"
0'
1(
0/
10
#699230000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#699240000000
0!
0'
0/
#699250000000
1!
1'
1/
#699260000000
0!
0'
0/
#699270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#699280000000
0!
0'
0/
#699290000000
1!
1'
1/
#699300000000
0!
1"
0'
1(
0/
10
#699310000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#699320000000
0!
1$
0'
1+
0/
#699330000000
1!
1'
1/
#699340000000
0!
0'
0/
#699350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#699360000000
0!
0'
0/
#699370000000
1!
1'
1/
#699380000000
0!
0'
0/
#699390000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#699400000000
0!
0'
0/
#699410000000
1!
1'
1/
#699420000000
0!
0'
0/
#699430000000
1!
1'
1/
#699440000000
0!
0'
0/
#699450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#699460000000
0!
0'
0/
#699470000000
1!
1'
1/
#699480000000
0!
0'
0/
#699490000000
1!
1'
1/
#699500000000
0!
0'
0/
#699510000000
1!
1'
1/
#699520000000
0!
0'
0/
#699530000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#699540000000
0!
0'
0/
#699550000000
1!
1'
1/
#699560000000
0!
0'
0/
#699570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#699580000000
0!
0'
0/
#699590000000
1!
1'
1/
#699600000000
0!
0'
0/
#699610000000
#699620000000
1!
1'
1/
#699630000000
0!
0'
0/
#699640000000
1!
1'
1/
#699650000000
0!
1"
0'
1(
0/
10
#699660000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#699670000000
0!
0'
0/
#699680000000
1!
1'
1/
#699690000000
0!
0'
0/
#699700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#699710000000
0!
0'
0/
#699720000000
1!
1'
1/
#699730000000
0!
1"
0'
1(
0/
10
#699740000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#699750000000
0!
1$
0'
1+
0/
#699760000000
1!
1'
1/
#699770000000
0!
0'
0/
#699780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#699790000000
0!
0'
0/
#699800000000
1!
1'
1/
#699810000000
0!
0'
0/
#699820000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#699830000000
0!
0'
0/
#699840000000
1!
1'
1/
#699850000000
0!
0'
0/
#699860000000
1!
1'
1/
#699870000000
0!
0'
0/
#699880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#699890000000
0!
0'
0/
#699900000000
1!
1'
1/
#699910000000
0!
0'
0/
#699920000000
1!
1'
1/
#699930000000
0!
0'
0/
#699940000000
1!
1'
1/
#699950000000
0!
0'
0/
#699960000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#699970000000
0!
0'
0/
#699980000000
1!
1'
1/
#699990000000
0!
0'
0/
#700000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#700010000000
0!
0'
0/
#700020000000
1!
1'
1/
#700030000000
0!
0'
0/
#700040000000
#700050000000
1!
1'
1/
#700060000000
0!
0'
0/
#700070000000
1!
1'
1/
#700080000000
0!
1"
0'
1(
0/
10
#700090000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#700100000000
0!
0'
0/
#700110000000
1!
1'
1/
#700120000000
0!
0'
0/
#700130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#700140000000
0!
0'
0/
#700150000000
1!
1'
1/
#700160000000
0!
1"
0'
1(
0/
10
#700170000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#700180000000
0!
1$
0'
1+
0/
#700190000000
1!
1'
1/
#700200000000
0!
0'
0/
#700210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#700220000000
0!
0'
0/
#700230000000
1!
1'
1/
#700240000000
0!
0'
0/
#700250000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#700260000000
0!
0'
0/
#700270000000
1!
1'
1/
#700280000000
0!
0'
0/
#700290000000
1!
1'
1/
#700300000000
0!
0'
0/
#700310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#700320000000
0!
0'
0/
#700330000000
1!
1'
1/
#700340000000
0!
0'
0/
#700350000000
1!
1'
1/
#700360000000
0!
0'
0/
#700370000000
1!
1'
1/
#700380000000
0!
0'
0/
#700390000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#700400000000
0!
0'
0/
#700410000000
1!
1'
1/
#700420000000
0!
0'
0/
#700430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#700440000000
0!
0'
0/
#700450000000
1!
1'
1/
#700460000000
0!
0'
0/
#700470000000
#700480000000
1!
1'
1/
#700490000000
0!
0'
0/
#700500000000
1!
1'
1/
#700510000000
0!
1"
0'
1(
0/
10
#700520000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#700530000000
0!
0'
0/
#700540000000
1!
1'
1/
#700550000000
0!
0'
0/
#700560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#700570000000
0!
0'
0/
#700580000000
1!
1'
1/
#700590000000
0!
1"
0'
1(
0/
10
#700600000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#700610000000
0!
1$
0'
1+
0/
#700620000000
1!
1'
1/
#700630000000
0!
0'
0/
#700640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#700650000000
0!
0'
0/
#700660000000
1!
1'
1/
#700670000000
0!
0'
0/
#700680000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#700690000000
0!
0'
0/
#700700000000
1!
1'
1/
#700710000000
0!
0'
0/
#700720000000
1!
1'
1/
#700730000000
0!
0'
0/
#700740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#700750000000
0!
0'
0/
#700760000000
1!
1'
1/
#700770000000
0!
0'
0/
#700780000000
1!
1'
1/
#700790000000
0!
0'
0/
#700800000000
1!
1'
1/
#700810000000
0!
0'
0/
#700820000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#700830000000
0!
0'
0/
#700840000000
1!
1'
1/
#700850000000
0!
0'
0/
#700860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#700870000000
0!
0'
0/
#700880000000
1!
1'
1/
#700890000000
0!
0'
0/
#700900000000
#700910000000
1!
1'
1/
#700920000000
0!
0'
0/
#700930000000
1!
1'
1/
#700940000000
0!
1"
0'
1(
0/
10
#700950000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#700960000000
0!
0'
0/
#700970000000
1!
1'
1/
#700980000000
0!
0'
0/
#700990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#701000000000
0!
0'
0/
#701010000000
1!
1'
1/
#701020000000
0!
1"
0'
1(
0/
10
#701030000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#701040000000
0!
1$
0'
1+
0/
#701050000000
1!
1'
1/
#701060000000
0!
0'
0/
#701070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#701080000000
0!
0'
0/
#701090000000
1!
1'
1/
#701100000000
0!
0'
0/
#701110000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#701120000000
0!
0'
0/
#701130000000
1!
1'
1/
#701140000000
0!
0'
0/
#701150000000
1!
1'
1/
#701160000000
0!
0'
0/
#701170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#701180000000
0!
0'
0/
#701190000000
1!
1'
1/
#701200000000
0!
0'
0/
#701210000000
1!
1'
1/
#701220000000
0!
0'
0/
#701230000000
1!
1'
1/
#701240000000
0!
0'
0/
#701250000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#701260000000
0!
0'
0/
#701270000000
1!
1'
1/
#701280000000
0!
0'
0/
#701290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#701300000000
0!
0'
0/
#701310000000
1!
1'
1/
#701320000000
0!
0'
0/
#701330000000
#701340000000
1!
1'
1/
#701350000000
0!
0'
0/
#701360000000
1!
1'
1/
#701370000000
0!
1"
0'
1(
0/
10
#701380000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#701390000000
0!
0'
0/
#701400000000
1!
1'
1/
#701410000000
0!
0'
0/
#701420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#701430000000
0!
0'
0/
#701440000000
1!
1'
1/
#701450000000
0!
1"
0'
1(
0/
10
#701460000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#701470000000
0!
1$
0'
1+
0/
#701480000000
1!
1'
1/
#701490000000
0!
0'
0/
#701500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#701510000000
0!
0'
0/
#701520000000
1!
1'
1/
#701530000000
0!
0'
0/
#701540000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#701550000000
0!
0'
0/
#701560000000
1!
1'
1/
#701570000000
0!
0'
0/
#701580000000
1!
1'
1/
#701590000000
0!
0'
0/
#701600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#701610000000
0!
0'
0/
#701620000000
1!
1'
1/
#701630000000
0!
0'
0/
#701640000000
1!
1'
1/
#701650000000
0!
0'
0/
#701660000000
1!
1'
1/
#701670000000
0!
0'
0/
#701680000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#701690000000
0!
0'
0/
#701700000000
1!
1'
1/
#701710000000
0!
0'
0/
#701720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#701730000000
0!
0'
0/
#701740000000
1!
1'
1/
#701750000000
0!
0'
0/
#701760000000
#701770000000
1!
1'
1/
#701780000000
0!
0'
0/
#701790000000
1!
1'
1/
#701800000000
0!
1"
0'
1(
0/
10
#701810000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#701820000000
0!
0'
0/
#701830000000
1!
1'
1/
#701840000000
0!
0'
0/
#701850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#701860000000
0!
0'
0/
#701870000000
1!
1'
1/
#701880000000
0!
1"
0'
1(
0/
10
#701890000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#701900000000
0!
1$
0'
1+
0/
#701910000000
1!
1'
1/
#701920000000
0!
0'
0/
#701930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#701940000000
0!
0'
0/
#701950000000
1!
1'
1/
#701960000000
0!
0'
0/
#701970000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#701980000000
0!
0'
0/
#701990000000
1!
1'
1/
#702000000000
0!
0'
0/
#702010000000
1!
1'
1/
#702020000000
0!
0'
0/
#702030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#702040000000
0!
0'
0/
#702050000000
1!
1'
1/
#702060000000
0!
0'
0/
#702070000000
1!
1'
1/
#702080000000
0!
0'
0/
#702090000000
1!
1'
1/
#702100000000
0!
0'
0/
#702110000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#702120000000
0!
0'
0/
#702130000000
1!
1'
1/
#702140000000
0!
0'
0/
#702150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#702160000000
0!
0'
0/
#702170000000
1!
1'
1/
#702180000000
0!
0'
0/
#702190000000
#702200000000
1!
1'
1/
#702210000000
0!
0'
0/
#702220000000
1!
1'
1/
#702230000000
0!
1"
0'
1(
0/
10
#702240000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#702250000000
0!
0'
0/
#702260000000
1!
1'
1/
#702270000000
0!
0'
0/
#702280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#702290000000
0!
0'
0/
#702300000000
1!
1'
1/
#702310000000
0!
1"
0'
1(
0/
10
#702320000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#702330000000
0!
1$
0'
1+
0/
#702340000000
1!
1'
1/
#702350000000
0!
0'
0/
#702360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#702370000000
0!
0'
0/
#702380000000
1!
1'
1/
#702390000000
0!
0'
0/
#702400000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#702410000000
0!
0'
0/
#702420000000
1!
1'
1/
#702430000000
0!
0'
0/
#702440000000
1!
1'
1/
#702450000000
0!
0'
0/
#702460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#702470000000
0!
0'
0/
#702480000000
1!
1'
1/
#702490000000
0!
0'
0/
#702500000000
1!
1'
1/
#702510000000
0!
0'
0/
#702520000000
1!
1'
1/
#702530000000
0!
0'
0/
#702540000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#702550000000
0!
0'
0/
#702560000000
1!
1'
1/
#702570000000
0!
0'
0/
#702580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#702590000000
0!
0'
0/
#702600000000
1!
1'
1/
#702610000000
0!
0'
0/
#702620000000
#702630000000
1!
1'
1/
#702640000000
0!
0'
0/
#702650000000
1!
1'
1/
#702660000000
0!
1"
0'
1(
0/
10
#702670000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#702680000000
0!
0'
0/
#702690000000
1!
1'
1/
#702700000000
0!
0'
0/
#702710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#702720000000
0!
0'
0/
#702730000000
1!
1'
1/
#702740000000
0!
1"
0'
1(
0/
10
#702750000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#702760000000
0!
1$
0'
1+
0/
#702770000000
1!
1'
1/
#702780000000
0!
0'
0/
#702790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#702800000000
0!
0'
0/
#702810000000
1!
1'
1/
#702820000000
0!
0'
0/
#702830000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#702840000000
0!
0'
0/
#702850000000
1!
1'
1/
#702860000000
0!
0'
0/
#702870000000
1!
1'
1/
#702880000000
0!
0'
0/
#702890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#702900000000
0!
0'
0/
#702910000000
1!
1'
1/
#702920000000
0!
0'
0/
#702930000000
1!
1'
1/
#702940000000
0!
0'
0/
#702950000000
1!
1'
1/
#702960000000
0!
0'
0/
#702970000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#702980000000
0!
0'
0/
#702990000000
1!
1'
1/
#703000000000
0!
0'
0/
#703010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#703020000000
0!
0'
0/
#703030000000
1!
1'
1/
#703040000000
0!
0'
0/
#703050000000
#703060000000
1!
1'
1/
#703070000000
0!
0'
0/
#703080000000
1!
1'
1/
#703090000000
0!
1"
0'
1(
0/
10
#703100000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#703110000000
0!
0'
0/
#703120000000
1!
1'
1/
#703130000000
0!
0'
0/
#703140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#703150000000
0!
0'
0/
#703160000000
1!
1'
1/
#703170000000
0!
1"
0'
1(
0/
10
#703180000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#703190000000
0!
1$
0'
1+
0/
#703200000000
1!
1'
1/
#703210000000
0!
0'
0/
#703220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#703230000000
0!
0'
0/
#703240000000
1!
1'
1/
#703250000000
0!
0'
0/
#703260000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#703270000000
0!
0'
0/
#703280000000
1!
1'
1/
#703290000000
0!
0'
0/
#703300000000
1!
1'
1/
#703310000000
0!
0'
0/
#703320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#703330000000
0!
0'
0/
#703340000000
1!
1'
1/
#703350000000
0!
0'
0/
#703360000000
1!
1'
1/
#703370000000
0!
0'
0/
#703380000000
1!
1'
1/
#703390000000
0!
0'
0/
#703400000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#703410000000
0!
0'
0/
#703420000000
1!
1'
1/
#703430000000
0!
0'
0/
#703440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#703450000000
0!
0'
0/
#703460000000
1!
1'
1/
#703470000000
0!
0'
0/
#703480000000
#703490000000
1!
1'
1/
#703500000000
0!
0'
0/
#703510000000
1!
1'
1/
#703520000000
0!
1"
0'
1(
0/
10
#703530000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#703540000000
0!
0'
0/
#703550000000
1!
1'
1/
#703560000000
0!
0'
0/
#703570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#703580000000
0!
0'
0/
#703590000000
1!
1'
1/
#703600000000
0!
1"
0'
1(
0/
10
#703610000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#703620000000
0!
1$
0'
1+
0/
#703630000000
1!
1'
1/
#703640000000
0!
0'
0/
#703650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#703660000000
0!
0'
0/
#703670000000
1!
1'
1/
#703680000000
0!
0'
0/
#703690000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#703700000000
0!
0'
0/
#703710000000
1!
1'
1/
#703720000000
0!
0'
0/
#703730000000
1!
1'
1/
#703740000000
0!
0'
0/
#703750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#703760000000
0!
0'
0/
#703770000000
1!
1'
1/
#703780000000
0!
0'
0/
#703790000000
1!
1'
1/
#703800000000
0!
0'
0/
#703810000000
1!
1'
1/
#703820000000
0!
0'
0/
#703830000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#703840000000
0!
0'
0/
#703850000000
1!
1'
1/
#703860000000
0!
0'
0/
#703870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#703880000000
0!
0'
0/
#703890000000
1!
1'
1/
#703900000000
0!
0'
0/
#703910000000
#703920000000
1!
1'
1/
#703930000000
0!
0'
0/
#703940000000
1!
1'
1/
#703950000000
0!
1"
0'
1(
0/
10
#703960000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#703970000000
0!
0'
0/
#703980000000
1!
1'
1/
#703990000000
0!
0'
0/
#704000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#704010000000
0!
0'
0/
#704020000000
1!
1'
1/
#704030000000
0!
1"
0'
1(
0/
10
#704040000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#704050000000
0!
1$
0'
1+
0/
#704060000000
1!
1'
1/
#704070000000
0!
0'
0/
#704080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#704090000000
0!
0'
0/
#704100000000
1!
1'
1/
#704110000000
0!
0'
0/
#704120000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#704130000000
0!
0'
0/
#704140000000
1!
1'
1/
#704150000000
0!
0'
0/
#704160000000
1!
1'
1/
#704170000000
0!
0'
0/
#704180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#704190000000
0!
0'
0/
#704200000000
1!
1'
1/
#704210000000
0!
0'
0/
#704220000000
1!
1'
1/
#704230000000
0!
0'
0/
#704240000000
1!
1'
1/
#704250000000
0!
0'
0/
#704260000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#704270000000
0!
0'
0/
#704280000000
1!
1'
1/
#704290000000
0!
0'
0/
#704300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#704310000000
0!
0'
0/
#704320000000
1!
1'
1/
#704330000000
0!
0'
0/
#704340000000
#704350000000
1!
1'
1/
#704360000000
0!
0'
0/
#704370000000
1!
1'
1/
#704380000000
0!
1"
0'
1(
0/
10
#704390000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#704400000000
0!
0'
0/
#704410000000
1!
1'
1/
#704420000000
0!
0'
0/
#704430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#704440000000
0!
0'
0/
#704450000000
1!
1'
1/
#704460000000
0!
1"
0'
1(
0/
10
#704470000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#704480000000
0!
1$
0'
1+
0/
#704490000000
1!
1'
1/
#704500000000
0!
0'
0/
#704510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#704520000000
0!
0'
0/
#704530000000
1!
1'
1/
#704540000000
0!
0'
0/
#704550000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#704560000000
0!
0'
0/
#704570000000
1!
1'
1/
#704580000000
0!
0'
0/
#704590000000
1!
1'
1/
#704600000000
0!
0'
0/
#704610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#704620000000
0!
0'
0/
#704630000000
1!
1'
1/
#704640000000
0!
0'
0/
#704650000000
1!
1'
1/
#704660000000
0!
0'
0/
#704670000000
1!
1'
1/
#704680000000
0!
0'
0/
#704690000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#704700000000
0!
0'
0/
#704710000000
1!
1'
1/
#704720000000
0!
0'
0/
#704730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#704740000000
0!
0'
0/
#704750000000
1!
1'
1/
#704760000000
0!
0'
0/
#704770000000
#704780000000
1!
1'
1/
#704790000000
0!
0'
0/
#704800000000
1!
1'
1/
#704810000000
0!
1"
0'
1(
0/
10
#704820000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#704830000000
0!
0'
0/
#704840000000
1!
1'
1/
#704850000000
0!
0'
0/
#704860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#704870000000
0!
0'
0/
#704880000000
1!
1'
1/
#704890000000
0!
1"
0'
1(
0/
10
#704900000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#704910000000
0!
1$
0'
1+
0/
#704920000000
1!
1'
1/
#704930000000
0!
0'
0/
#704940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#704950000000
0!
0'
0/
#704960000000
1!
1'
1/
#704970000000
0!
0'
0/
#704980000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#704990000000
0!
0'
0/
#705000000000
1!
1'
1/
#705010000000
0!
0'
0/
#705020000000
1!
1'
1/
#705030000000
0!
0'
0/
#705040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#705050000000
0!
0'
0/
#705060000000
1!
1'
1/
#705070000000
0!
0'
0/
#705080000000
1!
1'
1/
#705090000000
0!
0'
0/
#705100000000
1!
1'
1/
#705110000000
0!
0'
0/
#705120000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#705130000000
0!
0'
0/
#705140000000
1!
1'
1/
#705150000000
0!
0'
0/
#705160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#705170000000
0!
0'
0/
#705180000000
1!
1'
1/
#705190000000
0!
0'
0/
#705200000000
#705210000000
1!
1'
1/
#705220000000
0!
0'
0/
#705230000000
1!
1'
1/
#705240000000
0!
1"
0'
1(
0/
10
#705250000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#705260000000
0!
0'
0/
#705270000000
1!
1'
1/
#705280000000
0!
0'
0/
#705290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#705300000000
0!
0'
0/
#705310000000
1!
1'
1/
#705320000000
0!
1"
0'
1(
0/
10
#705330000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#705340000000
0!
1$
0'
1+
0/
#705350000000
1!
1'
1/
#705360000000
0!
0'
0/
#705370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#705380000000
0!
0'
0/
#705390000000
1!
1'
1/
#705400000000
0!
0'
0/
#705410000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#705420000000
0!
0'
0/
#705430000000
1!
1'
1/
#705440000000
0!
0'
0/
#705450000000
1!
1'
1/
#705460000000
0!
0'
0/
#705470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#705480000000
0!
0'
0/
#705490000000
1!
1'
1/
#705500000000
0!
0'
0/
#705510000000
1!
1'
1/
#705520000000
0!
0'
0/
#705530000000
1!
1'
1/
#705540000000
0!
0'
0/
#705550000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#705560000000
0!
0'
0/
#705570000000
1!
1'
1/
#705580000000
0!
0'
0/
#705590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#705600000000
0!
0'
0/
#705610000000
1!
1'
1/
#705620000000
0!
0'
0/
#705630000000
#705640000000
1!
1'
1/
#705650000000
0!
0'
0/
#705660000000
1!
1'
1/
#705670000000
0!
1"
0'
1(
0/
10
#705680000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#705690000000
0!
0'
0/
#705700000000
1!
1'
1/
#705710000000
0!
0'
0/
#705720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#705730000000
0!
0'
0/
#705740000000
1!
1'
1/
#705750000000
0!
1"
0'
1(
0/
10
#705760000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#705770000000
0!
1$
0'
1+
0/
#705780000000
1!
1'
1/
#705790000000
0!
0'
0/
#705800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#705810000000
0!
0'
0/
#705820000000
1!
1'
1/
#705830000000
0!
0'
0/
#705840000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#705850000000
0!
0'
0/
#705860000000
1!
1'
1/
#705870000000
0!
0'
0/
#705880000000
1!
1'
1/
#705890000000
0!
0'
0/
#705900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#705910000000
0!
0'
0/
#705920000000
1!
1'
1/
#705930000000
0!
0'
0/
#705940000000
1!
1'
1/
#705950000000
0!
0'
0/
#705960000000
1!
1'
1/
#705970000000
0!
0'
0/
#705980000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#705990000000
0!
0'
0/
#706000000000
1!
1'
1/
#706010000000
0!
0'
0/
#706020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#706030000000
0!
0'
0/
#706040000000
1!
1'
1/
#706050000000
0!
0'
0/
#706060000000
#706070000000
1!
1'
1/
#706080000000
0!
0'
0/
#706090000000
1!
1'
1/
#706100000000
0!
1"
0'
1(
0/
10
#706110000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#706120000000
0!
0'
0/
#706130000000
1!
1'
1/
#706140000000
0!
0'
0/
#706150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#706160000000
0!
0'
0/
#706170000000
1!
1'
1/
#706180000000
0!
1"
0'
1(
0/
10
#706190000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#706200000000
0!
1$
0'
1+
0/
#706210000000
1!
1'
1/
#706220000000
0!
0'
0/
#706230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#706240000000
0!
0'
0/
#706250000000
1!
1'
1/
#706260000000
0!
0'
0/
#706270000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#706280000000
0!
0'
0/
#706290000000
1!
1'
1/
#706300000000
0!
0'
0/
#706310000000
1!
1'
1/
#706320000000
0!
0'
0/
#706330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#706340000000
0!
0'
0/
#706350000000
1!
1'
1/
#706360000000
0!
0'
0/
#706370000000
1!
1'
1/
#706380000000
0!
0'
0/
#706390000000
1!
1'
1/
#706400000000
0!
0'
0/
#706410000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#706420000000
0!
0'
0/
#706430000000
1!
1'
1/
#706440000000
0!
0'
0/
#706450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#706460000000
0!
0'
0/
#706470000000
1!
1'
1/
#706480000000
0!
0'
0/
#706490000000
#706500000000
1!
1'
1/
#706510000000
0!
0'
0/
#706520000000
1!
1'
1/
#706530000000
0!
1"
0'
1(
0/
10
#706540000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#706550000000
0!
0'
0/
#706560000000
1!
1'
1/
#706570000000
0!
0'
0/
#706580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#706590000000
0!
0'
0/
#706600000000
1!
1'
1/
#706610000000
0!
1"
0'
1(
0/
10
#706620000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#706630000000
0!
1$
0'
1+
0/
#706640000000
1!
1'
1/
#706650000000
0!
0'
0/
#706660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#706670000000
0!
0'
0/
#706680000000
1!
1'
1/
#706690000000
0!
0'
0/
#706700000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#706710000000
0!
0'
0/
#706720000000
1!
1'
1/
#706730000000
0!
0'
0/
#706740000000
1!
1'
1/
#706750000000
0!
0'
0/
#706760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#706770000000
0!
0'
0/
#706780000000
1!
1'
1/
#706790000000
0!
0'
0/
#706800000000
1!
1'
1/
#706810000000
0!
0'
0/
#706820000000
1!
1'
1/
#706830000000
0!
0'
0/
#706840000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#706850000000
0!
0'
0/
#706860000000
1!
1'
1/
#706870000000
0!
0'
0/
#706880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#706890000000
0!
0'
0/
#706900000000
1!
1'
1/
#706910000000
0!
0'
0/
#706920000000
#706930000000
1!
1'
1/
#706940000000
0!
0'
0/
#706950000000
1!
1'
1/
#706960000000
0!
1"
0'
1(
0/
10
#706970000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#706980000000
0!
0'
0/
#706990000000
1!
1'
1/
#707000000000
0!
0'
0/
#707010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#707020000000
0!
0'
0/
#707030000000
1!
1'
1/
#707040000000
0!
1"
0'
1(
0/
10
#707050000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#707060000000
0!
1$
0'
1+
0/
#707070000000
1!
1'
1/
#707080000000
0!
0'
0/
#707090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#707100000000
0!
0'
0/
#707110000000
1!
1'
1/
#707120000000
0!
0'
0/
#707130000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#707140000000
0!
0'
0/
#707150000000
1!
1'
1/
#707160000000
0!
0'
0/
#707170000000
1!
1'
1/
#707180000000
0!
0'
0/
#707190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#707200000000
0!
0'
0/
#707210000000
1!
1'
1/
#707220000000
0!
0'
0/
#707230000000
1!
1'
1/
#707240000000
0!
0'
0/
#707250000000
1!
1'
1/
#707260000000
0!
0'
0/
#707270000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#707280000000
0!
0'
0/
#707290000000
1!
1'
1/
#707300000000
0!
0'
0/
#707310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#707320000000
0!
0'
0/
#707330000000
1!
1'
1/
#707340000000
0!
0'
0/
#707350000000
#707360000000
1!
1'
1/
#707370000000
0!
0'
0/
#707380000000
1!
1'
1/
#707390000000
0!
1"
0'
1(
0/
10
#707400000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#707410000000
0!
0'
0/
#707420000000
1!
1'
1/
#707430000000
0!
0'
0/
#707440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#707450000000
0!
0'
0/
#707460000000
1!
1'
1/
#707470000000
0!
1"
0'
1(
0/
10
#707480000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#707490000000
0!
1$
0'
1+
0/
#707500000000
1!
1'
1/
#707510000000
0!
0'
0/
#707520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#707530000000
0!
0'
0/
#707540000000
1!
1'
1/
#707550000000
0!
0'
0/
#707560000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#707570000000
0!
0'
0/
#707580000000
1!
1'
1/
#707590000000
0!
0'
0/
#707600000000
1!
1'
1/
#707610000000
0!
0'
0/
#707620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#707630000000
0!
0'
0/
#707640000000
1!
1'
1/
#707650000000
0!
0'
0/
#707660000000
1!
1'
1/
#707670000000
0!
0'
0/
#707680000000
1!
1'
1/
#707690000000
0!
0'
0/
#707700000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#707710000000
0!
0'
0/
#707720000000
1!
1'
1/
#707730000000
0!
0'
0/
#707740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#707750000000
0!
0'
0/
#707760000000
1!
1'
1/
#707770000000
0!
0'
0/
#707780000000
#707790000000
1!
1'
1/
#707800000000
0!
0'
0/
#707810000000
1!
1'
1/
#707820000000
0!
1"
0'
1(
0/
10
#707830000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#707840000000
0!
0'
0/
#707850000000
1!
1'
1/
#707860000000
0!
0'
0/
#707870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#707880000000
0!
0'
0/
#707890000000
1!
1'
1/
#707900000000
0!
1"
0'
1(
0/
10
#707910000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#707920000000
0!
1$
0'
1+
0/
#707930000000
1!
1'
1/
#707940000000
0!
0'
0/
#707950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#707960000000
0!
0'
0/
#707970000000
1!
1'
1/
#707980000000
0!
0'
0/
#707990000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#708000000000
0!
0'
0/
#708010000000
1!
1'
1/
#708020000000
0!
0'
0/
#708030000000
1!
1'
1/
#708040000000
0!
0'
0/
#708050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#708060000000
0!
0'
0/
#708070000000
1!
1'
1/
#708080000000
0!
0'
0/
#708090000000
1!
1'
1/
#708100000000
0!
0'
0/
#708110000000
1!
1'
1/
#708120000000
0!
0'
0/
#708130000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#708140000000
0!
0'
0/
#708150000000
1!
1'
1/
#708160000000
0!
0'
0/
#708170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#708180000000
0!
0'
0/
#708190000000
1!
1'
1/
#708200000000
0!
0'
0/
#708210000000
#708220000000
1!
1'
1/
#708230000000
0!
0'
0/
#708240000000
1!
1'
1/
#708250000000
0!
1"
0'
1(
0/
10
#708260000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#708270000000
0!
0'
0/
#708280000000
1!
1'
1/
#708290000000
0!
0'
0/
#708300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#708310000000
0!
0'
0/
#708320000000
1!
1'
1/
#708330000000
0!
1"
0'
1(
0/
10
#708340000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#708350000000
0!
1$
0'
1+
0/
#708360000000
1!
1'
1/
#708370000000
0!
0'
0/
#708380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#708390000000
0!
0'
0/
#708400000000
1!
1'
1/
#708410000000
0!
0'
0/
#708420000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#708430000000
0!
0'
0/
#708440000000
1!
1'
1/
#708450000000
0!
0'
0/
#708460000000
1!
1'
1/
#708470000000
0!
0'
0/
#708480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#708490000000
0!
0'
0/
#708500000000
1!
1'
1/
#708510000000
0!
0'
0/
#708520000000
1!
1'
1/
#708530000000
0!
0'
0/
#708540000000
1!
1'
1/
#708550000000
0!
0'
0/
#708560000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#708570000000
0!
0'
0/
#708580000000
1!
1'
1/
#708590000000
0!
0'
0/
#708600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#708610000000
0!
0'
0/
#708620000000
1!
1'
1/
#708630000000
0!
0'
0/
#708640000000
#708650000000
1!
1'
1/
#708660000000
0!
0'
0/
#708670000000
1!
1'
1/
#708680000000
0!
1"
0'
1(
0/
10
#708690000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#708700000000
0!
0'
0/
#708710000000
1!
1'
1/
#708720000000
0!
0'
0/
#708730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#708740000000
0!
0'
0/
#708750000000
1!
1'
1/
#708760000000
0!
1"
0'
1(
0/
10
#708770000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#708780000000
0!
1$
0'
1+
0/
#708790000000
1!
1'
1/
#708800000000
0!
0'
0/
#708810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#708820000000
0!
0'
0/
#708830000000
1!
1'
1/
#708840000000
0!
0'
0/
#708850000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#708860000000
0!
0'
0/
#708870000000
1!
1'
1/
#708880000000
0!
0'
0/
#708890000000
1!
1'
1/
#708900000000
0!
0'
0/
#708910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#708920000000
0!
0'
0/
#708930000000
1!
1'
1/
#708940000000
0!
0'
0/
#708950000000
1!
1'
1/
#708960000000
0!
0'
0/
#708970000000
1!
1'
1/
#708980000000
0!
0'
0/
#708990000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#709000000000
0!
0'
0/
#709010000000
1!
1'
1/
#709020000000
0!
0'
0/
#709030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#709040000000
0!
0'
0/
#709050000000
1!
1'
1/
#709060000000
0!
0'
0/
#709070000000
#709080000000
1!
1'
1/
#709090000000
0!
0'
0/
#709100000000
1!
1'
1/
#709110000000
0!
1"
0'
1(
0/
10
#709120000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#709130000000
0!
0'
0/
#709140000000
1!
1'
1/
#709150000000
0!
0'
0/
#709160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#709170000000
0!
0'
0/
#709180000000
1!
1'
1/
#709190000000
0!
1"
0'
1(
0/
10
#709200000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#709210000000
0!
1$
0'
1+
0/
#709220000000
1!
1'
1/
#709230000000
0!
0'
0/
#709240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#709250000000
0!
0'
0/
#709260000000
1!
1'
1/
#709270000000
0!
0'
0/
#709280000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#709290000000
0!
0'
0/
#709300000000
1!
1'
1/
#709310000000
0!
0'
0/
#709320000000
1!
1'
1/
#709330000000
0!
0'
0/
#709340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#709350000000
0!
0'
0/
#709360000000
1!
1'
1/
#709370000000
0!
0'
0/
#709380000000
1!
1'
1/
#709390000000
0!
0'
0/
#709400000000
1!
1'
1/
#709410000000
0!
0'
0/
#709420000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#709430000000
0!
0'
0/
#709440000000
1!
1'
1/
#709450000000
0!
0'
0/
#709460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#709470000000
0!
0'
0/
#709480000000
1!
1'
1/
#709490000000
0!
0'
0/
#709500000000
#709510000000
1!
1'
1/
#709520000000
0!
0'
0/
#709530000000
1!
1'
1/
#709540000000
0!
1"
0'
1(
0/
10
#709550000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#709560000000
0!
0'
0/
#709570000000
1!
1'
1/
#709580000000
0!
0'
0/
#709590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#709600000000
0!
0'
0/
#709610000000
1!
1'
1/
#709620000000
0!
1"
0'
1(
0/
10
#709630000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#709640000000
0!
1$
0'
1+
0/
#709650000000
1!
1'
1/
#709660000000
0!
0'
0/
#709670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#709680000000
0!
0'
0/
#709690000000
1!
1'
1/
#709700000000
0!
0'
0/
#709710000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#709720000000
0!
0'
0/
#709730000000
1!
1'
1/
#709740000000
0!
0'
0/
#709750000000
1!
1'
1/
#709760000000
0!
0'
0/
#709770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#709780000000
0!
0'
0/
#709790000000
1!
1'
1/
#709800000000
0!
0'
0/
#709810000000
1!
1'
1/
#709820000000
0!
0'
0/
#709830000000
1!
1'
1/
#709840000000
0!
0'
0/
#709850000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#709860000000
0!
0'
0/
#709870000000
1!
1'
1/
#709880000000
0!
0'
0/
#709890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#709900000000
0!
0'
0/
#709910000000
1!
1'
1/
#709920000000
0!
0'
0/
#709930000000
#709940000000
1!
1'
1/
#709950000000
0!
0'
0/
#709960000000
1!
1'
1/
#709970000000
0!
1"
0'
1(
0/
10
#709980000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#709990000000
0!
0'
0/
#710000000000
1!
1'
1/
#710010000000
0!
0'
0/
#710020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#710030000000
0!
0'
0/
#710040000000
1!
1'
1/
#710050000000
0!
1"
0'
1(
0/
10
#710060000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#710070000000
0!
1$
0'
1+
0/
#710080000000
1!
1'
1/
#710090000000
0!
0'
0/
#710100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#710110000000
0!
0'
0/
#710120000000
1!
1'
1/
#710130000000
0!
0'
0/
#710140000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#710150000000
0!
0'
0/
#710160000000
1!
1'
1/
#710170000000
0!
0'
0/
#710180000000
1!
1'
1/
#710190000000
0!
0'
0/
#710200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#710210000000
0!
0'
0/
#710220000000
1!
1'
1/
#710230000000
0!
0'
0/
#710240000000
1!
1'
1/
#710250000000
0!
0'
0/
#710260000000
1!
1'
1/
#710270000000
0!
0'
0/
#710280000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#710290000000
0!
0'
0/
#710300000000
1!
1'
1/
#710310000000
0!
0'
0/
#710320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#710330000000
0!
0'
0/
#710340000000
1!
1'
1/
#710350000000
0!
0'
0/
#710360000000
#710370000000
1!
1'
1/
#710380000000
0!
0'
0/
#710390000000
1!
1'
1/
#710400000000
0!
1"
0'
1(
0/
10
#710410000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#710420000000
0!
0'
0/
#710430000000
1!
1'
1/
#710440000000
0!
0'
0/
#710450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#710460000000
0!
0'
0/
#710470000000
1!
1'
1/
#710480000000
0!
1"
0'
1(
0/
10
#710490000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#710500000000
0!
1$
0'
1+
0/
#710510000000
1!
1'
1/
#710520000000
0!
0'
0/
#710530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#710540000000
0!
0'
0/
#710550000000
1!
1'
1/
#710560000000
0!
0'
0/
#710570000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#710580000000
0!
0'
0/
#710590000000
1!
1'
1/
#710600000000
0!
0'
0/
#710610000000
1!
1'
1/
#710620000000
0!
0'
0/
#710630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#710640000000
0!
0'
0/
#710650000000
1!
1'
1/
#710660000000
0!
0'
0/
#710670000000
1!
1'
1/
#710680000000
0!
0'
0/
#710690000000
1!
1'
1/
#710700000000
0!
0'
0/
#710710000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#710720000000
0!
0'
0/
#710730000000
1!
1'
1/
#710740000000
0!
0'
0/
#710750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#710760000000
0!
0'
0/
#710770000000
1!
1'
1/
#710780000000
0!
0'
0/
#710790000000
#710800000000
1!
1'
1/
#710810000000
0!
0'
0/
#710820000000
1!
1'
1/
#710830000000
0!
1"
0'
1(
0/
10
#710840000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#710850000000
0!
0'
0/
#710860000000
1!
1'
1/
#710870000000
0!
0'
0/
#710880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#710890000000
0!
0'
0/
#710900000000
1!
1'
1/
#710910000000
0!
1"
0'
1(
0/
10
#710920000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#710930000000
0!
1$
0'
1+
0/
#710940000000
1!
1'
1/
#710950000000
0!
0'
0/
#710960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#710970000000
0!
0'
0/
#710980000000
1!
1'
1/
#710990000000
0!
0'
0/
#711000000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#711010000000
0!
0'
0/
#711020000000
1!
1'
1/
#711030000000
0!
0'
0/
#711040000000
1!
1'
1/
#711050000000
0!
0'
0/
#711060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#711070000000
0!
0'
0/
#711080000000
1!
1'
1/
#711090000000
0!
0'
0/
#711100000000
1!
1'
1/
#711110000000
0!
0'
0/
#711120000000
1!
1'
1/
#711130000000
0!
0'
0/
#711140000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#711150000000
0!
0'
0/
#711160000000
1!
1'
1/
#711170000000
0!
0'
0/
#711180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#711190000000
0!
0'
0/
#711200000000
1!
1'
1/
#711210000000
0!
0'
0/
#711220000000
#711230000000
1!
1'
1/
#711240000000
0!
0'
0/
#711250000000
1!
1'
1/
#711260000000
0!
1"
0'
1(
0/
10
#711270000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#711280000000
0!
0'
0/
#711290000000
1!
1'
1/
#711300000000
0!
0'
0/
#711310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#711320000000
0!
0'
0/
#711330000000
1!
1'
1/
#711340000000
0!
1"
0'
1(
0/
10
#711350000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#711360000000
0!
1$
0'
1+
0/
#711370000000
1!
1'
1/
#711380000000
0!
0'
0/
#711390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#711400000000
0!
0'
0/
#711410000000
1!
1'
1/
#711420000000
0!
0'
0/
#711430000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#711440000000
0!
0'
0/
#711450000000
1!
1'
1/
#711460000000
0!
0'
0/
#711470000000
1!
1'
1/
#711480000000
0!
0'
0/
#711490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#711500000000
0!
0'
0/
#711510000000
1!
1'
1/
#711520000000
0!
0'
0/
#711530000000
1!
1'
1/
#711540000000
0!
0'
0/
#711550000000
1!
1'
1/
#711560000000
0!
0'
0/
#711570000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#711580000000
0!
0'
0/
#711590000000
1!
1'
1/
#711600000000
0!
0'
0/
#711610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#711620000000
0!
0'
0/
#711630000000
1!
1'
1/
#711640000000
0!
0'
0/
#711650000000
#711660000000
1!
1'
1/
#711670000000
0!
0'
0/
#711680000000
1!
1'
1/
#711690000000
0!
1"
0'
1(
0/
10
#711700000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#711710000000
0!
0'
0/
#711720000000
1!
1'
1/
#711730000000
0!
0'
0/
#711740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#711750000000
0!
0'
0/
#711760000000
1!
1'
1/
#711770000000
0!
1"
0'
1(
0/
10
#711780000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#711790000000
0!
1$
0'
1+
0/
#711800000000
1!
1'
1/
#711810000000
0!
0'
0/
#711820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#711830000000
0!
0'
0/
#711840000000
1!
1'
1/
#711850000000
0!
0'
0/
#711860000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#711870000000
0!
0'
0/
#711880000000
1!
1'
1/
#711890000000
0!
0'
0/
#711900000000
1!
1'
1/
#711910000000
0!
0'
0/
#711920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#711930000000
0!
0'
0/
#711940000000
1!
1'
1/
#711950000000
0!
0'
0/
#711960000000
1!
1'
1/
#711970000000
0!
0'
0/
#711980000000
1!
1'
1/
#711990000000
0!
0'
0/
#712000000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#712010000000
0!
0'
0/
#712020000000
1!
1'
1/
#712030000000
0!
0'
0/
#712040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#712050000000
0!
0'
0/
#712060000000
1!
1'
1/
#712070000000
0!
0'
0/
#712080000000
#712090000000
1!
1'
1/
#712100000000
0!
0'
0/
#712110000000
1!
1'
1/
#712120000000
0!
1"
0'
1(
0/
10
#712130000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#712140000000
0!
0'
0/
#712150000000
1!
1'
1/
#712160000000
0!
0'
0/
#712170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#712180000000
0!
0'
0/
#712190000000
1!
1'
1/
#712200000000
0!
1"
0'
1(
0/
10
#712210000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#712220000000
0!
1$
0'
1+
0/
#712230000000
1!
1'
1/
#712240000000
0!
0'
0/
#712250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#712260000000
0!
0'
0/
#712270000000
1!
1'
1/
#712280000000
0!
0'
0/
#712290000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#712300000000
0!
0'
0/
#712310000000
1!
1'
1/
#712320000000
0!
0'
0/
#712330000000
1!
1'
1/
#712340000000
0!
0'
0/
#712350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#712360000000
0!
0'
0/
#712370000000
1!
1'
1/
#712380000000
0!
0'
0/
#712390000000
1!
1'
1/
#712400000000
0!
0'
0/
#712410000000
1!
1'
1/
#712420000000
0!
0'
0/
#712430000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#712440000000
0!
0'
0/
#712450000000
1!
1'
1/
#712460000000
0!
0'
0/
#712470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#712480000000
0!
0'
0/
#712490000000
1!
1'
1/
#712500000000
0!
0'
0/
#712510000000
#712520000000
1!
1'
1/
#712530000000
0!
0'
0/
#712540000000
1!
1'
1/
#712550000000
0!
1"
0'
1(
0/
10
#712560000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#712570000000
0!
0'
0/
#712580000000
1!
1'
1/
#712590000000
0!
0'
0/
#712600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#712610000000
0!
0'
0/
#712620000000
1!
1'
1/
#712630000000
0!
1"
0'
1(
0/
10
#712640000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#712650000000
0!
1$
0'
1+
0/
#712660000000
1!
1'
1/
#712670000000
0!
0'
0/
#712680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#712690000000
0!
0'
0/
#712700000000
1!
1'
1/
#712710000000
0!
0'
0/
#712720000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#712730000000
0!
0'
0/
#712740000000
1!
1'
1/
#712750000000
0!
0'
0/
#712760000000
1!
1'
1/
#712770000000
0!
0'
0/
#712780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#712790000000
0!
0'
0/
#712800000000
1!
1'
1/
#712810000000
0!
0'
0/
#712820000000
1!
1'
1/
#712830000000
0!
0'
0/
#712840000000
1!
1'
1/
#712850000000
0!
0'
0/
#712860000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#712870000000
0!
0'
0/
#712880000000
1!
1'
1/
#712890000000
0!
0'
0/
#712900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#712910000000
0!
0'
0/
#712920000000
1!
1'
1/
#712930000000
0!
0'
0/
#712940000000
#712950000000
1!
1'
1/
#712960000000
0!
0'
0/
#712970000000
1!
1'
1/
#712980000000
0!
1"
0'
1(
0/
10
#712990000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#713000000000
0!
0'
0/
#713010000000
1!
1'
1/
#713020000000
0!
0'
0/
#713030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#713040000000
0!
0'
0/
#713050000000
1!
1'
1/
#713060000000
0!
1"
0'
1(
0/
10
#713070000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#713080000000
0!
1$
0'
1+
0/
#713090000000
1!
1'
1/
#713100000000
0!
0'
0/
#713110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#713120000000
0!
0'
0/
#713130000000
1!
1'
1/
#713140000000
0!
0'
0/
#713150000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#713160000000
0!
0'
0/
#713170000000
1!
1'
1/
#713180000000
0!
0'
0/
#713190000000
1!
1'
1/
#713200000000
0!
0'
0/
#713210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#713220000000
0!
0'
0/
#713230000000
1!
1'
1/
#713240000000
0!
0'
0/
#713250000000
1!
1'
1/
#713260000000
0!
0'
0/
#713270000000
1!
1'
1/
#713280000000
0!
0'
0/
#713290000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#713300000000
0!
0'
0/
#713310000000
1!
1'
1/
#713320000000
0!
0'
0/
#713330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#713340000000
0!
0'
0/
#713350000000
1!
1'
1/
#713360000000
0!
0'
0/
#713370000000
#713380000000
1!
1'
1/
#713390000000
0!
0'
0/
#713400000000
1!
1'
1/
#713410000000
0!
1"
0'
1(
0/
10
#713420000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#713430000000
0!
0'
0/
#713440000000
1!
1'
1/
#713450000000
0!
0'
0/
#713460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#713470000000
0!
0'
0/
#713480000000
1!
1'
1/
#713490000000
0!
1"
0'
1(
0/
10
#713500000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#713510000000
0!
1$
0'
1+
0/
#713520000000
1!
1'
1/
#713530000000
0!
0'
0/
#713540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#713550000000
0!
0'
0/
#713560000000
1!
1'
1/
#713570000000
0!
0'
0/
#713580000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#713590000000
0!
0'
0/
#713600000000
1!
1'
1/
#713610000000
0!
0'
0/
#713620000000
1!
1'
1/
#713630000000
0!
0'
0/
#713640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#713650000000
0!
0'
0/
#713660000000
1!
1'
1/
#713670000000
0!
0'
0/
#713680000000
1!
1'
1/
#713690000000
0!
0'
0/
#713700000000
1!
1'
1/
#713710000000
0!
0'
0/
#713720000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#713730000000
0!
0'
0/
#713740000000
1!
1'
1/
#713750000000
0!
0'
0/
#713760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#713770000000
0!
0'
0/
#713780000000
1!
1'
1/
#713790000000
0!
0'
0/
#713800000000
#713810000000
1!
1'
1/
#713820000000
0!
0'
0/
#713830000000
1!
1'
1/
#713840000000
0!
1"
0'
1(
0/
10
#713850000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#713860000000
0!
0'
0/
#713870000000
1!
1'
1/
#713880000000
0!
0'
0/
#713890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#713900000000
0!
0'
0/
#713910000000
1!
1'
1/
#713920000000
0!
1"
0'
1(
0/
10
#713930000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#713940000000
0!
1$
0'
1+
0/
#713950000000
1!
1'
1/
#713960000000
0!
0'
0/
#713970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#713980000000
0!
0'
0/
#713990000000
1!
1'
1/
#714000000000
0!
0'
0/
#714010000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#714020000000
0!
0'
0/
#714030000000
1!
1'
1/
#714040000000
0!
0'
0/
#714050000000
1!
1'
1/
#714060000000
0!
0'
0/
#714070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#714080000000
0!
0'
0/
#714090000000
1!
1'
1/
#714100000000
0!
0'
0/
#714110000000
1!
1'
1/
#714120000000
0!
0'
0/
#714130000000
1!
1'
1/
#714140000000
0!
0'
0/
#714150000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#714160000000
0!
0'
0/
#714170000000
1!
1'
1/
#714180000000
0!
0'
0/
#714190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#714200000000
0!
0'
0/
#714210000000
1!
1'
1/
#714220000000
0!
0'
0/
#714230000000
#714240000000
1!
1'
1/
#714250000000
0!
0'
0/
#714260000000
1!
1'
1/
#714270000000
0!
1"
0'
1(
0/
10
#714280000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#714290000000
0!
0'
0/
#714300000000
1!
1'
1/
#714310000000
0!
0'
0/
#714320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#714330000000
0!
0'
0/
#714340000000
1!
1'
1/
#714350000000
0!
1"
0'
1(
0/
10
#714360000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#714370000000
0!
1$
0'
1+
0/
#714380000000
1!
1'
1/
#714390000000
0!
0'
0/
#714400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#714410000000
0!
0'
0/
#714420000000
1!
1'
1/
#714430000000
0!
0'
0/
#714440000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#714450000000
0!
0'
0/
#714460000000
1!
1'
1/
#714470000000
0!
0'
0/
#714480000000
1!
1'
1/
#714490000000
0!
0'
0/
#714500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#714510000000
0!
0'
0/
#714520000000
1!
1'
1/
#714530000000
0!
0'
0/
#714540000000
1!
1'
1/
#714550000000
0!
0'
0/
#714560000000
1!
1'
1/
#714570000000
0!
0'
0/
#714580000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#714590000000
0!
0'
0/
#714600000000
1!
1'
1/
#714610000000
0!
0'
0/
#714620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#714630000000
0!
0'
0/
#714640000000
1!
1'
1/
#714650000000
0!
0'
0/
#714660000000
#714670000000
1!
1'
1/
#714680000000
0!
0'
0/
#714690000000
1!
1'
1/
#714700000000
0!
1"
0'
1(
0/
10
#714710000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#714720000000
0!
0'
0/
#714730000000
1!
1'
1/
#714740000000
0!
0'
0/
#714750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#714760000000
0!
0'
0/
#714770000000
1!
1'
1/
#714780000000
0!
1"
0'
1(
0/
10
#714790000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#714800000000
0!
1$
0'
1+
0/
#714810000000
1!
1'
1/
#714820000000
0!
0'
0/
#714830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#714840000000
0!
0'
0/
#714850000000
1!
1'
1/
#714860000000
0!
0'
0/
#714870000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#714880000000
0!
0'
0/
#714890000000
1!
1'
1/
#714900000000
0!
0'
0/
#714910000000
1!
1'
1/
#714920000000
0!
0'
0/
#714930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#714940000000
0!
0'
0/
#714950000000
1!
1'
1/
#714960000000
0!
0'
0/
#714970000000
1!
1'
1/
#714980000000
0!
0'
0/
#714990000000
1!
1'
1/
#715000000000
0!
0'
0/
#715010000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#715020000000
0!
0'
0/
#715030000000
1!
1'
1/
#715040000000
0!
0'
0/
#715050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#715060000000
0!
0'
0/
#715070000000
1!
1'
1/
#715080000000
0!
0'
0/
#715090000000
#715100000000
1!
1'
1/
#715110000000
0!
0'
0/
#715120000000
1!
1'
1/
#715130000000
0!
1"
0'
1(
0/
10
#715140000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#715150000000
0!
0'
0/
#715160000000
1!
1'
1/
#715170000000
0!
0'
0/
#715180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#715190000000
0!
0'
0/
#715200000000
1!
1'
1/
#715210000000
0!
1"
0'
1(
0/
10
#715220000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#715230000000
0!
1$
0'
1+
0/
#715240000000
1!
1'
1/
#715250000000
0!
0'
0/
#715260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#715270000000
0!
0'
0/
#715280000000
1!
1'
1/
#715290000000
0!
0'
0/
#715300000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#715310000000
0!
0'
0/
#715320000000
1!
1'
1/
#715330000000
0!
0'
0/
#715340000000
1!
1'
1/
#715350000000
0!
0'
0/
#715360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#715370000000
0!
0'
0/
#715380000000
1!
1'
1/
#715390000000
0!
0'
0/
#715400000000
1!
1'
1/
#715410000000
0!
0'
0/
#715420000000
1!
1'
1/
#715430000000
0!
0'
0/
#715440000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#715450000000
0!
0'
0/
#715460000000
1!
1'
1/
#715470000000
0!
0'
0/
#715480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#715490000000
0!
0'
0/
#715500000000
1!
1'
1/
#715510000000
0!
0'
0/
#715520000000
#715530000000
1!
1'
1/
#715540000000
0!
0'
0/
#715550000000
1!
1'
1/
#715560000000
0!
1"
0'
1(
0/
10
#715570000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#715580000000
0!
0'
0/
#715590000000
1!
1'
1/
#715600000000
0!
0'
0/
#715610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#715620000000
0!
0'
0/
#715630000000
1!
1'
1/
#715640000000
0!
1"
0'
1(
0/
10
#715650000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#715660000000
0!
1$
0'
1+
0/
#715670000000
1!
1'
1/
#715680000000
0!
0'
0/
#715690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#715700000000
0!
0'
0/
#715710000000
1!
1'
1/
#715720000000
0!
0'
0/
#715730000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#715740000000
0!
0'
0/
#715750000000
1!
1'
1/
#715760000000
0!
0'
0/
#715770000000
1!
1'
1/
#715780000000
0!
0'
0/
#715790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#715800000000
0!
0'
0/
#715810000000
1!
1'
1/
#715820000000
0!
0'
0/
#715830000000
1!
1'
1/
#715840000000
0!
0'
0/
#715850000000
1!
1'
1/
#715860000000
0!
0'
0/
#715870000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#715880000000
0!
0'
0/
#715890000000
1!
1'
1/
#715900000000
0!
0'
0/
#715910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#715920000000
0!
0'
0/
#715930000000
1!
1'
1/
#715940000000
0!
0'
0/
#715950000000
#715960000000
1!
1'
1/
#715970000000
0!
0'
0/
#715980000000
1!
1'
1/
#715990000000
0!
1"
0'
1(
0/
10
#716000000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#716010000000
0!
0'
0/
#716020000000
1!
1'
1/
#716030000000
0!
0'
0/
#716040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#716050000000
0!
0'
0/
#716060000000
1!
1'
1/
#716070000000
0!
1"
0'
1(
0/
10
#716080000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#716090000000
0!
1$
0'
1+
0/
#716100000000
1!
1'
1/
#716110000000
0!
0'
0/
#716120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#716130000000
0!
0'
0/
#716140000000
1!
1'
1/
#716150000000
0!
0'
0/
#716160000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#716170000000
0!
0'
0/
#716180000000
1!
1'
1/
#716190000000
0!
0'
0/
#716200000000
1!
1'
1/
#716210000000
0!
0'
0/
#716220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#716230000000
0!
0'
0/
#716240000000
1!
1'
1/
#716250000000
0!
0'
0/
#716260000000
1!
1'
1/
#716270000000
0!
0'
0/
#716280000000
1!
1'
1/
#716290000000
0!
0'
0/
#716300000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#716310000000
0!
0'
0/
#716320000000
1!
1'
1/
#716330000000
0!
0'
0/
#716340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#716350000000
0!
0'
0/
#716360000000
1!
1'
1/
#716370000000
0!
0'
0/
#716380000000
#716390000000
1!
1'
1/
#716400000000
0!
0'
0/
#716410000000
1!
1'
1/
#716420000000
0!
1"
0'
1(
0/
10
#716430000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#716440000000
0!
0'
0/
#716450000000
1!
1'
1/
#716460000000
0!
0'
0/
#716470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#716480000000
0!
0'
0/
#716490000000
1!
1'
1/
#716500000000
0!
1"
0'
1(
0/
10
#716510000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#716520000000
0!
1$
0'
1+
0/
#716530000000
1!
1'
1/
#716540000000
0!
0'
0/
#716550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#716560000000
0!
0'
0/
#716570000000
1!
1'
1/
#716580000000
0!
0'
0/
#716590000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#716600000000
0!
0'
0/
#716610000000
1!
1'
1/
#716620000000
0!
0'
0/
#716630000000
1!
1'
1/
#716640000000
0!
0'
0/
#716650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#716660000000
0!
0'
0/
#716670000000
1!
1'
1/
#716680000000
0!
0'
0/
#716690000000
1!
1'
1/
#716700000000
0!
0'
0/
#716710000000
1!
1'
1/
#716720000000
0!
0'
0/
#716730000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#716740000000
0!
0'
0/
#716750000000
1!
1'
1/
#716760000000
0!
0'
0/
#716770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#716780000000
0!
0'
0/
#716790000000
1!
1'
1/
#716800000000
0!
0'
0/
#716810000000
#716820000000
1!
1'
1/
#716830000000
0!
0'
0/
#716840000000
1!
1'
1/
#716850000000
0!
1"
0'
1(
0/
10
#716860000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#716870000000
0!
0'
0/
#716880000000
1!
1'
1/
#716890000000
0!
0'
0/
#716900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#716910000000
0!
0'
0/
#716920000000
1!
1'
1/
#716930000000
0!
1"
0'
1(
0/
10
#716940000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#716950000000
0!
1$
0'
1+
0/
#716960000000
1!
1'
1/
#716970000000
0!
0'
0/
#716980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#716990000000
0!
0'
0/
#717000000000
1!
1'
1/
#717010000000
0!
0'
0/
#717020000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#717030000000
0!
0'
0/
#717040000000
1!
1'
1/
#717050000000
0!
0'
0/
#717060000000
1!
1'
1/
#717070000000
0!
0'
0/
#717080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#717090000000
0!
0'
0/
#717100000000
1!
1'
1/
#717110000000
0!
0'
0/
#717120000000
1!
1'
1/
#717130000000
0!
0'
0/
#717140000000
1!
1'
1/
#717150000000
0!
0'
0/
#717160000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#717170000000
0!
0'
0/
#717180000000
1!
1'
1/
#717190000000
0!
0'
0/
#717200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#717210000000
0!
0'
0/
#717220000000
1!
1'
1/
#717230000000
0!
0'
0/
#717240000000
#717250000000
1!
1'
1/
#717260000000
0!
0'
0/
#717270000000
1!
1'
1/
#717280000000
0!
1"
0'
1(
0/
10
#717290000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#717300000000
0!
0'
0/
#717310000000
1!
1'
1/
#717320000000
0!
0'
0/
#717330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#717340000000
0!
0'
0/
#717350000000
1!
1'
1/
#717360000000
0!
1"
0'
1(
0/
10
#717370000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#717380000000
0!
1$
0'
1+
0/
#717390000000
1!
1'
1/
#717400000000
0!
0'
0/
#717410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#717420000000
0!
0'
0/
#717430000000
1!
1'
1/
#717440000000
0!
0'
0/
#717450000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#717460000000
0!
0'
0/
#717470000000
1!
1'
1/
#717480000000
0!
0'
0/
#717490000000
1!
1'
1/
#717500000000
0!
0'
0/
#717510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#717520000000
0!
0'
0/
#717530000000
1!
1'
1/
#717540000000
0!
0'
0/
#717550000000
1!
1'
1/
#717560000000
0!
0'
0/
#717570000000
1!
1'
1/
#717580000000
0!
0'
0/
#717590000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#717600000000
0!
0'
0/
#717610000000
1!
1'
1/
#717620000000
0!
0'
0/
#717630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#717640000000
0!
0'
0/
#717650000000
1!
1'
1/
#717660000000
0!
0'
0/
#717670000000
#717680000000
1!
1'
1/
#717690000000
0!
0'
0/
#717700000000
1!
1'
1/
#717710000000
0!
1"
0'
1(
0/
10
#717720000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#717730000000
0!
0'
0/
#717740000000
1!
1'
1/
#717750000000
0!
0'
0/
#717760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#717770000000
0!
0'
0/
#717780000000
1!
1'
1/
#717790000000
0!
1"
0'
1(
0/
10
#717800000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#717810000000
0!
1$
0'
1+
0/
#717820000000
1!
1'
1/
#717830000000
0!
0'
0/
#717840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#717850000000
0!
0'
0/
#717860000000
1!
1'
1/
#717870000000
0!
0'
0/
#717880000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#717890000000
0!
0'
0/
#717900000000
1!
1'
1/
#717910000000
0!
0'
0/
#717920000000
1!
1'
1/
#717930000000
0!
0'
0/
#717940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#717950000000
0!
0'
0/
#717960000000
1!
1'
1/
#717970000000
0!
0'
0/
#717980000000
1!
1'
1/
#717990000000
0!
0'
0/
#718000000000
1!
1'
1/
#718010000000
0!
0'
0/
#718020000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#718030000000
0!
0'
0/
#718040000000
1!
1'
1/
#718050000000
0!
0'
0/
#718060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#718070000000
0!
0'
0/
#718080000000
1!
1'
1/
#718090000000
0!
0'
0/
#718100000000
#718110000000
1!
1'
1/
#718120000000
0!
0'
0/
#718130000000
1!
1'
1/
#718140000000
0!
1"
0'
1(
0/
10
#718150000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#718160000000
0!
0'
0/
#718170000000
1!
1'
1/
#718180000000
0!
0'
0/
#718190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#718200000000
0!
0'
0/
#718210000000
1!
1'
1/
#718220000000
0!
1"
0'
1(
0/
10
#718230000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#718240000000
0!
1$
0'
1+
0/
#718250000000
1!
1'
1/
#718260000000
0!
0'
0/
#718270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#718280000000
0!
0'
0/
#718290000000
1!
1'
1/
#718300000000
0!
0'
0/
#718310000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#718320000000
0!
0'
0/
#718330000000
1!
1'
1/
#718340000000
0!
0'
0/
#718350000000
1!
1'
1/
#718360000000
0!
0'
0/
#718370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#718380000000
0!
0'
0/
#718390000000
1!
1'
1/
#718400000000
0!
0'
0/
#718410000000
1!
1'
1/
#718420000000
0!
0'
0/
#718430000000
1!
1'
1/
#718440000000
0!
0'
0/
#718450000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#718460000000
0!
0'
0/
#718470000000
1!
1'
1/
#718480000000
0!
0'
0/
#718490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#718500000000
0!
0'
0/
#718510000000
1!
1'
1/
#718520000000
0!
0'
0/
#718530000000
#718540000000
1!
1'
1/
#718550000000
0!
0'
0/
#718560000000
1!
1'
1/
#718570000000
0!
1"
0'
1(
0/
10
#718580000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#718590000000
0!
0'
0/
#718600000000
1!
1'
1/
#718610000000
0!
0'
0/
#718620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#718630000000
0!
0'
0/
#718640000000
1!
1'
1/
#718650000000
0!
1"
0'
1(
0/
10
#718660000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#718670000000
0!
1$
0'
1+
0/
#718680000000
1!
1'
1/
#718690000000
0!
0'
0/
#718700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#718710000000
0!
0'
0/
#718720000000
1!
1'
1/
#718730000000
0!
0'
0/
#718740000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#718750000000
0!
0'
0/
#718760000000
1!
1'
1/
#718770000000
0!
0'
0/
#718780000000
1!
1'
1/
#718790000000
0!
0'
0/
#718800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#718810000000
0!
0'
0/
#718820000000
1!
1'
1/
#718830000000
0!
0'
0/
#718840000000
1!
1'
1/
#718850000000
0!
0'
0/
#718860000000
1!
1'
1/
#718870000000
0!
0'
0/
#718880000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#718890000000
0!
0'
0/
#718900000000
1!
1'
1/
#718910000000
0!
0'
0/
#718920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#718930000000
0!
0'
0/
#718940000000
1!
1'
1/
#718950000000
0!
0'
0/
#718960000000
#718970000000
1!
1'
1/
#718980000000
0!
0'
0/
#718990000000
1!
1'
1/
#719000000000
0!
1"
0'
1(
0/
10
#719010000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#719020000000
0!
0'
0/
#719030000000
1!
1'
1/
#719040000000
0!
0'
0/
#719050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#719060000000
0!
0'
0/
#719070000000
1!
1'
1/
#719080000000
0!
1"
0'
1(
0/
10
#719090000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#719100000000
0!
1$
0'
1+
0/
#719110000000
1!
1'
1/
#719120000000
0!
0'
0/
#719130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#719140000000
0!
0'
0/
#719150000000
1!
1'
1/
#719160000000
0!
0'
0/
#719170000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#719180000000
0!
0'
0/
#719190000000
1!
1'
1/
#719200000000
0!
0'
0/
#719210000000
1!
1'
1/
#719220000000
0!
0'
0/
#719230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#719240000000
0!
0'
0/
#719250000000
1!
1'
1/
#719260000000
0!
0'
0/
#719270000000
1!
1'
1/
#719280000000
0!
0'
0/
#719290000000
1!
1'
1/
#719300000000
0!
0'
0/
#719310000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#719320000000
0!
0'
0/
#719330000000
1!
1'
1/
#719340000000
0!
0'
0/
#719350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#719360000000
0!
0'
0/
#719370000000
1!
1'
1/
#719380000000
0!
0'
0/
#719390000000
#719400000000
1!
1'
1/
#719410000000
0!
0'
0/
#719420000000
1!
1'
1/
#719430000000
0!
1"
0'
1(
0/
10
#719440000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#719450000000
0!
0'
0/
#719460000000
1!
1'
1/
#719470000000
0!
0'
0/
#719480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#719490000000
0!
0'
0/
#719500000000
1!
1'
1/
#719510000000
0!
1"
0'
1(
0/
10
#719520000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#719530000000
0!
1$
0'
1+
0/
#719540000000
1!
1'
1/
#719550000000
0!
0'
0/
#719560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#719570000000
0!
0'
0/
#719580000000
1!
1'
1/
#719590000000
0!
0'
0/
#719600000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#719610000000
0!
0'
0/
#719620000000
1!
1'
1/
#719630000000
0!
0'
0/
#719640000000
1!
1'
1/
#719650000000
0!
0'
0/
#719660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#719670000000
0!
0'
0/
#719680000000
1!
1'
1/
#719690000000
0!
0'
0/
#719700000000
1!
1'
1/
#719710000000
0!
0'
0/
#719720000000
1!
1'
1/
#719730000000
0!
0'
0/
#719740000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#719750000000
0!
0'
0/
#719760000000
1!
1'
1/
#719770000000
0!
0'
0/
#719780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#719790000000
0!
0'
0/
#719800000000
1!
1'
1/
#719810000000
0!
0'
0/
#719820000000
#719830000000
1!
1'
1/
#719840000000
0!
0'
0/
#719850000000
1!
1'
1/
#719860000000
0!
1"
0'
1(
0/
10
#719870000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#719880000000
0!
0'
0/
#719890000000
1!
1'
1/
#719900000000
0!
0'
0/
#719910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#719920000000
0!
0'
0/
#719930000000
1!
1'
1/
#719940000000
0!
1"
0'
1(
0/
10
#719950000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#719960000000
0!
1$
0'
1+
0/
#719970000000
1!
1'
1/
#719980000000
0!
0'
0/
#719990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#720000000000
0!
0'
0/
#720010000000
1!
1'
1/
#720020000000
0!
0'
0/
#720030000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#720040000000
0!
0'
0/
#720050000000
1!
1'
1/
#720060000000
0!
0'
0/
#720070000000
1!
1'
1/
#720080000000
0!
0'
0/
#720090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#720100000000
0!
0'
0/
#720110000000
1!
1'
1/
#720120000000
0!
0'
0/
#720130000000
1!
1'
1/
#720140000000
0!
0'
0/
#720150000000
1!
1'
1/
#720160000000
0!
0'
0/
#720170000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#720180000000
0!
0'
0/
#720190000000
1!
1'
1/
#720200000000
0!
0'
0/
#720210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#720220000000
0!
0'
0/
#720230000000
1!
1'
1/
#720240000000
0!
0'
0/
#720250000000
#720260000000
1!
1'
1/
#720270000000
0!
0'
0/
#720280000000
1!
1'
1/
#720290000000
0!
1"
0'
1(
0/
10
#720300000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#720310000000
0!
0'
0/
#720320000000
1!
1'
1/
#720330000000
0!
0'
0/
#720340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#720350000000
0!
0'
0/
#720360000000
1!
1'
1/
#720370000000
0!
1"
0'
1(
0/
10
#720380000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#720390000000
0!
1$
0'
1+
0/
#720400000000
1!
1'
1/
#720410000000
0!
0'
0/
#720420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#720430000000
0!
0'
0/
#720440000000
1!
1'
1/
#720450000000
0!
0'
0/
#720460000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#720470000000
0!
0'
0/
#720480000000
1!
1'
1/
#720490000000
0!
0'
0/
#720500000000
1!
1'
1/
#720510000000
0!
0'
0/
#720520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#720530000000
0!
0'
0/
#720540000000
1!
1'
1/
#720550000000
0!
0'
0/
#720560000000
1!
1'
1/
#720570000000
0!
0'
0/
#720580000000
1!
1'
1/
#720590000000
0!
0'
0/
#720600000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#720610000000
0!
0'
0/
#720620000000
1!
1'
1/
#720630000000
0!
0'
0/
#720640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#720650000000
0!
0'
0/
#720660000000
1!
1'
1/
#720670000000
0!
0'
0/
#720680000000
#720690000000
1!
1'
1/
#720700000000
0!
0'
0/
#720710000000
1!
1'
1/
#720720000000
0!
1"
0'
1(
0/
10
#720730000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#720740000000
0!
0'
0/
#720750000000
1!
1'
1/
#720760000000
0!
0'
0/
#720770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#720780000000
0!
0'
0/
#720790000000
1!
1'
1/
#720800000000
0!
1"
0'
1(
0/
10
#720810000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#720820000000
0!
1$
0'
1+
0/
#720830000000
1!
1'
1/
#720840000000
0!
0'
0/
#720850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#720860000000
0!
0'
0/
#720870000000
1!
1'
1/
#720880000000
0!
0'
0/
#720890000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#720900000000
0!
0'
0/
#720910000000
1!
1'
1/
#720920000000
0!
0'
0/
#720930000000
1!
1'
1/
#720940000000
0!
0'
0/
#720950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#720960000000
0!
0'
0/
#720970000000
1!
1'
1/
#720980000000
0!
0'
0/
#720990000000
1!
1'
1/
#721000000000
0!
0'
0/
#721010000000
1!
1'
1/
#721020000000
0!
0'
0/
#721030000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#721040000000
0!
0'
0/
#721050000000
1!
1'
1/
#721060000000
0!
0'
0/
#721070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#721080000000
0!
0'
0/
#721090000000
1!
1'
1/
#721100000000
0!
0'
0/
#721110000000
#721120000000
1!
1'
1/
#721130000000
0!
0'
0/
#721140000000
1!
1'
1/
#721150000000
0!
1"
0'
1(
0/
10
#721160000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#721170000000
0!
0'
0/
#721180000000
1!
1'
1/
#721190000000
0!
0'
0/
#721200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#721210000000
0!
0'
0/
#721220000000
1!
1'
1/
#721230000000
0!
1"
0'
1(
0/
10
#721240000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#721250000000
0!
1$
0'
1+
0/
#721260000000
1!
1'
1/
#721270000000
0!
0'
0/
#721280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#721290000000
0!
0'
0/
#721300000000
1!
1'
1/
#721310000000
0!
0'
0/
#721320000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#721330000000
0!
0'
0/
#721340000000
1!
1'
1/
#721350000000
0!
0'
0/
#721360000000
1!
1'
1/
#721370000000
0!
0'
0/
#721380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#721390000000
0!
0'
0/
#721400000000
1!
1'
1/
#721410000000
0!
0'
0/
#721420000000
1!
1'
1/
#721430000000
0!
0'
0/
#721440000000
1!
1'
1/
#721450000000
0!
0'
0/
#721460000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#721470000000
0!
0'
0/
#721480000000
1!
1'
1/
#721490000000
0!
0'
0/
#721500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#721510000000
0!
0'
0/
#721520000000
1!
1'
1/
#721530000000
0!
0'
0/
#721540000000
#721550000000
1!
1'
1/
#721560000000
0!
0'
0/
#721570000000
1!
1'
1/
#721580000000
0!
1"
0'
1(
0/
10
#721590000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#721600000000
0!
0'
0/
#721610000000
1!
1'
1/
#721620000000
0!
0'
0/
#721630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#721640000000
0!
0'
0/
#721650000000
1!
1'
1/
#721660000000
0!
1"
0'
1(
0/
10
#721670000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#721680000000
0!
1$
0'
1+
0/
#721690000000
1!
1'
1/
#721700000000
0!
0'
0/
#721710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#721720000000
0!
0'
0/
#721730000000
1!
1'
1/
#721740000000
0!
0'
0/
#721750000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#721760000000
0!
0'
0/
#721770000000
1!
1'
1/
#721780000000
0!
0'
0/
#721790000000
1!
1'
1/
#721800000000
0!
0'
0/
#721810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#721820000000
0!
0'
0/
#721830000000
1!
1'
1/
#721840000000
0!
0'
0/
#721850000000
1!
1'
1/
#721860000000
0!
0'
0/
#721870000000
1!
1'
1/
#721880000000
0!
0'
0/
#721890000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#721900000000
0!
0'
0/
#721910000000
1!
1'
1/
#721920000000
0!
0'
0/
#721930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#721940000000
0!
0'
0/
#721950000000
1!
1'
1/
#721960000000
0!
0'
0/
#721970000000
#721980000000
1!
1'
1/
#721990000000
0!
0'
0/
#722000000000
1!
1'
1/
#722010000000
0!
1"
0'
1(
0/
10
#722020000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#722030000000
0!
0'
0/
#722040000000
1!
1'
1/
#722050000000
0!
0'
0/
#722060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#722070000000
0!
0'
0/
#722080000000
1!
1'
1/
#722090000000
0!
1"
0'
1(
0/
10
#722100000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#722110000000
0!
1$
0'
1+
0/
#722120000000
1!
1'
1/
#722130000000
0!
0'
0/
#722140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#722150000000
0!
0'
0/
#722160000000
1!
1'
1/
#722170000000
0!
0'
0/
#722180000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#722190000000
0!
0'
0/
#722200000000
1!
1'
1/
#722210000000
0!
0'
0/
#722220000000
1!
1'
1/
#722230000000
0!
0'
0/
#722240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#722250000000
0!
0'
0/
#722260000000
1!
1'
1/
#722270000000
0!
0'
0/
#722280000000
1!
1'
1/
#722290000000
0!
0'
0/
#722300000000
1!
1'
1/
#722310000000
0!
0'
0/
#722320000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#722330000000
0!
0'
0/
#722340000000
1!
1'
1/
#722350000000
0!
0'
0/
#722360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#722370000000
0!
0'
0/
#722380000000
1!
1'
1/
#722390000000
0!
0'
0/
#722400000000
#722410000000
1!
1'
1/
#722420000000
0!
0'
0/
#722430000000
1!
1'
1/
#722440000000
0!
1"
0'
1(
0/
10
#722450000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#722460000000
0!
0'
0/
#722470000000
1!
1'
1/
#722480000000
0!
0'
0/
#722490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#722500000000
0!
0'
0/
#722510000000
1!
1'
1/
#722520000000
0!
1"
0'
1(
0/
10
#722530000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#722540000000
0!
1$
0'
1+
0/
#722550000000
1!
1'
1/
#722560000000
0!
0'
0/
#722570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#722580000000
0!
0'
0/
#722590000000
1!
1'
1/
#722600000000
0!
0'
0/
#722610000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#722620000000
0!
0'
0/
#722630000000
1!
1'
1/
#722640000000
0!
0'
0/
#722650000000
1!
1'
1/
#722660000000
0!
0'
0/
#722670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#722680000000
0!
0'
0/
#722690000000
1!
1'
1/
#722700000000
0!
0'
0/
#722710000000
1!
1'
1/
#722720000000
0!
0'
0/
#722730000000
1!
1'
1/
#722740000000
0!
0'
0/
#722750000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#722760000000
0!
0'
0/
#722770000000
1!
1'
1/
#722780000000
0!
0'
0/
#722790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#722800000000
0!
0'
0/
#722810000000
1!
1'
1/
#722820000000
0!
0'
0/
#722830000000
#722840000000
1!
1'
1/
#722850000000
0!
0'
0/
#722860000000
1!
1'
1/
#722870000000
0!
1"
0'
1(
0/
10
#722880000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#722890000000
0!
0'
0/
#722900000000
1!
1'
1/
#722910000000
0!
0'
0/
#722920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#722930000000
0!
0'
0/
#722940000000
1!
1'
1/
#722950000000
0!
1"
0'
1(
0/
10
#722960000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#722970000000
0!
1$
0'
1+
0/
#722980000000
1!
1'
1/
#722990000000
0!
0'
0/
#723000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#723010000000
0!
0'
0/
#723020000000
1!
1'
1/
#723030000000
0!
0'
0/
#723040000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#723050000000
0!
0'
0/
#723060000000
1!
1'
1/
#723070000000
0!
0'
0/
#723080000000
1!
1'
1/
#723090000000
0!
0'
0/
#723100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#723110000000
0!
0'
0/
#723120000000
1!
1'
1/
#723130000000
0!
0'
0/
#723140000000
1!
1'
1/
#723150000000
0!
0'
0/
#723160000000
1!
1'
1/
#723170000000
0!
0'
0/
#723180000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#723190000000
0!
0'
0/
#723200000000
1!
1'
1/
#723210000000
0!
0'
0/
#723220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#723230000000
0!
0'
0/
#723240000000
1!
1'
1/
#723250000000
0!
0'
0/
#723260000000
#723270000000
1!
1'
1/
#723280000000
0!
0'
0/
#723290000000
1!
1'
1/
#723300000000
0!
1"
0'
1(
0/
10
#723310000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#723320000000
0!
0'
0/
#723330000000
1!
1'
1/
#723340000000
0!
0'
0/
#723350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#723360000000
0!
0'
0/
#723370000000
1!
1'
1/
#723380000000
0!
1"
0'
1(
0/
10
#723390000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#723400000000
0!
1$
0'
1+
0/
#723410000000
1!
1'
1/
#723420000000
0!
0'
0/
#723430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#723440000000
0!
0'
0/
#723450000000
1!
1'
1/
#723460000000
0!
0'
0/
#723470000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#723480000000
0!
0'
0/
#723490000000
1!
1'
1/
#723500000000
0!
0'
0/
#723510000000
1!
1'
1/
#723520000000
0!
0'
0/
#723530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#723540000000
0!
0'
0/
#723550000000
1!
1'
1/
#723560000000
0!
0'
0/
#723570000000
1!
1'
1/
#723580000000
0!
0'
0/
#723590000000
1!
1'
1/
#723600000000
0!
0'
0/
#723610000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#723620000000
0!
0'
0/
#723630000000
1!
1'
1/
#723640000000
0!
0'
0/
#723650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#723660000000
0!
0'
0/
#723670000000
1!
1'
1/
#723680000000
0!
0'
0/
#723690000000
#723700000000
1!
1'
1/
#723710000000
0!
0'
0/
#723720000000
1!
1'
1/
#723730000000
0!
1"
0'
1(
0/
10
#723740000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#723750000000
0!
0'
0/
#723760000000
1!
1'
1/
#723770000000
0!
0'
0/
#723780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#723790000000
0!
0'
0/
#723800000000
1!
1'
1/
#723810000000
0!
1"
0'
1(
0/
10
#723820000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#723830000000
0!
1$
0'
1+
0/
#723840000000
1!
1'
1/
#723850000000
0!
0'
0/
#723860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#723870000000
0!
0'
0/
#723880000000
1!
1'
1/
#723890000000
0!
0'
0/
#723900000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#723910000000
0!
0'
0/
#723920000000
1!
1'
1/
#723930000000
0!
0'
0/
#723940000000
1!
1'
1/
#723950000000
0!
0'
0/
#723960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#723970000000
0!
0'
0/
#723980000000
1!
1'
1/
#723990000000
0!
0'
0/
#724000000000
1!
1'
1/
#724010000000
0!
0'
0/
#724020000000
1!
1'
1/
#724030000000
0!
0'
0/
#724040000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#724050000000
0!
0'
0/
#724060000000
1!
1'
1/
#724070000000
0!
0'
0/
#724080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#724090000000
0!
0'
0/
#724100000000
1!
1'
1/
#724110000000
0!
0'
0/
#724120000000
#724130000000
1!
1'
1/
#724140000000
0!
0'
0/
#724150000000
1!
1'
1/
#724160000000
0!
1"
0'
1(
0/
10
#724170000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#724180000000
0!
0'
0/
#724190000000
1!
1'
1/
#724200000000
0!
0'
0/
#724210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#724220000000
0!
0'
0/
#724230000000
1!
1'
1/
#724240000000
0!
1"
0'
1(
0/
10
#724250000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#724260000000
0!
1$
0'
1+
0/
#724270000000
1!
1'
1/
#724280000000
0!
0'
0/
#724290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#724300000000
0!
0'
0/
#724310000000
1!
1'
1/
#724320000000
0!
0'
0/
#724330000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#724340000000
0!
0'
0/
#724350000000
1!
1'
1/
#724360000000
0!
0'
0/
#724370000000
1!
1'
1/
#724380000000
0!
0'
0/
#724390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#724400000000
0!
0'
0/
#724410000000
1!
1'
1/
#724420000000
0!
0'
0/
#724430000000
1!
1'
1/
#724440000000
0!
0'
0/
#724450000000
1!
1'
1/
#724460000000
0!
0'
0/
#724470000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#724480000000
0!
0'
0/
#724490000000
1!
1'
1/
#724500000000
0!
0'
0/
#724510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#724520000000
0!
0'
0/
#724530000000
1!
1'
1/
#724540000000
0!
0'
0/
#724550000000
#724560000000
1!
1'
1/
#724570000000
0!
0'
0/
#724580000000
1!
1'
1/
#724590000000
0!
1"
0'
1(
0/
10
#724600000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#724610000000
0!
0'
0/
#724620000000
1!
1'
1/
#724630000000
0!
0'
0/
#724640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#724650000000
0!
0'
0/
#724660000000
1!
1'
1/
#724670000000
0!
1"
0'
1(
0/
10
#724680000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#724690000000
0!
1$
0'
1+
0/
#724700000000
1!
1'
1/
#724710000000
0!
0'
0/
#724720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#724730000000
0!
0'
0/
#724740000000
1!
1'
1/
#724750000000
0!
0'
0/
#724760000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#724770000000
0!
0'
0/
#724780000000
1!
1'
1/
#724790000000
0!
0'
0/
#724800000000
1!
1'
1/
#724810000000
0!
0'
0/
#724820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#724830000000
0!
0'
0/
#724840000000
1!
1'
1/
#724850000000
0!
0'
0/
#724860000000
1!
1'
1/
#724870000000
0!
0'
0/
#724880000000
1!
1'
1/
#724890000000
0!
0'
0/
#724900000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#724910000000
0!
0'
0/
#724920000000
1!
1'
1/
#724930000000
0!
0'
0/
#724940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#724950000000
0!
0'
0/
#724960000000
1!
1'
1/
#724970000000
0!
0'
0/
#724980000000
#724990000000
1!
1'
1/
#725000000000
0!
0'
0/
#725010000000
1!
1'
1/
#725020000000
0!
1"
0'
1(
0/
10
#725030000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#725040000000
0!
0'
0/
#725050000000
1!
1'
1/
#725060000000
0!
0'
0/
#725070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#725080000000
0!
0'
0/
#725090000000
1!
1'
1/
#725100000000
0!
1"
0'
1(
0/
10
#725110000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#725120000000
0!
1$
0'
1+
0/
#725130000000
1!
1'
1/
#725140000000
0!
0'
0/
#725150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#725160000000
0!
0'
0/
#725170000000
1!
1'
1/
#725180000000
0!
0'
0/
#725190000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#725200000000
0!
0'
0/
#725210000000
1!
1'
1/
#725220000000
0!
0'
0/
#725230000000
1!
1'
1/
#725240000000
0!
0'
0/
#725250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#725260000000
0!
0'
0/
#725270000000
1!
1'
1/
#725280000000
0!
0'
0/
#725290000000
1!
1'
1/
#725300000000
0!
0'
0/
#725310000000
1!
1'
1/
#725320000000
0!
0'
0/
#725330000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#725340000000
0!
0'
0/
#725350000000
1!
1'
1/
#725360000000
0!
0'
0/
#725370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#725380000000
0!
0'
0/
#725390000000
1!
1'
1/
#725400000000
0!
0'
0/
#725410000000
#725420000000
1!
1'
1/
#725430000000
0!
0'
0/
#725440000000
1!
1'
1/
#725450000000
0!
1"
0'
1(
0/
10
#725460000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#725470000000
0!
0'
0/
#725480000000
1!
1'
1/
#725490000000
0!
0'
0/
#725500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#725510000000
0!
0'
0/
#725520000000
1!
1'
1/
#725530000000
0!
1"
0'
1(
0/
10
#725540000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#725550000000
0!
1$
0'
1+
0/
#725560000000
1!
1'
1/
#725570000000
0!
0'
0/
#725580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#725590000000
0!
0'
0/
#725600000000
1!
1'
1/
#725610000000
0!
0'
0/
#725620000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#725630000000
0!
0'
0/
#725640000000
1!
1'
1/
#725650000000
0!
0'
0/
#725660000000
1!
1'
1/
#725670000000
0!
0'
0/
#725680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#725690000000
0!
0'
0/
#725700000000
1!
1'
1/
#725710000000
0!
0'
0/
#725720000000
1!
1'
1/
#725730000000
0!
0'
0/
#725740000000
1!
1'
1/
#725750000000
0!
0'
0/
#725760000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#725770000000
0!
0'
0/
#725780000000
1!
1'
1/
#725790000000
0!
0'
0/
#725800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#725810000000
0!
0'
0/
#725820000000
1!
1'
1/
#725830000000
0!
0'
0/
#725840000000
#725850000000
1!
1'
1/
#725860000000
0!
0'
0/
#725870000000
1!
1'
1/
#725880000000
0!
1"
0'
1(
0/
10
#725890000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#725900000000
0!
0'
0/
#725910000000
1!
1'
1/
#725920000000
0!
0'
0/
#725930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#725940000000
0!
0'
0/
#725950000000
1!
1'
1/
#725960000000
0!
1"
0'
1(
0/
10
#725970000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#725980000000
0!
1$
0'
1+
0/
#725990000000
1!
1'
1/
#726000000000
0!
0'
0/
#726010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#726020000000
0!
0'
0/
#726030000000
1!
1'
1/
#726040000000
0!
0'
0/
#726050000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#726060000000
0!
0'
0/
#726070000000
1!
1'
1/
#726080000000
0!
0'
0/
#726090000000
1!
1'
1/
#726100000000
0!
0'
0/
#726110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#726120000000
0!
0'
0/
#726130000000
1!
1'
1/
#726140000000
0!
0'
0/
#726150000000
1!
1'
1/
#726160000000
0!
0'
0/
#726170000000
1!
1'
1/
#726180000000
0!
0'
0/
#726190000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#726200000000
0!
0'
0/
#726210000000
1!
1'
1/
#726220000000
0!
0'
0/
#726230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#726240000000
0!
0'
0/
#726250000000
1!
1'
1/
#726260000000
0!
0'
0/
#726270000000
#726280000000
1!
1'
1/
#726290000000
0!
0'
0/
#726300000000
1!
1'
1/
#726310000000
0!
1"
0'
1(
0/
10
#726320000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#726330000000
0!
0'
0/
#726340000000
1!
1'
1/
#726350000000
0!
0'
0/
#726360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#726370000000
0!
0'
0/
#726380000000
1!
1'
1/
#726390000000
0!
1"
0'
1(
0/
10
#726400000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#726410000000
0!
1$
0'
1+
0/
#726420000000
1!
1'
1/
#726430000000
0!
0'
0/
#726440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#726450000000
0!
0'
0/
#726460000000
1!
1'
1/
#726470000000
0!
0'
0/
#726480000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#726490000000
0!
0'
0/
#726500000000
1!
1'
1/
#726510000000
0!
0'
0/
#726520000000
1!
1'
1/
#726530000000
0!
0'
0/
#726540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#726550000000
0!
0'
0/
#726560000000
1!
1'
1/
#726570000000
0!
0'
0/
#726580000000
1!
1'
1/
#726590000000
0!
0'
0/
#726600000000
1!
1'
1/
#726610000000
0!
0'
0/
#726620000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#726630000000
0!
0'
0/
#726640000000
1!
1'
1/
#726650000000
0!
0'
0/
#726660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#726670000000
0!
0'
0/
#726680000000
1!
1'
1/
#726690000000
0!
0'
0/
#726700000000
#726710000000
1!
1'
1/
#726720000000
0!
0'
0/
#726730000000
1!
1'
1/
#726740000000
0!
1"
0'
1(
0/
10
#726750000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#726760000000
0!
0'
0/
#726770000000
1!
1'
1/
#726780000000
0!
0'
0/
#726790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#726800000000
0!
0'
0/
#726810000000
1!
1'
1/
#726820000000
0!
1"
0'
1(
0/
10
#726830000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#726840000000
0!
1$
0'
1+
0/
#726850000000
1!
1'
1/
#726860000000
0!
0'
0/
#726870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#726880000000
0!
0'
0/
#726890000000
1!
1'
1/
#726900000000
0!
0'
0/
#726910000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#726920000000
0!
0'
0/
#726930000000
1!
1'
1/
#726940000000
0!
0'
0/
#726950000000
1!
1'
1/
#726960000000
0!
0'
0/
#726970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#726980000000
0!
0'
0/
#726990000000
1!
1'
1/
#727000000000
0!
0'
0/
#727010000000
1!
1'
1/
#727020000000
0!
0'
0/
#727030000000
1!
1'
1/
#727040000000
0!
0'
0/
#727050000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#727060000000
0!
0'
0/
#727070000000
1!
1'
1/
#727080000000
0!
0'
0/
#727090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#727100000000
0!
0'
0/
#727110000000
1!
1'
1/
#727120000000
0!
0'
0/
#727130000000
#727140000000
1!
1'
1/
#727150000000
0!
0'
0/
#727160000000
1!
1'
1/
#727170000000
0!
1"
0'
1(
0/
10
#727180000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#727190000000
0!
0'
0/
#727200000000
1!
1'
1/
#727210000000
0!
0'
0/
#727220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#727230000000
0!
0'
0/
#727240000000
1!
1'
1/
#727250000000
0!
1"
0'
1(
0/
10
#727260000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#727270000000
0!
1$
0'
1+
0/
#727280000000
1!
1'
1/
#727290000000
0!
0'
0/
#727300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#727310000000
0!
0'
0/
#727320000000
1!
1'
1/
#727330000000
0!
0'
0/
#727340000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#727350000000
0!
0'
0/
#727360000000
1!
1'
1/
#727370000000
0!
0'
0/
#727380000000
1!
1'
1/
#727390000000
0!
0'
0/
#727400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#727410000000
0!
0'
0/
#727420000000
1!
1'
1/
#727430000000
0!
0'
0/
#727440000000
1!
1'
1/
#727450000000
0!
0'
0/
#727460000000
1!
1'
1/
#727470000000
0!
0'
0/
#727480000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#727490000000
0!
0'
0/
#727500000000
1!
1'
1/
#727510000000
0!
0'
0/
#727520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#727530000000
0!
0'
0/
#727540000000
1!
1'
1/
#727550000000
0!
0'
0/
#727560000000
#727570000000
1!
1'
1/
#727580000000
0!
0'
0/
#727590000000
1!
1'
1/
#727600000000
0!
1"
0'
1(
0/
10
#727610000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#727620000000
0!
0'
0/
#727630000000
1!
1'
1/
#727640000000
0!
0'
0/
#727650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#727660000000
0!
0'
0/
#727670000000
1!
1'
1/
#727680000000
0!
1"
0'
1(
0/
10
#727690000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#727700000000
0!
1$
0'
1+
0/
#727710000000
1!
1'
1/
#727720000000
0!
0'
0/
#727730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#727740000000
0!
0'
0/
#727750000000
1!
1'
1/
#727760000000
0!
0'
0/
#727770000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#727780000000
0!
0'
0/
#727790000000
1!
1'
1/
#727800000000
0!
0'
0/
#727810000000
1!
1'
1/
#727820000000
0!
0'
0/
#727830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#727840000000
0!
0'
0/
#727850000000
1!
1'
1/
#727860000000
0!
0'
0/
#727870000000
1!
1'
1/
#727880000000
0!
0'
0/
#727890000000
1!
1'
1/
#727900000000
0!
0'
0/
#727910000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#727920000000
0!
0'
0/
#727930000000
1!
1'
1/
#727940000000
0!
0'
0/
#727950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#727960000000
0!
0'
0/
#727970000000
1!
1'
1/
#727980000000
0!
0'
0/
#727990000000
#728000000000
1!
1'
1/
#728010000000
0!
0'
0/
#728020000000
1!
1'
1/
#728030000000
0!
1"
0'
1(
0/
10
#728040000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#728050000000
0!
0'
0/
#728060000000
1!
1'
1/
#728070000000
0!
0'
0/
#728080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#728090000000
0!
0'
0/
#728100000000
1!
1'
1/
#728110000000
0!
1"
0'
1(
0/
10
#728120000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#728130000000
0!
1$
0'
1+
0/
#728140000000
1!
1'
1/
#728150000000
0!
0'
0/
#728160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#728170000000
0!
0'
0/
#728180000000
1!
1'
1/
#728190000000
0!
0'
0/
#728200000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#728210000000
0!
0'
0/
#728220000000
1!
1'
1/
#728230000000
0!
0'
0/
#728240000000
1!
1'
1/
#728250000000
0!
0'
0/
#728260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#728270000000
0!
0'
0/
#728280000000
1!
1'
1/
#728290000000
0!
0'
0/
#728300000000
1!
1'
1/
#728310000000
0!
0'
0/
#728320000000
1!
1'
1/
#728330000000
0!
0'
0/
#728340000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#728350000000
0!
0'
0/
#728360000000
1!
1'
1/
#728370000000
0!
0'
0/
#728380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#728390000000
0!
0'
0/
#728400000000
1!
1'
1/
#728410000000
0!
0'
0/
#728420000000
#728430000000
1!
1'
1/
#728440000000
0!
0'
0/
#728450000000
1!
1'
1/
#728460000000
0!
1"
0'
1(
0/
10
#728470000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#728480000000
0!
0'
0/
#728490000000
1!
1'
1/
#728500000000
0!
0'
0/
#728510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#728520000000
0!
0'
0/
#728530000000
1!
1'
1/
#728540000000
0!
1"
0'
1(
0/
10
#728550000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#728560000000
0!
1$
0'
1+
0/
#728570000000
1!
1'
1/
#728580000000
0!
0'
0/
#728590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#728600000000
0!
0'
0/
#728610000000
1!
1'
1/
#728620000000
0!
0'
0/
#728630000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#728640000000
0!
0'
0/
#728650000000
1!
1'
1/
#728660000000
0!
0'
0/
#728670000000
1!
1'
1/
#728680000000
0!
0'
0/
#728690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#728700000000
0!
0'
0/
#728710000000
1!
1'
1/
#728720000000
0!
0'
0/
#728730000000
1!
1'
1/
#728740000000
0!
0'
0/
#728750000000
1!
1'
1/
#728760000000
0!
0'
0/
#728770000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#728780000000
0!
0'
0/
#728790000000
1!
1'
1/
#728800000000
0!
0'
0/
#728810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#728820000000
0!
0'
0/
#728830000000
1!
1'
1/
#728840000000
0!
0'
0/
#728850000000
#728860000000
1!
1'
1/
#728870000000
0!
0'
0/
#728880000000
1!
1'
1/
#728890000000
0!
1"
0'
1(
0/
10
#728900000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#728910000000
0!
0'
0/
#728920000000
1!
1'
1/
#728930000000
0!
0'
0/
#728940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#728950000000
0!
0'
0/
#728960000000
1!
1'
1/
#728970000000
0!
1"
0'
1(
0/
10
#728980000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#728990000000
0!
1$
0'
1+
0/
#729000000000
1!
1'
1/
#729010000000
0!
0'
0/
#729020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#729030000000
0!
0'
0/
#729040000000
1!
1'
1/
#729050000000
0!
0'
0/
#729060000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#729070000000
0!
0'
0/
#729080000000
1!
1'
1/
#729090000000
0!
0'
0/
#729100000000
1!
1'
1/
#729110000000
0!
0'
0/
#729120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#729130000000
0!
0'
0/
#729140000000
1!
1'
1/
#729150000000
0!
0'
0/
#729160000000
1!
1'
1/
#729170000000
0!
0'
0/
#729180000000
1!
1'
1/
#729190000000
0!
0'
0/
#729200000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#729210000000
0!
0'
0/
#729220000000
1!
1'
1/
#729230000000
0!
0'
0/
#729240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#729250000000
0!
0'
0/
#729260000000
1!
1'
1/
#729270000000
0!
0'
0/
#729280000000
#729290000000
1!
1'
1/
#729300000000
0!
0'
0/
#729310000000
1!
1'
1/
#729320000000
0!
1"
0'
1(
0/
10
#729330000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#729340000000
0!
0'
0/
#729350000000
1!
1'
1/
#729360000000
0!
0'
0/
#729370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#729380000000
0!
0'
0/
#729390000000
1!
1'
1/
#729400000000
0!
1"
0'
1(
0/
10
#729410000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#729420000000
0!
1$
0'
1+
0/
#729430000000
1!
1'
1/
#729440000000
0!
0'
0/
#729450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#729460000000
0!
0'
0/
#729470000000
1!
1'
1/
#729480000000
0!
0'
0/
#729490000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#729500000000
0!
0'
0/
#729510000000
1!
1'
1/
#729520000000
0!
0'
0/
#729530000000
1!
1'
1/
#729540000000
0!
0'
0/
#729550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#729560000000
0!
0'
0/
#729570000000
1!
1'
1/
#729580000000
0!
0'
0/
#729590000000
1!
1'
1/
#729600000000
0!
0'
0/
#729610000000
1!
1'
1/
#729620000000
0!
0'
0/
#729630000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#729640000000
0!
0'
0/
#729650000000
1!
1'
1/
#729660000000
0!
0'
0/
#729670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#729680000000
0!
0'
0/
#729690000000
1!
1'
1/
#729700000000
0!
0'
0/
#729710000000
#729720000000
1!
1'
1/
#729730000000
0!
0'
0/
#729740000000
1!
1'
1/
#729750000000
0!
1"
0'
1(
0/
10
#729760000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#729770000000
0!
0'
0/
#729780000000
1!
1'
1/
#729790000000
0!
0'
0/
#729800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#729810000000
0!
0'
0/
#729820000000
1!
1'
1/
#729830000000
0!
1"
0'
1(
0/
10
#729840000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#729850000000
0!
1$
0'
1+
0/
#729860000000
1!
1'
1/
#729870000000
0!
0'
0/
#729880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#729890000000
0!
0'
0/
#729900000000
1!
1'
1/
#729910000000
0!
0'
0/
#729920000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#729930000000
0!
0'
0/
#729940000000
1!
1'
1/
#729950000000
0!
0'
0/
#729960000000
1!
1'
1/
#729970000000
0!
0'
0/
#729980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#729990000000
0!
0'
0/
#730000000000
1!
1'
1/
#730010000000
0!
0'
0/
#730020000000
1!
1'
1/
#730030000000
0!
0'
0/
#730040000000
1!
1'
1/
#730050000000
0!
0'
0/
#730060000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#730070000000
0!
0'
0/
#730080000000
1!
1'
1/
#730090000000
0!
0'
0/
#730100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#730110000000
0!
0'
0/
#730120000000
1!
1'
1/
#730130000000
0!
0'
0/
#730140000000
#730150000000
1!
1'
1/
#730160000000
0!
0'
0/
#730170000000
1!
1'
1/
#730180000000
0!
1"
0'
1(
0/
10
#730190000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#730200000000
0!
0'
0/
#730210000000
1!
1'
1/
#730220000000
0!
0'
0/
#730230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#730240000000
0!
0'
0/
#730250000000
1!
1'
1/
#730260000000
0!
1"
0'
1(
0/
10
#730270000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#730280000000
0!
1$
0'
1+
0/
#730290000000
1!
1'
1/
#730300000000
0!
0'
0/
#730310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#730320000000
0!
0'
0/
#730330000000
1!
1'
1/
#730340000000
0!
0'
0/
#730350000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#730360000000
0!
0'
0/
#730370000000
1!
1'
1/
#730380000000
0!
0'
0/
#730390000000
1!
1'
1/
#730400000000
0!
0'
0/
#730410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#730420000000
0!
0'
0/
#730430000000
1!
1'
1/
#730440000000
0!
0'
0/
#730450000000
1!
1'
1/
#730460000000
0!
0'
0/
#730470000000
1!
1'
1/
#730480000000
0!
0'
0/
#730490000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#730500000000
0!
0'
0/
#730510000000
1!
1'
1/
#730520000000
0!
0'
0/
#730530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#730540000000
0!
0'
0/
#730550000000
1!
1'
1/
#730560000000
0!
0'
0/
#730570000000
#730580000000
1!
1'
1/
#730590000000
0!
0'
0/
#730600000000
1!
1'
1/
#730610000000
0!
1"
0'
1(
0/
10
#730620000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#730630000000
0!
0'
0/
#730640000000
1!
1'
1/
#730650000000
0!
0'
0/
#730660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#730670000000
0!
0'
0/
#730680000000
1!
1'
1/
#730690000000
0!
1"
0'
1(
0/
10
#730700000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#730710000000
0!
1$
0'
1+
0/
#730720000000
1!
1'
1/
#730730000000
0!
0'
0/
#730740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#730750000000
0!
0'
0/
#730760000000
1!
1'
1/
#730770000000
0!
0'
0/
#730780000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#730790000000
0!
0'
0/
#730800000000
1!
1'
1/
#730810000000
0!
0'
0/
#730820000000
1!
1'
1/
#730830000000
0!
0'
0/
#730840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#730850000000
0!
0'
0/
#730860000000
1!
1'
1/
#730870000000
0!
0'
0/
#730880000000
1!
1'
1/
#730890000000
0!
0'
0/
#730900000000
1!
1'
1/
#730910000000
0!
0'
0/
#730920000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#730930000000
0!
0'
0/
#730940000000
1!
1'
1/
#730950000000
0!
0'
0/
#730960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#730970000000
0!
0'
0/
#730980000000
1!
1'
1/
#730990000000
0!
0'
0/
#731000000000
#731010000000
1!
1'
1/
#731020000000
0!
0'
0/
#731030000000
1!
1'
1/
#731040000000
0!
1"
0'
1(
0/
10
#731050000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#731060000000
0!
0'
0/
#731070000000
1!
1'
1/
#731080000000
0!
0'
0/
#731090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#731100000000
0!
0'
0/
#731110000000
1!
1'
1/
#731120000000
0!
1"
0'
1(
0/
10
#731130000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#731140000000
0!
1$
0'
1+
0/
#731150000000
1!
1'
1/
#731160000000
0!
0'
0/
#731170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#731180000000
0!
0'
0/
#731190000000
1!
1'
1/
#731200000000
0!
0'
0/
#731210000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#731220000000
0!
0'
0/
#731230000000
1!
1'
1/
#731240000000
0!
0'
0/
#731250000000
1!
1'
1/
#731260000000
0!
0'
0/
#731270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#731280000000
0!
0'
0/
#731290000000
1!
1'
1/
#731300000000
0!
0'
0/
#731310000000
1!
1'
1/
#731320000000
0!
0'
0/
#731330000000
1!
1'
1/
#731340000000
0!
0'
0/
#731350000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#731360000000
0!
0'
0/
#731370000000
1!
1'
1/
#731380000000
0!
0'
0/
#731390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#731400000000
0!
0'
0/
#731410000000
1!
1'
1/
#731420000000
0!
0'
0/
#731430000000
#731440000000
1!
1'
1/
#731450000000
0!
0'
0/
#731460000000
1!
1'
1/
#731470000000
0!
1"
0'
1(
0/
10
#731480000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#731490000000
0!
0'
0/
#731500000000
1!
1'
1/
#731510000000
0!
0'
0/
#731520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#731530000000
0!
0'
0/
#731540000000
1!
1'
1/
#731550000000
0!
1"
0'
1(
0/
10
#731560000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#731570000000
0!
1$
0'
1+
0/
#731580000000
1!
1'
1/
#731590000000
0!
0'
0/
#731600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#731610000000
0!
0'
0/
#731620000000
1!
1'
1/
#731630000000
0!
0'
0/
#731640000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#731650000000
0!
0'
0/
#731660000000
1!
1'
1/
#731670000000
0!
0'
0/
#731680000000
1!
1'
1/
#731690000000
0!
0'
0/
#731700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#731710000000
0!
0'
0/
#731720000000
1!
1'
1/
#731730000000
0!
0'
0/
#731740000000
1!
1'
1/
#731750000000
0!
0'
0/
#731760000000
1!
1'
1/
#731770000000
0!
0'
0/
#731780000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#731790000000
0!
0'
0/
#731800000000
1!
1'
1/
#731810000000
0!
0'
0/
#731820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#731830000000
0!
0'
0/
#731840000000
1!
1'
1/
#731850000000
0!
0'
0/
#731860000000
#731870000000
1!
1'
1/
#731880000000
0!
0'
0/
#731890000000
1!
1'
1/
#731900000000
0!
1"
0'
1(
0/
10
#731910000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#731920000000
0!
0'
0/
#731930000000
1!
1'
1/
#731940000000
0!
0'
0/
#731950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#731960000000
0!
0'
0/
#731970000000
1!
1'
1/
#731980000000
0!
1"
0'
1(
0/
10
#731990000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#732000000000
0!
1$
0'
1+
0/
#732010000000
1!
1'
1/
#732020000000
0!
0'
0/
#732030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#732040000000
0!
0'
0/
#732050000000
1!
1'
1/
#732060000000
0!
0'
0/
#732070000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#732080000000
0!
0'
0/
#732090000000
1!
1'
1/
#732100000000
0!
0'
0/
#732110000000
1!
1'
1/
#732120000000
0!
0'
0/
#732130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#732140000000
0!
0'
0/
#732150000000
1!
1'
1/
#732160000000
0!
0'
0/
#732170000000
1!
1'
1/
#732180000000
0!
0'
0/
#732190000000
1!
1'
1/
#732200000000
0!
0'
0/
#732210000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#732220000000
0!
0'
0/
#732230000000
1!
1'
1/
#732240000000
0!
0'
0/
#732250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#732260000000
0!
0'
0/
#732270000000
1!
1'
1/
#732280000000
0!
0'
0/
#732290000000
#732300000000
1!
1'
1/
#732310000000
0!
0'
0/
#732320000000
1!
1'
1/
#732330000000
0!
1"
0'
1(
0/
10
#732340000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#732350000000
0!
0'
0/
#732360000000
1!
1'
1/
#732370000000
0!
0'
0/
#732380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#732390000000
0!
0'
0/
#732400000000
1!
1'
1/
#732410000000
0!
1"
0'
1(
0/
10
#732420000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#732430000000
0!
1$
0'
1+
0/
#732440000000
1!
1'
1/
#732450000000
0!
0'
0/
#732460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#732470000000
0!
0'
0/
#732480000000
1!
1'
1/
#732490000000
0!
0'
0/
#732500000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#732510000000
0!
0'
0/
#732520000000
1!
1'
1/
#732530000000
0!
0'
0/
#732540000000
1!
1'
1/
#732550000000
0!
0'
0/
#732560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#732570000000
0!
0'
0/
#732580000000
1!
1'
1/
#732590000000
0!
0'
0/
#732600000000
1!
1'
1/
#732610000000
0!
0'
0/
#732620000000
1!
1'
1/
#732630000000
0!
0'
0/
#732640000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#732650000000
0!
0'
0/
#732660000000
1!
1'
1/
#732670000000
0!
0'
0/
#732680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#732690000000
0!
0'
0/
#732700000000
1!
1'
1/
#732710000000
0!
0'
0/
#732720000000
#732730000000
1!
1'
1/
#732740000000
0!
0'
0/
#732750000000
1!
1'
1/
#732760000000
0!
1"
0'
1(
0/
10
#732770000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#732780000000
0!
0'
0/
#732790000000
1!
1'
1/
#732800000000
0!
0'
0/
#732810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#732820000000
0!
0'
0/
#732830000000
1!
1'
1/
#732840000000
0!
1"
0'
1(
0/
10
#732850000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#732860000000
0!
1$
0'
1+
0/
#732870000000
1!
1'
1/
#732880000000
0!
0'
0/
#732890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#732900000000
0!
0'
0/
#732910000000
1!
1'
1/
#732920000000
0!
0'
0/
#732930000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#732940000000
0!
0'
0/
#732950000000
1!
1'
1/
#732960000000
0!
0'
0/
#732970000000
1!
1'
1/
#732980000000
0!
0'
0/
#732990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#733000000000
0!
0'
0/
#733010000000
1!
1'
1/
#733020000000
0!
0'
0/
#733030000000
1!
1'
1/
#733040000000
0!
0'
0/
#733050000000
1!
1'
1/
#733060000000
0!
0'
0/
#733070000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#733080000000
0!
0'
0/
#733090000000
1!
1'
1/
#733100000000
0!
0'
0/
#733110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#733120000000
0!
0'
0/
#733130000000
1!
1'
1/
#733140000000
0!
0'
0/
#733150000000
#733160000000
1!
1'
1/
#733170000000
0!
0'
0/
#733180000000
1!
1'
1/
#733190000000
0!
1"
0'
1(
0/
10
#733200000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#733210000000
0!
0'
0/
#733220000000
1!
1'
1/
#733230000000
0!
0'
0/
#733240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#733250000000
0!
0'
0/
#733260000000
1!
1'
1/
#733270000000
0!
1"
0'
1(
0/
10
#733280000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#733290000000
0!
1$
0'
1+
0/
#733300000000
1!
1'
1/
#733310000000
0!
0'
0/
#733320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#733330000000
0!
0'
0/
#733340000000
1!
1'
1/
#733350000000
0!
0'
0/
#733360000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#733370000000
0!
0'
0/
#733380000000
1!
1'
1/
#733390000000
0!
0'
0/
#733400000000
1!
1'
1/
#733410000000
0!
0'
0/
#733420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#733430000000
0!
0'
0/
#733440000000
1!
1'
1/
#733450000000
0!
0'
0/
#733460000000
1!
1'
1/
#733470000000
0!
0'
0/
#733480000000
1!
1'
1/
#733490000000
0!
0'
0/
#733500000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#733510000000
0!
0'
0/
#733520000000
1!
1'
1/
#733530000000
0!
0'
0/
#733540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#733550000000
0!
0'
0/
#733560000000
1!
1'
1/
#733570000000
0!
0'
0/
#733580000000
#733590000000
1!
1'
1/
#733600000000
0!
0'
0/
#733610000000
1!
1'
1/
#733620000000
0!
1"
0'
1(
0/
10
#733630000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#733640000000
0!
0'
0/
#733650000000
1!
1'
1/
#733660000000
0!
0'
0/
#733670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#733680000000
0!
0'
0/
#733690000000
1!
1'
1/
#733700000000
0!
1"
0'
1(
0/
10
#733710000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#733720000000
0!
1$
0'
1+
0/
#733730000000
1!
1'
1/
#733740000000
0!
0'
0/
#733750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#733760000000
0!
0'
0/
#733770000000
1!
1'
1/
#733780000000
0!
0'
0/
#733790000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#733800000000
0!
0'
0/
#733810000000
1!
1'
1/
#733820000000
0!
0'
0/
#733830000000
1!
1'
1/
#733840000000
0!
0'
0/
#733850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#733860000000
0!
0'
0/
#733870000000
1!
1'
1/
#733880000000
0!
0'
0/
#733890000000
1!
1'
1/
#733900000000
0!
0'
0/
#733910000000
1!
1'
1/
#733920000000
0!
0'
0/
#733930000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#733940000000
0!
0'
0/
#733950000000
1!
1'
1/
#733960000000
0!
0'
0/
#733970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#733980000000
0!
0'
0/
#733990000000
1!
1'
1/
#734000000000
0!
0'
0/
#734010000000
#734020000000
1!
1'
1/
#734030000000
0!
0'
0/
#734040000000
1!
1'
1/
#734050000000
0!
1"
0'
1(
0/
10
#734060000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#734070000000
0!
0'
0/
#734080000000
1!
1'
1/
#734090000000
0!
0'
0/
#734100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#734110000000
0!
0'
0/
#734120000000
1!
1'
1/
#734130000000
0!
1"
0'
1(
0/
10
#734140000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#734150000000
0!
1$
0'
1+
0/
#734160000000
1!
1'
1/
#734170000000
0!
0'
0/
#734180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#734190000000
0!
0'
0/
#734200000000
1!
1'
1/
#734210000000
0!
0'
0/
#734220000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#734230000000
0!
0'
0/
#734240000000
1!
1'
1/
#734250000000
0!
0'
0/
#734260000000
1!
1'
1/
#734270000000
0!
0'
0/
#734280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#734290000000
0!
0'
0/
#734300000000
1!
1'
1/
#734310000000
0!
0'
0/
#734320000000
1!
1'
1/
#734330000000
0!
0'
0/
#734340000000
1!
1'
1/
#734350000000
0!
0'
0/
#734360000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#734370000000
0!
0'
0/
#734380000000
1!
1'
1/
#734390000000
0!
0'
0/
#734400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#734410000000
0!
0'
0/
#734420000000
1!
1'
1/
#734430000000
0!
0'
0/
#734440000000
#734450000000
1!
1'
1/
#734460000000
0!
0'
0/
#734470000000
1!
1'
1/
#734480000000
0!
1"
0'
1(
0/
10
#734490000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#734500000000
0!
0'
0/
#734510000000
1!
1'
1/
#734520000000
0!
0'
0/
#734530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#734540000000
0!
0'
0/
#734550000000
1!
1'
1/
#734560000000
0!
1"
0'
1(
0/
10
#734570000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#734580000000
0!
1$
0'
1+
0/
#734590000000
1!
1'
1/
#734600000000
0!
0'
0/
#734610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#734620000000
0!
0'
0/
#734630000000
1!
1'
1/
#734640000000
0!
0'
0/
#734650000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#734660000000
0!
0'
0/
#734670000000
1!
1'
1/
#734680000000
0!
0'
0/
#734690000000
1!
1'
1/
#734700000000
0!
0'
0/
#734710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#734720000000
0!
0'
0/
#734730000000
1!
1'
1/
#734740000000
0!
0'
0/
#734750000000
1!
1'
1/
#734760000000
0!
0'
0/
#734770000000
1!
1'
1/
#734780000000
0!
0'
0/
#734790000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#734800000000
0!
0'
0/
#734810000000
1!
1'
1/
#734820000000
0!
0'
0/
#734830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#734840000000
0!
0'
0/
#734850000000
1!
1'
1/
#734860000000
0!
0'
0/
#734870000000
#734880000000
1!
1'
1/
#734890000000
0!
0'
0/
#734900000000
1!
1'
1/
#734910000000
0!
1"
0'
1(
0/
10
#734920000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#734930000000
0!
0'
0/
#734940000000
1!
1'
1/
#734950000000
0!
0'
0/
#734960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#734970000000
0!
0'
0/
#734980000000
1!
1'
1/
#734990000000
0!
1"
0'
1(
0/
10
#735000000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#735010000000
0!
1$
0'
1+
0/
#735020000000
1!
1'
1/
#735030000000
0!
0'
0/
#735040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#735050000000
0!
0'
0/
#735060000000
1!
1'
1/
#735070000000
0!
0'
0/
#735080000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#735090000000
0!
0'
0/
#735100000000
1!
1'
1/
#735110000000
0!
0'
0/
#735120000000
1!
1'
1/
#735130000000
0!
0'
0/
#735140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#735150000000
0!
0'
0/
#735160000000
1!
1'
1/
#735170000000
0!
0'
0/
#735180000000
1!
1'
1/
#735190000000
0!
0'
0/
#735200000000
1!
1'
1/
#735210000000
0!
0'
0/
#735220000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#735230000000
0!
0'
0/
#735240000000
1!
1'
1/
#735250000000
0!
0'
0/
#735260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#735270000000
0!
0'
0/
#735280000000
1!
1'
1/
#735290000000
0!
0'
0/
#735300000000
#735310000000
1!
1'
1/
#735320000000
0!
0'
0/
#735330000000
1!
1'
1/
#735340000000
0!
1"
0'
1(
0/
10
#735350000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#735360000000
0!
0'
0/
#735370000000
1!
1'
1/
#735380000000
0!
0'
0/
#735390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#735400000000
0!
0'
0/
#735410000000
1!
1'
1/
#735420000000
0!
1"
0'
1(
0/
10
#735430000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#735440000000
0!
1$
0'
1+
0/
#735450000000
1!
1'
1/
#735460000000
0!
0'
0/
#735470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#735480000000
0!
0'
0/
#735490000000
1!
1'
1/
#735500000000
0!
0'
0/
#735510000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#735520000000
0!
0'
0/
#735530000000
1!
1'
1/
#735540000000
0!
0'
0/
#735550000000
1!
1'
1/
#735560000000
0!
0'
0/
#735570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#735580000000
0!
0'
0/
#735590000000
1!
1'
1/
#735600000000
0!
0'
0/
#735610000000
1!
1'
1/
#735620000000
0!
0'
0/
#735630000000
1!
1'
1/
#735640000000
0!
0'
0/
#735650000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#735660000000
0!
0'
0/
#735670000000
1!
1'
1/
#735680000000
0!
0'
0/
#735690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#735700000000
0!
0'
0/
#735710000000
1!
1'
1/
#735720000000
0!
0'
0/
#735730000000
#735740000000
1!
1'
1/
#735750000000
0!
0'
0/
#735760000000
1!
1'
1/
#735770000000
0!
1"
0'
1(
0/
10
#735780000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#735790000000
0!
0'
0/
#735800000000
1!
1'
1/
#735810000000
0!
0'
0/
#735820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#735830000000
0!
0'
0/
#735840000000
1!
1'
1/
#735850000000
0!
1"
0'
1(
0/
10
#735860000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#735870000000
0!
1$
0'
1+
0/
#735880000000
1!
1'
1/
#735890000000
0!
0'
0/
#735900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#735910000000
0!
0'
0/
#735920000000
1!
1'
1/
#735930000000
0!
0'
0/
#735940000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#735950000000
0!
0'
0/
#735960000000
1!
1'
1/
#735970000000
0!
0'
0/
#735980000000
1!
1'
1/
#735990000000
0!
0'
0/
#736000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#736010000000
0!
0'
0/
#736020000000
1!
1'
1/
#736030000000
0!
0'
0/
#736040000000
1!
1'
1/
#736050000000
0!
0'
0/
#736060000000
1!
1'
1/
#736070000000
0!
0'
0/
#736080000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#736090000000
0!
0'
0/
#736100000000
1!
1'
1/
#736110000000
0!
0'
0/
#736120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#736130000000
0!
0'
0/
#736140000000
1!
1'
1/
#736150000000
0!
0'
0/
#736160000000
#736170000000
1!
1'
1/
#736180000000
0!
0'
0/
#736190000000
1!
1'
1/
#736200000000
0!
1"
0'
1(
0/
10
#736210000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#736220000000
0!
0'
0/
#736230000000
1!
1'
1/
#736240000000
0!
0'
0/
#736250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#736260000000
0!
0'
0/
#736270000000
1!
1'
1/
#736280000000
0!
1"
0'
1(
0/
10
#736290000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#736300000000
0!
1$
0'
1+
0/
#736310000000
1!
1'
1/
#736320000000
0!
0'
0/
#736330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#736340000000
0!
0'
0/
#736350000000
1!
1'
1/
#736360000000
0!
0'
0/
#736370000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#736380000000
0!
0'
0/
#736390000000
1!
1'
1/
#736400000000
0!
0'
0/
#736410000000
1!
1'
1/
#736420000000
0!
0'
0/
#736430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#736440000000
0!
0'
0/
#736450000000
1!
1'
1/
#736460000000
0!
0'
0/
#736470000000
1!
1'
1/
#736480000000
0!
0'
0/
#736490000000
1!
1'
1/
#736500000000
0!
0'
0/
#736510000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#736520000000
0!
0'
0/
#736530000000
1!
1'
1/
#736540000000
0!
0'
0/
#736550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#736560000000
0!
0'
0/
#736570000000
1!
1'
1/
#736580000000
0!
0'
0/
#736590000000
#736600000000
1!
1'
1/
#736610000000
0!
0'
0/
#736620000000
1!
1'
1/
#736630000000
0!
1"
0'
1(
0/
10
#736640000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#736650000000
0!
0'
0/
#736660000000
1!
1'
1/
#736670000000
0!
0'
0/
#736680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#736690000000
0!
0'
0/
#736700000000
1!
1'
1/
#736710000000
0!
1"
0'
1(
0/
10
#736720000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#736730000000
0!
1$
0'
1+
0/
#736740000000
1!
1'
1/
#736750000000
0!
0'
0/
#736760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#736770000000
0!
0'
0/
#736780000000
1!
1'
1/
#736790000000
0!
0'
0/
#736800000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#736810000000
0!
0'
0/
#736820000000
1!
1'
1/
#736830000000
0!
0'
0/
#736840000000
1!
1'
1/
#736850000000
0!
0'
0/
#736860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#736870000000
0!
0'
0/
#736880000000
1!
1'
1/
#736890000000
0!
0'
0/
#736900000000
1!
1'
1/
#736910000000
0!
0'
0/
#736920000000
1!
1'
1/
#736930000000
0!
0'
0/
#736940000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#736950000000
0!
0'
0/
#736960000000
1!
1'
1/
#736970000000
0!
0'
0/
#736980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#736990000000
0!
0'
0/
#737000000000
1!
1'
1/
#737010000000
0!
0'
0/
#737020000000
#737030000000
1!
1'
1/
#737040000000
0!
0'
0/
#737050000000
1!
1'
1/
#737060000000
0!
1"
0'
1(
0/
10
#737070000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#737080000000
0!
0'
0/
#737090000000
1!
1'
1/
#737100000000
0!
0'
0/
#737110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#737120000000
0!
0'
0/
#737130000000
1!
1'
1/
#737140000000
0!
1"
0'
1(
0/
10
#737150000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#737160000000
0!
1$
0'
1+
0/
#737170000000
1!
1'
1/
#737180000000
0!
0'
0/
#737190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#737200000000
0!
0'
0/
#737210000000
1!
1'
1/
#737220000000
0!
0'
0/
#737230000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#737240000000
0!
0'
0/
#737250000000
1!
1'
1/
#737260000000
0!
0'
0/
#737270000000
1!
1'
1/
#737280000000
0!
0'
0/
#737290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#737300000000
0!
0'
0/
#737310000000
1!
1'
1/
#737320000000
0!
0'
0/
#737330000000
1!
1'
1/
#737340000000
0!
0'
0/
#737350000000
1!
1'
1/
#737360000000
0!
0'
0/
#737370000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#737380000000
0!
0'
0/
#737390000000
1!
1'
1/
#737400000000
0!
0'
0/
#737410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#737420000000
0!
0'
0/
#737430000000
1!
1'
1/
#737440000000
0!
0'
0/
#737450000000
#737460000000
1!
1'
1/
#737470000000
0!
0'
0/
#737480000000
1!
1'
1/
#737490000000
0!
1"
0'
1(
0/
10
#737500000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#737510000000
0!
0'
0/
#737520000000
1!
1'
1/
#737530000000
0!
0'
0/
#737540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#737550000000
0!
0'
0/
#737560000000
1!
1'
1/
#737570000000
0!
1"
0'
1(
0/
10
#737580000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#737590000000
0!
1$
0'
1+
0/
#737600000000
1!
1'
1/
#737610000000
0!
0'
0/
#737620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#737630000000
0!
0'
0/
#737640000000
1!
1'
1/
#737650000000
0!
0'
0/
#737660000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#737670000000
0!
0'
0/
#737680000000
1!
1'
1/
#737690000000
0!
0'
0/
#737700000000
1!
1'
1/
#737710000000
0!
0'
0/
#737720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#737730000000
0!
0'
0/
#737740000000
1!
1'
1/
#737750000000
0!
0'
0/
#737760000000
1!
1'
1/
#737770000000
0!
0'
0/
#737780000000
1!
1'
1/
#737790000000
0!
0'
0/
#737800000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#737810000000
0!
0'
0/
#737820000000
1!
1'
1/
#737830000000
0!
0'
0/
#737840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#737850000000
0!
0'
0/
#737860000000
1!
1'
1/
#737870000000
0!
0'
0/
#737880000000
#737890000000
1!
1'
1/
#737900000000
0!
0'
0/
#737910000000
1!
1'
1/
#737920000000
0!
1"
0'
1(
0/
10
#737930000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#737940000000
0!
0'
0/
#737950000000
1!
1'
1/
#737960000000
0!
0'
0/
#737970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#737980000000
0!
0'
0/
#737990000000
1!
1'
1/
#738000000000
0!
1"
0'
1(
0/
10
#738010000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#738020000000
0!
1$
0'
1+
0/
#738030000000
1!
1'
1/
#738040000000
0!
0'
0/
#738050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#738060000000
0!
0'
0/
#738070000000
1!
1'
1/
#738080000000
0!
0'
0/
#738090000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#738100000000
0!
0'
0/
#738110000000
1!
1'
1/
#738120000000
0!
0'
0/
#738130000000
1!
1'
1/
#738140000000
0!
0'
0/
#738150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#738160000000
0!
0'
0/
#738170000000
1!
1'
1/
#738180000000
0!
0'
0/
#738190000000
1!
1'
1/
#738200000000
0!
0'
0/
#738210000000
1!
1'
1/
#738220000000
0!
0'
0/
#738230000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#738240000000
0!
0'
0/
#738250000000
1!
1'
1/
#738260000000
0!
0'
0/
#738270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#738280000000
0!
0'
0/
#738290000000
1!
1'
1/
#738300000000
0!
0'
0/
#738310000000
#738320000000
1!
1'
1/
#738330000000
0!
0'
0/
#738340000000
1!
1'
1/
#738350000000
0!
1"
0'
1(
0/
10
#738360000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#738370000000
0!
0'
0/
#738380000000
1!
1'
1/
#738390000000
0!
0'
0/
#738400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#738410000000
0!
0'
0/
#738420000000
1!
1'
1/
#738430000000
0!
1"
0'
1(
0/
10
#738440000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#738450000000
0!
1$
0'
1+
0/
#738460000000
1!
1'
1/
#738470000000
0!
0'
0/
#738480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#738490000000
0!
0'
0/
#738500000000
1!
1'
1/
#738510000000
0!
0'
0/
#738520000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#738530000000
0!
0'
0/
#738540000000
1!
1'
1/
#738550000000
0!
0'
0/
#738560000000
1!
1'
1/
#738570000000
0!
0'
0/
#738580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#738590000000
0!
0'
0/
#738600000000
1!
1'
1/
#738610000000
0!
0'
0/
#738620000000
1!
1'
1/
#738630000000
0!
0'
0/
#738640000000
1!
1'
1/
#738650000000
0!
0'
0/
#738660000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#738670000000
0!
0'
0/
#738680000000
1!
1'
1/
#738690000000
0!
0'
0/
#738700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#738710000000
0!
0'
0/
#738720000000
1!
1'
1/
#738730000000
0!
0'
0/
#738740000000
#738750000000
1!
1'
1/
#738760000000
0!
0'
0/
#738770000000
1!
1'
1/
#738780000000
0!
1"
0'
1(
0/
10
#738790000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#738800000000
0!
0'
0/
#738810000000
1!
1'
1/
#738820000000
0!
0'
0/
#738830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#738840000000
0!
0'
0/
#738850000000
1!
1'
1/
#738860000000
0!
1"
0'
1(
0/
10
#738870000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#738880000000
0!
1$
0'
1+
0/
#738890000000
1!
1'
1/
#738900000000
0!
0'
0/
#738910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#738920000000
0!
0'
0/
#738930000000
1!
1'
1/
#738940000000
0!
0'
0/
#738950000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#738960000000
0!
0'
0/
#738970000000
1!
1'
1/
#738980000000
0!
0'
0/
#738990000000
1!
1'
1/
#739000000000
0!
0'
0/
#739010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#739020000000
0!
0'
0/
#739030000000
1!
1'
1/
#739040000000
0!
0'
0/
#739050000000
1!
1'
1/
#739060000000
0!
0'
0/
#739070000000
1!
1'
1/
#739080000000
0!
0'
0/
#739090000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#739100000000
0!
0'
0/
#739110000000
1!
1'
1/
#739120000000
0!
0'
0/
#739130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#739140000000
0!
0'
0/
#739150000000
1!
1'
1/
#739160000000
0!
0'
0/
#739170000000
#739180000000
1!
1'
1/
#739190000000
0!
0'
0/
#739200000000
1!
1'
1/
#739210000000
0!
1"
0'
1(
0/
10
#739220000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#739230000000
0!
0'
0/
#739240000000
1!
1'
1/
#739250000000
0!
0'
0/
#739260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#739270000000
0!
0'
0/
#739280000000
1!
1'
1/
#739290000000
0!
1"
0'
1(
0/
10
#739300000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#739310000000
0!
1$
0'
1+
0/
#739320000000
1!
1'
1/
#739330000000
0!
0'
0/
#739340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#739350000000
0!
0'
0/
#739360000000
1!
1'
1/
#739370000000
0!
0'
0/
#739380000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#739390000000
0!
0'
0/
#739400000000
1!
1'
1/
#739410000000
0!
0'
0/
#739420000000
1!
1'
1/
#739430000000
0!
0'
0/
#739440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#739450000000
0!
0'
0/
#739460000000
1!
1'
1/
#739470000000
0!
0'
0/
#739480000000
1!
1'
1/
#739490000000
0!
0'
0/
#739500000000
1!
1'
1/
#739510000000
0!
0'
0/
#739520000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#739530000000
0!
0'
0/
#739540000000
1!
1'
1/
#739550000000
0!
0'
0/
#739560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#739570000000
0!
0'
0/
#739580000000
1!
1'
1/
#739590000000
0!
0'
0/
#739600000000
#739610000000
1!
1'
1/
#739620000000
0!
0'
0/
#739630000000
1!
1'
1/
#739640000000
0!
1"
0'
1(
0/
10
#739650000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#739660000000
0!
0'
0/
#739670000000
1!
1'
1/
#739680000000
0!
0'
0/
#739690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#739700000000
0!
0'
0/
#739710000000
1!
1'
1/
#739720000000
0!
1"
0'
1(
0/
10
#739730000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#739740000000
0!
1$
0'
1+
0/
#739750000000
1!
1'
1/
#739760000000
0!
0'
0/
#739770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#739780000000
0!
0'
0/
#739790000000
1!
1'
1/
#739800000000
0!
0'
0/
#739810000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#739820000000
0!
0'
0/
#739830000000
1!
1'
1/
#739840000000
0!
0'
0/
#739850000000
1!
1'
1/
#739860000000
0!
0'
0/
#739870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#739880000000
0!
0'
0/
#739890000000
1!
1'
1/
#739900000000
0!
0'
0/
#739910000000
1!
1'
1/
#739920000000
0!
0'
0/
#739930000000
1!
1'
1/
#739940000000
0!
0'
0/
#739950000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#739960000000
0!
0'
0/
#739970000000
1!
1'
1/
#739980000000
0!
0'
0/
#739990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#740000000000
0!
0'
0/
#740010000000
1!
1'
1/
#740020000000
0!
0'
0/
#740030000000
#740040000000
1!
1'
1/
#740050000000
0!
0'
0/
#740060000000
1!
1'
1/
#740070000000
0!
1"
0'
1(
0/
10
#740080000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#740090000000
0!
0'
0/
#740100000000
1!
1'
1/
#740110000000
0!
0'
0/
#740120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#740130000000
0!
0'
0/
#740140000000
1!
1'
1/
#740150000000
0!
1"
0'
1(
0/
10
#740160000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#740170000000
0!
1$
0'
1+
0/
#740180000000
1!
1'
1/
#740190000000
0!
0'
0/
#740200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#740210000000
0!
0'
0/
#740220000000
1!
1'
1/
#740230000000
0!
0'
0/
#740240000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#740250000000
0!
0'
0/
#740260000000
1!
1'
1/
#740270000000
0!
0'
0/
#740280000000
1!
1'
1/
#740290000000
0!
0'
0/
#740300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#740310000000
0!
0'
0/
#740320000000
1!
1'
1/
#740330000000
0!
0'
0/
#740340000000
1!
1'
1/
#740350000000
0!
0'
0/
#740360000000
1!
1'
1/
#740370000000
0!
0'
0/
#740380000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#740390000000
0!
0'
0/
#740400000000
1!
1'
1/
#740410000000
0!
0'
0/
#740420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#740430000000
0!
0'
0/
#740440000000
1!
1'
1/
#740450000000
0!
0'
0/
#740460000000
#740470000000
1!
1'
1/
#740480000000
0!
0'
0/
#740490000000
1!
1'
1/
#740500000000
0!
1"
0'
1(
0/
10
#740510000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#740520000000
0!
0'
0/
#740530000000
1!
1'
1/
#740540000000
0!
0'
0/
#740550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#740560000000
0!
0'
0/
#740570000000
1!
1'
1/
#740580000000
0!
1"
0'
1(
0/
10
#740590000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#740600000000
0!
1$
0'
1+
0/
#740610000000
1!
1'
1/
#740620000000
0!
0'
0/
#740630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#740640000000
0!
0'
0/
#740650000000
1!
1'
1/
#740660000000
0!
0'
0/
#740670000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#740680000000
0!
0'
0/
#740690000000
1!
1'
1/
#740700000000
0!
0'
0/
#740710000000
1!
1'
1/
#740720000000
0!
0'
0/
#740730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#740740000000
0!
0'
0/
#740750000000
1!
1'
1/
#740760000000
0!
0'
0/
#740770000000
1!
1'
1/
#740780000000
0!
0'
0/
#740790000000
1!
1'
1/
#740800000000
0!
0'
0/
#740810000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#740820000000
0!
0'
0/
#740830000000
1!
1'
1/
#740840000000
0!
0'
0/
#740850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#740860000000
0!
0'
0/
#740870000000
1!
1'
1/
#740880000000
0!
0'
0/
#740890000000
#740900000000
1!
1'
1/
#740910000000
0!
0'
0/
#740920000000
1!
1'
1/
#740930000000
0!
1"
0'
1(
0/
10
#740940000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#740950000000
0!
0'
0/
#740960000000
1!
1'
1/
#740970000000
0!
0'
0/
#740980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#740990000000
0!
0'
0/
#741000000000
1!
1'
1/
#741010000000
0!
1"
0'
1(
0/
10
#741020000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#741030000000
0!
1$
0'
1+
0/
#741040000000
1!
1'
1/
#741050000000
0!
0'
0/
#741060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#741070000000
0!
0'
0/
#741080000000
1!
1'
1/
#741090000000
0!
0'
0/
#741100000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#741110000000
0!
0'
0/
#741120000000
1!
1'
1/
#741130000000
0!
0'
0/
#741140000000
1!
1'
1/
#741150000000
0!
0'
0/
#741160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#741170000000
0!
0'
0/
#741180000000
1!
1'
1/
#741190000000
0!
0'
0/
#741200000000
1!
1'
1/
#741210000000
0!
0'
0/
#741220000000
1!
1'
1/
#741230000000
0!
0'
0/
#741240000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#741250000000
0!
0'
0/
#741260000000
1!
1'
1/
#741270000000
0!
0'
0/
#741280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#741290000000
0!
0'
0/
#741300000000
1!
1'
1/
#741310000000
0!
0'
0/
#741320000000
#741330000000
1!
1'
1/
#741340000000
0!
0'
0/
#741350000000
1!
1'
1/
#741360000000
0!
1"
0'
1(
0/
10
#741370000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#741380000000
0!
0'
0/
#741390000000
1!
1'
1/
#741400000000
0!
0'
0/
#741410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#741420000000
0!
0'
0/
#741430000000
1!
1'
1/
#741440000000
0!
1"
0'
1(
0/
10
#741450000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#741460000000
0!
1$
0'
1+
0/
#741470000000
1!
1'
1/
#741480000000
0!
0'
0/
#741490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#741500000000
0!
0'
0/
#741510000000
1!
1'
1/
#741520000000
0!
0'
0/
#741530000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#741540000000
0!
0'
0/
#741550000000
1!
1'
1/
#741560000000
0!
0'
0/
#741570000000
1!
1'
1/
#741580000000
0!
0'
0/
#741590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#741600000000
0!
0'
0/
#741610000000
1!
1'
1/
#741620000000
0!
0'
0/
#741630000000
1!
1'
1/
#741640000000
0!
0'
0/
#741650000000
1!
1'
1/
#741660000000
0!
0'
0/
#741670000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#741680000000
0!
0'
0/
#741690000000
1!
1'
1/
#741700000000
0!
0'
0/
#741710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#741720000000
0!
0'
0/
#741730000000
1!
1'
1/
#741740000000
0!
0'
0/
#741750000000
#741760000000
1!
1'
1/
#741770000000
0!
0'
0/
#741780000000
1!
1'
1/
#741790000000
0!
1"
0'
1(
0/
10
#741800000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#741810000000
0!
0'
0/
#741820000000
1!
1'
1/
#741830000000
0!
0'
0/
#741840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#741850000000
0!
0'
0/
#741860000000
1!
1'
1/
#741870000000
0!
1"
0'
1(
0/
10
#741880000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#741890000000
0!
1$
0'
1+
0/
#741900000000
1!
1'
1/
#741910000000
0!
0'
0/
#741920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#741930000000
0!
0'
0/
#741940000000
1!
1'
1/
#741950000000
0!
0'
0/
#741960000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#741970000000
0!
0'
0/
#741980000000
1!
1'
1/
#741990000000
0!
0'
0/
#742000000000
1!
1'
1/
#742010000000
0!
0'
0/
#742020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#742030000000
0!
0'
0/
#742040000000
1!
1'
1/
#742050000000
0!
0'
0/
#742060000000
1!
1'
1/
#742070000000
0!
0'
0/
#742080000000
1!
1'
1/
#742090000000
0!
0'
0/
#742100000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#742110000000
0!
0'
0/
#742120000000
1!
1'
1/
#742130000000
0!
0'
0/
#742140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#742150000000
0!
0'
0/
#742160000000
1!
1'
1/
#742170000000
0!
0'
0/
#742180000000
#742190000000
1!
1'
1/
#742200000000
0!
0'
0/
#742210000000
1!
1'
1/
#742220000000
0!
1"
0'
1(
0/
10
#742230000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#742240000000
0!
0'
0/
#742250000000
1!
1'
1/
#742260000000
0!
0'
0/
#742270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#742280000000
0!
0'
0/
#742290000000
1!
1'
1/
#742300000000
0!
1"
0'
1(
0/
10
#742310000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#742320000000
0!
1$
0'
1+
0/
#742330000000
1!
1'
1/
#742340000000
0!
0'
0/
#742350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#742360000000
0!
0'
0/
#742370000000
1!
1'
1/
#742380000000
0!
0'
0/
#742390000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#742400000000
0!
0'
0/
#742410000000
1!
1'
1/
#742420000000
0!
0'
0/
#742430000000
1!
1'
1/
#742440000000
0!
0'
0/
#742450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#742460000000
0!
0'
0/
#742470000000
1!
1'
1/
#742480000000
0!
0'
0/
#742490000000
1!
1'
1/
#742500000000
0!
0'
0/
#742510000000
1!
1'
1/
#742520000000
0!
0'
0/
#742530000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#742540000000
0!
0'
0/
#742550000000
1!
1'
1/
#742560000000
0!
0'
0/
#742570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#742580000000
0!
0'
0/
#742590000000
1!
1'
1/
#742600000000
0!
0'
0/
#742610000000
#742620000000
1!
1'
1/
#742630000000
0!
0'
0/
#742640000000
1!
1'
1/
#742650000000
0!
1"
0'
1(
0/
10
#742660000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#742670000000
0!
0'
0/
#742680000000
1!
1'
1/
#742690000000
0!
0'
0/
#742700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#742710000000
0!
0'
0/
#742720000000
1!
1'
1/
#742730000000
0!
1"
0'
1(
0/
10
#742740000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#742750000000
0!
1$
0'
1+
0/
#742760000000
1!
1'
1/
#742770000000
0!
0'
0/
#742780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#742790000000
0!
0'
0/
#742800000000
1!
1'
1/
#742810000000
0!
0'
0/
#742820000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#742830000000
0!
0'
0/
#742840000000
1!
1'
1/
#742850000000
0!
0'
0/
#742860000000
1!
1'
1/
#742870000000
0!
0'
0/
#742880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#742890000000
0!
0'
0/
#742900000000
1!
1'
1/
#742910000000
0!
0'
0/
#742920000000
1!
1'
1/
#742930000000
0!
0'
0/
#742940000000
1!
1'
1/
#742950000000
0!
0'
0/
#742960000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#742970000000
0!
0'
0/
#742980000000
1!
1'
1/
#742990000000
0!
0'
0/
#743000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#743010000000
0!
0'
0/
#743020000000
1!
1'
1/
#743030000000
0!
0'
0/
#743040000000
#743050000000
1!
1'
1/
#743060000000
0!
0'
0/
#743070000000
1!
1'
1/
#743080000000
0!
1"
0'
1(
0/
10
#743090000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#743100000000
0!
0'
0/
#743110000000
1!
1'
1/
#743120000000
0!
0'
0/
#743130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#743140000000
0!
0'
0/
#743150000000
1!
1'
1/
#743160000000
0!
1"
0'
1(
0/
10
#743170000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#743180000000
0!
1$
0'
1+
0/
#743190000000
1!
1'
1/
#743200000000
0!
0'
0/
#743210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#743220000000
0!
0'
0/
#743230000000
1!
1'
1/
#743240000000
0!
0'
0/
#743250000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#743260000000
0!
0'
0/
#743270000000
1!
1'
1/
#743280000000
0!
0'
0/
#743290000000
1!
1'
1/
#743300000000
0!
0'
0/
#743310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#743320000000
0!
0'
0/
#743330000000
1!
1'
1/
#743340000000
0!
0'
0/
#743350000000
1!
1'
1/
#743360000000
0!
0'
0/
#743370000000
1!
1'
1/
#743380000000
0!
0'
0/
#743390000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#743400000000
0!
0'
0/
#743410000000
1!
1'
1/
#743420000000
0!
0'
0/
#743430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#743440000000
0!
0'
0/
#743450000000
1!
1'
1/
#743460000000
0!
0'
0/
#743470000000
#743480000000
1!
1'
1/
#743490000000
0!
0'
0/
#743500000000
1!
1'
1/
#743510000000
0!
1"
0'
1(
0/
10
#743520000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#743530000000
0!
0'
0/
#743540000000
1!
1'
1/
#743550000000
0!
0'
0/
#743560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#743570000000
0!
0'
0/
#743580000000
1!
1'
1/
#743590000000
0!
1"
0'
1(
0/
10
#743600000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#743610000000
0!
1$
0'
1+
0/
#743620000000
1!
1'
1/
#743630000000
0!
0'
0/
#743640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#743650000000
0!
0'
0/
#743660000000
1!
1'
1/
#743670000000
0!
0'
0/
#743680000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#743690000000
0!
0'
0/
#743700000000
1!
1'
1/
#743710000000
0!
0'
0/
#743720000000
1!
1'
1/
#743730000000
0!
0'
0/
#743740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#743750000000
0!
0'
0/
#743760000000
1!
1'
1/
#743770000000
0!
0'
0/
#743780000000
1!
1'
1/
#743790000000
0!
0'
0/
#743800000000
1!
1'
1/
#743810000000
0!
0'
0/
#743820000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#743830000000
0!
0'
0/
#743840000000
1!
1'
1/
#743850000000
0!
0'
0/
#743860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#743870000000
0!
0'
0/
#743880000000
1!
1'
1/
#743890000000
0!
0'
0/
#743900000000
#743910000000
1!
1'
1/
#743920000000
0!
0'
0/
#743930000000
1!
1'
1/
#743940000000
0!
1"
0'
1(
0/
10
#743950000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#743960000000
0!
0'
0/
#743970000000
1!
1'
1/
#743980000000
0!
0'
0/
#743990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#744000000000
0!
0'
0/
#744010000000
1!
1'
1/
#744020000000
0!
1"
0'
1(
0/
10
#744030000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#744040000000
0!
1$
0'
1+
0/
#744050000000
1!
1'
1/
#744060000000
0!
0'
0/
#744070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#744080000000
0!
0'
0/
#744090000000
1!
1'
1/
#744100000000
0!
0'
0/
#744110000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#744120000000
0!
0'
0/
#744130000000
1!
1'
1/
#744140000000
0!
0'
0/
#744150000000
1!
1'
1/
#744160000000
0!
0'
0/
#744170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#744180000000
0!
0'
0/
#744190000000
1!
1'
1/
#744200000000
0!
0'
0/
#744210000000
1!
1'
1/
#744220000000
0!
0'
0/
#744230000000
1!
1'
1/
#744240000000
0!
0'
0/
#744250000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#744260000000
0!
0'
0/
#744270000000
1!
1'
1/
#744280000000
0!
0'
0/
#744290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#744300000000
0!
0'
0/
#744310000000
1!
1'
1/
#744320000000
0!
0'
0/
#744330000000
#744340000000
1!
1'
1/
#744350000000
0!
0'
0/
#744360000000
1!
1'
1/
#744370000000
0!
1"
0'
1(
0/
10
#744380000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#744390000000
0!
0'
0/
#744400000000
1!
1'
1/
#744410000000
0!
0'
0/
#744420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#744430000000
0!
0'
0/
#744440000000
1!
1'
1/
#744450000000
0!
1"
0'
1(
0/
10
#744460000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#744470000000
0!
1$
0'
1+
0/
#744480000000
1!
1'
1/
#744490000000
0!
0'
0/
#744500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#744510000000
0!
0'
0/
#744520000000
1!
1'
1/
#744530000000
0!
0'
0/
#744540000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#744550000000
0!
0'
0/
#744560000000
1!
1'
1/
#744570000000
0!
0'
0/
#744580000000
1!
1'
1/
#744590000000
0!
0'
0/
#744600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#744610000000
0!
0'
0/
#744620000000
1!
1'
1/
#744630000000
0!
0'
0/
#744640000000
1!
1'
1/
#744650000000
0!
0'
0/
#744660000000
1!
1'
1/
#744670000000
0!
0'
0/
#744680000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#744690000000
0!
0'
0/
#744700000000
1!
1'
1/
#744710000000
0!
0'
0/
#744720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#744730000000
0!
0'
0/
#744740000000
1!
1'
1/
#744750000000
0!
0'
0/
#744760000000
#744770000000
1!
1'
1/
#744780000000
0!
0'
0/
#744790000000
1!
1'
1/
#744800000000
0!
1"
0'
1(
0/
10
#744810000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#744820000000
0!
0'
0/
#744830000000
1!
1'
1/
#744840000000
0!
0'
0/
#744850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#744860000000
0!
0'
0/
#744870000000
1!
1'
1/
#744880000000
0!
1"
0'
1(
0/
10
#744890000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#744900000000
0!
1$
0'
1+
0/
#744910000000
1!
1'
1/
#744920000000
0!
0'
0/
#744930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#744940000000
0!
0'
0/
#744950000000
1!
1'
1/
#744960000000
0!
0'
0/
#744970000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#744980000000
0!
0'
0/
#744990000000
1!
1'
1/
#745000000000
0!
0'
0/
#745010000000
1!
1'
1/
#745020000000
0!
0'
0/
#745030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#745040000000
0!
0'
0/
#745050000000
1!
1'
1/
#745060000000
0!
0'
0/
#745070000000
1!
1'
1/
#745080000000
0!
0'
0/
#745090000000
1!
1'
1/
#745100000000
0!
0'
0/
#745110000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#745120000000
0!
0'
0/
#745130000000
1!
1'
1/
#745140000000
0!
0'
0/
#745150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#745160000000
0!
0'
0/
#745170000000
1!
1'
1/
#745180000000
0!
0'
0/
#745190000000
#745200000000
1!
1'
1/
#745210000000
0!
0'
0/
#745220000000
1!
1'
1/
#745230000000
0!
1"
0'
1(
0/
10
#745240000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#745250000000
0!
0'
0/
#745260000000
1!
1'
1/
#745270000000
0!
0'
0/
#745280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#745290000000
0!
0'
0/
#745300000000
1!
1'
1/
#745310000000
0!
1"
0'
1(
0/
10
#745320000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#745330000000
0!
1$
0'
1+
0/
#745340000000
1!
1'
1/
#745350000000
0!
0'
0/
#745360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#745370000000
0!
0'
0/
#745380000000
1!
1'
1/
#745390000000
0!
0'
0/
#745400000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#745410000000
0!
0'
0/
#745420000000
1!
1'
1/
#745430000000
0!
0'
0/
#745440000000
1!
1'
1/
#745450000000
0!
0'
0/
#745460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#745470000000
0!
0'
0/
#745480000000
1!
1'
1/
#745490000000
0!
0'
0/
#745500000000
1!
1'
1/
#745510000000
0!
0'
0/
#745520000000
1!
1'
1/
#745530000000
0!
0'
0/
#745540000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#745550000000
0!
0'
0/
#745560000000
1!
1'
1/
#745570000000
0!
0'
0/
#745580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#745590000000
0!
0'
0/
#745600000000
1!
1'
1/
#745610000000
0!
0'
0/
#745620000000
#745630000000
1!
1'
1/
#745640000000
0!
0'
0/
#745650000000
1!
1'
1/
#745660000000
0!
1"
0'
1(
0/
10
#745670000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#745680000000
0!
0'
0/
#745690000000
1!
1'
1/
#745700000000
0!
0'
0/
#745710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#745720000000
0!
0'
0/
#745730000000
1!
1'
1/
#745740000000
0!
1"
0'
1(
0/
10
#745750000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#745760000000
0!
1$
0'
1+
0/
#745770000000
1!
1'
1/
#745780000000
0!
0'
0/
#745790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#745800000000
0!
0'
0/
#745810000000
1!
1'
1/
#745820000000
0!
0'
0/
#745830000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#745840000000
0!
0'
0/
#745850000000
1!
1'
1/
#745860000000
0!
0'
0/
#745870000000
1!
1'
1/
#745880000000
0!
0'
0/
#745890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#745900000000
0!
0'
0/
#745910000000
1!
1'
1/
#745920000000
0!
0'
0/
#745930000000
1!
1'
1/
#745940000000
0!
0'
0/
#745950000000
1!
1'
1/
#745960000000
0!
0'
0/
#745970000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#745980000000
0!
0'
0/
#745990000000
1!
1'
1/
#746000000000
0!
0'
0/
#746010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#746020000000
0!
0'
0/
#746030000000
1!
1'
1/
#746040000000
0!
0'
0/
#746050000000
#746060000000
1!
1'
1/
#746070000000
0!
0'
0/
#746080000000
1!
1'
1/
#746090000000
0!
1"
0'
1(
0/
10
#746100000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#746110000000
0!
0'
0/
#746120000000
1!
1'
1/
#746130000000
0!
0'
0/
#746140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#746150000000
0!
0'
0/
#746160000000
1!
1'
1/
#746170000000
0!
1"
0'
1(
0/
10
#746180000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#746190000000
0!
1$
0'
1+
0/
#746200000000
1!
1'
1/
#746210000000
0!
0'
0/
#746220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#746230000000
0!
0'
0/
#746240000000
1!
1'
1/
#746250000000
0!
0'
0/
#746260000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#746270000000
0!
0'
0/
#746280000000
1!
1'
1/
#746290000000
0!
0'
0/
#746300000000
1!
1'
1/
#746310000000
0!
0'
0/
#746320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#746330000000
0!
0'
0/
#746340000000
1!
1'
1/
#746350000000
0!
0'
0/
#746360000000
1!
1'
1/
#746370000000
0!
0'
0/
#746380000000
1!
1'
1/
#746390000000
0!
0'
0/
#746400000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#746410000000
0!
0'
0/
#746420000000
1!
1'
1/
#746430000000
0!
0'
0/
#746440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#746450000000
0!
0'
0/
#746460000000
1!
1'
1/
#746470000000
0!
0'
0/
#746480000000
#746490000000
1!
1'
1/
#746500000000
0!
0'
0/
#746510000000
1!
1'
1/
#746520000000
0!
1"
0'
1(
0/
10
#746530000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#746540000000
0!
0'
0/
#746550000000
1!
1'
1/
#746560000000
0!
0'
0/
#746570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#746580000000
0!
0'
0/
#746590000000
1!
1'
1/
#746600000000
0!
1"
0'
1(
0/
10
#746610000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#746620000000
0!
1$
0'
1+
0/
#746630000000
1!
1'
1/
#746640000000
0!
0'
0/
#746650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#746660000000
0!
0'
0/
#746670000000
1!
1'
1/
#746680000000
0!
0'
0/
#746690000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#746700000000
0!
0'
0/
#746710000000
1!
1'
1/
#746720000000
0!
0'
0/
#746730000000
1!
1'
1/
#746740000000
0!
0'
0/
#746750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#746760000000
0!
0'
0/
#746770000000
1!
1'
1/
#746780000000
0!
0'
0/
#746790000000
1!
1'
1/
#746800000000
0!
0'
0/
#746810000000
1!
1'
1/
#746820000000
0!
0'
0/
#746830000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#746840000000
0!
0'
0/
#746850000000
1!
1'
1/
#746860000000
0!
0'
0/
#746870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#746880000000
0!
0'
0/
#746890000000
1!
1'
1/
#746900000000
0!
0'
0/
#746910000000
#746920000000
1!
1'
1/
#746930000000
0!
0'
0/
#746940000000
1!
1'
1/
#746950000000
0!
1"
0'
1(
0/
10
#746960000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#746970000000
0!
0'
0/
#746980000000
1!
1'
1/
#746990000000
0!
0'
0/
#747000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#747010000000
0!
0'
0/
#747020000000
1!
1'
1/
#747030000000
0!
1"
0'
1(
0/
10
#747040000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#747050000000
0!
1$
0'
1+
0/
#747060000000
1!
1'
1/
#747070000000
0!
0'
0/
#747080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#747090000000
0!
0'
0/
#747100000000
1!
1'
1/
#747110000000
0!
0'
0/
#747120000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#747130000000
0!
0'
0/
#747140000000
1!
1'
1/
#747150000000
0!
0'
0/
#747160000000
1!
1'
1/
#747170000000
0!
0'
0/
#747180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#747190000000
0!
0'
0/
#747200000000
1!
1'
1/
#747210000000
0!
0'
0/
#747220000000
1!
1'
1/
#747230000000
0!
0'
0/
#747240000000
1!
1'
1/
#747250000000
0!
0'
0/
#747260000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#747270000000
0!
0'
0/
#747280000000
1!
1'
1/
#747290000000
0!
0'
0/
#747300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#747310000000
0!
0'
0/
#747320000000
1!
1'
1/
#747330000000
0!
0'
0/
#747340000000
#747350000000
1!
1'
1/
#747360000000
0!
0'
0/
#747370000000
1!
1'
1/
#747380000000
0!
1"
0'
1(
0/
10
#747390000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#747400000000
0!
0'
0/
#747410000000
1!
1'
1/
#747420000000
0!
0'
0/
#747430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#747440000000
0!
0'
0/
#747450000000
1!
1'
1/
#747460000000
0!
1"
0'
1(
0/
10
#747470000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#747480000000
0!
1$
0'
1+
0/
#747490000000
1!
1'
1/
#747500000000
0!
0'
0/
#747510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#747520000000
0!
0'
0/
#747530000000
1!
1'
1/
#747540000000
0!
0'
0/
#747550000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#747560000000
0!
0'
0/
#747570000000
1!
1'
1/
#747580000000
0!
0'
0/
#747590000000
1!
1'
1/
#747600000000
0!
0'
0/
#747610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#747620000000
0!
0'
0/
#747630000000
1!
1'
1/
#747640000000
0!
0'
0/
#747650000000
1!
1'
1/
#747660000000
0!
0'
0/
#747670000000
1!
1'
1/
#747680000000
0!
0'
0/
#747690000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#747700000000
0!
0'
0/
#747710000000
1!
1'
1/
#747720000000
0!
0'
0/
#747730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#747740000000
0!
0'
0/
#747750000000
1!
1'
1/
#747760000000
0!
0'
0/
#747770000000
#747780000000
1!
1'
1/
#747790000000
0!
0'
0/
#747800000000
1!
1'
1/
#747810000000
0!
1"
0'
1(
0/
10
#747820000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#747830000000
0!
0'
0/
#747840000000
1!
1'
1/
#747850000000
0!
0'
0/
#747860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#747870000000
0!
0'
0/
#747880000000
1!
1'
1/
#747890000000
0!
1"
0'
1(
0/
10
#747900000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#747910000000
0!
1$
0'
1+
0/
#747920000000
1!
1'
1/
#747930000000
0!
0'
0/
#747940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#747950000000
0!
0'
0/
#747960000000
1!
1'
1/
#747970000000
0!
0'
0/
#747980000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#747990000000
0!
0'
0/
#748000000000
1!
1'
1/
#748010000000
0!
0'
0/
#748020000000
1!
1'
1/
#748030000000
0!
0'
0/
#748040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#748050000000
0!
0'
0/
#748060000000
1!
1'
1/
#748070000000
0!
0'
0/
#748080000000
1!
1'
1/
#748090000000
0!
0'
0/
#748100000000
1!
1'
1/
#748110000000
0!
0'
0/
#748120000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#748130000000
0!
0'
0/
#748140000000
1!
1'
1/
#748150000000
0!
0'
0/
#748160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#748170000000
0!
0'
0/
#748180000000
1!
1'
1/
#748190000000
0!
0'
0/
#748200000000
#748210000000
1!
1'
1/
#748220000000
0!
0'
0/
#748230000000
1!
1'
1/
#748240000000
0!
1"
0'
1(
0/
10
#748250000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#748260000000
0!
0'
0/
#748270000000
1!
1'
1/
#748280000000
0!
0'
0/
#748290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#748300000000
0!
0'
0/
#748310000000
1!
1'
1/
#748320000000
0!
1"
0'
1(
0/
10
#748330000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#748340000000
0!
1$
0'
1+
0/
#748350000000
1!
1'
1/
#748360000000
0!
0'
0/
#748370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#748380000000
0!
0'
0/
#748390000000
1!
1'
1/
#748400000000
0!
0'
0/
#748410000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#748420000000
0!
0'
0/
#748430000000
1!
1'
1/
#748440000000
0!
0'
0/
#748450000000
1!
1'
1/
#748460000000
0!
0'
0/
#748470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#748480000000
0!
0'
0/
#748490000000
1!
1'
1/
#748500000000
0!
0'
0/
#748510000000
1!
1'
1/
#748520000000
0!
0'
0/
#748530000000
1!
1'
1/
#748540000000
0!
0'
0/
#748550000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#748560000000
0!
0'
0/
#748570000000
1!
1'
1/
#748580000000
0!
0'
0/
#748590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#748600000000
0!
0'
0/
#748610000000
1!
1'
1/
#748620000000
0!
0'
0/
#748630000000
#748640000000
1!
1'
1/
#748650000000
0!
0'
0/
#748660000000
1!
1'
1/
#748670000000
0!
1"
0'
1(
0/
10
#748680000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#748690000000
0!
0'
0/
#748700000000
1!
1'
1/
#748710000000
0!
0'
0/
#748720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#748730000000
0!
0'
0/
#748740000000
1!
1'
1/
#748750000000
0!
1"
0'
1(
0/
10
#748760000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#748770000000
0!
1$
0'
1+
0/
#748780000000
1!
1'
1/
#748790000000
0!
0'
0/
#748800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#748810000000
0!
0'
0/
#748820000000
1!
1'
1/
#748830000000
0!
0'
0/
#748840000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#748850000000
0!
0'
0/
#748860000000
1!
1'
1/
#748870000000
0!
0'
0/
#748880000000
1!
1'
1/
#748890000000
0!
0'
0/
#748900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#748910000000
0!
0'
0/
#748920000000
1!
1'
1/
#748930000000
0!
0'
0/
#748940000000
1!
1'
1/
#748950000000
0!
0'
0/
#748960000000
1!
1'
1/
#748970000000
0!
0'
0/
#748980000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#748990000000
0!
0'
0/
#749000000000
1!
1'
1/
#749010000000
0!
0'
0/
#749020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#749030000000
0!
0'
0/
#749040000000
1!
1'
1/
#749050000000
0!
0'
0/
#749060000000
#749070000000
1!
1'
1/
#749080000000
0!
0'
0/
#749090000000
1!
1'
1/
#749100000000
0!
1"
0'
1(
0/
10
#749110000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#749120000000
0!
0'
0/
#749130000000
1!
1'
1/
#749140000000
0!
0'
0/
#749150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#749160000000
0!
0'
0/
#749170000000
1!
1'
1/
#749180000000
0!
1"
0'
1(
0/
10
#749190000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#749200000000
0!
1$
0'
1+
0/
#749210000000
1!
1'
1/
#749220000000
0!
0'
0/
#749230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#749240000000
0!
0'
0/
#749250000000
1!
1'
1/
#749260000000
0!
0'
0/
#749270000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#749280000000
0!
0'
0/
#749290000000
1!
1'
1/
#749300000000
0!
0'
0/
#749310000000
1!
1'
1/
#749320000000
0!
0'
0/
#749330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#749340000000
0!
0'
0/
#749350000000
1!
1'
1/
#749360000000
0!
0'
0/
#749370000000
1!
1'
1/
#749380000000
0!
0'
0/
#749390000000
1!
1'
1/
#749400000000
0!
0'
0/
#749410000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#749420000000
0!
0'
0/
#749430000000
1!
1'
1/
#749440000000
0!
0'
0/
#749450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#749460000000
0!
0'
0/
#749470000000
1!
1'
1/
#749480000000
0!
0'
0/
#749490000000
#749500000000
1!
1'
1/
#749510000000
0!
0'
0/
#749520000000
1!
1'
1/
#749530000000
0!
1"
0'
1(
0/
10
#749540000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#749550000000
0!
0'
0/
#749560000000
1!
1'
1/
#749570000000
0!
0'
0/
#749580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#749590000000
0!
0'
0/
#749600000000
1!
1'
1/
#749610000000
0!
1"
0'
1(
0/
10
#749620000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#749630000000
0!
1$
0'
1+
0/
#749640000000
1!
1'
1/
#749650000000
0!
0'
0/
#749660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#749670000000
0!
0'
0/
#749680000000
1!
1'
1/
#749690000000
0!
0'
0/
#749700000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#749710000000
0!
0'
0/
#749720000000
1!
1'
1/
#749730000000
0!
0'
0/
#749740000000
1!
1'
1/
#749750000000
0!
0'
0/
#749760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#749770000000
0!
0'
0/
#749780000000
1!
1'
1/
#749790000000
0!
0'
0/
#749800000000
1!
1'
1/
#749810000000
0!
0'
0/
#749820000000
1!
1'
1/
#749830000000
0!
0'
0/
#749840000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#749850000000
0!
0'
0/
#749860000000
1!
1'
1/
#749870000000
0!
0'
0/
#749880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#749890000000
0!
0'
0/
#749900000000
1!
1'
1/
#749910000000
0!
0'
0/
#749920000000
#749930000000
1!
1'
1/
#749940000000
0!
0'
0/
#749950000000
1!
1'
1/
#749960000000
0!
1"
0'
1(
0/
10
#749970000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#749980000000
0!
0'
0/
#749990000000
1!
1'
1/
#750000000000
0!
0'
0/
#750010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#750020000000
0!
0'
0/
#750030000000
1!
1'
1/
#750040000000
0!
1"
0'
1(
0/
10
#750050000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#750060000000
0!
1$
0'
1+
0/
#750070000000
1!
1'
1/
#750080000000
0!
0'
0/
#750090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#750100000000
0!
0'
0/
#750110000000
1!
1'
1/
#750120000000
0!
0'
0/
#750130000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#750140000000
0!
0'
0/
#750150000000
1!
1'
1/
#750160000000
0!
0'
0/
#750170000000
1!
1'
1/
#750180000000
0!
0'
0/
#750190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#750200000000
0!
0'
0/
#750210000000
1!
1'
1/
#750220000000
0!
0'
0/
#750230000000
1!
1'
1/
#750240000000
0!
0'
0/
#750250000000
1!
1'
1/
#750260000000
0!
0'
0/
#750270000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#750280000000
0!
0'
0/
#750290000000
1!
1'
1/
#750300000000
0!
0'
0/
#750310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#750320000000
0!
0'
0/
#750330000000
1!
1'
1/
#750340000000
0!
0'
0/
#750350000000
#750360000000
1!
1'
1/
#750370000000
0!
0'
0/
#750380000000
1!
1'
1/
#750390000000
0!
1"
0'
1(
0/
10
#750400000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#750410000000
0!
0'
0/
#750420000000
1!
1'
1/
#750430000000
0!
0'
0/
#750440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#750450000000
0!
0'
0/
#750460000000
1!
1'
1/
#750470000000
0!
1"
0'
1(
0/
10
#750480000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#750490000000
0!
1$
0'
1+
0/
#750500000000
1!
1'
1/
#750510000000
0!
0'
0/
#750520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#750530000000
0!
0'
0/
#750540000000
1!
1'
1/
#750550000000
0!
0'
0/
#750560000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#750570000000
0!
0'
0/
#750580000000
1!
1'
1/
#750590000000
0!
0'
0/
#750600000000
1!
1'
1/
#750610000000
0!
0'
0/
#750620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#750630000000
0!
0'
0/
#750640000000
1!
1'
1/
#750650000000
0!
0'
0/
#750660000000
1!
1'
1/
#750670000000
0!
0'
0/
#750680000000
1!
1'
1/
#750690000000
0!
0'
0/
#750700000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#750710000000
0!
0'
0/
#750720000000
1!
1'
1/
#750730000000
0!
0'
0/
#750740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#750750000000
0!
0'
0/
#750760000000
1!
1'
1/
#750770000000
0!
0'
0/
#750780000000
#750790000000
1!
1'
1/
#750800000000
0!
0'
0/
#750810000000
1!
1'
1/
#750820000000
0!
1"
0'
1(
0/
10
#750830000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#750840000000
0!
0'
0/
#750850000000
1!
1'
1/
#750860000000
0!
0'
0/
#750870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#750880000000
0!
0'
0/
#750890000000
1!
1'
1/
#750900000000
0!
1"
0'
1(
0/
10
#750910000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#750920000000
0!
1$
0'
1+
0/
#750930000000
1!
1'
1/
#750940000000
0!
0'
0/
#750950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#750960000000
0!
0'
0/
#750970000000
1!
1'
1/
#750980000000
0!
0'
0/
#750990000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#751000000000
0!
0'
0/
#751010000000
1!
1'
1/
#751020000000
0!
0'
0/
#751030000000
1!
1'
1/
#751040000000
0!
0'
0/
#751050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#751060000000
0!
0'
0/
#751070000000
1!
1'
1/
#751080000000
0!
0'
0/
#751090000000
1!
1'
1/
#751100000000
0!
0'
0/
#751110000000
1!
1'
1/
#751120000000
0!
0'
0/
#751130000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#751140000000
0!
0'
0/
#751150000000
1!
1'
1/
#751160000000
0!
0'
0/
#751170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#751180000000
0!
0'
0/
#751190000000
1!
1'
1/
#751200000000
0!
0'
0/
#751210000000
#751220000000
1!
1'
1/
#751230000000
0!
0'
0/
#751240000000
1!
1'
1/
#751250000000
0!
1"
0'
1(
0/
10
#751260000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#751270000000
0!
0'
0/
#751280000000
1!
1'
1/
#751290000000
0!
0'
0/
#751300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#751310000000
0!
0'
0/
#751320000000
1!
1'
1/
#751330000000
0!
1"
0'
1(
0/
10
#751340000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#751350000000
0!
1$
0'
1+
0/
#751360000000
1!
1'
1/
#751370000000
0!
0'
0/
#751380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#751390000000
0!
0'
0/
#751400000000
1!
1'
1/
#751410000000
0!
0'
0/
#751420000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#751430000000
0!
0'
0/
#751440000000
1!
1'
1/
#751450000000
0!
0'
0/
#751460000000
1!
1'
1/
#751470000000
0!
0'
0/
#751480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#751490000000
0!
0'
0/
#751500000000
1!
1'
1/
#751510000000
0!
0'
0/
#751520000000
1!
1'
1/
#751530000000
0!
0'
0/
#751540000000
1!
1'
1/
#751550000000
0!
0'
0/
#751560000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#751570000000
0!
0'
0/
#751580000000
1!
1'
1/
#751590000000
0!
0'
0/
#751600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#751610000000
0!
0'
0/
#751620000000
1!
1'
1/
#751630000000
0!
0'
0/
#751640000000
#751650000000
1!
1'
1/
#751660000000
0!
0'
0/
#751670000000
1!
1'
1/
#751680000000
0!
1"
0'
1(
0/
10
#751690000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#751700000000
0!
0'
0/
#751710000000
1!
1'
1/
#751720000000
0!
0'
0/
#751730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#751740000000
0!
0'
0/
#751750000000
1!
1'
1/
#751760000000
0!
1"
0'
1(
0/
10
#751770000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#751780000000
0!
1$
0'
1+
0/
#751790000000
1!
1'
1/
#751800000000
0!
0'
0/
#751810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#751820000000
0!
0'
0/
#751830000000
1!
1'
1/
#751840000000
0!
0'
0/
#751850000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#751860000000
0!
0'
0/
#751870000000
1!
1'
1/
#751880000000
0!
0'
0/
#751890000000
1!
1'
1/
#751900000000
0!
0'
0/
#751910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#751920000000
0!
0'
0/
#751930000000
1!
1'
1/
#751940000000
0!
0'
0/
#751950000000
1!
1'
1/
#751960000000
0!
0'
0/
#751970000000
1!
1'
1/
#751980000000
0!
0'
0/
#751990000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#752000000000
0!
0'
0/
#752010000000
1!
1'
1/
#752020000000
0!
0'
0/
#752030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#752040000000
0!
0'
0/
#752050000000
1!
1'
1/
#752060000000
0!
0'
0/
#752070000000
#752080000000
1!
1'
1/
#752090000000
0!
0'
0/
#752100000000
1!
1'
1/
#752110000000
0!
1"
0'
1(
0/
10
#752120000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#752130000000
0!
0'
0/
#752140000000
1!
1'
1/
#752150000000
0!
0'
0/
#752160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#752170000000
0!
0'
0/
#752180000000
1!
1'
1/
#752190000000
0!
1"
0'
1(
0/
10
#752200000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#752210000000
0!
1$
0'
1+
0/
#752220000000
1!
1'
1/
#752230000000
0!
0'
0/
#752240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#752250000000
0!
0'
0/
#752260000000
1!
1'
1/
#752270000000
0!
0'
0/
#752280000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#752290000000
0!
0'
0/
#752300000000
1!
1'
1/
#752310000000
0!
0'
0/
#752320000000
1!
1'
1/
#752330000000
0!
0'
0/
#752340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#752350000000
0!
0'
0/
#752360000000
1!
1'
1/
#752370000000
0!
0'
0/
#752380000000
1!
1'
1/
#752390000000
0!
0'
0/
#752400000000
1!
1'
1/
#752410000000
0!
0'
0/
#752420000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#752430000000
0!
0'
0/
#752440000000
1!
1'
1/
#752450000000
0!
0'
0/
#752460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#752470000000
0!
0'
0/
#752480000000
1!
1'
1/
#752490000000
0!
0'
0/
#752500000000
#752510000000
1!
1'
1/
#752520000000
0!
0'
0/
#752530000000
1!
1'
1/
#752540000000
0!
1"
0'
1(
0/
10
#752550000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#752560000000
0!
0'
0/
#752570000000
1!
1'
1/
#752580000000
0!
0'
0/
#752590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#752600000000
0!
0'
0/
#752610000000
1!
1'
1/
#752620000000
0!
1"
0'
1(
0/
10
#752630000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#752640000000
0!
1$
0'
1+
0/
#752650000000
1!
1'
1/
#752660000000
0!
0'
0/
#752670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#752680000000
0!
0'
0/
#752690000000
1!
1'
1/
#752700000000
0!
0'
0/
#752710000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#752720000000
0!
0'
0/
#752730000000
1!
1'
1/
#752740000000
0!
0'
0/
#752750000000
1!
1'
1/
#752760000000
0!
0'
0/
#752770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#752780000000
0!
0'
0/
#752790000000
1!
1'
1/
#752800000000
0!
0'
0/
#752810000000
1!
1'
1/
#752820000000
0!
0'
0/
#752830000000
1!
1'
1/
#752840000000
0!
0'
0/
#752850000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#752860000000
0!
0'
0/
#752870000000
1!
1'
1/
#752880000000
0!
0'
0/
#752890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#752900000000
0!
0'
0/
#752910000000
1!
1'
1/
#752920000000
0!
0'
0/
#752930000000
#752940000000
1!
1'
1/
#752950000000
0!
0'
0/
#752960000000
1!
1'
1/
#752970000000
0!
1"
0'
1(
0/
10
#752980000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#752990000000
0!
0'
0/
#753000000000
1!
1'
1/
#753010000000
0!
0'
0/
#753020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#753030000000
0!
0'
0/
#753040000000
1!
1'
1/
#753050000000
0!
1"
0'
1(
0/
10
#753060000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#753070000000
0!
1$
0'
1+
0/
#753080000000
1!
1'
1/
#753090000000
0!
0'
0/
#753100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#753110000000
0!
0'
0/
#753120000000
1!
1'
1/
#753130000000
0!
0'
0/
#753140000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#753150000000
0!
0'
0/
#753160000000
1!
1'
1/
#753170000000
0!
0'
0/
#753180000000
1!
1'
1/
#753190000000
0!
0'
0/
#753200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#753210000000
0!
0'
0/
#753220000000
1!
1'
1/
#753230000000
0!
0'
0/
#753240000000
1!
1'
1/
#753250000000
0!
0'
0/
#753260000000
1!
1'
1/
#753270000000
0!
0'
0/
#753280000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#753290000000
0!
0'
0/
#753300000000
1!
1'
1/
#753310000000
0!
0'
0/
#753320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#753330000000
0!
0'
0/
#753340000000
1!
1'
1/
#753350000000
0!
0'
0/
#753360000000
#753370000000
1!
1'
1/
#753380000000
0!
0'
0/
#753390000000
1!
1'
1/
#753400000000
0!
1"
0'
1(
0/
10
#753410000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#753420000000
0!
0'
0/
#753430000000
1!
1'
1/
#753440000000
0!
0'
0/
#753450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#753460000000
0!
0'
0/
#753470000000
1!
1'
1/
#753480000000
0!
1"
0'
1(
0/
10
#753490000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#753500000000
0!
1$
0'
1+
0/
#753510000000
1!
1'
1/
#753520000000
0!
0'
0/
#753530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#753540000000
0!
0'
0/
#753550000000
1!
1'
1/
#753560000000
0!
0'
0/
#753570000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#753580000000
0!
0'
0/
#753590000000
1!
1'
1/
#753600000000
0!
0'
0/
#753610000000
1!
1'
1/
#753620000000
0!
0'
0/
#753630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#753640000000
0!
0'
0/
#753650000000
1!
1'
1/
#753660000000
0!
0'
0/
#753670000000
1!
1'
1/
#753680000000
0!
0'
0/
#753690000000
1!
1'
1/
#753700000000
0!
0'
0/
#753710000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#753720000000
0!
0'
0/
#753730000000
1!
1'
1/
#753740000000
0!
0'
0/
#753750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#753760000000
0!
0'
0/
#753770000000
1!
1'
1/
#753780000000
0!
0'
0/
#753790000000
#753800000000
1!
1'
1/
#753810000000
0!
0'
0/
#753820000000
1!
1'
1/
#753830000000
0!
1"
0'
1(
0/
10
#753840000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#753850000000
0!
0'
0/
#753860000000
1!
1'
1/
#753870000000
0!
0'
0/
#753880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#753890000000
0!
0'
0/
#753900000000
1!
1'
1/
#753910000000
0!
1"
0'
1(
0/
10
#753920000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#753930000000
0!
1$
0'
1+
0/
#753940000000
1!
1'
1/
#753950000000
0!
0'
0/
#753960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#753970000000
0!
0'
0/
#753980000000
1!
1'
1/
#753990000000
0!
0'
0/
#754000000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#754010000000
0!
0'
0/
#754020000000
1!
1'
1/
#754030000000
0!
0'
0/
#754040000000
1!
1'
1/
#754050000000
0!
0'
0/
#754060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#754070000000
0!
0'
0/
#754080000000
1!
1'
1/
#754090000000
0!
0'
0/
#754100000000
1!
1'
1/
#754110000000
0!
0'
0/
#754120000000
1!
1'
1/
#754130000000
0!
0'
0/
#754140000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#754150000000
0!
0'
0/
#754160000000
1!
1'
1/
#754170000000
0!
0'
0/
#754180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#754190000000
0!
0'
0/
#754200000000
1!
1'
1/
#754210000000
0!
0'
0/
#754220000000
#754230000000
1!
1'
1/
#754240000000
0!
0'
0/
#754250000000
1!
1'
1/
#754260000000
0!
1"
0'
1(
0/
10
#754270000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#754280000000
0!
0'
0/
#754290000000
1!
1'
1/
#754300000000
0!
0'
0/
#754310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#754320000000
0!
0'
0/
#754330000000
1!
1'
1/
#754340000000
0!
1"
0'
1(
0/
10
#754350000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#754360000000
0!
1$
0'
1+
0/
#754370000000
1!
1'
1/
#754380000000
0!
0'
0/
#754390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#754400000000
0!
0'
0/
#754410000000
1!
1'
1/
#754420000000
0!
0'
0/
#754430000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#754440000000
0!
0'
0/
#754450000000
1!
1'
1/
#754460000000
0!
0'
0/
#754470000000
1!
1'
1/
#754480000000
0!
0'
0/
#754490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#754500000000
0!
0'
0/
#754510000000
1!
1'
1/
#754520000000
0!
0'
0/
#754530000000
1!
1'
1/
#754540000000
0!
0'
0/
#754550000000
1!
1'
1/
#754560000000
0!
0'
0/
#754570000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#754580000000
0!
0'
0/
#754590000000
1!
1'
1/
#754600000000
0!
0'
0/
#754610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#754620000000
0!
0'
0/
#754630000000
1!
1'
1/
#754640000000
0!
0'
0/
#754650000000
#754660000000
1!
1'
1/
#754670000000
0!
0'
0/
#754680000000
1!
1'
1/
#754690000000
0!
1"
0'
1(
0/
10
#754700000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#754710000000
0!
0'
0/
#754720000000
1!
1'
1/
#754730000000
0!
0'
0/
#754740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#754750000000
0!
0'
0/
#754760000000
1!
1'
1/
#754770000000
0!
1"
0'
1(
0/
10
#754780000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#754790000000
0!
1$
0'
1+
0/
#754800000000
1!
1'
1/
#754810000000
0!
0'
0/
#754820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#754830000000
0!
0'
0/
#754840000000
1!
1'
1/
#754850000000
0!
0'
0/
#754860000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#754870000000
0!
0'
0/
#754880000000
1!
1'
1/
#754890000000
0!
0'
0/
#754900000000
1!
1'
1/
#754910000000
0!
0'
0/
#754920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#754930000000
0!
0'
0/
#754940000000
1!
1'
1/
#754950000000
0!
0'
0/
#754960000000
1!
1'
1/
#754970000000
0!
0'
0/
#754980000000
1!
1'
1/
#754990000000
0!
0'
0/
#755000000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#755010000000
0!
0'
0/
#755020000000
1!
1'
1/
#755030000000
0!
0'
0/
#755040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#755050000000
0!
0'
0/
#755060000000
1!
1'
1/
#755070000000
0!
0'
0/
#755080000000
#755090000000
1!
1'
1/
#755100000000
0!
0'
0/
#755110000000
1!
1'
1/
#755120000000
0!
1"
0'
1(
0/
10
#755130000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#755140000000
0!
0'
0/
#755150000000
1!
1'
1/
#755160000000
0!
0'
0/
#755170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#755180000000
0!
0'
0/
#755190000000
1!
1'
1/
#755200000000
0!
1"
0'
1(
0/
10
#755210000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#755220000000
0!
1$
0'
1+
0/
#755230000000
1!
1'
1/
#755240000000
0!
0'
0/
#755250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#755260000000
0!
0'
0/
#755270000000
1!
1'
1/
#755280000000
0!
0'
0/
#755290000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#755300000000
0!
0'
0/
#755310000000
1!
1'
1/
#755320000000
0!
0'
0/
#755330000000
1!
1'
1/
#755340000000
0!
0'
0/
#755350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#755360000000
0!
0'
0/
#755370000000
1!
1'
1/
#755380000000
0!
0'
0/
#755390000000
1!
1'
1/
#755400000000
0!
0'
0/
#755410000000
1!
1'
1/
#755420000000
0!
0'
0/
#755430000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#755440000000
0!
0'
0/
#755450000000
1!
1'
1/
#755460000000
0!
0'
0/
#755470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#755480000000
0!
0'
0/
#755490000000
1!
1'
1/
#755500000000
0!
0'
0/
#755510000000
#755520000000
1!
1'
1/
#755530000000
0!
0'
0/
#755540000000
1!
1'
1/
#755550000000
0!
1"
0'
1(
0/
10
#755560000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#755570000000
0!
0'
0/
#755580000000
1!
1'
1/
#755590000000
0!
0'
0/
#755600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#755610000000
0!
0'
0/
#755620000000
1!
1'
1/
#755630000000
0!
1"
0'
1(
0/
10
#755640000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#755650000000
0!
1$
0'
1+
0/
#755660000000
1!
1'
1/
#755670000000
0!
0'
0/
#755680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#755690000000
0!
0'
0/
#755700000000
1!
1'
1/
#755710000000
0!
0'
0/
#755720000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#755730000000
0!
0'
0/
#755740000000
1!
1'
1/
#755750000000
0!
0'
0/
#755760000000
1!
1'
1/
#755770000000
0!
0'
0/
#755780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#755790000000
0!
0'
0/
#755800000000
1!
1'
1/
#755810000000
0!
0'
0/
#755820000000
1!
1'
1/
#755830000000
0!
0'
0/
#755840000000
1!
1'
1/
#755850000000
0!
0'
0/
#755860000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#755870000000
0!
0'
0/
#755880000000
1!
1'
1/
#755890000000
0!
0'
0/
#755900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#755910000000
0!
0'
0/
#755920000000
1!
1'
1/
#755930000000
0!
0'
0/
#755940000000
#755950000000
1!
1'
1/
#755960000000
0!
0'
0/
#755970000000
1!
1'
1/
#755980000000
0!
1"
0'
1(
0/
10
#755990000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#756000000000
0!
0'
0/
#756010000000
1!
1'
1/
#756020000000
0!
0'
0/
#756030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#756040000000
0!
0'
0/
#756050000000
1!
1'
1/
#756060000000
0!
1"
0'
1(
0/
10
#756070000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#756080000000
0!
1$
0'
1+
0/
#756090000000
1!
1'
1/
#756100000000
0!
0'
0/
#756110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#756120000000
0!
0'
0/
#756130000000
1!
1'
1/
#756140000000
0!
0'
0/
#756150000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#756160000000
0!
0'
0/
#756170000000
1!
1'
1/
#756180000000
0!
0'
0/
#756190000000
1!
1'
1/
#756200000000
0!
0'
0/
#756210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#756220000000
0!
0'
0/
#756230000000
1!
1'
1/
#756240000000
0!
0'
0/
#756250000000
1!
1'
1/
#756260000000
0!
0'
0/
#756270000000
1!
1'
1/
#756280000000
0!
0'
0/
#756290000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#756300000000
0!
0'
0/
#756310000000
1!
1'
1/
#756320000000
0!
0'
0/
#756330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#756340000000
0!
0'
0/
#756350000000
1!
1'
1/
#756360000000
0!
0'
0/
#756370000000
#756380000000
1!
1'
1/
#756390000000
0!
0'
0/
#756400000000
1!
1'
1/
#756410000000
0!
1"
0'
1(
0/
10
#756420000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#756430000000
0!
0'
0/
#756440000000
1!
1'
1/
#756450000000
0!
0'
0/
#756460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#756470000000
0!
0'
0/
#756480000000
1!
1'
1/
#756490000000
0!
1"
0'
1(
0/
10
#756500000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#756510000000
0!
1$
0'
1+
0/
#756520000000
1!
1'
1/
#756530000000
0!
0'
0/
#756540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#756550000000
0!
0'
0/
#756560000000
1!
1'
1/
#756570000000
0!
0'
0/
#756580000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#756590000000
0!
0'
0/
#756600000000
1!
1'
1/
#756610000000
0!
0'
0/
#756620000000
1!
1'
1/
#756630000000
0!
0'
0/
#756640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#756650000000
0!
0'
0/
#756660000000
1!
1'
1/
#756670000000
0!
0'
0/
#756680000000
1!
1'
1/
#756690000000
0!
0'
0/
#756700000000
1!
1'
1/
#756710000000
0!
0'
0/
#756720000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#756730000000
0!
0'
0/
#756740000000
1!
1'
1/
#756750000000
0!
0'
0/
#756760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#756770000000
0!
0'
0/
#756780000000
1!
1'
1/
#756790000000
0!
0'
0/
#756800000000
#756810000000
1!
1'
1/
#756820000000
0!
0'
0/
#756830000000
1!
1'
1/
#756840000000
0!
1"
0'
1(
0/
10
#756850000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#756860000000
0!
0'
0/
#756870000000
1!
1'
1/
#756880000000
0!
0'
0/
#756890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#756900000000
0!
0'
0/
#756910000000
1!
1'
1/
#756920000000
0!
1"
0'
1(
0/
10
#756930000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#756940000000
0!
1$
0'
1+
0/
#756950000000
1!
1'
1/
#756960000000
0!
0'
0/
#756970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#756980000000
0!
0'
0/
#756990000000
1!
1'
1/
#757000000000
0!
0'
0/
#757010000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#757020000000
0!
0'
0/
#757030000000
1!
1'
1/
#757040000000
0!
0'
0/
#757050000000
1!
1'
1/
#757060000000
0!
0'
0/
#757070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#757080000000
0!
0'
0/
#757090000000
1!
1'
1/
#757100000000
0!
0'
0/
#757110000000
1!
1'
1/
#757120000000
0!
0'
0/
#757130000000
1!
1'
1/
#757140000000
0!
0'
0/
#757150000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#757160000000
0!
0'
0/
#757170000000
1!
1'
1/
#757180000000
0!
0'
0/
#757190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#757200000000
0!
0'
0/
#757210000000
1!
1'
1/
#757220000000
0!
0'
0/
#757230000000
#757240000000
1!
1'
1/
#757250000000
0!
0'
0/
#757260000000
1!
1'
1/
#757270000000
0!
1"
0'
1(
0/
10
#757280000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#757290000000
0!
0'
0/
#757300000000
1!
1'
1/
#757310000000
0!
0'
0/
#757320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#757330000000
0!
0'
0/
#757340000000
1!
1'
1/
#757350000000
0!
1"
0'
1(
0/
10
#757360000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#757370000000
0!
1$
0'
1+
0/
#757380000000
1!
1'
1/
#757390000000
0!
0'
0/
#757400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#757410000000
0!
0'
0/
#757420000000
1!
1'
1/
#757430000000
0!
0'
0/
#757440000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#757450000000
0!
0'
0/
#757460000000
1!
1'
1/
#757470000000
0!
0'
0/
#757480000000
1!
1'
1/
#757490000000
0!
0'
0/
#757500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#757510000000
0!
0'
0/
#757520000000
1!
1'
1/
#757530000000
0!
0'
0/
#757540000000
1!
1'
1/
#757550000000
0!
0'
0/
#757560000000
1!
1'
1/
#757570000000
0!
0'
0/
#757580000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#757590000000
0!
0'
0/
#757600000000
1!
1'
1/
#757610000000
0!
0'
0/
#757620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#757630000000
0!
0'
0/
#757640000000
1!
1'
1/
#757650000000
0!
0'
0/
#757660000000
#757670000000
1!
1'
1/
#757680000000
0!
0'
0/
#757690000000
1!
1'
1/
#757700000000
0!
1"
0'
1(
0/
10
#757710000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#757720000000
0!
0'
0/
#757730000000
1!
1'
1/
#757740000000
0!
0'
0/
#757750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#757760000000
0!
0'
0/
#757770000000
1!
1'
1/
#757780000000
0!
1"
0'
1(
0/
10
#757790000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#757800000000
0!
1$
0'
1+
0/
#757810000000
1!
1'
1/
#757820000000
0!
0'
0/
#757830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#757840000000
0!
0'
0/
#757850000000
1!
1'
1/
#757860000000
0!
0'
0/
#757870000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#757880000000
0!
0'
0/
#757890000000
1!
1'
1/
#757900000000
0!
0'
0/
#757910000000
1!
1'
1/
#757920000000
0!
0'
0/
#757930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#757940000000
0!
0'
0/
#757950000000
1!
1'
1/
#757960000000
0!
0'
0/
#757970000000
1!
1'
1/
#757980000000
0!
0'
0/
#757990000000
1!
1'
1/
#758000000000
0!
0'
0/
#758010000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#758020000000
0!
0'
0/
#758030000000
1!
1'
1/
#758040000000
0!
0'
0/
#758050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#758060000000
0!
0'
0/
#758070000000
1!
1'
1/
#758080000000
0!
0'
0/
#758090000000
#758100000000
1!
1'
1/
#758110000000
0!
0'
0/
#758120000000
1!
1'
1/
#758130000000
0!
1"
0'
1(
0/
10
#758140000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#758150000000
0!
0'
0/
#758160000000
1!
1'
1/
#758170000000
0!
0'
0/
#758180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#758190000000
0!
0'
0/
#758200000000
1!
1'
1/
#758210000000
0!
1"
0'
1(
0/
10
#758220000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#758230000000
0!
1$
0'
1+
0/
#758240000000
1!
1'
1/
#758250000000
0!
0'
0/
#758260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#758270000000
0!
0'
0/
#758280000000
1!
1'
1/
#758290000000
0!
0'
0/
#758300000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#758310000000
0!
0'
0/
#758320000000
1!
1'
1/
#758330000000
0!
0'
0/
#758340000000
1!
1'
1/
#758350000000
0!
0'
0/
#758360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#758370000000
0!
0'
0/
#758380000000
1!
1'
1/
#758390000000
0!
0'
0/
#758400000000
1!
1'
1/
#758410000000
0!
0'
0/
#758420000000
1!
1'
1/
#758430000000
0!
0'
0/
#758440000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#758450000000
0!
0'
0/
#758460000000
1!
1'
1/
#758470000000
0!
0'
0/
#758480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#758490000000
0!
0'
0/
#758500000000
1!
1'
1/
#758510000000
0!
0'
0/
#758520000000
#758530000000
1!
1'
1/
#758540000000
0!
0'
0/
#758550000000
1!
1'
1/
#758560000000
0!
1"
0'
1(
0/
10
#758570000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#758580000000
0!
0'
0/
#758590000000
1!
1'
1/
#758600000000
0!
0'
0/
#758610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#758620000000
0!
0'
0/
#758630000000
1!
1'
1/
#758640000000
0!
1"
0'
1(
0/
10
#758650000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#758660000000
0!
1$
0'
1+
0/
#758670000000
1!
1'
1/
#758680000000
0!
0'
0/
#758690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#758700000000
0!
0'
0/
#758710000000
1!
1'
1/
#758720000000
0!
0'
0/
#758730000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#758740000000
0!
0'
0/
#758750000000
1!
1'
1/
#758760000000
0!
0'
0/
#758770000000
1!
1'
1/
#758780000000
0!
0'
0/
#758790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#758800000000
0!
0'
0/
#758810000000
1!
1'
1/
#758820000000
0!
0'
0/
#758830000000
1!
1'
1/
#758840000000
0!
0'
0/
#758850000000
1!
1'
1/
#758860000000
0!
0'
0/
#758870000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#758880000000
0!
0'
0/
#758890000000
1!
1'
1/
#758900000000
0!
0'
0/
#758910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#758920000000
0!
0'
0/
#758930000000
1!
1'
1/
#758940000000
0!
0'
0/
#758950000000
#758960000000
1!
1'
1/
#758970000000
0!
0'
0/
#758980000000
1!
1'
1/
#758990000000
0!
1"
0'
1(
0/
10
#759000000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#759010000000
0!
0'
0/
#759020000000
1!
1'
1/
#759030000000
0!
0'
0/
#759040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#759050000000
0!
0'
0/
#759060000000
1!
1'
1/
#759070000000
0!
1"
0'
1(
0/
10
#759080000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#759090000000
0!
1$
0'
1+
0/
#759100000000
1!
1'
1/
#759110000000
0!
0'
0/
#759120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#759130000000
0!
0'
0/
#759140000000
1!
1'
1/
#759150000000
0!
0'
0/
#759160000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#759170000000
0!
0'
0/
#759180000000
1!
1'
1/
#759190000000
0!
0'
0/
#759200000000
1!
1'
1/
#759210000000
0!
0'
0/
#759220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#759230000000
0!
0'
0/
#759240000000
1!
1'
1/
#759250000000
0!
0'
0/
#759260000000
1!
1'
1/
#759270000000
0!
0'
0/
#759280000000
1!
1'
1/
#759290000000
0!
0'
0/
#759300000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#759310000000
0!
0'
0/
#759320000000
1!
1'
1/
#759330000000
0!
0'
0/
#759340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#759350000000
0!
0'
0/
#759360000000
1!
1'
1/
#759370000000
0!
0'
0/
#759380000000
#759390000000
1!
1'
1/
#759400000000
0!
0'
0/
#759410000000
1!
1'
1/
#759420000000
0!
1"
0'
1(
0/
10
#759430000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#759440000000
0!
0'
0/
#759450000000
1!
1'
1/
#759460000000
0!
0'
0/
#759470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#759480000000
0!
0'
0/
#759490000000
1!
1'
1/
#759500000000
0!
1"
0'
1(
0/
10
#759510000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#759520000000
0!
1$
0'
1+
0/
#759530000000
1!
1'
1/
#759540000000
0!
0'
0/
#759550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#759560000000
0!
0'
0/
#759570000000
1!
1'
1/
#759580000000
0!
0'
0/
#759590000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#759600000000
0!
0'
0/
#759610000000
1!
1'
1/
#759620000000
0!
0'
0/
#759630000000
1!
1'
1/
#759640000000
0!
0'
0/
#759650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#759660000000
0!
0'
0/
#759670000000
1!
1'
1/
#759680000000
0!
0'
0/
#759690000000
1!
1'
1/
#759700000000
0!
0'
0/
#759710000000
1!
1'
1/
#759720000000
0!
0'
0/
#759730000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#759740000000
0!
0'
0/
#759750000000
1!
1'
1/
#759760000000
0!
0'
0/
#759770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#759780000000
0!
0'
0/
#759790000000
1!
1'
1/
#759800000000
0!
0'
0/
#759810000000
#759820000000
1!
1'
1/
#759830000000
0!
0'
0/
#759840000000
1!
1'
1/
#759850000000
0!
1"
0'
1(
0/
10
#759860000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#759870000000
0!
0'
0/
#759880000000
1!
1'
1/
#759890000000
0!
0'
0/
#759900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#759910000000
0!
0'
0/
#759920000000
1!
1'
1/
#759930000000
0!
1"
0'
1(
0/
10
#759940000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#759950000000
0!
1$
0'
1+
0/
#759960000000
1!
1'
1/
#759970000000
0!
0'
0/
#759980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#759990000000
0!
0'
0/
#760000000000
1!
1'
1/
#760010000000
0!
0'
0/
#760020000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#760030000000
0!
0'
0/
#760040000000
1!
1'
1/
#760050000000
0!
0'
0/
#760060000000
1!
1'
1/
#760070000000
0!
0'
0/
#760080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#760090000000
0!
0'
0/
#760100000000
1!
1'
1/
#760110000000
0!
0'
0/
#760120000000
1!
1'
1/
#760130000000
0!
0'
0/
#760140000000
1!
1'
1/
#760150000000
0!
0'
0/
#760160000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#760170000000
0!
0'
0/
#760180000000
1!
1'
1/
#760190000000
0!
0'
0/
#760200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#760210000000
0!
0'
0/
#760220000000
1!
1'
1/
#760230000000
0!
0'
0/
#760240000000
#760250000000
1!
1'
1/
#760260000000
0!
0'
0/
#760270000000
1!
1'
1/
#760280000000
0!
1"
0'
1(
0/
10
#760290000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#760300000000
0!
0'
0/
#760310000000
1!
1'
1/
#760320000000
0!
0'
0/
#760330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#760340000000
0!
0'
0/
#760350000000
1!
1'
1/
#760360000000
0!
1"
0'
1(
0/
10
#760370000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#760380000000
0!
1$
0'
1+
0/
#760390000000
1!
1'
1/
#760400000000
0!
0'
0/
#760410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#760420000000
0!
0'
0/
#760430000000
1!
1'
1/
#760440000000
0!
0'
0/
#760450000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#760460000000
0!
0'
0/
#760470000000
1!
1'
1/
#760480000000
0!
0'
0/
#760490000000
1!
1'
1/
#760500000000
0!
0'
0/
#760510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#760520000000
0!
0'
0/
#760530000000
1!
1'
1/
#760540000000
0!
0'
0/
#760550000000
1!
1'
1/
#760560000000
0!
0'
0/
#760570000000
1!
1'
1/
#760580000000
0!
0'
0/
#760590000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#760600000000
0!
0'
0/
#760610000000
1!
1'
1/
#760620000000
0!
0'
0/
#760630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#760640000000
0!
0'
0/
#760650000000
1!
1'
1/
#760660000000
0!
0'
0/
#760670000000
#760680000000
1!
1'
1/
#760690000000
0!
0'
0/
#760700000000
1!
1'
1/
#760710000000
0!
1"
0'
1(
0/
10
#760720000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#760730000000
0!
0'
0/
#760740000000
1!
1'
1/
#760750000000
0!
0'
0/
#760760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#760770000000
0!
0'
0/
#760780000000
1!
1'
1/
#760790000000
0!
1"
0'
1(
0/
10
#760800000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#760810000000
0!
1$
0'
1+
0/
#760820000000
1!
1'
1/
#760830000000
0!
0'
0/
#760840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#760850000000
0!
0'
0/
#760860000000
1!
1'
1/
#760870000000
0!
0'
0/
#760880000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#760890000000
0!
0'
0/
#760900000000
1!
1'
1/
#760910000000
0!
0'
0/
#760920000000
1!
1'
1/
#760930000000
0!
0'
0/
#760940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#760950000000
0!
0'
0/
#760960000000
1!
1'
1/
#760970000000
0!
0'
0/
#760980000000
1!
1'
1/
#760990000000
0!
0'
0/
#761000000000
1!
1'
1/
#761010000000
0!
0'
0/
#761020000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#761030000000
0!
0'
0/
#761040000000
1!
1'
1/
#761050000000
0!
0'
0/
#761060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#761070000000
0!
0'
0/
#761080000000
1!
1'
1/
#761090000000
0!
0'
0/
#761100000000
#761110000000
1!
1'
1/
#761120000000
0!
0'
0/
#761130000000
1!
1'
1/
#761140000000
0!
1"
0'
1(
0/
10
#761150000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#761160000000
0!
0'
0/
#761170000000
1!
1'
1/
#761180000000
0!
0'
0/
#761190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#761200000000
0!
0'
0/
#761210000000
1!
1'
1/
#761220000000
0!
1"
0'
1(
0/
10
#761230000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#761240000000
0!
1$
0'
1+
0/
#761250000000
1!
1'
1/
#761260000000
0!
0'
0/
#761270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#761280000000
0!
0'
0/
#761290000000
1!
1'
1/
#761300000000
0!
0'
0/
#761310000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#761320000000
0!
0'
0/
#761330000000
1!
1'
1/
#761340000000
0!
0'
0/
#761350000000
1!
1'
1/
#761360000000
0!
0'
0/
#761370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#761380000000
0!
0'
0/
#761390000000
1!
1'
1/
#761400000000
0!
0'
0/
#761410000000
1!
1'
1/
#761420000000
0!
0'
0/
#761430000000
1!
1'
1/
#761440000000
0!
0'
0/
#761450000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#761460000000
0!
0'
0/
#761470000000
1!
1'
1/
#761480000000
0!
0'
0/
#761490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#761500000000
0!
0'
0/
#761510000000
1!
1'
1/
#761520000000
0!
0'
0/
#761530000000
#761540000000
1!
1'
1/
#761550000000
0!
0'
0/
#761560000000
1!
1'
1/
#761570000000
0!
1"
0'
1(
0/
10
#761580000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#761590000000
0!
0'
0/
#761600000000
1!
1'
1/
#761610000000
0!
0'
0/
#761620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#761630000000
0!
0'
0/
#761640000000
1!
1'
1/
#761650000000
0!
1"
0'
1(
0/
10
#761660000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#761670000000
0!
1$
0'
1+
0/
#761680000000
1!
1'
1/
#761690000000
0!
0'
0/
#761700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#761710000000
0!
0'
0/
#761720000000
1!
1'
1/
#761730000000
0!
0'
0/
#761740000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#761750000000
0!
0'
0/
#761760000000
1!
1'
1/
#761770000000
0!
0'
0/
#761780000000
1!
1'
1/
#761790000000
0!
0'
0/
#761800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#761810000000
0!
0'
0/
#761820000000
1!
1'
1/
#761830000000
0!
0'
0/
#761840000000
1!
1'
1/
#761850000000
0!
0'
0/
#761860000000
1!
1'
1/
#761870000000
0!
0'
0/
#761880000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#761890000000
0!
0'
0/
#761900000000
1!
1'
1/
#761910000000
0!
0'
0/
#761920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#761930000000
0!
0'
0/
#761940000000
1!
1'
1/
#761950000000
0!
0'
0/
#761960000000
#761970000000
1!
1'
1/
#761980000000
0!
0'
0/
#761990000000
1!
1'
1/
#762000000000
0!
1"
0'
1(
0/
10
#762010000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#762020000000
0!
0'
0/
#762030000000
1!
1'
1/
#762040000000
0!
0'
0/
#762050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#762060000000
0!
0'
0/
#762070000000
1!
1'
1/
#762080000000
0!
1"
0'
1(
0/
10
#762090000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#762100000000
0!
1$
0'
1+
0/
#762110000000
1!
1'
1/
#762120000000
0!
0'
0/
#762130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#762140000000
0!
0'
0/
#762150000000
1!
1'
1/
#762160000000
0!
0'
0/
#762170000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#762180000000
0!
0'
0/
#762190000000
1!
1'
1/
#762200000000
0!
0'
0/
#762210000000
1!
1'
1/
#762220000000
0!
0'
0/
#762230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#762240000000
0!
0'
0/
#762250000000
1!
1'
1/
#762260000000
0!
0'
0/
#762270000000
1!
1'
1/
#762280000000
0!
0'
0/
#762290000000
1!
1'
1/
#762300000000
0!
0'
0/
#762310000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#762320000000
0!
0'
0/
#762330000000
1!
1'
1/
#762340000000
0!
0'
0/
#762350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#762360000000
0!
0'
0/
#762370000000
1!
1'
1/
#762380000000
0!
0'
0/
#762390000000
#762400000000
1!
1'
1/
#762410000000
0!
0'
0/
#762420000000
1!
1'
1/
#762430000000
0!
1"
0'
1(
0/
10
#762440000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#762450000000
0!
0'
0/
#762460000000
1!
1'
1/
#762470000000
0!
0'
0/
#762480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#762490000000
0!
0'
0/
#762500000000
1!
1'
1/
#762510000000
0!
1"
0'
1(
0/
10
#762520000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#762530000000
0!
1$
0'
1+
0/
#762540000000
1!
1'
1/
#762550000000
0!
0'
0/
#762560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#762570000000
0!
0'
0/
#762580000000
1!
1'
1/
#762590000000
0!
0'
0/
#762600000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#762610000000
0!
0'
0/
#762620000000
1!
1'
1/
#762630000000
0!
0'
0/
#762640000000
1!
1'
1/
#762650000000
0!
0'
0/
#762660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#762670000000
0!
0'
0/
#762680000000
1!
1'
1/
#762690000000
0!
0'
0/
#762700000000
1!
1'
1/
#762710000000
0!
0'
0/
#762720000000
1!
1'
1/
#762730000000
0!
0'
0/
#762740000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#762750000000
0!
0'
0/
#762760000000
1!
1'
1/
#762770000000
0!
0'
0/
#762780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#762790000000
0!
0'
0/
#762800000000
1!
1'
1/
#762810000000
0!
0'
0/
#762820000000
#762830000000
1!
1'
1/
#762840000000
0!
0'
0/
#762850000000
1!
1'
1/
#762860000000
0!
1"
0'
1(
0/
10
#762870000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#762880000000
0!
0'
0/
#762890000000
1!
1'
1/
#762900000000
0!
0'
0/
#762910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#762920000000
0!
0'
0/
#762930000000
1!
1'
1/
#762940000000
0!
1"
0'
1(
0/
10
#762950000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#762960000000
0!
1$
0'
1+
0/
#762970000000
1!
1'
1/
#762980000000
0!
0'
0/
#762990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#763000000000
0!
0'
0/
#763010000000
1!
1'
1/
#763020000000
0!
0'
0/
#763030000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#763040000000
0!
0'
0/
#763050000000
1!
1'
1/
#763060000000
0!
0'
0/
#763070000000
1!
1'
1/
#763080000000
0!
0'
0/
#763090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#763100000000
0!
0'
0/
#763110000000
1!
1'
1/
#763120000000
0!
0'
0/
#763130000000
1!
1'
1/
#763140000000
0!
0'
0/
#763150000000
1!
1'
1/
#763160000000
0!
0'
0/
#763170000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#763180000000
0!
0'
0/
#763190000000
1!
1'
1/
#763200000000
0!
0'
0/
#763210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#763220000000
0!
0'
0/
#763230000000
1!
1'
1/
#763240000000
0!
0'
0/
#763250000000
#763260000000
1!
1'
1/
#763270000000
0!
0'
0/
#763280000000
1!
1'
1/
#763290000000
0!
1"
0'
1(
0/
10
#763300000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#763310000000
0!
0'
0/
#763320000000
1!
1'
1/
#763330000000
0!
0'
0/
#763340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#763350000000
0!
0'
0/
#763360000000
1!
1'
1/
#763370000000
0!
1"
0'
1(
0/
10
#763380000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#763390000000
0!
1$
0'
1+
0/
#763400000000
1!
1'
1/
#763410000000
0!
0'
0/
#763420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#763430000000
0!
0'
0/
#763440000000
1!
1'
1/
#763450000000
0!
0'
0/
#763460000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#763470000000
0!
0'
0/
#763480000000
1!
1'
1/
#763490000000
0!
0'
0/
#763500000000
1!
1'
1/
#763510000000
0!
0'
0/
#763520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#763530000000
0!
0'
0/
#763540000000
1!
1'
1/
#763550000000
0!
0'
0/
#763560000000
1!
1'
1/
#763570000000
0!
0'
0/
#763580000000
1!
1'
1/
#763590000000
0!
0'
0/
#763600000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#763610000000
0!
0'
0/
#763620000000
1!
1'
1/
#763630000000
0!
0'
0/
#763640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#763650000000
0!
0'
0/
#763660000000
1!
1'
1/
#763670000000
0!
0'
0/
#763680000000
#763690000000
1!
1'
1/
#763700000000
0!
0'
0/
#763710000000
1!
1'
1/
#763720000000
0!
1"
0'
1(
0/
10
#763730000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#763740000000
0!
0'
0/
#763750000000
1!
1'
1/
#763760000000
0!
0'
0/
#763770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#763780000000
0!
0'
0/
#763790000000
1!
1'
1/
#763800000000
0!
1"
0'
1(
0/
10
#763810000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#763820000000
0!
1$
0'
1+
0/
#763830000000
1!
1'
1/
#763840000000
0!
0'
0/
#763850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#763860000000
0!
0'
0/
#763870000000
1!
1'
1/
#763880000000
0!
0'
0/
#763890000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#763900000000
0!
0'
0/
#763910000000
1!
1'
1/
#763920000000
0!
0'
0/
#763930000000
1!
1'
1/
#763940000000
0!
0'
0/
#763950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#763960000000
0!
0'
0/
#763970000000
1!
1'
1/
#763980000000
0!
0'
0/
#763990000000
1!
1'
1/
#764000000000
0!
0'
0/
#764010000000
1!
1'
1/
#764020000000
0!
0'
0/
#764030000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#764040000000
0!
0'
0/
#764050000000
1!
1'
1/
#764060000000
0!
0'
0/
#764070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#764080000000
0!
0'
0/
#764090000000
1!
1'
1/
#764100000000
0!
0'
0/
#764110000000
#764120000000
1!
1'
1/
#764130000000
0!
0'
0/
#764140000000
1!
1'
1/
#764150000000
0!
1"
0'
1(
0/
10
#764160000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#764170000000
0!
0'
0/
#764180000000
1!
1'
1/
#764190000000
0!
0'
0/
#764200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#764210000000
0!
0'
0/
#764220000000
1!
1'
1/
#764230000000
0!
1"
0'
1(
0/
10
#764240000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#764250000000
0!
1$
0'
1+
0/
#764260000000
1!
1'
1/
#764270000000
0!
0'
0/
#764280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#764290000000
0!
0'
0/
#764300000000
1!
1'
1/
#764310000000
0!
0'
0/
#764320000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#764330000000
0!
0'
0/
#764340000000
1!
1'
1/
#764350000000
0!
0'
0/
#764360000000
1!
1'
1/
#764370000000
0!
0'
0/
#764380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#764390000000
0!
0'
0/
#764400000000
1!
1'
1/
#764410000000
0!
0'
0/
#764420000000
1!
1'
1/
#764430000000
0!
0'
0/
#764440000000
1!
1'
1/
#764450000000
0!
0'
0/
#764460000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#764470000000
0!
0'
0/
#764480000000
1!
1'
1/
#764490000000
0!
0'
0/
#764500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#764510000000
0!
0'
0/
#764520000000
1!
1'
1/
#764530000000
0!
0'
0/
#764540000000
#764550000000
1!
1'
1/
#764560000000
0!
0'
0/
#764570000000
1!
1'
1/
#764580000000
0!
1"
0'
1(
0/
10
#764590000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#764600000000
0!
0'
0/
#764610000000
1!
1'
1/
#764620000000
0!
0'
0/
#764630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#764640000000
0!
0'
0/
#764650000000
1!
1'
1/
#764660000000
0!
1"
0'
1(
0/
10
#764670000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#764680000000
0!
1$
0'
1+
0/
#764690000000
1!
1'
1/
#764700000000
0!
0'
0/
#764710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#764720000000
0!
0'
0/
#764730000000
1!
1'
1/
#764740000000
0!
0'
0/
#764750000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#764760000000
0!
0'
0/
#764770000000
1!
1'
1/
#764780000000
0!
0'
0/
#764790000000
1!
1'
1/
#764800000000
0!
0'
0/
#764810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#764820000000
0!
0'
0/
#764830000000
1!
1'
1/
#764840000000
0!
0'
0/
#764850000000
1!
1'
1/
#764860000000
0!
0'
0/
#764870000000
1!
1'
1/
#764880000000
0!
0'
0/
#764890000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#764900000000
0!
0'
0/
#764910000000
1!
1'
1/
#764920000000
0!
0'
0/
#764930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#764940000000
0!
0'
0/
#764950000000
1!
1'
1/
#764960000000
0!
0'
0/
#764970000000
#764980000000
1!
1'
1/
#764990000000
0!
0'
0/
#765000000000
1!
1'
1/
#765010000000
0!
1"
0'
1(
0/
10
#765020000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#765030000000
0!
0'
0/
#765040000000
1!
1'
1/
#765050000000
0!
0'
0/
#765060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#765070000000
0!
0'
0/
#765080000000
1!
1'
1/
#765090000000
0!
1"
0'
1(
0/
10
#765100000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#765110000000
0!
1$
0'
1+
0/
#765120000000
1!
1'
1/
#765130000000
0!
0'
0/
#765140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#765150000000
0!
0'
0/
#765160000000
1!
1'
1/
#765170000000
0!
0'
0/
#765180000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#765190000000
0!
0'
0/
#765200000000
1!
1'
1/
#765210000000
0!
0'
0/
#765220000000
1!
1'
1/
#765230000000
0!
0'
0/
#765240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#765250000000
0!
0'
0/
#765260000000
1!
1'
1/
#765270000000
0!
0'
0/
#765280000000
1!
1'
1/
#765290000000
0!
0'
0/
#765300000000
1!
1'
1/
#765310000000
0!
0'
0/
#765320000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#765330000000
0!
0'
0/
#765340000000
1!
1'
1/
#765350000000
0!
0'
0/
#765360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#765370000000
0!
0'
0/
#765380000000
1!
1'
1/
#765390000000
0!
0'
0/
#765400000000
#765410000000
1!
1'
1/
#765420000000
0!
0'
0/
#765430000000
1!
1'
1/
#765440000000
0!
1"
0'
1(
0/
10
#765450000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#765460000000
0!
0'
0/
#765470000000
1!
1'
1/
#765480000000
0!
0'
0/
#765490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#765500000000
0!
0'
0/
#765510000000
1!
1'
1/
#765520000000
0!
1"
0'
1(
0/
10
#765530000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#765540000000
0!
1$
0'
1+
0/
#765550000000
1!
1'
1/
#765560000000
0!
0'
0/
#765570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#765580000000
0!
0'
0/
#765590000000
1!
1'
1/
#765600000000
0!
0'
0/
#765610000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#765620000000
0!
0'
0/
#765630000000
1!
1'
1/
#765640000000
0!
0'
0/
#765650000000
1!
1'
1/
#765660000000
0!
0'
0/
#765670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#765680000000
0!
0'
0/
#765690000000
1!
1'
1/
#765700000000
0!
0'
0/
#765710000000
1!
1'
1/
#765720000000
0!
0'
0/
#765730000000
1!
1'
1/
#765740000000
0!
0'
0/
#765750000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#765760000000
0!
0'
0/
#765770000000
1!
1'
1/
#765780000000
0!
0'
0/
#765790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#765800000000
0!
0'
0/
#765810000000
1!
1'
1/
#765820000000
0!
0'
0/
#765830000000
#765840000000
1!
1'
1/
#765850000000
0!
0'
0/
#765860000000
1!
1'
1/
#765870000000
0!
1"
0'
1(
0/
10
#765880000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#765890000000
0!
0'
0/
#765900000000
1!
1'
1/
#765910000000
0!
0'
0/
#765920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#765930000000
0!
0'
0/
#765940000000
1!
1'
1/
#765950000000
0!
1"
0'
1(
0/
10
#765960000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#765970000000
0!
1$
0'
1+
0/
#765980000000
1!
1'
1/
#765990000000
0!
0'
0/
#766000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#766010000000
0!
0'
0/
#766020000000
1!
1'
1/
#766030000000
0!
0'
0/
#766040000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#766050000000
0!
0'
0/
#766060000000
1!
1'
1/
#766070000000
0!
0'
0/
#766080000000
1!
1'
1/
#766090000000
0!
0'
0/
#766100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#766110000000
0!
0'
0/
#766120000000
1!
1'
1/
#766130000000
0!
0'
0/
#766140000000
1!
1'
1/
#766150000000
0!
0'
0/
#766160000000
1!
1'
1/
#766170000000
0!
0'
0/
#766180000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#766190000000
0!
0'
0/
#766200000000
1!
1'
1/
#766210000000
0!
0'
0/
#766220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#766230000000
0!
0'
0/
#766240000000
1!
1'
1/
#766250000000
0!
0'
0/
#766260000000
#766270000000
1!
1'
1/
#766280000000
0!
0'
0/
#766290000000
1!
1'
1/
#766300000000
0!
1"
0'
1(
0/
10
#766310000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#766320000000
0!
0'
0/
#766330000000
1!
1'
1/
#766340000000
0!
0'
0/
#766350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#766360000000
0!
0'
0/
#766370000000
1!
1'
1/
#766380000000
0!
1"
0'
1(
0/
10
#766390000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#766400000000
0!
1$
0'
1+
0/
#766410000000
1!
1'
1/
#766420000000
0!
0'
0/
#766430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#766440000000
0!
0'
0/
#766450000000
1!
1'
1/
#766460000000
0!
0'
0/
#766470000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#766480000000
0!
0'
0/
#766490000000
1!
1'
1/
#766500000000
0!
0'
0/
#766510000000
1!
1'
1/
#766520000000
0!
0'
0/
#766530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#766540000000
0!
0'
0/
#766550000000
1!
1'
1/
#766560000000
0!
0'
0/
#766570000000
1!
1'
1/
#766580000000
0!
0'
0/
#766590000000
1!
1'
1/
#766600000000
0!
0'
0/
#766610000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#766620000000
0!
0'
0/
#766630000000
1!
1'
1/
#766640000000
0!
0'
0/
#766650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#766660000000
0!
0'
0/
#766670000000
1!
1'
1/
#766680000000
0!
0'
0/
#766690000000
#766700000000
1!
1'
1/
#766710000000
0!
0'
0/
#766720000000
1!
1'
1/
#766730000000
0!
1"
0'
1(
0/
10
#766740000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#766750000000
0!
0'
0/
#766760000000
1!
1'
1/
#766770000000
0!
0'
0/
#766780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#766790000000
0!
0'
0/
#766800000000
1!
1'
1/
#766810000000
0!
1"
0'
1(
0/
10
#766820000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#766830000000
0!
1$
0'
1+
0/
#766840000000
1!
1'
1/
#766850000000
0!
0'
0/
#766860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#766870000000
0!
0'
0/
#766880000000
1!
1'
1/
#766890000000
0!
0'
0/
#766900000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#766910000000
0!
0'
0/
#766920000000
1!
1'
1/
#766930000000
0!
0'
0/
#766940000000
1!
1'
1/
#766950000000
0!
0'
0/
#766960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#766970000000
0!
0'
0/
#766980000000
1!
1'
1/
#766990000000
0!
0'
0/
#767000000000
1!
1'
1/
#767010000000
0!
0'
0/
#767020000000
1!
1'
1/
#767030000000
0!
0'
0/
#767040000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#767050000000
0!
0'
0/
#767060000000
1!
1'
1/
#767070000000
0!
0'
0/
#767080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#767090000000
0!
0'
0/
#767100000000
1!
1'
1/
#767110000000
0!
0'
0/
#767120000000
#767130000000
1!
1'
1/
#767140000000
0!
0'
0/
#767150000000
1!
1'
1/
#767160000000
0!
1"
0'
1(
0/
10
#767170000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#767180000000
0!
0'
0/
#767190000000
1!
1'
1/
#767200000000
0!
0'
0/
#767210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#767220000000
0!
0'
0/
#767230000000
1!
1'
1/
#767240000000
0!
1"
0'
1(
0/
10
#767250000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#767260000000
0!
1$
0'
1+
0/
#767270000000
1!
1'
1/
#767280000000
0!
0'
0/
#767290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#767300000000
0!
0'
0/
#767310000000
1!
1'
1/
#767320000000
0!
0'
0/
#767330000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#767340000000
0!
0'
0/
#767350000000
1!
1'
1/
#767360000000
0!
0'
0/
#767370000000
1!
1'
1/
#767380000000
0!
0'
0/
#767390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#767400000000
0!
0'
0/
#767410000000
1!
1'
1/
#767420000000
0!
0'
0/
#767430000000
1!
1'
1/
#767440000000
0!
0'
0/
#767450000000
1!
1'
1/
#767460000000
0!
0'
0/
#767470000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#767480000000
0!
0'
0/
#767490000000
1!
1'
1/
#767500000000
0!
0'
0/
#767510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#767520000000
0!
0'
0/
#767530000000
1!
1'
1/
#767540000000
0!
0'
0/
#767550000000
#767560000000
1!
1'
1/
#767570000000
0!
0'
0/
#767580000000
1!
1'
1/
#767590000000
0!
1"
0'
1(
0/
10
#767600000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#767610000000
0!
0'
0/
#767620000000
1!
1'
1/
#767630000000
0!
0'
0/
#767640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#767650000000
0!
0'
0/
#767660000000
1!
1'
1/
#767670000000
0!
1"
0'
1(
0/
10
#767680000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#767690000000
0!
1$
0'
1+
0/
#767700000000
1!
1'
1/
#767710000000
0!
0'
0/
#767720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#767730000000
0!
0'
0/
#767740000000
1!
1'
1/
#767750000000
0!
0'
0/
#767760000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#767770000000
0!
0'
0/
#767780000000
1!
1'
1/
#767790000000
0!
0'
0/
#767800000000
1!
1'
1/
#767810000000
0!
0'
0/
#767820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#767830000000
0!
0'
0/
#767840000000
1!
1'
1/
#767850000000
0!
0'
0/
#767860000000
1!
1'
1/
#767870000000
0!
0'
0/
#767880000000
1!
1'
1/
#767890000000
0!
0'
0/
#767900000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#767910000000
0!
0'
0/
#767920000000
1!
1'
1/
#767930000000
0!
0'
0/
#767940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#767950000000
0!
0'
0/
#767960000000
1!
1'
1/
#767970000000
0!
0'
0/
#767980000000
#767990000000
1!
1'
1/
#768000000000
0!
0'
0/
#768010000000
1!
1'
1/
#768020000000
0!
1"
0'
1(
0/
10
#768030000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#768040000000
0!
0'
0/
#768050000000
1!
1'
1/
#768060000000
0!
0'
0/
#768070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#768080000000
0!
0'
0/
#768090000000
1!
1'
1/
#768100000000
0!
1"
0'
1(
0/
10
#768110000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#768120000000
0!
1$
0'
1+
0/
#768130000000
1!
1'
1/
#768140000000
0!
0'
0/
#768150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#768160000000
0!
0'
0/
#768170000000
1!
1'
1/
#768180000000
0!
0'
0/
#768190000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#768200000000
0!
0'
0/
#768210000000
1!
1'
1/
#768220000000
0!
0'
0/
#768230000000
1!
1'
1/
#768240000000
0!
0'
0/
#768250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#768260000000
0!
0'
0/
#768270000000
1!
1'
1/
#768280000000
0!
0'
0/
#768290000000
1!
1'
1/
#768300000000
0!
0'
0/
#768310000000
1!
1'
1/
#768320000000
0!
0'
0/
#768330000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#768340000000
0!
0'
0/
#768350000000
1!
1'
1/
#768360000000
0!
0'
0/
#768370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#768380000000
0!
0'
0/
#768390000000
1!
1'
1/
#768400000000
0!
0'
0/
#768410000000
#768420000000
1!
1'
1/
#768430000000
0!
0'
0/
#768440000000
1!
1'
1/
#768450000000
0!
1"
0'
1(
0/
10
#768460000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#768470000000
0!
0'
0/
#768480000000
1!
1'
1/
#768490000000
0!
0'
0/
#768500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#768510000000
0!
0'
0/
#768520000000
1!
1'
1/
#768530000000
0!
1"
0'
1(
0/
10
#768540000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#768550000000
0!
1$
0'
1+
0/
#768560000000
1!
1'
1/
#768570000000
0!
0'
0/
#768580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#768590000000
0!
0'
0/
#768600000000
1!
1'
1/
#768610000000
0!
0'
0/
#768620000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#768630000000
0!
0'
0/
#768640000000
1!
1'
1/
#768650000000
0!
0'
0/
#768660000000
1!
1'
1/
#768670000000
0!
0'
0/
#768680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#768690000000
0!
0'
0/
#768700000000
1!
1'
1/
#768710000000
0!
0'
0/
#768720000000
1!
1'
1/
#768730000000
0!
0'
0/
#768740000000
1!
1'
1/
#768750000000
0!
0'
0/
#768760000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#768770000000
0!
0'
0/
#768780000000
1!
1'
1/
#768790000000
0!
0'
0/
#768800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#768810000000
0!
0'
0/
#768820000000
1!
1'
1/
#768830000000
0!
0'
0/
#768840000000
#768850000000
1!
1'
1/
#768860000000
0!
0'
0/
#768870000000
1!
1'
1/
#768880000000
0!
1"
0'
1(
0/
10
#768890000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#768900000000
0!
0'
0/
#768910000000
1!
1'
1/
#768920000000
0!
0'
0/
#768930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#768940000000
0!
0'
0/
#768950000000
1!
1'
1/
#768960000000
0!
1"
0'
1(
0/
10
#768970000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#768980000000
0!
1$
0'
1+
0/
#768990000000
1!
1'
1/
#769000000000
0!
0'
0/
#769010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#769020000000
0!
0'
0/
#769030000000
1!
1'
1/
#769040000000
0!
0'
0/
#769050000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#769060000000
0!
0'
0/
#769070000000
1!
1'
1/
#769080000000
0!
0'
0/
#769090000000
1!
1'
1/
#769100000000
0!
0'
0/
#769110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#769120000000
0!
0'
0/
#769130000000
1!
1'
1/
#769140000000
0!
0'
0/
#769150000000
1!
1'
1/
#769160000000
0!
0'
0/
#769170000000
1!
1'
1/
#769180000000
0!
0'
0/
#769190000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#769200000000
0!
0'
0/
#769210000000
1!
1'
1/
#769220000000
0!
0'
0/
#769230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#769240000000
0!
0'
0/
#769250000000
1!
1'
1/
#769260000000
0!
0'
0/
#769270000000
#769280000000
1!
1'
1/
#769290000000
0!
0'
0/
#769300000000
1!
1'
1/
#769310000000
0!
1"
0'
1(
0/
10
#769320000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#769330000000
0!
0'
0/
#769340000000
1!
1'
1/
#769350000000
0!
0'
0/
#769360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#769370000000
0!
0'
0/
#769380000000
1!
1'
1/
#769390000000
0!
1"
0'
1(
0/
10
#769400000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#769410000000
0!
1$
0'
1+
0/
#769420000000
1!
1'
1/
#769430000000
0!
0'
0/
#769440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#769450000000
0!
0'
0/
#769460000000
1!
1'
1/
#769470000000
0!
0'
0/
#769480000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#769490000000
0!
0'
0/
#769500000000
1!
1'
1/
#769510000000
0!
0'
0/
#769520000000
1!
1'
1/
#769530000000
0!
0'
0/
#769540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#769550000000
0!
0'
0/
#769560000000
1!
1'
1/
#769570000000
0!
0'
0/
#769580000000
1!
1'
1/
#769590000000
0!
0'
0/
#769600000000
1!
1'
1/
#769610000000
0!
0'
0/
#769620000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#769630000000
0!
0'
0/
#769640000000
1!
1'
1/
#769650000000
0!
0'
0/
#769660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#769670000000
0!
0'
0/
#769680000000
1!
1'
1/
#769690000000
0!
0'
0/
#769700000000
#769710000000
1!
1'
1/
#769720000000
0!
0'
0/
#769730000000
1!
1'
1/
#769740000000
0!
1"
0'
1(
0/
10
#769750000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#769760000000
0!
0'
0/
#769770000000
1!
1'
1/
#769780000000
0!
0'
0/
#769790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#769800000000
0!
0'
0/
#769810000000
1!
1'
1/
#769820000000
0!
1"
0'
1(
0/
10
#769830000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#769840000000
0!
1$
0'
1+
0/
#769850000000
1!
1'
1/
#769860000000
0!
0'
0/
#769870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#769880000000
0!
0'
0/
#769890000000
1!
1'
1/
#769900000000
0!
0'
0/
#769910000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#769920000000
0!
0'
0/
#769930000000
1!
1'
1/
#769940000000
0!
0'
0/
#769950000000
1!
1'
1/
#769960000000
0!
0'
0/
#769970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#769980000000
0!
0'
0/
#769990000000
1!
1'
1/
#770000000000
0!
0'
0/
#770010000000
1!
1'
1/
#770020000000
0!
0'
0/
#770030000000
1!
1'
1/
#770040000000
0!
0'
0/
#770050000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#770060000000
0!
0'
0/
#770070000000
1!
1'
1/
#770080000000
0!
0'
0/
#770090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#770100000000
0!
0'
0/
#770110000000
1!
1'
1/
#770120000000
0!
0'
0/
#770130000000
#770140000000
1!
1'
1/
#770150000000
0!
0'
0/
#770160000000
1!
1'
1/
#770170000000
0!
1"
0'
1(
0/
10
#770180000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#770190000000
0!
0'
0/
#770200000000
1!
1'
1/
#770210000000
0!
0'
0/
#770220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#770230000000
0!
0'
0/
#770240000000
1!
1'
1/
#770250000000
0!
1"
0'
1(
0/
10
#770260000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#770270000000
0!
1$
0'
1+
0/
#770280000000
1!
1'
1/
#770290000000
0!
0'
0/
#770300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#770310000000
0!
0'
0/
#770320000000
1!
1'
1/
#770330000000
0!
0'
0/
#770340000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#770350000000
0!
0'
0/
#770360000000
1!
1'
1/
#770370000000
0!
0'
0/
#770380000000
1!
1'
1/
#770390000000
0!
0'
0/
#770400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#770410000000
0!
0'
0/
#770420000000
1!
1'
1/
#770430000000
0!
0'
0/
#770440000000
1!
1'
1/
#770450000000
0!
0'
0/
#770460000000
1!
1'
1/
#770470000000
0!
0'
0/
#770480000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#770490000000
0!
0'
0/
#770500000000
1!
1'
1/
#770510000000
0!
0'
0/
#770520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#770530000000
0!
0'
0/
#770540000000
1!
1'
1/
#770550000000
0!
0'
0/
#770560000000
#770570000000
1!
1'
1/
#770580000000
0!
0'
0/
#770590000000
1!
1'
1/
#770600000000
0!
1"
0'
1(
0/
10
#770610000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#770620000000
0!
0'
0/
#770630000000
1!
1'
1/
#770640000000
0!
0'
0/
#770650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#770660000000
0!
0'
0/
#770670000000
1!
1'
1/
#770680000000
0!
1"
0'
1(
0/
10
#770690000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#770700000000
0!
1$
0'
1+
0/
#770710000000
1!
1'
1/
#770720000000
0!
0'
0/
#770730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#770740000000
0!
0'
0/
#770750000000
1!
1'
1/
#770760000000
0!
0'
0/
#770770000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#770780000000
0!
0'
0/
#770790000000
1!
1'
1/
#770800000000
0!
0'
0/
#770810000000
1!
1'
1/
#770820000000
0!
0'
0/
#770830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#770840000000
0!
0'
0/
#770850000000
1!
1'
1/
#770860000000
0!
0'
0/
#770870000000
1!
1'
1/
#770880000000
0!
0'
0/
#770890000000
1!
1'
1/
#770900000000
0!
0'
0/
#770910000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#770920000000
0!
0'
0/
#770930000000
1!
1'
1/
#770940000000
0!
0'
0/
#770950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#770960000000
0!
0'
0/
#770970000000
1!
1'
1/
#770980000000
0!
0'
0/
#770990000000
#771000000000
1!
1'
1/
#771010000000
0!
0'
0/
#771020000000
1!
1'
1/
#771030000000
0!
1"
0'
1(
0/
10
#771040000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#771050000000
0!
0'
0/
#771060000000
1!
1'
1/
#771070000000
0!
0'
0/
#771080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#771090000000
0!
0'
0/
#771100000000
1!
1'
1/
#771110000000
0!
1"
0'
1(
0/
10
#771120000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#771130000000
0!
1$
0'
1+
0/
#771140000000
1!
1'
1/
#771150000000
0!
0'
0/
#771160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#771170000000
0!
0'
0/
#771180000000
1!
1'
1/
#771190000000
0!
0'
0/
#771200000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#771210000000
0!
0'
0/
#771220000000
1!
1'
1/
#771230000000
0!
0'
0/
#771240000000
1!
1'
1/
#771250000000
0!
0'
0/
#771260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#771270000000
0!
0'
0/
#771280000000
1!
1'
1/
#771290000000
0!
0'
0/
#771300000000
1!
1'
1/
#771310000000
0!
0'
0/
#771320000000
1!
1'
1/
#771330000000
0!
0'
0/
#771340000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#771350000000
0!
0'
0/
#771360000000
1!
1'
1/
#771370000000
0!
0'
0/
#771380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#771390000000
0!
0'
0/
#771400000000
1!
1'
1/
#771410000000
0!
0'
0/
#771420000000
#771430000000
1!
1'
1/
#771440000000
0!
0'
0/
#771450000000
1!
1'
1/
#771460000000
0!
1"
0'
1(
0/
10
#771470000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#771480000000
0!
0'
0/
#771490000000
1!
1'
1/
#771500000000
0!
0'
0/
#771510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#771520000000
0!
0'
0/
#771530000000
1!
1'
1/
#771540000000
0!
1"
0'
1(
0/
10
#771550000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#771560000000
0!
1$
0'
1+
0/
#771570000000
1!
1'
1/
#771580000000
0!
0'
0/
#771590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#771600000000
0!
0'
0/
#771610000000
1!
1'
1/
#771620000000
0!
0'
0/
#771630000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#771640000000
0!
0'
0/
#771650000000
1!
1'
1/
#771660000000
0!
0'
0/
#771670000000
1!
1'
1/
#771680000000
0!
0'
0/
#771690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#771700000000
0!
0'
0/
#771710000000
1!
1'
1/
#771720000000
0!
0'
0/
#771730000000
1!
1'
1/
#771740000000
0!
0'
0/
#771750000000
1!
1'
1/
#771760000000
0!
0'
0/
#771770000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#771780000000
0!
0'
0/
#771790000000
1!
1'
1/
#771800000000
0!
0'
0/
#771810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#771820000000
0!
0'
0/
#771830000000
1!
1'
1/
#771840000000
0!
0'
0/
#771850000000
#771860000000
1!
1'
1/
#771870000000
0!
0'
0/
#771880000000
1!
1'
1/
#771890000000
0!
1"
0'
1(
0/
10
#771900000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#771910000000
0!
0'
0/
#771920000000
1!
1'
1/
#771930000000
0!
0'
0/
#771940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#771950000000
0!
0'
0/
#771960000000
1!
1'
1/
#771970000000
0!
1"
0'
1(
0/
10
#771980000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#771990000000
0!
1$
0'
1+
0/
#772000000000
1!
1'
1/
#772010000000
0!
0'
0/
#772020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#772030000000
0!
0'
0/
#772040000000
1!
1'
1/
#772050000000
0!
0'
0/
#772060000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#772070000000
0!
0'
0/
#772080000000
1!
1'
1/
#772090000000
0!
0'
0/
#772100000000
1!
1'
1/
#772110000000
0!
0'
0/
#772120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#772130000000
0!
0'
0/
#772140000000
1!
1'
1/
#772150000000
0!
0'
0/
#772160000000
1!
1'
1/
#772170000000
0!
0'
0/
#772180000000
1!
1'
1/
#772190000000
0!
0'
0/
#772200000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#772210000000
0!
0'
0/
#772220000000
1!
1'
1/
#772230000000
0!
0'
0/
#772240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#772250000000
0!
0'
0/
#772260000000
1!
1'
1/
#772270000000
0!
0'
0/
#772280000000
#772290000000
1!
1'
1/
#772300000000
0!
0'
0/
#772310000000
1!
1'
1/
#772320000000
0!
1"
0'
1(
0/
10
#772330000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#772340000000
0!
0'
0/
#772350000000
1!
1'
1/
#772360000000
0!
0'
0/
#772370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#772380000000
0!
0'
0/
#772390000000
1!
1'
1/
#772400000000
0!
1"
0'
1(
0/
10
#772410000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#772420000000
0!
1$
0'
1+
0/
#772430000000
1!
1'
1/
#772440000000
0!
0'
0/
#772450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#772460000000
0!
0'
0/
#772470000000
1!
1'
1/
#772480000000
0!
0'
0/
#772490000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#772500000000
0!
0'
0/
#772510000000
1!
1'
1/
#772520000000
0!
0'
0/
#772530000000
1!
1'
1/
#772540000000
0!
0'
0/
#772550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#772560000000
0!
0'
0/
#772570000000
1!
1'
1/
#772580000000
0!
0'
0/
#772590000000
1!
1'
1/
#772600000000
0!
0'
0/
#772610000000
1!
1'
1/
#772620000000
0!
0'
0/
#772630000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#772640000000
0!
0'
0/
#772650000000
1!
1'
1/
#772660000000
0!
0'
0/
#772670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#772680000000
0!
0'
0/
#772690000000
1!
1'
1/
#772700000000
0!
0'
0/
#772710000000
#772720000000
1!
1'
1/
#772730000000
0!
0'
0/
#772740000000
1!
1'
1/
#772750000000
0!
1"
0'
1(
0/
10
#772760000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#772770000000
0!
0'
0/
#772780000000
1!
1'
1/
#772790000000
0!
0'
0/
#772800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#772810000000
0!
0'
0/
#772820000000
1!
1'
1/
#772830000000
0!
1"
0'
1(
0/
10
#772840000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#772850000000
0!
1$
0'
1+
0/
#772860000000
1!
1'
1/
#772870000000
0!
0'
0/
#772880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#772890000000
0!
0'
0/
#772900000000
1!
1'
1/
#772910000000
0!
0'
0/
#772920000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#772930000000
0!
0'
0/
#772940000000
1!
1'
1/
#772950000000
0!
0'
0/
#772960000000
1!
1'
1/
#772970000000
0!
0'
0/
#772980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#772990000000
0!
0'
0/
#773000000000
1!
1'
1/
#773010000000
0!
0'
0/
#773020000000
1!
1'
1/
#773030000000
0!
0'
0/
#773040000000
1!
1'
1/
#773050000000
0!
0'
0/
#773060000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#773070000000
0!
0'
0/
#773080000000
1!
1'
1/
#773090000000
0!
0'
0/
#773100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#773110000000
0!
0'
0/
#773120000000
1!
1'
1/
#773130000000
0!
0'
0/
#773140000000
#773150000000
1!
1'
1/
#773160000000
0!
0'
0/
#773170000000
1!
1'
1/
#773180000000
0!
1"
0'
1(
0/
10
#773190000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#773200000000
0!
0'
0/
#773210000000
1!
1'
1/
#773220000000
0!
0'
0/
#773230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#773240000000
0!
0'
0/
#773250000000
1!
1'
1/
#773260000000
0!
1"
0'
1(
0/
10
#773270000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#773280000000
0!
1$
0'
1+
0/
#773290000000
1!
1'
1/
#773300000000
0!
0'
0/
#773310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#773320000000
0!
0'
0/
#773330000000
1!
1'
1/
#773340000000
0!
0'
0/
#773350000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#773360000000
0!
0'
0/
#773370000000
1!
1'
1/
#773380000000
0!
0'
0/
#773390000000
1!
1'
1/
#773400000000
0!
0'
0/
#773410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#773420000000
0!
0'
0/
#773430000000
1!
1'
1/
#773440000000
0!
0'
0/
#773450000000
1!
1'
1/
#773460000000
0!
0'
0/
#773470000000
1!
1'
1/
#773480000000
0!
0'
0/
#773490000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#773500000000
0!
0'
0/
#773510000000
1!
1'
1/
#773520000000
0!
0'
0/
#773530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#773540000000
0!
0'
0/
#773550000000
1!
1'
1/
#773560000000
0!
0'
0/
#773570000000
#773580000000
1!
1'
1/
#773590000000
0!
0'
0/
#773600000000
1!
1'
1/
#773610000000
0!
1"
0'
1(
0/
10
#773620000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#773630000000
0!
0'
0/
#773640000000
1!
1'
1/
#773650000000
0!
0'
0/
#773660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#773670000000
0!
0'
0/
#773680000000
1!
1'
1/
#773690000000
0!
1"
0'
1(
0/
10
#773700000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#773710000000
0!
1$
0'
1+
0/
#773720000000
1!
1'
1/
#773730000000
0!
0'
0/
#773740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#773750000000
0!
0'
0/
#773760000000
1!
1'
1/
#773770000000
0!
0'
0/
#773780000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#773790000000
0!
0'
0/
#773800000000
1!
1'
1/
#773810000000
0!
0'
0/
#773820000000
1!
1'
1/
#773830000000
0!
0'
0/
#773840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#773850000000
0!
0'
0/
#773860000000
1!
1'
1/
#773870000000
0!
0'
0/
#773880000000
1!
1'
1/
#773890000000
0!
0'
0/
#773900000000
1!
1'
1/
#773910000000
0!
0'
0/
#773920000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#773930000000
0!
0'
0/
#773940000000
1!
1'
1/
#773950000000
0!
0'
0/
#773960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#773970000000
0!
0'
0/
#773980000000
1!
1'
1/
#773990000000
0!
0'
0/
#774000000000
#774010000000
1!
1'
1/
#774020000000
0!
0'
0/
#774030000000
1!
1'
1/
#774040000000
0!
1"
0'
1(
0/
10
#774050000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#774060000000
0!
0'
0/
#774070000000
1!
1'
1/
#774080000000
0!
0'
0/
#774090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#774100000000
0!
0'
0/
#774110000000
1!
1'
1/
#774120000000
0!
1"
0'
1(
0/
10
#774130000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#774140000000
0!
1$
0'
1+
0/
#774150000000
1!
1'
1/
#774160000000
0!
0'
0/
#774170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#774180000000
0!
0'
0/
#774190000000
1!
1'
1/
#774200000000
0!
0'
0/
#774210000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#774220000000
0!
0'
0/
#774230000000
1!
1'
1/
#774240000000
0!
0'
0/
#774250000000
1!
1'
1/
#774260000000
0!
0'
0/
#774270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#774280000000
0!
0'
0/
#774290000000
1!
1'
1/
#774300000000
0!
0'
0/
#774310000000
1!
1'
1/
#774320000000
0!
0'
0/
#774330000000
1!
1'
1/
#774340000000
0!
0'
0/
#774350000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#774360000000
0!
0'
0/
#774370000000
1!
1'
1/
#774380000000
0!
0'
0/
#774390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#774400000000
0!
0'
0/
#774410000000
1!
1'
1/
#774420000000
0!
0'
0/
#774430000000
#774440000000
1!
1'
1/
#774450000000
0!
0'
0/
#774460000000
1!
1'
1/
#774470000000
0!
1"
0'
1(
0/
10
#774480000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#774490000000
0!
0'
0/
#774500000000
1!
1'
1/
#774510000000
0!
0'
0/
#774520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#774530000000
0!
0'
0/
#774540000000
1!
1'
1/
#774550000000
0!
1"
0'
1(
0/
10
#774560000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#774570000000
0!
1$
0'
1+
0/
#774580000000
1!
1'
1/
#774590000000
0!
0'
0/
#774600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#774610000000
0!
0'
0/
#774620000000
1!
1'
1/
#774630000000
0!
0'
0/
#774640000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#774650000000
0!
0'
0/
#774660000000
1!
1'
1/
#774670000000
0!
0'
0/
#774680000000
1!
1'
1/
#774690000000
0!
0'
0/
#774700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#774710000000
0!
0'
0/
#774720000000
1!
1'
1/
#774730000000
0!
0'
0/
#774740000000
1!
1'
1/
#774750000000
0!
0'
0/
#774760000000
1!
1'
1/
#774770000000
0!
0'
0/
#774780000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#774790000000
0!
0'
0/
#774800000000
1!
1'
1/
#774810000000
0!
0'
0/
#774820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#774830000000
0!
0'
0/
#774840000000
1!
1'
1/
#774850000000
0!
0'
0/
#774860000000
#774870000000
1!
1'
1/
#774880000000
0!
0'
0/
#774890000000
1!
1'
1/
#774900000000
0!
1"
0'
1(
0/
10
#774910000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#774920000000
0!
0'
0/
#774930000000
1!
1'
1/
#774940000000
0!
0'
0/
#774950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#774960000000
0!
0'
0/
#774970000000
1!
1'
1/
#774980000000
0!
1"
0'
1(
0/
10
#774990000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#775000000000
0!
1$
0'
1+
0/
#775010000000
1!
1'
1/
#775020000000
0!
0'
0/
#775030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#775040000000
0!
0'
0/
#775050000000
1!
1'
1/
#775060000000
0!
0'
0/
#775070000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#775080000000
0!
0'
0/
#775090000000
1!
1'
1/
#775100000000
0!
0'
0/
#775110000000
1!
1'
1/
#775120000000
0!
0'
0/
#775130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#775140000000
0!
0'
0/
#775150000000
1!
1'
1/
#775160000000
0!
0'
0/
#775170000000
1!
1'
1/
#775180000000
0!
0'
0/
#775190000000
1!
1'
1/
#775200000000
0!
0'
0/
#775210000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#775220000000
0!
0'
0/
#775230000000
1!
1'
1/
#775240000000
0!
0'
0/
#775250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#775260000000
0!
0'
0/
#775270000000
1!
1'
1/
#775280000000
0!
0'
0/
#775290000000
#775300000000
1!
1'
1/
#775310000000
0!
0'
0/
#775320000000
1!
1'
1/
#775330000000
0!
1"
0'
1(
0/
10
#775340000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#775350000000
0!
0'
0/
#775360000000
1!
1'
1/
#775370000000
0!
0'
0/
#775380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#775390000000
0!
0'
0/
#775400000000
1!
1'
1/
#775410000000
0!
1"
0'
1(
0/
10
#775420000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#775430000000
0!
1$
0'
1+
0/
#775440000000
1!
1'
1/
#775450000000
0!
0'
0/
#775460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#775470000000
0!
0'
0/
#775480000000
1!
1'
1/
#775490000000
0!
0'
0/
#775500000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#775510000000
0!
0'
0/
#775520000000
1!
1'
1/
#775530000000
0!
0'
0/
#775540000000
1!
1'
1/
#775550000000
0!
0'
0/
#775560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#775570000000
0!
0'
0/
#775580000000
1!
1'
1/
#775590000000
0!
0'
0/
#775600000000
1!
1'
1/
#775610000000
0!
0'
0/
#775620000000
1!
1'
1/
#775630000000
0!
0'
0/
#775640000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#775650000000
0!
0'
0/
#775660000000
1!
1'
1/
#775670000000
0!
0'
0/
#775680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#775690000000
0!
0'
0/
#775700000000
1!
1'
1/
#775710000000
0!
0'
0/
#775720000000
#775730000000
1!
1'
1/
#775740000000
0!
0'
0/
#775750000000
1!
1'
1/
#775760000000
0!
1"
0'
1(
0/
10
#775770000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#775780000000
0!
0'
0/
#775790000000
1!
1'
1/
#775800000000
0!
0'
0/
#775810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#775820000000
0!
0'
0/
#775830000000
1!
1'
1/
#775840000000
0!
1"
0'
1(
0/
10
#775850000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#775860000000
0!
1$
0'
1+
0/
#775870000000
1!
1'
1/
#775880000000
0!
0'
0/
#775890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#775900000000
0!
0'
0/
#775910000000
1!
1'
1/
#775920000000
0!
0'
0/
#775930000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#775940000000
0!
0'
0/
#775950000000
1!
1'
1/
#775960000000
0!
0'
0/
#775970000000
1!
1'
1/
#775980000000
0!
0'
0/
#775990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#776000000000
0!
0'
0/
#776010000000
1!
1'
1/
#776020000000
0!
0'
0/
#776030000000
1!
1'
1/
#776040000000
0!
0'
0/
#776050000000
1!
1'
1/
#776060000000
0!
0'
0/
#776070000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#776080000000
0!
0'
0/
#776090000000
1!
1'
1/
#776100000000
0!
0'
0/
#776110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#776120000000
0!
0'
0/
#776130000000
1!
1'
1/
#776140000000
0!
0'
0/
#776150000000
#776160000000
1!
1'
1/
#776170000000
0!
0'
0/
#776180000000
1!
1'
1/
#776190000000
0!
1"
0'
1(
0/
10
#776200000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#776210000000
0!
0'
0/
#776220000000
1!
1'
1/
#776230000000
0!
0'
0/
#776240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#776250000000
0!
0'
0/
#776260000000
1!
1'
1/
#776270000000
0!
1"
0'
1(
0/
10
#776280000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#776290000000
0!
1$
0'
1+
0/
#776300000000
1!
1'
1/
#776310000000
0!
0'
0/
#776320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#776330000000
0!
0'
0/
#776340000000
1!
1'
1/
#776350000000
0!
0'
0/
#776360000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#776370000000
0!
0'
0/
#776380000000
1!
1'
1/
#776390000000
0!
0'
0/
#776400000000
1!
1'
1/
#776410000000
0!
0'
0/
#776420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#776430000000
0!
0'
0/
#776440000000
1!
1'
1/
#776450000000
0!
0'
0/
#776460000000
1!
1'
1/
#776470000000
0!
0'
0/
#776480000000
1!
1'
1/
#776490000000
0!
0'
0/
#776500000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#776510000000
0!
0'
0/
#776520000000
1!
1'
1/
#776530000000
0!
0'
0/
#776540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#776550000000
0!
0'
0/
#776560000000
1!
1'
1/
#776570000000
0!
0'
0/
#776580000000
#776590000000
1!
1'
1/
#776600000000
0!
0'
0/
#776610000000
1!
1'
1/
#776620000000
0!
1"
0'
1(
0/
10
#776630000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#776640000000
0!
0'
0/
#776650000000
1!
1'
1/
#776660000000
0!
0'
0/
#776670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#776680000000
0!
0'
0/
#776690000000
1!
1'
1/
#776700000000
0!
1"
0'
1(
0/
10
#776710000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#776720000000
0!
1$
0'
1+
0/
#776730000000
1!
1'
1/
#776740000000
0!
0'
0/
#776750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#776760000000
0!
0'
0/
#776770000000
1!
1'
1/
#776780000000
0!
0'
0/
#776790000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#776800000000
0!
0'
0/
#776810000000
1!
1'
1/
#776820000000
0!
0'
0/
#776830000000
1!
1'
1/
#776840000000
0!
0'
0/
#776850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#776860000000
0!
0'
0/
#776870000000
1!
1'
1/
#776880000000
0!
0'
0/
#776890000000
1!
1'
1/
#776900000000
0!
0'
0/
#776910000000
1!
1'
1/
#776920000000
0!
0'
0/
#776930000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#776940000000
0!
0'
0/
#776950000000
1!
1'
1/
#776960000000
0!
0'
0/
#776970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#776980000000
0!
0'
0/
#776990000000
1!
1'
1/
#777000000000
0!
0'
0/
#777010000000
#777020000000
1!
1'
1/
#777030000000
0!
0'
0/
#777040000000
1!
1'
1/
#777050000000
0!
1"
0'
1(
0/
10
#777060000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#777070000000
0!
0'
0/
#777080000000
1!
1'
1/
#777090000000
0!
0'
0/
#777100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#777110000000
0!
0'
0/
#777120000000
1!
1'
1/
#777130000000
0!
1"
0'
1(
0/
10
#777140000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#777150000000
0!
1$
0'
1+
0/
#777160000000
1!
1'
1/
#777170000000
0!
0'
0/
#777180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#777190000000
0!
0'
0/
#777200000000
1!
1'
1/
#777210000000
0!
0'
0/
#777220000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#777230000000
0!
0'
0/
#777240000000
1!
1'
1/
#777250000000
0!
0'
0/
#777260000000
1!
1'
1/
#777270000000
0!
0'
0/
#777280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#777290000000
0!
0'
0/
#777300000000
1!
1'
1/
#777310000000
0!
0'
0/
#777320000000
1!
1'
1/
#777330000000
0!
0'
0/
#777340000000
1!
1'
1/
#777350000000
0!
0'
0/
#777360000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#777370000000
0!
0'
0/
#777380000000
1!
1'
1/
#777390000000
0!
0'
0/
#777400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#777410000000
0!
0'
0/
#777420000000
1!
1'
1/
#777430000000
0!
0'
0/
#777440000000
#777450000000
1!
1'
1/
#777460000000
0!
0'
0/
#777470000000
1!
1'
1/
#777480000000
0!
1"
0'
1(
0/
10
#777490000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#777500000000
0!
0'
0/
#777510000000
1!
1'
1/
#777520000000
0!
0'
0/
#777530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#777540000000
0!
0'
0/
#777550000000
1!
1'
1/
#777560000000
0!
1"
0'
1(
0/
10
#777570000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#777580000000
0!
1$
0'
1+
0/
#777590000000
1!
1'
1/
#777600000000
0!
0'
0/
#777610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#777620000000
0!
0'
0/
#777630000000
1!
1'
1/
#777640000000
0!
0'
0/
#777650000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#777660000000
0!
0'
0/
#777670000000
1!
1'
1/
#777680000000
0!
0'
0/
#777690000000
1!
1'
1/
#777700000000
0!
0'
0/
#777710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#777720000000
0!
0'
0/
#777730000000
1!
1'
1/
#777740000000
0!
0'
0/
#777750000000
1!
1'
1/
#777760000000
0!
0'
0/
#777770000000
1!
1'
1/
#777780000000
0!
0'
0/
#777790000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#777800000000
0!
0'
0/
#777810000000
1!
1'
1/
#777820000000
0!
0'
0/
#777830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#777840000000
0!
0'
0/
#777850000000
1!
1'
1/
#777860000000
0!
0'
0/
#777870000000
#777880000000
1!
1'
1/
#777890000000
0!
0'
0/
#777900000000
1!
1'
1/
#777910000000
0!
1"
0'
1(
0/
10
#777920000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#777930000000
0!
0'
0/
#777940000000
1!
1'
1/
#777950000000
0!
0'
0/
#777960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#777970000000
0!
0'
0/
#777980000000
1!
1'
1/
#777990000000
0!
1"
0'
1(
0/
10
#778000000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#778010000000
0!
1$
0'
1+
0/
#778020000000
1!
1'
1/
#778030000000
0!
0'
0/
#778040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#778050000000
0!
0'
0/
#778060000000
1!
1'
1/
#778070000000
0!
0'
0/
#778080000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#778090000000
0!
0'
0/
#778100000000
1!
1'
1/
#778110000000
0!
0'
0/
#778120000000
1!
1'
1/
#778130000000
0!
0'
0/
#778140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#778150000000
0!
0'
0/
#778160000000
1!
1'
1/
#778170000000
0!
0'
0/
#778180000000
1!
1'
1/
#778190000000
0!
0'
0/
#778200000000
1!
1'
1/
#778210000000
0!
0'
0/
#778220000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#778230000000
0!
0'
0/
#778240000000
1!
1'
1/
#778250000000
0!
0'
0/
#778260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#778270000000
0!
0'
0/
#778280000000
1!
1'
1/
#778290000000
0!
0'
0/
#778300000000
#778310000000
1!
1'
1/
#778320000000
0!
0'
0/
#778330000000
1!
1'
1/
#778340000000
0!
1"
0'
1(
0/
10
#778350000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#778360000000
0!
0'
0/
#778370000000
1!
1'
1/
#778380000000
0!
0'
0/
#778390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#778400000000
0!
0'
0/
#778410000000
1!
1'
1/
#778420000000
0!
1"
0'
1(
0/
10
#778430000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#778440000000
0!
1$
0'
1+
0/
#778450000000
1!
1'
1/
#778460000000
0!
0'
0/
#778470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#778480000000
0!
0'
0/
#778490000000
1!
1'
1/
#778500000000
0!
0'
0/
#778510000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#778520000000
0!
0'
0/
#778530000000
1!
1'
1/
#778540000000
0!
0'
0/
#778550000000
1!
1'
1/
#778560000000
0!
0'
0/
#778570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#778580000000
0!
0'
0/
#778590000000
1!
1'
1/
#778600000000
0!
0'
0/
#778610000000
1!
1'
1/
#778620000000
0!
0'
0/
#778630000000
1!
1'
1/
#778640000000
0!
0'
0/
#778650000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#778660000000
0!
0'
0/
#778670000000
1!
1'
1/
#778680000000
0!
0'
0/
#778690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#778700000000
0!
0'
0/
#778710000000
1!
1'
1/
#778720000000
0!
0'
0/
#778730000000
#778740000000
1!
1'
1/
#778750000000
0!
0'
0/
#778760000000
1!
1'
1/
#778770000000
0!
1"
0'
1(
0/
10
#778780000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#778790000000
0!
0'
0/
#778800000000
1!
1'
1/
#778810000000
0!
0'
0/
#778820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#778830000000
0!
0'
0/
#778840000000
1!
1'
1/
#778850000000
0!
1"
0'
1(
0/
10
#778860000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#778870000000
0!
1$
0'
1+
0/
#778880000000
1!
1'
1/
#778890000000
0!
0'
0/
#778900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#778910000000
0!
0'
0/
#778920000000
1!
1'
1/
#778930000000
0!
0'
0/
#778940000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#778950000000
0!
0'
0/
#778960000000
1!
1'
1/
#778970000000
0!
0'
0/
#778980000000
1!
1'
1/
#778990000000
0!
0'
0/
#779000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#779010000000
0!
0'
0/
#779020000000
1!
1'
1/
#779030000000
0!
0'
0/
#779040000000
1!
1'
1/
#779050000000
0!
0'
0/
#779060000000
1!
1'
1/
#779070000000
0!
0'
0/
#779080000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#779090000000
0!
0'
0/
#779100000000
1!
1'
1/
#779110000000
0!
0'
0/
#779120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#779130000000
0!
0'
0/
#779140000000
1!
1'
1/
#779150000000
0!
0'
0/
#779160000000
#779170000000
1!
1'
1/
#779180000000
0!
0'
0/
#779190000000
1!
1'
1/
#779200000000
0!
1"
0'
1(
0/
10
#779210000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#779220000000
0!
0'
0/
#779230000000
1!
1'
1/
#779240000000
0!
0'
0/
#779250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#779260000000
0!
0'
0/
#779270000000
1!
1'
1/
#779280000000
0!
1"
0'
1(
0/
10
#779290000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#779300000000
0!
1$
0'
1+
0/
#779310000000
1!
1'
1/
#779320000000
0!
0'
0/
#779330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#779340000000
0!
0'
0/
#779350000000
1!
1'
1/
#779360000000
0!
0'
0/
#779370000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#779380000000
0!
0'
0/
#779390000000
1!
1'
1/
#779400000000
0!
0'
0/
#779410000000
1!
1'
1/
#779420000000
0!
0'
0/
#779430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#779440000000
0!
0'
0/
#779450000000
1!
1'
1/
#779460000000
0!
0'
0/
#779470000000
1!
1'
1/
#779480000000
0!
0'
0/
#779490000000
1!
1'
1/
#779500000000
0!
0'
0/
#779510000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#779520000000
0!
0'
0/
#779530000000
1!
1'
1/
#779540000000
0!
0'
0/
#779550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#779560000000
0!
0'
0/
#779570000000
1!
1'
1/
#779580000000
0!
0'
0/
#779590000000
#779600000000
1!
1'
1/
#779610000000
0!
0'
0/
#779620000000
1!
1'
1/
#779630000000
0!
1"
0'
1(
0/
10
#779640000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#779650000000
0!
0'
0/
#779660000000
1!
1'
1/
#779670000000
0!
0'
0/
#779680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#779690000000
0!
0'
0/
#779700000000
1!
1'
1/
#779710000000
0!
1"
0'
1(
0/
10
#779720000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#779730000000
0!
1$
0'
1+
0/
#779740000000
1!
1'
1/
#779750000000
0!
0'
0/
#779760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#779770000000
0!
0'
0/
#779780000000
1!
1'
1/
#779790000000
0!
0'
0/
#779800000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#779810000000
0!
0'
0/
#779820000000
1!
1'
1/
#779830000000
0!
0'
0/
#779840000000
1!
1'
1/
#779850000000
0!
0'
0/
#779860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#779870000000
0!
0'
0/
#779880000000
1!
1'
1/
#779890000000
0!
0'
0/
#779900000000
1!
1'
1/
#779910000000
0!
0'
0/
#779920000000
1!
1'
1/
#779930000000
0!
0'
0/
#779940000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#779950000000
0!
0'
0/
#779960000000
1!
1'
1/
#779970000000
0!
0'
0/
#779980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#779990000000
0!
0'
0/
#780000000000
1!
1'
1/
#780010000000
0!
0'
0/
#780020000000
#780030000000
1!
1'
1/
#780040000000
0!
0'
0/
#780050000000
1!
1'
1/
#780060000000
0!
1"
0'
1(
0/
10
#780070000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#780080000000
0!
0'
0/
#780090000000
1!
1'
1/
#780100000000
0!
0'
0/
#780110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#780120000000
0!
0'
0/
#780130000000
1!
1'
1/
#780140000000
0!
1"
0'
1(
0/
10
#780150000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#780160000000
0!
1$
0'
1+
0/
#780170000000
1!
1'
1/
#780180000000
0!
0'
0/
#780190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#780200000000
0!
0'
0/
#780210000000
1!
1'
1/
#780220000000
0!
0'
0/
#780230000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#780240000000
0!
0'
0/
#780250000000
1!
1'
1/
#780260000000
0!
0'
0/
#780270000000
1!
1'
1/
#780280000000
0!
0'
0/
#780290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#780300000000
0!
0'
0/
#780310000000
1!
1'
1/
#780320000000
0!
0'
0/
#780330000000
1!
1'
1/
#780340000000
0!
0'
0/
#780350000000
1!
1'
1/
#780360000000
0!
0'
0/
#780370000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#780380000000
0!
0'
0/
#780390000000
1!
1'
1/
#780400000000
0!
0'
0/
#780410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#780420000000
0!
0'
0/
#780430000000
1!
1'
1/
#780440000000
0!
0'
0/
#780450000000
#780460000000
1!
1'
1/
#780470000000
0!
0'
0/
#780480000000
1!
1'
1/
#780490000000
0!
1"
0'
1(
0/
10
#780500000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#780510000000
0!
0'
0/
#780520000000
1!
1'
1/
#780530000000
0!
0'
0/
#780540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#780550000000
0!
0'
0/
#780560000000
1!
1'
1/
#780570000000
0!
1"
0'
1(
0/
10
#780580000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#780590000000
0!
1$
0'
1+
0/
#780600000000
1!
1'
1/
#780610000000
0!
0'
0/
#780620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#780630000000
0!
0'
0/
#780640000000
1!
1'
1/
#780650000000
0!
0'
0/
#780660000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#780670000000
0!
0'
0/
#780680000000
1!
1'
1/
#780690000000
0!
0'
0/
#780700000000
1!
1'
1/
#780710000000
0!
0'
0/
#780720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#780730000000
0!
0'
0/
#780740000000
1!
1'
1/
#780750000000
0!
0'
0/
#780760000000
1!
1'
1/
#780770000000
0!
0'
0/
#780780000000
1!
1'
1/
#780790000000
0!
0'
0/
#780800000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#780810000000
0!
0'
0/
#780820000000
1!
1'
1/
#780830000000
0!
0'
0/
#780840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#780850000000
0!
0'
0/
#780860000000
1!
1'
1/
#780870000000
0!
0'
0/
#780880000000
#780890000000
1!
1'
1/
#780900000000
0!
0'
0/
#780910000000
1!
1'
1/
#780920000000
0!
1"
0'
1(
0/
10
#780930000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#780940000000
0!
0'
0/
#780950000000
1!
1'
1/
#780960000000
0!
0'
0/
#780970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#780980000000
0!
0'
0/
#780990000000
1!
1'
1/
#781000000000
0!
1"
0'
1(
0/
10
#781010000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#781020000000
0!
1$
0'
1+
0/
#781030000000
1!
1'
1/
#781040000000
0!
0'
0/
#781050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#781060000000
0!
0'
0/
#781070000000
1!
1'
1/
#781080000000
0!
0'
0/
#781090000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#781100000000
0!
0'
0/
#781110000000
1!
1'
1/
#781120000000
0!
0'
0/
#781130000000
1!
1'
1/
#781140000000
0!
0'
0/
#781150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#781160000000
0!
0'
0/
#781170000000
1!
1'
1/
#781180000000
0!
0'
0/
#781190000000
1!
1'
1/
#781200000000
0!
0'
0/
#781210000000
1!
1'
1/
#781220000000
0!
0'
0/
#781230000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#781240000000
0!
0'
0/
#781250000000
1!
1'
1/
#781260000000
0!
0'
0/
#781270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#781280000000
0!
0'
0/
#781290000000
1!
1'
1/
#781300000000
0!
0'
0/
#781310000000
#781320000000
1!
1'
1/
#781330000000
0!
0'
0/
#781340000000
1!
1'
1/
#781350000000
0!
1"
0'
1(
0/
10
#781360000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#781370000000
0!
0'
0/
#781380000000
1!
1'
1/
#781390000000
0!
0'
0/
#781400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#781410000000
0!
0'
0/
#781420000000
1!
1'
1/
#781430000000
0!
1"
0'
1(
0/
10
#781440000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#781450000000
0!
1$
0'
1+
0/
#781460000000
1!
1'
1/
#781470000000
0!
0'
0/
#781480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#781490000000
0!
0'
0/
#781500000000
1!
1'
1/
#781510000000
0!
0'
0/
#781520000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#781530000000
0!
0'
0/
#781540000000
1!
1'
1/
#781550000000
0!
0'
0/
#781560000000
1!
1'
1/
#781570000000
0!
0'
0/
#781580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#781590000000
0!
0'
0/
#781600000000
1!
1'
1/
#781610000000
0!
0'
0/
#781620000000
1!
1'
1/
#781630000000
0!
0'
0/
#781640000000
1!
1'
1/
#781650000000
0!
0'
0/
#781660000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#781670000000
0!
0'
0/
#781680000000
1!
1'
1/
#781690000000
0!
0'
0/
#781700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#781710000000
0!
0'
0/
#781720000000
1!
1'
1/
#781730000000
0!
0'
0/
#781740000000
#781750000000
1!
1'
1/
#781760000000
0!
0'
0/
#781770000000
1!
1'
1/
#781780000000
0!
1"
0'
1(
0/
10
#781790000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#781800000000
0!
0'
0/
#781810000000
1!
1'
1/
#781820000000
0!
0'
0/
#781830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#781840000000
0!
0'
0/
#781850000000
1!
1'
1/
#781860000000
0!
1"
0'
1(
0/
10
#781870000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#781880000000
0!
1$
0'
1+
0/
#781890000000
1!
1'
1/
#781900000000
0!
0'
0/
#781910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#781920000000
0!
0'
0/
#781930000000
1!
1'
1/
#781940000000
0!
0'
0/
#781950000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#781960000000
0!
0'
0/
#781970000000
1!
1'
1/
#781980000000
0!
0'
0/
#781990000000
1!
1'
1/
#782000000000
0!
0'
0/
#782010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#782020000000
0!
0'
0/
#782030000000
1!
1'
1/
#782040000000
0!
0'
0/
#782050000000
1!
1'
1/
#782060000000
0!
0'
0/
#782070000000
1!
1'
1/
#782080000000
0!
0'
0/
#782090000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#782100000000
0!
0'
0/
#782110000000
1!
1'
1/
#782120000000
0!
0'
0/
#782130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#782140000000
0!
0'
0/
#782150000000
1!
1'
1/
#782160000000
0!
0'
0/
#782170000000
#782180000000
1!
1'
1/
#782190000000
0!
0'
0/
#782200000000
1!
1'
1/
#782210000000
0!
1"
0'
1(
0/
10
#782220000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#782230000000
0!
0'
0/
#782240000000
1!
1'
1/
#782250000000
0!
0'
0/
#782260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#782270000000
0!
0'
0/
#782280000000
1!
1'
1/
#782290000000
0!
1"
0'
1(
0/
10
#782300000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#782310000000
0!
1$
0'
1+
0/
#782320000000
1!
1'
1/
#782330000000
0!
0'
0/
#782340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#782350000000
0!
0'
0/
#782360000000
1!
1'
1/
#782370000000
0!
0'
0/
#782380000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#782390000000
0!
0'
0/
#782400000000
1!
1'
1/
#782410000000
0!
0'
0/
#782420000000
1!
1'
1/
#782430000000
0!
0'
0/
#782440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#782450000000
0!
0'
0/
#782460000000
1!
1'
1/
#782470000000
0!
0'
0/
#782480000000
1!
1'
1/
#782490000000
0!
0'
0/
#782500000000
1!
1'
1/
#782510000000
0!
0'
0/
#782520000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#782530000000
0!
0'
0/
#782540000000
1!
1'
1/
#782550000000
0!
0'
0/
#782560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#782570000000
0!
0'
0/
#782580000000
1!
1'
1/
#782590000000
0!
0'
0/
#782600000000
#782610000000
1!
1'
1/
#782620000000
0!
0'
0/
#782630000000
1!
1'
1/
#782640000000
0!
1"
0'
1(
0/
10
#782650000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#782660000000
0!
0'
0/
#782670000000
1!
1'
1/
#782680000000
0!
0'
0/
#782690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#782700000000
0!
0'
0/
#782710000000
1!
1'
1/
#782720000000
0!
1"
0'
1(
0/
10
#782730000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#782740000000
0!
1$
0'
1+
0/
#782750000000
1!
1'
1/
#782760000000
0!
0'
0/
#782770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#782780000000
0!
0'
0/
#782790000000
1!
1'
1/
#782800000000
0!
0'
0/
#782810000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#782820000000
0!
0'
0/
#782830000000
1!
1'
1/
#782840000000
0!
0'
0/
#782850000000
1!
1'
1/
#782860000000
0!
0'
0/
#782870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#782880000000
0!
0'
0/
#782890000000
1!
1'
1/
#782900000000
0!
0'
0/
#782910000000
1!
1'
1/
#782920000000
0!
0'
0/
#782930000000
1!
1'
1/
#782940000000
0!
0'
0/
#782950000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#782960000000
0!
0'
0/
#782970000000
1!
1'
1/
#782980000000
0!
0'
0/
#782990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#783000000000
0!
0'
0/
#783010000000
1!
1'
1/
#783020000000
0!
0'
0/
#783030000000
#783040000000
1!
1'
1/
#783050000000
0!
0'
0/
#783060000000
1!
1'
1/
#783070000000
0!
1"
0'
1(
0/
10
#783080000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#783090000000
0!
0'
0/
#783100000000
1!
1'
1/
#783110000000
0!
0'
0/
#783120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#783130000000
0!
0'
0/
#783140000000
1!
1'
1/
#783150000000
0!
1"
0'
1(
0/
10
#783160000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#783170000000
0!
1$
0'
1+
0/
#783180000000
1!
1'
1/
#783190000000
0!
0'
0/
#783200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#783210000000
0!
0'
0/
#783220000000
1!
1'
1/
#783230000000
0!
0'
0/
#783240000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#783250000000
0!
0'
0/
#783260000000
1!
1'
1/
#783270000000
0!
0'
0/
#783280000000
1!
1'
1/
#783290000000
0!
0'
0/
#783300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#783310000000
0!
0'
0/
#783320000000
1!
1'
1/
#783330000000
0!
0'
0/
#783340000000
1!
1'
1/
#783350000000
0!
0'
0/
#783360000000
1!
1'
1/
#783370000000
0!
0'
0/
#783380000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#783390000000
0!
0'
0/
#783400000000
1!
1'
1/
#783410000000
0!
0'
0/
#783420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#783430000000
0!
0'
0/
#783440000000
1!
1'
1/
#783450000000
0!
0'
0/
#783460000000
#783470000000
1!
1'
1/
#783480000000
0!
0'
0/
#783490000000
1!
1'
1/
#783500000000
0!
1"
0'
1(
0/
10
#783510000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#783520000000
0!
0'
0/
#783530000000
1!
1'
1/
#783540000000
0!
0'
0/
#783550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#783560000000
0!
0'
0/
#783570000000
1!
1'
1/
#783580000000
0!
1"
0'
1(
0/
10
#783590000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#783600000000
0!
1$
0'
1+
0/
#783610000000
1!
1'
1/
#783620000000
0!
0'
0/
#783630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#783640000000
0!
0'
0/
#783650000000
1!
1'
1/
#783660000000
0!
0'
0/
#783670000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#783680000000
0!
0'
0/
#783690000000
1!
1'
1/
#783700000000
0!
0'
0/
#783710000000
1!
1'
1/
#783720000000
0!
0'
0/
#783730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#783740000000
0!
0'
0/
#783750000000
1!
1'
1/
#783760000000
0!
0'
0/
#783770000000
1!
1'
1/
#783780000000
0!
0'
0/
#783790000000
1!
1'
1/
#783800000000
0!
0'
0/
#783810000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#783820000000
0!
0'
0/
#783830000000
1!
1'
1/
#783840000000
0!
0'
0/
#783850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#783860000000
0!
0'
0/
#783870000000
1!
1'
1/
#783880000000
0!
0'
0/
#783890000000
#783900000000
1!
1'
1/
#783910000000
0!
0'
0/
#783920000000
1!
1'
1/
#783930000000
0!
1"
0'
1(
0/
10
#783940000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#783950000000
0!
0'
0/
#783960000000
1!
1'
1/
#783970000000
0!
0'
0/
#783980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#783990000000
0!
0'
0/
#784000000000
1!
1'
1/
#784010000000
0!
1"
0'
1(
0/
10
#784020000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#784030000000
0!
1$
0'
1+
0/
#784040000000
1!
1'
1/
#784050000000
0!
0'
0/
#784060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#784070000000
0!
0'
0/
#784080000000
1!
1'
1/
#784090000000
0!
0'
0/
#784100000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#784110000000
0!
0'
0/
#784120000000
1!
1'
1/
#784130000000
0!
0'
0/
#784140000000
1!
1'
1/
#784150000000
0!
0'
0/
#784160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#784170000000
0!
0'
0/
#784180000000
1!
1'
1/
#784190000000
0!
0'
0/
#784200000000
1!
1'
1/
#784210000000
0!
0'
0/
#784220000000
1!
1'
1/
#784230000000
0!
0'
0/
#784240000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#784250000000
0!
0'
0/
#784260000000
1!
1'
1/
#784270000000
0!
0'
0/
#784280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#784290000000
0!
0'
0/
#784300000000
1!
1'
1/
#784310000000
0!
0'
0/
#784320000000
#784330000000
1!
1'
1/
#784340000000
0!
0'
0/
#784350000000
1!
1'
1/
#784360000000
0!
1"
0'
1(
0/
10
#784370000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#784380000000
0!
0'
0/
#784390000000
1!
1'
1/
#784400000000
0!
0'
0/
#784410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#784420000000
0!
0'
0/
#784430000000
1!
1'
1/
#784440000000
0!
1"
0'
1(
0/
10
#784450000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#784460000000
0!
1$
0'
1+
0/
#784470000000
1!
1'
1/
#784480000000
0!
0'
0/
#784490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#784500000000
0!
0'
0/
#784510000000
1!
1'
1/
#784520000000
0!
0'
0/
#784530000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#784540000000
0!
0'
0/
#784550000000
1!
1'
1/
#784560000000
0!
0'
0/
#784570000000
1!
1'
1/
#784580000000
0!
0'
0/
#784590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#784600000000
0!
0'
0/
#784610000000
1!
1'
1/
#784620000000
0!
0'
0/
#784630000000
1!
1'
1/
#784640000000
0!
0'
0/
#784650000000
1!
1'
1/
#784660000000
0!
0'
0/
#784670000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#784680000000
0!
0'
0/
#784690000000
1!
1'
1/
#784700000000
0!
0'
0/
#784710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#784720000000
0!
0'
0/
#784730000000
1!
1'
1/
#784740000000
0!
0'
0/
#784750000000
#784760000000
1!
1'
1/
#784770000000
0!
0'
0/
#784780000000
1!
1'
1/
#784790000000
0!
1"
0'
1(
0/
10
#784800000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#784810000000
0!
0'
0/
#784820000000
1!
1'
1/
#784830000000
0!
0'
0/
#784840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#784850000000
0!
0'
0/
#784860000000
1!
1'
1/
#784870000000
0!
1"
0'
1(
0/
10
#784880000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#784890000000
0!
1$
0'
1+
0/
#784900000000
1!
1'
1/
#784910000000
0!
0'
0/
#784920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#784930000000
0!
0'
0/
#784940000000
1!
1'
1/
#784950000000
0!
0'
0/
#784960000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#784970000000
0!
0'
0/
#784980000000
1!
1'
1/
#784990000000
0!
0'
0/
#785000000000
1!
1'
1/
#785010000000
0!
0'
0/
#785020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#785030000000
0!
0'
0/
#785040000000
1!
1'
1/
#785050000000
0!
0'
0/
#785060000000
1!
1'
1/
#785070000000
0!
0'
0/
#785080000000
1!
1'
1/
#785090000000
0!
0'
0/
#785100000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#785110000000
0!
0'
0/
#785120000000
1!
1'
1/
#785130000000
0!
0'
0/
#785140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#785150000000
0!
0'
0/
#785160000000
1!
1'
1/
#785170000000
0!
0'
0/
#785180000000
#785190000000
1!
1'
1/
#785200000000
0!
0'
0/
#785210000000
1!
1'
1/
#785220000000
0!
1"
0'
1(
0/
10
#785230000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#785240000000
0!
0'
0/
#785250000000
1!
1'
1/
#785260000000
0!
0'
0/
#785270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#785280000000
0!
0'
0/
#785290000000
1!
1'
1/
#785300000000
0!
1"
0'
1(
0/
10
#785310000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#785320000000
0!
1$
0'
1+
0/
#785330000000
1!
1'
1/
#785340000000
0!
0'
0/
#785350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#785360000000
0!
0'
0/
#785370000000
1!
1'
1/
#785380000000
0!
0'
0/
#785390000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#785400000000
0!
0'
0/
#785410000000
1!
1'
1/
#785420000000
0!
0'
0/
#785430000000
1!
1'
1/
#785440000000
0!
0'
0/
#785450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#785460000000
0!
0'
0/
#785470000000
1!
1'
1/
#785480000000
0!
0'
0/
#785490000000
1!
1'
1/
#785500000000
0!
0'
0/
#785510000000
1!
1'
1/
#785520000000
0!
0'
0/
#785530000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#785540000000
0!
0'
0/
#785550000000
1!
1'
1/
#785560000000
0!
0'
0/
#785570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#785580000000
0!
0'
0/
#785590000000
1!
1'
1/
#785600000000
0!
0'
0/
#785610000000
#785620000000
1!
1'
1/
#785630000000
0!
0'
0/
#785640000000
1!
1'
1/
#785650000000
0!
1"
0'
1(
0/
10
#785660000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#785670000000
0!
0'
0/
#785680000000
1!
1'
1/
#785690000000
0!
0'
0/
#785700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#785710000000
0!
0'
0/
#785720000000
1!
1'
1/
#785730000000
0!
1"
0'
1(
0/
10
#785740000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#785750000000
0!
1$
0'
1+
0/
#785760000000
1!
1'
1/
#785770000000
0!
0'
0/
#785780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#785790000000
0!
0'
0/
#785800000000
1!
1'
1/
#785810000000
0!
0'
0/
#785820000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#785830000000
0!
0'
0/
#785840000000
1!
1'
1/
#785850000000
0!
0'
0/
#785860000000
1!
1'
1/
#785870000000
0!
0'
0/
#785880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#785890000000
0!
0'
0/
#785900000000
1!
1'
1/
#785910000000
0!
0'
0/
#785920000000
1!
1'
1/
#785930000000
0!
0'
0/
#785940000000
1!
1'
1/
#785950000000
0!
0'
0/
#785960000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#785970000000
0!
0'
0/
#785980000000
1!
1'
1/
#785990000000
0!
0'
0/
#786000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#786010000000
0!
0'
0/
#786020000000
1!
1'
1/
#786030000000
0!
0'
0/
#786040000000
#786050000000
1!
1'
1/
#786060000000
0!
0'
0/
#786070000000
1!
1'
1/
#786080000000
0!
1"
0'
1(
0/
10
#786090000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#786100000000
0!
0'
0/
#786110000000
1!
1'
1/
#786120000000
0!
0'
0/
#786130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#786140000000
0!
0'
0/
#786150000000
1!
1'
1/
#786160000000
0!
1"
0'
1(
0/
10
#786170000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#786180000000
0!
1$
0'
1+
0/
#786190000000
1!
1'
1/
#786200000000
0!
0'
0/
#786210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#786220000000
0!
0'
0/
#786230000000
1!
1'
1/
#786240000000
0!
0'
0/
#786250000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#786260000000
0!
0'
0/
#786270000000
1!
1'
1/
#786280000000
0!
0'
0/
#786290000000
1!
1'
1/
#786300000000
0!
0'
0/
#786310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#786320000000
0!
0'
0/
#786330000000
1!
1'
1/
#786340000000
0!
0'
0/
#786350000000
1!
1'
1/
#786360000000
0!
0'
0/
#786370000000
1!
1'
1/
#786380000000
0!
0'
0/
#786390000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#786400000000
0!
0'
0/
#786410000000
1!
1'
1/
#786420000000
0!
0'
0/
#786430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#786440000000
0!
0'
0/
#786450000000
1!
1'
1/
#786460000000
0!
0'
0/
#786470000000
#786480000000
1!
1'
1/
#786490000000
0!
0'
0/
#786500000000
1!
1'
1/
#786510000000
0!
1"
0'
1(
0/
10
#786520000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#786530000000
0!
0'
0/
#786540000000
1!
1'
1/
#786550000000
0!
0'
0/
#786560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#786570000000
0!
0'
0/
#786580000000
1!
1'
1/
#786590000000
0!
1"
0'
1(
0/
10
#786600000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#786610000000
0!
1$
0'
1+
0/
#786620000000
1!
1'
1/
#786630000000
0!
0'
0/
#786640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#786650000000
0!
0'
0/
#786660000000
1!
1'
1/
#786670000000
0!
0'
0/
#786680000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#786690000000
0!
0'
0/
#786700000000
1!
1'
1/
#786710000000
0!
0'
0/
#786720000000
1!
1'
1/
#786730000000
0!
0'
0/
#786740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#786750000000
0!
0'
0/
#786760000000
1!
1'
1/
#786770000000
0!
0'
0/
#786780000000
1!
1'
1/
#786790000000
0!
0'
0/
#786800000000
1!
1'
1/
#786810000000
0!
0'
0/
#786820000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#786830000000
0!
0'
0/
#786840000000
1!
1'
1/
#786850000000
0!
0'
0/
#786860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#786870000000
0!
0'
0/
#786880000000
1!
1'
1/
#786890000000
0!
0'
0/
#786900000000
#786910000000
1!
1'
1/
#786920000000
0!
0'
0/
#786930000000
1!
1'
1/
#786940000000
0!
1"
0'
1(
0/
10
#786950000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#786960000000
0!
0'
0/
#786970000000
1!
1'
1/
#786980000000
0!
0'
0/
#786990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#787000000000
0!
0'
0/
#787010000000
1!
1'
1/
#787020000000
0!
1"
0'
1(
0/
10
#787030000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#787040000000
0!
1$
0'
1+
0/
#787050000000
1!
1'
1/
#787060000000
0!
0'
0/
#787070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#787080000000
0!
0'
0/
#787090000000
1!
1'
1/
#787100000000
0!
0'
0/
#787110000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#787120000000
0!
0'
0/
#787130000000
1!
1'
1/
#787140000000
0!
0'
0/
#787150000000
1!
1'
1/
#787160000000
0!
0'
0/
#787170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#787180000000
0!
0'
0/
#787190000000
1!
1'
1/
#787200000000
0!
0'
0/
#787210000000
1!
1'
1/
#787220000000
0!
0'
0/
#787230000000
1!
1'
1/
#787240000000
0!
0'
0/
#787250000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#787260000000
0!
0'
0/
#787270000000
1!
1'
1/
#787280000000
0!
0'
0/
#787290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#787300000000
0!
0'
0/
#787310000000
1!
1'
1/
#787320000000
0!
0'
0/
#787330000000
#787340000000
1!
1'
1/
#787350000000
0!
0'
0/
#787360000000
1!
1'
1/
#787370000000
0!
1"
0'
1(
0/
10
#787380000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#787390000000
0!
0'
0/
#787400000000
1!
1'
1/
#787410000000
0!
0'
0/
#787420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#787430000000
0!
0'
0/
#787440000000
1!
1'
1/
#787450000000
0!
1"
0'
1(
0/
10
#787460000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#787470000000
0!
1$
0'
1+
0/
#787480000000
1!
1'
1/
#787490000000
0!
0'
0/
#787500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#787510000000
0!
0'
0/
#787520000000
1!
1'
1/
#787530000000
0!
0'
0/
#787540000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#787550000000
0!
0'
0/
#787560000000
1!
1'
1/
#787570000000
0!
0'
0/
#787580000000
1!
1'
1/
#787590000000
0!
0'
0/
#787600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#787610000000
0!
0'
0/
#787620000000
1!
1'
1/
#787630000000
0!
0'
0/
#787640000000
1!
1'
1/
#787650000000
0!
0'
0/
#787660000000
1!
1'
1/
#787670000000
0!
0'
0/
#787680000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#787690000000
0!
0'
0/
#787700000000
1!
1'
1/
#787710000000
0!
0'
0/
#787720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#787730000000
0!
0'
0/
#787740000000
1!
1'
1/
#787750000000
0!
0'
0/
#787760000000
#787770000000
1!
1'
1/
#787780000000
0!
0'
0/
#787790000000
1!
1'
1/
#787800000000
0!
1"
0'
1(
0/
10
#787810000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#787820000000
0!
0'
0/
#787830000000
1!
1'
1/
#787840000000
0!
0'
0/
#787850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#787860000000
0!
0'
0/
#787870000000
1!
1'
1/
#787880000000
0!
1"
0'
1(
0/
10
#787890000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#787900000000
0!
1$
0'
1+
0/
#787910000000
1!
1'
1/
#787920000000
0!
0'
0/
#787930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#787940000000
0!
0'
0/
#787950000000
1!
1'
1/
#787960000000
0!
0'
0/
#787970000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#787980000000
0!
0'
0/
#787990000000
1!
1'
1/
#788000000000
0!
0'
0/
#788010000000
1!
1'
1/
#788020000000
0!
0'
0/
#788030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#788040000000
0!
0'
0/
#788050000000
1!
1'
1/
#788060000000
0!
0'
0/
#788070000000
1!
1'
1/
#788080000000
0!
0'
0/
#788090000000
1!
1'
1/
#788100000000
0!
0'
0/
#788110000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#788120000000
0!
0'
0/
#788130000000
1!
1'
1/
#788140000000
0!
0'
0/
#788150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#788160000000
0!
0'
0/
#788170000000
1!
1'
1/
#788180000000
0!
0'
0/
#788190000000
#788200000000
1!
1'
1/
#788210000000
0!
0'
0/
#788220000000
1!
1'
1/
#788230000000
0!
1"
0'
1(
0/
10
#788240000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#788250000000
0!
0'
0/
#788260000000
1!
1'
1/
#788270000000
0!
0'
0/
#788280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#788290000000
0!
0'
0/
#788300000000
1!
1'
1/
#788310000000
0!
1"
0'
1(
0/
10
#788320000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#788330000000
0!
1$
0'
1+
0/
#788340000000
1!
1'
1/
#788350000000
0!
0'
0/
#788360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#788370000000
0!
0'
0/
#788380000000
1!
1'
1/
#788390000000
0!
0'
0/
#788400000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#788410000000
0!
0'
0/
#788420000000
1!
1'
1/
#788430000000
0!
0'
0/
#788440000000
1!
1'
1/
#788450000000
0!
0'
0/
#788460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#788470000000
0!
0'
0/
#788480000000
1!
1'
1/
#788490000000
0!
0'
0/
#788500000000
1!
1'
1/
#788510000000
0!
0'
0/
#788520000000
1!
1'
1/
#788530000000
0!
0'
0/
#788540000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#788550000000
0!
0'
0/
#788560000000
1!
1'
1/
#788570000000
0!
0'
0/
#788580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#788590000000
0!
0'
0/
#788600000000
1!
1'
1/
#788610000000
0!
0'
0/
#788620000000
#788630000000
1!
1'
1/
#788640000000
0!
0'
0/
#788650000000
1!
1'
1/
#788660000000
0!
1"
0'
1(
0/
10
#788670000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#788680000000
0!
0'
0/
#788690000000
1!
1'
1/
#788700000000
0!
0'
0/
#788710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#788720000000
0!
0'
0/
#788730000000
1!
1'
1/
#788740000000
0!
1"
0'
1(
0/
10
#788750000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#788760000000
0!
1$
0'
1+
0/
#788770000000
1!
1'
1/
#788780000000
0!
0'
0/
#788790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#788800000000
0!
0'
0/
#788810000000
1!
1'
1/
#788820000000
0!
0'
0/
#788830000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#788840000000
0!
0'
0/
#788850000000
1!
1'
1/
#788860000000
0!
0'
0/
#788870000000
1!
1'
1/
#788880000000
0!
0'
0/
#788890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#788900000000
0!
0'
0/
#788910000000
1!
1'
1/
#788920000000
0!
0'
0/
#788930000000
1!
1'
1/
#788940000000
0!
0'
0/
#788950000000
1!
1'
1/
#788960000000
0!
0'
0/
#788970000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#788980000000
0!
0'
0/
#788990000000
1!
1'
1/
#789000000000
0!
0'
0/
#789010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#789020000000
0!
0'
0/
#789030000000
1!
1'
1/
#789040000000
0!
0'
0/
#789050000000
#789060000000
1!
1'
1/
#789070000000
0!
0'
0/
#789080000000
1!
1'
1/
#789090000000
0!
1"
0'
1(
0/
10
#789100000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#789110000000
0!
0'
0/
#789120000000
1!
1'
1/
#789130000000
0!
0'
0/
#789140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#789150000000
0!
0'
0/
#789160000000
1!
1'
1/
#789170000000
0!
1"
0'
1(
0/
10
#789180000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#789190000000
0!
1$
0'
1+
0/
#789200000000
1!
1'
1/
#789210000000
0!
0'
0/
#789220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#789230000000
0!
0'
0/
#789240000000
1!
1'
1/
#789250000000
0!
0'
0/
#789260000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#789270000000
0!
0'
0/
#789280000000
1!
1'
1/
#789290000000
0!
0'
0/
#789300000000
1!
1'
1/
#789310000000
0!
0'
0/
#789320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#789330000000
0!
0'
0/
#789340000000
1!
1'
1/
#789350000000
0!
0'
0/
#789360000000
1!
1'
1/
#789370000000
0!
0'
0/
#789380000000
1!
1'
1/
#789390000000
0!
0'
0/
#789400000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#789410000000
0!
0'
0/
#789420000000
1!
1'
1/
#789430000000
0!
0'
0/
#789440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#789450000000
0!
0'
0/
#789460000000
1!
1'
1/
#789470000000
0!
0'
0/
#789480000000
#789490000000
1!
1'
1/
#789500000000
0!
0'
0/
#789510000000
1!
1'
1/
#789520000000
0!
1"
0'
1(
0/
10
#789530000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#789540000000
0!
0'
0/
#789550000000
1!
1'
1/
#789560000000
0!
0'
0/
#789570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#789580000000
0!
0'
0/
#789590000000
1!
1'
1/
#789600000000
0!
1"
0'
1(
0/
10
#789610000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#789620000000
0!
1$
0'
1+
0/
#789630000000
1!
1'
1/
#789640000000
0!
0'
0/
#789650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#789660000000
0!
0'
0/
#789670000000
1!
1'
1/
#789680000000
0!
0'
0/
#789690000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#789700000000
0!
0'
0/
#789710000000
1!
1'
1/
#789720000000
0!
0'
0/
#789730000000
1!
1'
1/
#789740000000
0!
0'
0/
#789750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#789760000000
0!
0'
0/
#789770000000
1!
1'
1/
#789780000000
0!
0'
0/
#789790000000
1!
1'
1/
#789800000000
0!
0'
0/
#789810000000
1!
1'
1/
#789820000000
0!
0'
0/
#789830000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#789840000000
0!
0'
0/
#789850000000
1!
1'
1/
#789860000000
0!
0'
0/
#789870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#789880000000
0!
0'
0/
#789890000000
1!
1'
1/
#789900000000
0!
0'
0/
#789910000000
#789920000000
1!
1'
1/
#789930000000
0!
0'
0/
#789940000000
1!
1'
1/
#789950000000
0!
1"
0'
1(
0/
10
#789960000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#789970000000
0!
0'
0/
#789980000000
1!
1'
1/
#789990000000
0!
0'
0/
#790000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#790010000000
0!
0'
0/
#790020000000
1!
1'
1/
#790030000000
0!
1"
0'
1(
0/
10
#790040000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#790050000000
0!
1$
0'
1+
0/
#790060000000
1!
1'
1/
#790070000000
0!
0'
0/
#790080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#790090000000
0!
0'
0/
#790100000000
1!
1'
1/
#790110000000
0!
0'
0/
#790120000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#790130000000
0!
0'
0/
#790140000000
1!
1'
1/
#790150000000
0!
0'
0/
#790160000000
1!
1'
1/
#790170000000
0!
0'
0/
#790180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#790190000000
0!
0'
0/
#790200000000
1!
1'
1/
#790210000000
0!
0'
0/
#790220000000
1!
1'
1/
#790230000000
0!
0'
0/
#790240000000
1!
1'
1/
#790250000000
0!
0'
0/
#790260000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#790270000000
0!
0'
0/
#790280000000
1!
1'
1/
#790290000000
0!
0'
0/
#790300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#790310000000
0!
0'
0/
#790320000000
1!
1'
1/
#790330000000
0!
0'
0/
#790340000000
#790350000000
1!
1'
1/
#790360000000
0!
0'
0/
#790370000000
1!
1'
1/
#790380000000
0!
1"
0'
1(
0/
10
#790390000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#790400000000
0!
0'
0/
#790410000000
1!
1'
1/
#790420000000
0!
0'
0/
#790430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#790440000000
0!
0'
0/
#790450000000
1!
1'
1/
#790460000000
0!
1"
0'
1(
0/
10
#790470000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#790480000000
0!
1$
0'
1+
0/
#790490000000
1!
1'
1/
#790500000000
0!
0'
0/
#790510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#790520000000
0!
0'
0/
#790530000000
1!
1'
1/
#790540000000
0!
0'
0/
#790550000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#790560000000
0!
0'
0/
#790570000000
1!
1'
1/
#790580000000
0!
0'
0/
#790590000000
1!
1'
1/
#790600000000
0!
0'
0/
#790610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#790620000000
0!
0'
0/
#790630000000
1!
1'
1/
#790640000000
0!
0'
0/
#790650000000
1!
1'
1/
#790660000000
0!
0'
0/
#790670000000
1!
1'
1/
#790680000000
0!
0'
0/
#790690000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#790700000000
0!
0'
0/
#790710000000
1!
1'
1/
#790720000000
0!
0'
0/
#790730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#790740000000
0!
0'
0/
#790750000000
1!
1'
1/
#790760000000
0!
0'
0/
#790770000000
#790780000000
1!
1'
1/
#790790000000
0!
0'
0/
#790800000000
1!
1'
1/
#790810000000
0!
1"
0'
1(
0/
10
#790820000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#790830000000
0!
0'
0/
#790840000000
1!
1'
1/
#790850000000
0!
0'
0/
#790860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#790870000000
0!
0'
0/
#790880000000
1!
1'
1/
#790890000000
0!
1"
0'
1(
0/
10
#790900000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#790910000000
0!
1$
0'
1+
0/
#790920000000
1!
1'
1/
#790930000000
0!
0'
0/
#790940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#790950000000
0!
0'
0/
#790960000000
1!
1'
1/
#790970000000
0!
0'
0/
#790980000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#790990000000
0!
0'
0/
#791000000000
1!
1'
1/
#791010000000
0!
0'
0/
#791020000000
1!
1'
1/
#791030000000
0!
0'
0/
#791040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#791050000000
0!
0'
0/
#791060000000
1!
1'
1/
#791070000000
0!
0'
0/
#791080000000
1!
1'
1/
#791090000000
0!
0'
0/
#791100000000
1!
1'
1/
#791110000000
0!
0'
0/
#791120000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#791130000000
0!
0'
0/
#791140000000
1!
1'
1/
#791150000000
0!
0'
0/
#791160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#791170000000
0!
0'
0/
#791180000000
1!
1'
1/
#791190000000
0!
0'
0/
#791200000000
#791210000000
1!
1'
1/
#791220000000
0!
0'
0/
#791230000000
1!
1'
1/
#791240000000
0!
1"
0'
1(
0/
10
#791250000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#791260000000
0!
0'
0/
#791270000000
1!
1'
1/
#791280000000
0!
0'
0/
#791290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#791300000000
0!
0'
0/
#791310000000
1!
1'
1/
#791320000000
0!
1"
0'
1(
0/
10
#791330000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#791340000000
0!
1$
0'
1+
0/
#791350000000
1!
1'
1/
#791360000000
0!
0'
0/
#791370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#791380000000
0!
0'
0/
#791390000000
1!
1'
1/
#791400000000
0!
0'
0/
#791410000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#791420000000
0!
0'
0/
#791430000000
1!
1'
1/
#791440000000
0!
0'
0/
#791450000000
1!
1'
1/
#791460000000
0!
0'
0/
#791470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#791480000000
0!
0'
0/
#791490000000
1!
1'
1/
#791500000000
0!
0'
0/
#791510000000
1!
1'
1/
#791520000000
0!
0'
0/
#791530000000
1!
1'
1/
#791540000000
0!
0'
0/
#791550000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#791560000000
0!
0'
0/
#791570000000
1!
1'
1/
#791580000000
0!
0'
0/
#791590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#791600000000
0!
0'
0/
#791610000000
1!
1'
1/
#791620000000
0!
0'
0/
#791630000000
#791640000000
1!
1'
1/
#791650000000
0!
0'
0/
#791660000000
1!
1'
1/
#791670000000
0!
1"
0'
1(
0/
10
#791680000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#791690000000
0!
0'
0/
#791700000000
1!
1'
1/
#791710000000
0!
0'
0/
#791720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#791730000000
0!
0'
0/
#791740000000
1!
1'
1/
#791750000000
0!
1"
0'
1(
0/
10
#791760000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#791770000000
0!
1$
0'
1+
0/
#791780000000
1!
1'
1/
#791790000000
0!
0'
0/
#791800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#791810000000
0!
0'
0/
#791820000000
1!
1'
1/
#791830000000
0!
0'
0/
#791840000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#791850000000
0!
0'
0/
#791860000000
1!
1'
1/
#791870000000
0!
0'
0/
#791880000000
1!
1'
1/
#791890000000
0!
0'
0/
#791900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#791910000000
0!
0'
0/
#791920000000
1!
1'
1/
#791930000000
0!
0'
0/
#791940000000
1!
1'
1/
#791950000000
0!
0'
0/
#791960000000
1!
1'
1/
#791970000000
0!
0'
0/
#791980000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#791990000000
0!
0'
0/
#792000000000
1!
1'
1/
#792010000000
0!
0'
0/
#792020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#792030000000
0!
0'
0/
#792040000000
1!
1'
1/
#792050000000
0!
0'
0/
#792060000000
#792070000000
1!
1'
1/
#792080000000
0!
0'
0/
#792090000000
1!
1'
1/
#792100000000
0!
1"
0'
1(
0/
10
#792110000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#792120000000
0!
0'
0/
#792130000000
1!
1'
1/
#792140000000
0!
0'
0/
#792150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#792160000000
0!
0'
0/
#792170000000
1!
1'
1/
#792180000000
0!
1"
0'
1(
0/
10
#792190000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#792200000000
0!
1$
0'
1+
0/
#792210000000
1!
1'
1/
#792220000000
0!
0'
0/
#792230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#792240000000
0!
0'
0/
#792250000000
1!
1'
1/
#792260000000
0!
0'
0/
#792270000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#792280000000
0!
0'
0/
#792290000000
1!
1'
1/
#792300000000
0!
0'
0/
#792310000000
1!
1'
1/
#792320000000
0!
0'
0/
#792330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#792340000000
0!
0'
0/
#792350000000
1!
1'
1/
#792360000000
0!
0'
0/
#792370000000
1!
1'
1/
#792380000000
0!
0'
0/
#792390000000
1!
1'
1/
#792400000000
0!
0'
0/
#792410000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#792420000000
0!
0'
0/
#792430000000
1!
1'
1/
#792440000000
0!
0'
0/
#792450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#792460000000
0!
0'
0/
#792470000000
1!
1'
1/
#792480000000
0!
0'
0/
#792490000000
#792500000000
1!
1'
1/
#792510000000
0!
0'
0/
#792520000000
1!
1'
1/
#792530000000
0!
1"
0'
1(
0/
10
#792540000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#792550000000
0!
0'
0/
#792560000000
1!
1'
1/
#792570000000
0!
0'
0/
#792580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#792590000000
0!
0'
0/
#792600000000
1!
1'
1/
#792610000000
0!
1"
0'
1(
0/
10
#792620000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#792630000000
0!
1$
0'
1+
0/
#792640000000
1!
1'
1/
#792650000000
0!
0'
0/
#792660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#792670000000
0!
0'
0/
#792680000000
1!
1'
1/
#792690000000
0!
0'
0/
#792700000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#792710000000
0!
0'
0/
#792720000000
1!
1'
1/
#792730000000
0!
0'
0/
#792740000000
1!
1'
1/
#792750000000
0!
0'
0/
#792760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#792770000000
0!
0'
0/
#792780000000
1!
1'
1/
#792790000000
0!
0'
0/
#792800000000
1!
1'
1/
#792810000000
0!
0'
0/
#792820000000
1!
1'
1/
#792830000000
0!
0'
0/
#792840000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#792850000000
0!
0'
0/
#792860000000
1!
1'
1/
#792870000000
0!
0'
0/
#792880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#792890000000
0!
0'
0/
#792900000000
1!
1'
1/
#792910000000
0!
0'
0/
#792920000000
#792930000000
1!
1'
1/
#792940000000
0!
0'
0/
#792950000000
1!
1'
1/
#792960000000
0!
1"
0'
1(
0/
10
#792970000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#792980000000
0!
0'
0/
#792990000000
1!
1'
1/
#793000000000
0!
0'
0/
#793010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#793020000000
0!
0'
0/
#793030000000
1!
1'
1/
#793040000000
0!
1"
0'
1(
0/
10
#793050000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#793060000000
0!
1$
0'
1+
0/
#793070000000
1!
1'
1/
#793080000000
0!
0'
0/
#793090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#793100000000
0!
0'
0/
#793110000000
1!
1'
1/
#793120000000
0!
0'
0/
#793130000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#793140000000
0!
0'
0/
#793150000000
1!
1'
1/
#793160000000
0!
0'
0/
#793170000000
1!
1'
1/
#793180000000
0!
0'
0/
#793190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#793200000000
0!
0'
0/
#793210000000
1!
1'
1/
#793220000000
0!
0'
0/
#793230000000
1!
1'
1/
#793240000000
0!
0'
0/
#793250000000
1!
1'
1/
#793260000000
0!
0'
0/
#793270000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#793280000000
0!
0'
0/
#793290000000
1!
1'
1/
#793300000000
0!
0'
0/
#793310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#793320000000
0!
0'
0/
#793330000000
1!
1'
1/
#793340000000
0!
0'
0/
#793350000000
#793360000000
1!
1'
1/
#793370000000
0!
0'
0/
#793380000000
1!
1'
1/
#793390000000
0!
1"
0'
1(
0/
10
#793400000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#793410000000
0!
0'
0/
#793420000000
1!
1'
1/
#793430000000
0!
0'
0/
#793440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#793450000000
0!
0'
0/
#793460000000
1!
1'
1/
#793470000000
0!
1"
0'
1(
0/
10
#793480000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#793490000000
0!
1$
0'
1+
0/
#793500000000
1!
1'
1/
#793510000000
0!
0'
0/
#793520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#793530000000
0!
0'
0/
#793540000000
1!
1'
1/
#793550000000
0!
0'
0/
#793560000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#793570000000
0!
0'
0/
#793580000000
1!
1'
1/
#793590000000
0!
0'
0/
#793600000000
1!
1'
1/
#793610000000
0!
0'
0/
#793620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#793630000000
0!
0'
0/
#793640000000
1!
1'
1/
#793650000000
0!
0'
0/
#793660000000
1!
1'
1/
#793670000000
0!
0'
0/
#793680000000
1!
1'
1/
#793690000000
0!
0'
0/
#793700000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#793710000000
0!
0'
0/
#793720000000
1!
1'
1/
#793730000000
0!
0'
0/
#793740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#793750000000
0!
0'
0/
#793760000000
1!
1'
1/
#793770000000
0!
0'
0/
#793780000000
#793790000000
1!
1'
1/
#793800000000
0!
0'
0/
#793810000000
1!
1'
1/
#793820000000
0!
1"
0'
1(
0/
10
#793830000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#793840000000
0!
0'
0/
#793850000000
1!
1'
1/
#793860000000
0!
0'
0/
#793870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#793880000000
0!
0'
0/
#793890000000
1!
1'
1/
#793900000000
0!
1"
0'
1(
0/
10
#793910000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#793920000000
0!
1$
0'
1+
0/
#793930000000
1!
1'
1/
#793940000000
0!
0'
0/
#793950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#793960000000
0!
0'
0/
#793970000000
1!
1'
1/
#793980000000
0!
0'
0/
#793990000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#794000000000
0!
0'
0/
#794010000000
1!
1'
1/
#794020000000
0!
0'
0/
#794030000000
1!
1'
1/
#794040000000
0!
0'
0/
#794050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#794060000000
0!
0'
0/
#794070000000
1!
1'
1/
#794080000000
0!
0'
0/
#794090000000
1!
1'
1/
#794100000000
0!
0'
0/
#794110000000
1!
1'
1/
#794120000000
0!
0'
0/
#794130000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#794140000000
0!
0'
0/
#794150000000
1!
1'
1/
#794160000000
0!
0'
0/
#794170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#794180000000
0!
0'
0/
#794190000000
1!
1'
1/
#794200000000
0!
0'
0/
#794210000000
#794220000000
1!
1'
1/
#794230000000
0!
0'
0/
#794240000000
1!
1'
1/
#794250000000
0!
1"
0'
1(
0/
10
#794260000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#794270000000
0!
0'
0/
#794280000000
1!
1'
1/
#794290000000
0!
0'
0/
#794300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#794310000000
0!
0'
0/
#794320000000
1!
1'
1/
#794330000000
0!
1"
0'
1(
0/
10
#794340000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#794350000000
0!
1$
0'
1+
0/
#794360000000
1!
1'
1/
#794370000000
0!
0'
0/
#794380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#794390000000
0!
0'
0/
#794400000000
1!
1'
1/
#794410000000
0!
0'
0/
#794420000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#794430000000
0!
0'
0/
#794440000000
1!
1'
1/
#794450000000
0!
0'
0/
#794460000000
1!
1'
1/
#794470000000
0!
0'
0/
#794480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#794490000000
0!
0'
0/
#794500000000
1!
1'
1/
#794510000000
0!
0'
0/
#794520000000
1!
1'
1/
#794530000000
0!
0'
0/
#794540000000
1!
1'
1/
#794550000000
0!
0'
0/
#794560000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#794570000000
0!
0'
0/
#794580000000
1!
1'
1/
#794590000000
0!
0'
0/
#794600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#794610000000
0!
0'
0/
#794620000000
1!
1'
1/
#794630000000
0!
0'
0/
#794640000000
#794650000000
1!
1'
1/
#794660000000
0!
0'
0/
#794670000000
1!
1'
1/
#794680000000
0!
1"
0'
1(
0/
10
#794690000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#794700000000
0!
0'
0/
#794710000000
1!
1'
1/
#794720000000
0!
0'
0/
#794730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#794740000000
0!
0'
0/
#794750000000
1!
1'
1/
#794760000000
0!
1"
0'
1(
0/
10
#794770000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#794780000000
0!
1$
0'
1+
0/
#794790000000
1!
1'
1/
#794800000000
0!
0'
0/
#794810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#794820000000
0!
0'
0/
#794830000000
1!
1'
1/
#794840000000
0!
0'
0/
#794850000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#794860000000
0!
0'
0/
#794870000000
1!
1'
1/
#794880000000
0!
0'
0/
#794890000000
1!
1'
1/
#794900000000
0!
0'
0/
#794910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#794920000000
0!
0'
0/
#794930000000
1!
1'
1/
#794940000000
0!
0'
0/
#794950000000
1!
1'
1/
#794960000000
0!
0'
0/
#794970000000
1!
1'
1/
#794980000000
0!
0'
0/
#794990000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#795000000000
0!
0'
0/
#795010000000
1!
1'
1/
#795020000000
0!
0'
0/
#795030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#795040000000
0!
0'
0/
#795050000000
1!
1'
1/
#795060000000
0!
0'
0/
#795070000000
#795080000000
1!
1'
1/
#795090000000
0!
0'
0/
#795100000000
1!
1'
1/
#795110000000
0!
1"
0'
1(
0/
10
#795120000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#795130000000
0!
0'
0/
#795140000000
1!
1'
1/
#795150000000
0!
0'
0/
#795160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#795170000000
0!
0'
0/
#795180000000
1!
1'
1/
#795190000000
0!
1"
0'
1(
0/
10
#795200000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#795210000000
0!
1$
0'
1+
0/
#795220000000
1!
1'
1/
#795230000000
0!
0'
0/
#795240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#795250000000
0!
0'
0/
#795260000000
1!
1'
1/
#795270000000
0!
0'
0/
#795280000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#795290000000
0!
0'
0/
#795300000000
1!
1'
1/
#795310000000
0!
0'
0/
#795320000000
1!
1'
1/
#795330000000
0!
0'
0/
#795340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#795350000000
0!
0'
0/
#795360000000
1!
1'
1/
#795370000000
0!
0'
0/
#795380000000
1!
1'
1/
#795390000000
0!
0'
0/
#795400000000
1!
1'
1/
#795410000000
0!
0'
0/
#795420000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#795430000000
0!
0'
0/
#795440000000
1!
1'
1/
#795450000000
0!
0'
0/
#795460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#795470000000
0!
0'
0/
#795480000000
1!
1'
1/
#795490000000
0!
0'
0/
#795500000000
#795510000000
1!
1'
1/
#795520000000
0!
0'
0/
#795530000000
1!
1'
1/
#795540000000
0!
1"
0'
1(
0/
10
#795550000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#795560000000
0!
0'
0/
#795570000000
1!
1'
1/
#795580000000
0!
0'
0/
#795590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#795600000000
0!
0'
0/
#795610000000
1!
1'
1/
#795620000000
0!
1"
0'
1(
0/
10
#795630000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#795640000000
0!
1$
0'
1+
0/
#795650000000
1!
1'
1/
#795660000000
0!
0'
0/
#795670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#795680000000
0!
0'
0/
#795690000000
1!
1'
1/
#795700000000
0!
0'
0/
#795710000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#795720000000
0!
0'
0/
#795730000000
1!
1'
1/
#795740000000
0!
0'
0/
#795750000000
1!
1'
1/
#795760000000
0!
0'
0/
#795770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#795780000000
0!
0'
0/
#795790000000
1!
1'
1/
#795800000000
0!
0'
0/
#795810000000
1!
1'
1/
#795820000000
0!
0'
0/
#795830000000
1!
1'
1/
#795840000000
0!
0'
0/
#795850000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#795860000000
0!
0'
0/
#795870000000
1!
1'
1/
#795880000000
0!
0'
0/
#795890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#795900000000
0!
0'
0/
#795910000000
1!
1'
1/
#795920000000
0!
0'
0/
#795930000000
#795940000000
1!
1'
1/
#795950000000
0!
0'
0/
#795960000000
1!
1'
1/
#795970000000
0!
1"
0'
1(
0/
10
#795980000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#795990000000
0!
0'
0/
#796000000000
1!
1'
1/
#796010000000
0!
0'
0/
#796020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#796030000000
0!
0'
0/
#796040000000
1!
1'
1/
#796050000000
0!
1"
0'
1(
0/
10
#796060000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#796070000000
0!
1$
0'
1+
0/
#796080000000
1!
1'
1/
#796090000000
0!
0'
0/
#796100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#796110000000
0!
0'
0/
#796120000000
1!
1'
1/
#796130000000
0!
0'
0/
#796140000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#796150000000
0!
0'
0/
#796160000000
1!
1'
1/
#796170000000
0!
0'
0/
#796180000000
1!
1'
1/
#796190000000
0!
0'
0/
#796200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#796210000000
0!
0'
0/
#796220000000
1!
1'
1/
#796230000000
0!
0'
0/
#796240000000
1!
1'
1/
#796250000000
0!
0'
0/
#796260000000
1!
1'
1/
#796270000000
0!
0'
0/
#796280000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#796290000000
0!
0'
0/
#796300000000
1!
1'
1/
#796310000000
0!
0'
0/
#796320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#796330000000
0!
0'
0/
#796340000000
1!
1'
1/
#796350000000
0!
0'
0/
#796360000000
#796370000000
1!
1'
1/
#796380000000
0!
0'
0/
#796390000000
1!
1'
1/
#796400000000
0!
1"
0'
1(
0/
10
#796410000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#796420000000
0!
0'
0/
#796430000000
1!
1'
1/
#796440000000
0!
0'
0/
#796450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#796460000000
0!
0'
0/
#796470000000
1!
1'
1/
#796480000000
0!
1"
0'
1(
0/
10
#796490000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#796500000000
0!
1$
0'
1+
0/
#796510000000
1!
1'
1/
#796520000000
0!
0'
0/
#796530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#796540000000
0!
0'
0/
#796550000000
1!
1'
1/
#796560000000
0!
0'
0/
#796570000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#796580000000
0!
0'
0/
#796590000000
1!
1'
1/
#796600000000
0!
0'
0/
#796610000000
1!
1'
1/
#796620000000
0!
0'
0/
#796630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#796640000000
0!
0'
0/
#796650000000
1!
1'
1/
#796660000000
0!
0'
0/
#796670000000
1!
1'
1/
#796680000000
0!
0'
0/
#796690000000
1!
1'
1/
#796700000000
0!
0'
0/
#796710000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#796720000000
0!
0'
0/
#796730000000
1!
1'
1/
#796740000000
0!
0'
0/
#796750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#796760000000
0!
0'
0/
#796770000000
1!
1'
1/
#796780000000
0!
0'
0/
#796790000000
#796800000000
1!
1'
1/
#796810000000
0!
0'
0/
#796820000000
1!
1'
1/
#796830000000
0!
1"
0'
1(
0/
10
#796840000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#796850000000
0!
0'
0/
#796860000000
1!
1'
1/
#796870000000
0!
0'
0/
#796880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#796890000000
0!
0'
0/
#796900000000
1!
1'
1/
#796910000000
0!
1"
0'
1(
0/
10
#796920000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#796930000000
0!
1$
0'
1+
0/
#796940000000
1!
1'
1/
#796950000000
0!
0'
0/
#796960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#796970000000
0!
0'
0/
#796980000000
1!
1'
1/
#796990000000
0!
0'
0/
#797000000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#797010000000
0!
0'
0/
#797020000000
1!
1'
1/
#797030000000
0!
0'
0/
#797040000000
1!
1'
1/
#797050000000
0!
0'
0/
#797060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#797070000000
0!
0'
0/
#797080000000
1!
1'
1/
#797090000000
0!
0'
0/
#797100000000
1!
1'
1/
#797110000000
0!
0'
0/
#797120000000
1!
1'
1/
#797130000000
0!
0'
0/
#797140000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#797150000000
0!
0'
0/
#797160000000
1!
1'
1/
#797170000000
0!
0'
0/
#797180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#797190000000
0!
0'
0/
#797200000000
1!
1'
1/
#797210000000
0!
0'
0/
#797220000000
#797230000000
1!
1'
1/
#797240000000
0!
0'
0/
#797250000000
1!
1'
1/
#797260000000
0!
1"
0'
1(
0/
10
#797270000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#797280000000
0!
0'
0/
#797290000000
1!
1'
1/
#797300000000
0!
0'
0/
#797310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#797320000000
0!
0'
0/
#797330000000
1!
1'
1/
#797340000000
0!
1"
0'
1(
0/
10
#797350000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#797360000000
0!
1$
0'
1+
0/
#797370000000
1!
1'
1/
#797380000000
0!
0'
0/
#797390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#797400000000
0!
0'
0/
#797410000000
1!
1'
1/
#797420000000
0!
0'
0/
#797430000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#797440000000
0!
0'
0/
#797450000000
1!
1'
1/
#797460000000
0!
0'
0/
#797470000000
1!
1'
1/
#797480000000
0!
0'
0/
#797490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#797500000000
0!
0'
0/
#797510000000
1!
1'
1/
#797520000000
0!
0'
0/
#797530000000
1!
1'
1/
#797540000000
0!
0'
0/
#797550000000
1!
1'
1/
#797560000000
0!
0'
0/
#797570000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#797580000000
0!
0'
0/
#797590000000
1!
1'
1/
#797600000000
0!
0'
0/
#797610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#797620000000
0!
0'
0/
#797630000000
1!
1'
1/
#797640000000
0!
0'
0/
#797650000000
#797660000000
1!
1'
1/
#797670000000
0!
0'
0/
#797680000000
1!
1'
1/
#797690000000
0!
1"
0'
1(
0/
10
#797700000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#797710000000
0!
0'
0/
#797720000000
1!
1'
1/
#797730000000
0!
0'
0/
#797740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#797750000000
0!
0'
0/
#797760000000
1!
1'
1/
#797770000000
0!
1"
0'
1(
0/
10
#797780000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#797790000000
0!
1$
0'
1+
0/
#797800000000
1!
1'
1/
#797810000000
0!
0'
0/
#797820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#797830000000
0!
0'
0/
#797840000000
1!
1'
1/
#797850000000
0!
0'
0/
#797860000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#797870000000
0!
0'
0/
#797880000000
1!
1'
1/
#797890000000
0!
0'
0/
#797900000000
1!
1'
1/
#797910000000
0!
0'
0/
#797920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#797930000000
0!
0'
0/
#797940000000
1!
1'
1/
#797950000000
0!
0'
0/
#797960000000
1!
1'
1/
#797970000000
0!
0'
0/
#797980000000
1!
1'
1/
#797990000000
0!
0'
0/
#798000000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#798010000000
0!
0'
0/
#798020000000
1!
1'
1/
#798030000000
0!
0'
0/
#798040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#798050000000
0!
0'
0/
#798060000000
1!
1'
1/
#798070000000
0!
0'
0/
#798080000000
#798090000000
1!
1'
1/
#798100000000
0!
0'
0/
#798110000000
1!
1'
1/
#798120000000
0!
1"
0'
1(
0/
10
#798130000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#798140000000
0!
0'
0/
#798150000000
1!
1'
1/
#798160000000
0!
0'
0/
#798170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#798180000000
0!
0'
0/
#798190000000
1!
1'
1/
#798200000000
0!
1"
0'
1(
0/
10
#798210000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#798220000000
0!
1$
0'
1+
0/
#798230000000
1!
1'
1/
#798240000000
0!
0'
0/
#798250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#798260000000
0!
0'
0/
#798270000000
1!
1'
1/
#798280000000
0!
0'
0/
#798290000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#798300000000
0!
0'
0/
#798310000000
1!
1'
1/
#798320000000
0!
0'
0/
#798330000000
1!
1'
1/
#798340000000
0!
0'
0/
#798350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#798360000000
0!
0'
0/
#798370000000
1!
1'
1/
#798380000000
0!
0'
0/
#798390000000
1!
1'
1/
#798400000000
0!
0'
0/
#798410000000
1!
1'
1/
#798420000000
0!
0'
0/
#798430000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#798440000000
0!
0'
0/
#798450000000
1!
1'
1/
#798460000000
0!
0'
0/
#798470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#798480000000
0!
0'
0/
#798490000000
1!
1'
1/
#798500000000
0!
0'
0/
#798510000000
#798520000000
1!
1'
1/
#798530000000
0!
0'
0/
#798540000000
1!
1'
1/
#798550000000
0!
1"
0'
1(
0/
10
#798560000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#798570000000
0!
0'
0/
#798580000000
1!
1'
1/
#798590000000
0!
0'
0/
#798600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#798610000000
0!
0'
0/
#798620000000
1!
1'
1/
#798630000000
0!
1"
0'
1(
0/
10
#798640000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#798650000000
0!
1$
0'
1+
0/
#798660000000
1!
1'
1/
#798670000000
0!
0'
0/
#798680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#798690000000
0!
0'
0/
#798700000000
1!
1'
1/
#798710000000
0!
0'
0/
#798720000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#798730000000
0!
0'
0/
#798740000000
1!
1'
1/
#798750000000
0!
0'
0/
#798760000000
1!
1'
1/
#798770000000
0!
0'
0/
#798780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#798790000000
0!
0'
0/
#798800000000
1!
1'
1/
#798810000000
0!
0'
0/
#798820000000
1!
1'
1/
#798830000000
0!
0'
0/
#798840000000
1!
1'
1/
#798850000000
0!
0'
0/
#798860000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#798870000000
0!
0'
0/
#798880000000
1!
1'
1/
#798890000000
0!
0'
0/
#798900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#798910000000
0!
0'
0/
#798920000000
1!
1'
1/
#798930000000
0!
0'
0/
#798940000000
#798950000000
1!
1'
1/
#798960000000
0!
0'
0/
#798970000000
1!
1'
1/
#798980000000
0!
1"
0'
1(
0/
10
#798990000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#799000000000
0!
0'
0/
#799010000000
1!
1'
1/
#799020000000
0!
0'
0/
#799030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#799040000000
0!
0'
0/
#799050000000
1!
1'
1/
#799060000000
0!
1"
0'
1(
0/
10
#799070000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#799080000000
0!
1$
0'
1+
0/
#799090000000
1!
1'
1/
#799100000000
0!
0'
0/
#799110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#799120000000
0!
0'
0/
#799130000000
1!
1'
1/
#799140000000
0!
0'
0/
#799150000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#799160000000
0!
0'
0/
#799170000000
1!
1'
1/
#799180000000
0!
0'
0/
#799190000000
1!
1'
1/
#799200000000
0!
0'
0/
#799210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#799220000000
0!
0'
0/
#799230000000
1!
1'
1/
#799240000000
0!
0'
0/
#799250000000
1!
1'
1/
#799260000000
0!
0'
0/
#799270000000
1!
1'
1/
#799280000000
0!
0'
0/
#799290000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#799300000000
0!
0'
0/
#799310000000
1!
1'
1/
#799320000000
0!
0'
0/
#799330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#799340000000
0!
0'
0/
#799350000000
1!
1'
1/
#799360000000
0!
0'
0/
#799370000000
#799380000000
1!
1'
1/
#799390000000
0!
0'
0/
#799400000000
1!
1'
1/
#799410000000
0!
1"
0'
1(
0/
10
#799420000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#799430000000
0!
0'
0/
#799440000000
1!
1'
1/
#799450000000
0!
0'
0/
#799460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#799470000000
0!
0'
0/
#799480000000
1!
1'
1/
#799490000000
0!
1"
0'
1(
0/
10
#799500000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#799510000000
0!
1$
0'
1+
0/
#799520000000
1!
1'
1/
#799530000000
0!
0'
0/
#799540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#799550000000
0!
0'
0/
#799560000000
1!
1'
1/
#799570000000
0!
0'
0/
#799580000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#799590000000
0!
0'
0/
#799600000000
1!
1'
1/
#799610000000
0!
0'
0/
#799620000000
1!
1'
1/
#799630000000
0!
0'
0/
#799640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#799650000000
0!
0'
0/
#799660000000
1!
1'
1/
#799670000000
0!
0'
0/
#799680000000
1!
1'
1/
#799690000000
0!
0'
0/
#799700000000
1!
1'
1/
#799710000000
0!
0'
0/
#799720000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#799730000000
0!
0'
0/
#799740000000
1!
1'
1/
#799750000000
0!
0'
0/
#799760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#799770000000
0!
0'
0/
#799780000000
1!
1'
1/
#799790000000
0!
0'
0/
#799800000000
#799810000000
1!
1'
1/
#799820000000
0!
0'
0/
#799830000000
1!
1'
1/
#799840000000
0!
1"
0'
1(
0/
10
#799850000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#799860000000
0!
0'
0/
#799870000000
1!
1'
1/
#799880000000
0!
0'
0/
#799890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#799900000000
0!
0'
0/
#799910000000
1!
1'
1/
#799920000000
0!
1"
0'
1(
0/
10
#799930000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#799940000000
0!
1$
0'
1+
0/
#799950000000
1!
1'
1/
#799960000000
0!
0'
0/
#799970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#799980000000
0!
0'
0/
#799990000000
1!
1'
1/
#800000000000
0!
0'
0/
#800010000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#800020000000
0!
0'
0/
#800030000000
1!
1'
1/
#800040000000
0!
0'
0/
#800050000000
1!
1'
1/
#800060000000
0!
0'
0/
#800070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#800080000000
0!
0'
0/
#800090000000
1!
1'
1/
#800100000000
0!
0'
0/
#800110000000
1!
1'
1/
#800120000000
0!
0'
0/
#800130000000
1!
1'
1/
#800140000000
0!
0'
0/
#800150000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#800160000000
0!
0'
0/
#800170000000
1!
1'
1/
#800180000000
0!
0'
0/
#800190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#800200000000
0!
0'
0/
#800210000000
1!
1'
1/
#800220000000
0!
0'
0/
#800230000000
#800240000000
1!
1'
1/
#800250000000
0!
0'
0/
#800260000000
1!
1'
1/
#800270000000
0!
1"
0'
1(
0/
10
#800280000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#800290000000
0!
0'
0/
#800300000000
1!
1'
1/
#800310000000
0!
0'
0/
#800320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#800330000000
0!
0'
0/
#800340000000
1!
1'
1/
#800350000000
0!
1"
0'
1(
0/
10
#800360000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#800370000000
0!
1$
0'
1+
0/
#800380000000
1!
1'
1/
#800390000000
0!
0'
0/
#800400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#800410000000
0!
0'
0/
#800420000000
1!
1'
1/
#800430000000
0!
0'
0/
#800440000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#800450000000
0!
0'
0/
#800460000000
1!
1'
1/
#800470000000
0!
0'
0/
#800480000000
1!
1'
1/
#800490000000
0!
0'
0/
#800500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#800510000000
0!
0'
0/
#800520000000
1!
1'
1/
#800530000000
0!
0'
0/
#800540000000
1!
1'
1/
#800550000000
0!
0'
0/
#800560000000
1!
1'
1/
#800570000000
0!
0'
0/
#800580000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#800590000000
0!
0'
0/
#800600000000
1!
1'
1/
#800610000000
0!
0'
0/
#800620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#800630000000
0!
0'
0/
#800640000000
1!
1'
1/
#800650000000
0!
0'
0/
#800660000000
#800670000000
1!
1'
1/
#800680000000
0!
0'
0/
#800690000000
1!
1'
1/
#800700000000
0!
1"
0'
1(
0/
10
#800710000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#800720000000
0!
0'
0/
#800730000000
1!
1'
1/
#800740000000
0!
0'
0/
#800750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#800760000000
0!
0'
0/
#800770000000
1!
1'
1/
#800780000000
0!
1"
0'
1(
0/
10
#800790000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#800800000000
0!
1$
0'
1+
0/
#800810000000
1!
1'
1/
#800820000000
0!
0'
0/
#800830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#800840000000
0!
0'
0/
#800850000000
1!
1'
1/
#800860000000
0!
0'
0/
#800870000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#800880000000
0!
0'
0/
#800890000000
1!
1'
1/
#800900000000
0!
0'
0/
#800910000000
1!
1'
1/
#800920000000
0!
0'
0/
#800930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#800940000000
0!
0'
0/
#800950000000
1!
1'
1/
#800960000000
0!
0'
0/
#800970000000
1!
1'
1/
#800980000000
0!
0'
0/
#800990000000
1!
1'
1/
#801000000000
0!
0'
0/
#801010000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#801020000000
0!
0'
0/
#801030000000
1!
1'
1/
#801040000000
0!
0'
0/
#801050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#801060000000
0!
0'
0/
#801070000000
1!
1'
1/
#801080000000
0!
0'
0/
#801090000000
#801100000000
1!
1'
1/
#801110000000
0!
0'
0/
#801120000000
1!
1'
1/
#801130000000
0!
1"
0'
1(
0/
10
#801140000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#801150000000
0!
0'
0/
#801160000000
1!
1'
1/
#801170000000
0!
0'
0/
#801180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#801190000000
0!
0'
0/
#801200000000
1!
1'
1/
#801210000000
0!
1"
0'
1(
0/
10
#801220000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#801230000000
0!
1$
0'
1+
0/
#801240000000
1!
1'
1/
#801250000000
0!
0'
0/
#801260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#801270000000
0!
0'
0/
#801280000000
1!
1'
1/
#801290000000
0!
0'
0/
#801300000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#801310000000
0!
0'
0/
#801320000000
1!
1'
1/
#801330000000
0!
0'
0/
#801340000000
1!
1'
1/
#801350000000
0!
0'
0/
#801360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#801370000000
0!
0'
0/
#801380000000
1!
1'
1/
#801390000000
0!
0'
0/
#801400000000
1!
1'
1/
#801410000000
0!
0'
0/
#801420000000
1!
1'
1/
#801430000000
0!
0'
0/
#801440000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#801450000000
0!
0'
0/
#801460000000
1!
1'
1/
#801470000000
0!
0'
0/
#801480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#801490000000
0!
0'
0/
#801500000000
1!
1'
1/
#801510000000
0!
0'
0/
#801520000000
#801530000000
1!
1'
1/
#801540000000
0!
0'
0/
#801550000000
1!
1'
1/
#801560000000
0!
1"
0'
1(
0/
10
#801570000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#801580000000
0!
0'
0/
#801590000000
1!
1'
1/
#801600000000
0!
0'
0/
#801610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#801620000000
0!
0'
0/
#801630000000
1!
1'
1/
#801640000000
0!
1"
0'
1(
0/
10
#801650000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#801660000000
0!
1$
0'
1+
0/
#801670000000
1!
1'
1/
#801680000000
0!
0'
0/
#801690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#801700000000
0!
0'
0/
#801710000000
1!
1'
1/
#801720000000
0!
0'
0/
#801730000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#801740000000
0!
0'
0/
#801750000000
1!
1'
1/
#801760000000
0!
0'
0/
#801770000000
1!
1'
1/
#801780000000
0!
0'
0/
#801790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#801800000000
0!
0'
0/
#801810000000
1!
1'
1/
#801820000000
0!
0'
0/
#801830000000
1!
1'
1/
#801840000000
0!
0'
0/
#801850000000
1!
1'
1/
#801860000000
0!
0'
0/
#801870000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#801880000000
0!
0'
0/
#801890000000
1!
1'
1/
#801900000000
0!
0'
0/
#801910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#801920000000
0!
0'
0/
#801930000000
1!
1'
1/
#801940000000
0!
0'
0/
#801950000000
#801960000000
1!
1'
1/
#801970000000
0!
0'
0/
#801980000000
1!
1'
1/
#801990000000
0!
1"
0'
1(
0/
10
#802000000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#802010000000
0!
0'
0/
#802020000000
1!
1'
1/
#802030000000
0!
0'
0/
#802040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#802050000000
0!
0'
0/
#802060000000
1!
1'
1/
#802070000000
0!
1"
0'
1(
0/
10
#802080000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#802090000000
0!
1$
0'
1+
0/
#802100000000
1!
1'
1/
#802110000000
0!
0'
0/
#802120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#802130000000
0!
0'
0/
#802140000000
1!
1'
1/
#802150000000
0!
0'
0/
#802160000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#802170000000
0!
0'
0/
#802180000000
1!
1'
1/
#802190000000
0!
0'
0/
#802200000000
1!
1'
1/
#802210000000
0!
0'
0/
#802220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#802230000000
0!
0'
0/
#802240000000
1!
1'
1/
#802250000000
0!
0'
0/
#802260000000
1!
1'
1/
#802270000000
0!
0'
0/
#802280000000
1!
1'
1/
#802290000000
0!
0'
0/
#802300000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#802310000000
0!
0'
0/
#802320000000
1!
1'
1/
#802330000000
0!
0'
0/
#802340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#802350000000
0!
0'
0/
#802360000000
1!
1'
1/
#802370000000
0!
0'
0/
#802380000000
#802390000000
1!
1'
1/
#802400000000
0!
0'
0/
#802410000000
1!
1'
1/
#802420000000
0!
1"
0'
1(
0/
10
#802430000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#802440000000
0!
0'
0/
#802450000000
1!
1'
1/
#802460000000
0!
0'
0/
#802470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#802480000000
0!
0'
0/
#802490000000
1!
1'
1/
#802500000000
0!
1"
0'
1(
0/
10
#802510000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#802520000000
0!
1$
0'
1+
0/
#802530000000
1!
1'
1/
#802540000000
0!
0'
0/
#802550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#802560000000
0!
0'
0/
#802570000000
1!
1'
1/
#802580000000
0!
0'
0/
#802590000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#802600000000
0!
0'
0/
#802610000000
1!
1'
1/
#802620000000
0!
0'
0/
#802630000000
1!
1'
1/
#802640000000
0!
0'
0/
#802650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#802660000000
0!
0'
0/
#802670000000
1!
1'
1/
#802680000000
0!
0'
0/
#802690000000
1!
1'
1/
#802700000000
0!
0'
0/
#802710000000
1!
1'
1/
#802720000000
0!
0'
0/
#802730000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#802740000000
0!
0'
0/
#802750000000
1!
1'
1/
#802760000000
0!
0'
0/
#802770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#802780000000
0!
0'
0/
#802790000000
1!
1'
1/
#802800000000
0!
0'
0/
#802810000000
#802820000000
1!
1'
1/
#802830000000
0!
0'
0/
#802840000000
1!
1'
1/
#802850000000
0!
1"
0'
1(
0/
10
#802860000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#802870000000
0!
0'
0/
#802880000000
1!
1'
1/
#802890000000
0!
0'
0/
#802900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#802910000000
0!
0'
0/
#802920000000
1!
1'
1/
#802930000000
0!
1"
0'
1(
0/
10
#802940000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#802950000000
0!
1$
0'
1+
0/
#802960000000
1!
1'
1/
#802970000000
0!
0'
0/
#802980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#802990000000
0!
0'
0/
#803000000000
1!
1'
1/
#803010000000
0!
0'
0/
#803020000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#803030000000
0!
0'
0/
#803040000000
1!
1'
1/
#803050000000
0!
0'
0/
#803060000000
1!
1'
1/
#803070000000
0!
0'
0/
#803080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#803090000000
0!
0'
0/
#803100000000
1!
1'
1/
#803110000000
0!
0'
0/
#803120000000
1!
1'
1/
#803130000000
0!
0'
0/
#803140000000
1!
1'
1/
#803150000000
0!
0'
0/
#803160000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#803170000000
0!
0'
0/
#803180000000
1!
1'
1/
#803190000000
0!
0'
0/
#803200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#803210000000
0!
0'
0/
#803220000000
1!
1'
1/
#803230000000
0!
0'
0/
#803240000000
#803250000000
1!
1'
1/
#803260000000
0!
0'
0/
#803270000000
1!
1'
1/
#803280000000
0!
1"
0'
1(
0/
10
#803290000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#803300000000
0!
0'
0/
#803310000000
1!
1'
1/
#803320000000
0!
0'
0/
#803330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#803340000000
0!
0'
0/
#803350000000
1!
1'
1/
#803360000000
0!
1"
0'
1(
0/
10
#803370000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#803380000000
0!
1$
0'
1+
0/
#803390000000
1!
1'
1/
#803400000000
0!
0'
0/
#803410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#803420000000
0!
0'
0/
#803430000000
1!
1'
1/
#803440000000
0!
0'
0/
#803450000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#803460000000
0!
0'
0/
#803470000000
1!
1'
1/
#803480000000
0!
0'
0/
#803490000000
1!
1'
1/
#803500000000
0!
0'
0/
#803510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#803520000000
0!
0'
0/
#803530000000
1!
1'
1/
#803540000000
0!
0'
0/
#803550000000
1!
1'
1/
#803560000000
0!
0'
0/
#803570000000
1!
1'
1/
#803580000000
0!
0'
0/
#803590000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#803600000000
0!
0'
0/
#803610000000
1!
1'
1/
#803620000000
0!
0'
0/
#803630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#803640000000
0!
0'
0/
#803650000000
1!
1'
1/
#803660000000
0!
0'
0/
#803670000000
#803680000000
1!
1'
1/
#803690000000
0!
0'
0/
#803700000000
1!
1'
1/
#803710000000
0!
1"
0'
1(
0/
10
#803720000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#803730000000
0!
0'
0/
#803740000000
1!
1'
1/
#803750000000
0!
0'
0/
#803760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#803770000000
0!
0'
0/
#803780000000
1!
1'
1/
#803790000000
0!
1"
0'
1(
0/
10
#803800000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#803810000000
0!
1$
0'
1+
0/
#803820000000
1!
1'
1/
#803830000000
0!
0'
0/
#803840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#803850000000
0!
0'
0/
#803860000000
1!
1'
1/
#803870000000
0!
0'
0/
#803880000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#803890000000
0!
0'
0/
#803900000000
1!
1'
1/
#803910000000
0!
0'
0/
#803920000000
1!
1'
1/
#803930000000
0!
0'
0/
#803940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#803950000000
0!
0'
0/
#803960000000
1!
1'
1/
#803970000000
0!
0'
0/
#803980000000
1!
1'
1/
#803990000000
0!
0'
0/
#804000000000
1!
1'
1/
#804010000000
0!
0'
0/
#804020000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#804030000000
0!
0'
0/
#804040000000
1!
1'
1/
#804050000000
0!
0'
0/
#804060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#804070000000
0!
0'
0/
#804080000000
1!
1'
1/
#804090000000
0!
0'
0/
#804100000000
#804110000000
1!
1'
1/
#804120000000
0!
0'
0/
#804130000000
1!
1'
1/
#804140000000
0!
1"
0'
1(
0/
10
#804150000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#804160000000
0!
0'
0/
#804170000000
1!
1'
1/
#804180000000
0!
0'
0/
#804190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#804200000000
0!
0'
0/
#804210000000
1!
1'
1/
#804220000000
0!
1"
0'
1(
0/
10
#804230000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#804240000000
0!
1$
0'
1+
0/
#804250000000
1!
1'
1/
#804260000000
0!
0'
0/
#804270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#804280000000
0!
0'
0/
#804290000000
1!
1'
1/
#804300000000
0!
0'
0/
#804310000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#804320000000
0!
0'
0/
#804330000000
1!
1'
1/
#804340000000
0!
0'
0/
#804350000000
1!
1'
1/
#804360000000
0!
0'
0/
#804370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#804380000000
0!
0'
0/
#804390000000
1!
1'
1/
#804400000000
0!
0'
0/
#804410000000
1!
1'
1/
#804420000000
0!
0'
0/
#804430000000
1!
1'
1/
#804440000000
0!
0'
0/
#804450000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#804460000000
0!
0'
0/
#804470000000
1!
1'
1/
#804480000000
0!
0'
0/
#804490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#804500000000
0!
0'
0/
#804510000000
1!
1'
1/
#804520000000
0!
0'
0/
#804530000000
#804540000000
1!
1'
1/
#804550000000
0!
0'
0/
#804560000000
1!
1'
1/
#804570000000
0!
1"
0'
1(
0/
10
#804580000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#804590000000
0!
0'
0/
#804600000000
1!
1'
1/
#804610000000
0!
0'
0/
#804620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#804630000000
0!
0'
0/
#804640000000
1!
1'
1/
#804650000000
0!
1"
0'
1(
0/
10
#804660000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#804670000000
0!
1$
0'
1+
0/
#804680000000
1!
1'
1/
#804690000000
0!
0'
0/
#804700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#804710000000
0!
0'
0/
#804720000000
1!
1'
1/
#804730000000
0!
0'
0/
#804740000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#804750000000
0!
0'
0/
#804760000000
1!
1'
1/
#804770000000
0!
0'
0/
#804780000000
1!
1'
1/
#804790000000
0!
0'
0/
#804800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#804810000000
0!
0'
0/
#804820000000
1!
1'
1/
#804830000000
0!
0'
0/
#804840000000
1!
1'
1/
#804850000000
0!
0'
0/
#804860000000
1!
1'
1/
#804870000000
0!
0'
0/
#804880000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#804890000000
0!
0'
0/
#804900000000
1!
1'
1/
#804910000000
0!
0'
0/
#804920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#804930000000
0!
0'
0/
#804940000000
1!
1'
1/
#804950000000
0!
0'
0/
#804960000000
#804970000000
1!
1'
1/
#804980000000
0!
0'
0/
#804990000000
1!
1'
1/
#805000000000
0!
1"
0'
1(
0/
10
#805010000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#805020000000
0!
0'
0/
#805030000000
1!
1'
1/
#805040000000
0!
0'
0/
#805050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#805060000000
0!
0'
0/
#805070000000
1!
1'
1/
#805080000000
0!
1"
0'
1(
0/
10
#805090000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#805100000000
0!
1$
0'
1+
0/
#805110000000
1!
1'
1/
#805120000000
0!
0'
0/
#805130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#805140000000
0!
0'
0/
#805150000000
1!
1'
1/
#805160000000
0!
0'
0/
#805170000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#805180000000
0!
0'
0/
#805190000000
1!
1'
1/
#805200000000
0!
0'
0/
#805210000000
1!
1'
1/
#805220000000
0!
0'
0/
#805230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#805240000000
0!
0'
0/
#805250000000
1!
1'
1/
#805260000000
0!
0'
0/
#805270000000
1!
1'
1/
#805280000000
0!
0'
0/
#805290000000
1!
1'
1/
#805300000000
0!
0'
0/
#805310000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#805320000000
0!
0'
0/
#805330000000
1!
1'
1/
#805340000000
0!
0'
0/
#805350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#805360000000
0!
0'
0/
#805370000000
1!
1'
1/
#805380000000
0!
0'
0/
#805390000000
#805400000000
1!
1'
1/
#805410000000
0!
0'
0/
#805420000000
1!
1'
1/
#805430000000
0!
1"
0'
1(
0/
10
#805440000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#805450000000
0!
0'
0/
#805460000000
1!
1'
1/
#805470000000
0!
0'
0/
#805480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#805490000000
0!
0'
0/
#805500000000
1!
1'
1/
#805510000000
0!
1"
0'
1(
0/
10
#805520000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#805530000000
0!
1$
0'
1+
0/
#805540000000
1!
1'
1/
#805550000000
0!
0'
0/
#805560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#805570000000
0!
0'
0/
#805580000000
1!
1'
1/
#805590000000
0!
0'
0/
#805600000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#805610000000
0!
0'
0/
#805620000000
1!
1'
1/
#805630000000
0!
0'
0/
#805640000000
1!
1'
1/
#805650000000
0!
0'
0/
#805660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#805670000000
0!
0'
0/
#805680000000
1!
1'
1/
#805690000000
0!
0'
0/
#805700000000
1!
1'
1/
#805710000000
0!
0'
0/
#805720000000
1!
1'
1/
#805730000000
0!
0'
0/
#805740000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#805750000000
0!
0'
0/
#805760000000
1!
1'
1/
#805770000000
0!
0'
0/
#805780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#805790000000
0!
0'
0/
#805800000000
1!
1'
1/
#805810000000
0!
0'
0/
#805820000000
#805830000000
1!
1'
1/
#805840000000
0!
0'
0/
#805850000000
1!
1'
1/
#805860000000
0!
1"
0'
1(
0/
10
#805870000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#805880000000
0!
0'
0/
#805890000000
1!
1'
1/
#805900000000
0!
0'
0/
#805910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#805920000000
0!
0'
0/
#805930000000
1!
1'
1/
#805940000000
0!
1"
0'
1(
0/
10
#805950000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#805960000000
0!
1$
0'
1+
0/
#805970000000
1!
1'
1/
#805980000000
0!
0'
0/
#805990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#806000000000
0!
0'
0/
#806010000000
1!
1'
1/
#806020000000
0!
0'
0/
#806030000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#806040000000
0!
0'
0/
#806050000000
1!
1'
1/
#806060000000
0!
0'
0/
#806070000000
1!
1'
1/
#806080000000
0!
0'
0/
#806090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#806100000000
0!
0'
0/
#806110000000
1!
1'
1/
#806120000000
0!
0'
0/
#806130000000
1!
1'
1/
#806140000000
0!
0'
0/
#806150000000
1!
1'
1/
#806160000000
0!
0'
0/
#806170000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#806180000000
0!
0'
0/
#806190000000
1!
1'
1/
#806200000000
0!
0'
0/
#806210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#806220000000
0!
0'
0/
#806230000000
1!
1'
1/
#806240000000
0!
0'
0/
#806250000000
#806260000000
1!
1'
1/
#806270000000
0!
0'
0/
#806280000000
1!
1'
1/
#806290000000
0!
1"
0'
1(
0/
10
#806300000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#806310000000
0!
0'
0/
#806320000000
1!
1'
1/
#806330000000
0!
0'
0/
#806340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#806350000000
0!
0'
0/
#806360000000
1!
1'
1/
#806370000000
0!
1"
0'
1(
0/
10
#806380000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#806390000000
0!
1$
0'
1+
0/
#806400000000
1!
1'
1/
#806410000000
0!
0'
0/
#806420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#806430000000
0!
0'
0/
#806440000000
1!
1'
1/
#806450000000
0!
0'
0/
#806460000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#806470000000
0!
0'
0/
#806480000000
1!
1'
1/
#806490000000
0!
0'
0/
#806500000000
1!
1'
1/
#806510000000
0!
0'
0/
#806520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#806530000000
0!
0'
0/
#806540000000
1!
1'
1/
#806550000000
0!
0'
0/
#806560000000
1!
1'
1/
#806570000000
0!
0'
0/
#806580000000
1!
1'
1/
#806590000000
0!
0'
0/
#806600000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#806610000000
0!
0'
0/
#806620000000
1!
1'
1/
#806630000000
0!
0'
0/
#806640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#806650000000
0!
0'
0/
#806660000000
1!
1'
1/
#806670000000
0!
0'
0/
#806680000000
#806690000000
1!
1'
1/
#806700000000
0!
0'
0/
#806710000000
1!
1'
1/
#806720000000
0!
1"
0'
1(
0/
10
#806730000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#806740000000
0!
0'
0/
#806750000000
1!
1'
1/
#806760000000
0!
0'
0/
#806770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#806780000000
0!
0'
0/
#806790000000
1!
1'
1/
#806800000000
0!
1"
0'
1(
0/
10
#806810000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#806820000000
0!
1$
0'
1+
0/
#806830000000
1!
1'
1/
#806840000000
0!
0'
0/
#806850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#806860000000
0!
0'
0/
#806870000000
1!
1'
1/
#806880000000
0!
0'
0/
#806890000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#806900000000
0!
0'
0/
#806910000000
1!
1'
1/
#806920000000
0!
0'
0/
#806930000000
1!
1'
1/
#806940000000
0!
0'
0/
#806950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#806960000000
0!
0'
0/
#806970000000
1!
1'
1/
#806980000000
0!
0'
0/
#806990000000
1!
1'
1/
#807000000000
0!
0'
0/
#807010000000
1!
1'
1/
#807020000000
0!
0'
0/
#807030000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#807040000000
0!
0'
0/
#807050000000
1!
1'
1/
#807060000000
0!
0'
0/
#807070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#807080000000
0!
0'
0/
#807090000000
1!
1'
1/
#807100000000
0!
0'
0/
#807110000000
#807120000000
1!
1'
1/
#807130000000
0!
0'
0/
#807140000000
1!
1'
1/
#807150000000
0!
1"
0'
1(
0/
10
#807160000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#807170000000
0!
0'
0/
#807180000000
1!
1'
1/
#807190000000
0!
0'
0/
#807200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#807210000000
0!
0'
0/
#807220000000
1!
1'
1/
#807230000000
0!
1"
0'
1(
0/
10
#807240000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#807250000000
0!
1$
0'
1+
0/
#807260000000
1!
1'
1/
#807270000000
0!
0'
0/
#807280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#807290000000
0!
0'
0/
#807300000000
1!
1'
1/
#807310000000
0!
0'
0/
#807320000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#807330000000
0!
0'
0/
#807340000000
1!
1'
1/
#807350000000
0!
0'
0/
#807360000000
1!
1'
1/
#807370000000
0!
0'
0/
#807380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#807390000000
0!
0'
0/
#807400000000
1!
1'
1/
#807410000000
0!
0'
0/
#807420000000
1!
1'
1/
#807430000000
0!
0'
0/
#807440000000
1!
1'
1/
#807450000000
0!
0'
0/
#807460000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#807470000000
0!
0'
0/
#807480000000
1!
1'
1/
#807490000000
0!
0'
0/
#807500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#807510000000
0!
0'
0/
#807520000000
1!
1'
1/
#807530000000
0!
0'
0/
#807540000000
#807550000000
1!
1'
1/
#807560000000
0!
0'
0/
#807570000000
1!
1'
1/
#807580000000
0!
1"
0'
1(
0/
10
#807590000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#807600000000
0!
0'
0/
#807610000000
1!
1'
1/
#807620000000
0!
0'
0/
#807630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#807640000000
0!
0'
0/
#807650000000
1!
1'
1/
#807660000000
0!
1"
0'
1(
0/
10
#807670000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#807680000000
0!
1$
0'
1+
0/
#807690000000
1!
1'
1/
#807700000000
0!
0'
0/
#807710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#807720000000
0!
0'
0/
#807730000000
1!
1'
1/
#807740000000
0!
0'
0/
#807750000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#807760000000
0!
0'
0/
#807770000000
1!
1'
1/
#807780000000
0!
0'
0/
#807790000000
1!
1'
1/
#807800000000
0!
0'
0/
#807810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#807820000000
0!
0'
0/
#807830000000
1!
1'
1/
#807840000000
0!
0'
0/
#807850000000
1!
1'
1/
#807860000000
0!
0'
0/
#807870000000
1!
1'
1/
#807880000000
0!
0'
0/
#807890000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#807900000000
0!
0'
0/
#807910000000
1!
1'
1/
#807920000000
0!
0'
0/
#807930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#807940000000
0!
0'
0/
#807950000000
1!
1'
1/
#807960000000
0!
0'
0/
#807970000000
#807980000000
1!
1'
1/
#807990000000
0!
0'
0/
#808000000000
1!
1'
1/
#808010000000
0!
1"
0'
1(
0/
10
#808020000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#808030000000
0!
0'
0/
#808040000000
1!
1'
1/
#808050000000
0!
0'
0/
#808060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#808070000000
0!
0'
0/
#808080000000
1!
1'
1/
#808090000000
0!
1"
0'
1(
0/
10
#808100000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#808110000000
0!
1$
0'
1+
0/
#808120000000
1!
1'
1/
#808130000000
0!
0'
0/
#808140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#808150000000
0!
0'
0/
#808160000000
1!
1'
1/
#808170000000
0!
0'
0/
#808180000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#808190000000
0!
0'
0/
#808200000000
1!
1'
1/
#808210000000
0!
0'
0/
#808220000000
1!
1'
1/
#808230000000
0!
0'
0/
#808240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#808250000000
0!
0'
0/
#808260000000
1!
1'
1/
#808270000000
0!
0'
0/
#808280000000
1!
1'
1/
#808290000000
0!
0'
0/
#808300000000
1!
1'
1/
#808310000000
0!
0'
0/
#808320000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#808330000000
0!
0'
0/
#808340000000
1!
1'
1/
#808350000000
0!
0'
0/
#808360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#808370000000
0!
0'
0/
#808380000000
1!
1'
1/
#808390000000
0!
0'
0/
#808400000000
#808410000000
1!
1'
1/
#808420000000
0!
0'
0/
#808430000000
1!
1'
1/
#808440000000
0!
1"
0'
1(
0/
10
#808450000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#808460000000
0!
0'
0/
#808470000000
1!
1'
1/
#808480000000
0!
0'
0/
#808490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#808500000000
0!
0'
0/
#808510000000
1!
1'
1/
#808520000000
0!
1"
0'
1(
0/
10
#808530000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#808540000000
0!
1$
0'
1+
0/
#808550000000
1!
1'
1/
#808560000000
0!
0'
0/
#808570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#808580000000
0!
0'
0/
#808590000000
1!
1'
1/
#808600000000
0!
0'
0/
#808610000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#808620000000
0!
0'
0/
#808630000000
1!
1'
1/
#808640000000
0!
0'
0/
#808650000000
1!
1'
1/
#808660000000
0!
0'
0/
#808670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#808680000000
0!
0'
0/
#808690000000
1!
1'
1/
#808700000000
0!
0'
0/
#808710000000
1!
1'
1/
#808720000000
0!
0'
0/
#808730000000
1!
1'
1/
#808740000000
0!
0'
0/
#808750000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#808760000000
0!
0'
0/
#808770000000
1!
1'
1/
#808780000000
0!
0'
0/
#808790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#808800000000
0!
0'
0/
#808810000000
1!
1'
1/
#808820000000
0!
0'
0/
#808830000000
#808840000000
1!
1'
1/
#808850000000
0!
0'
0/
#808860000000
1!
1'
1/
#808870000000
0!
1"
0'
1(
0/
10
#808880000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#808890000000
0!
0'
0/
#808900000000
1!
1'
1/
#808910000000
0!
0'
0/
#808920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#808930000000
0!
0'
0/
#808940000000
1!
1'
1/
#808950000000
0!
1"
0'
1(
0/
10
#808960000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#808970000000
0!
1$
0'
1+
0/
#808980000000
1!
1'
1/
#808990000000
0!
0'
0/
#809000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#809010000000
0!
0'
0/
#809020000000
1!
1'
1/
#809030000000
0!
0'
0/
#809040000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#809050000000
0!
0'
0/
#809060000000
1!
1'
1/
#809070000000
0!
0'
0/
#809080000000
1!
1'
1/
#809090000000
0!
0'
0/
#809100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#809110000000
0!
0'
0/
#809120000000
1!
1'
1/
#809130000000
0!
0'
0/
#809140000000
1!
1'
1/
#809150000000
0!
0'
0/
#809160000000
1!
1'
1/
#809170000000
0!
0'
0/
#809180000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#809190000000
0!
0'
0/
#809200000000
1!
1'
1/
#809210000000
0!
0'
0/
#809220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#809230000000
0!
0'
0/
#809240000000
1!
1'
1/
#809250000000
0!
0'
0/
#809260000000
#809270000000
1!
1'
1/
#809280000000
0!
0'
0/
#809290000000
1!
1'
1/
#809300000000
0!
1"
0'
1(
0/
10
#809310000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#809320000000
0!
0'
0/
#809330000000
1!
1'
1/
#809340000000
0!
0'
0/
#809350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#809360000000
0!
0'
0/
#809370000000
1!
1'
1/
#809380000000
0!
1"
0'
1(
0/
10
#809390000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#809400000000
0!
1$
0'
1+
0/
#809410000000
1!
1'
1/
#809420000000
0!
0'
0/
#809430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#809440000000
0!
0'
0/
#809450000000
1!
1'
1/
#809460000000
0!
0'
0/
#809470000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#809480000000
0!
0'
0/
#809490000000
1!
1'
1/
#809500000000
0!
0'
0/
#809510000000
1!
1'
1/
#809520000000
0!
0'
0/
#809530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#809540000000
0!
0'
0/
#809550000000
1!
1'
1/
#809560000000
0!
0'
0/
#809570000000
1!
1'
1/
#809580000000
0!
0'
0/
#809590000000
1!
1'
1/
#809600000000
0!
0'
0/
#809610000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#809620000000
0!
0'
0/
#809630000000
1!
1'
1/
#809640000000
0!
0'
0/
#809650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#809660000000
0!
0'
0/
#809670000000
1!
1'
1/
#809680000000
0!
0'
0/
#809690000000
#809700000000
1!
1'
1/
#809710000000
0!
0'
0/
#809720000000
1!
1'
1/
#809730000000
0!
1"
0'
1(
0/
10
#809740000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#809750000000
0!
0'
0/
#809760000000
1!
1'
1/
#809770000000
0!
0'
0/
#809780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#809790000000
0!
0'
0/
#809800000000
1!
1'
1/
#809810000000
0!
1"
0'
1(
0/
10
#809820000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#809830000000
0!
1$
0'
1+
0/
#809840000000
1!
1'
1/
#809850000000
0!
0'
0/
#809860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#809870000000
0!
0'
0/
#809880000000
1!
1'
1/
#809890000000
0!
0'
0/
#809900000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#809910000000
0!
0'
0/
#809920000000
1!
1'
1/
#809930000000
0!
0'
0/
#809940000000
1!
1'
1/
#809950000000
0!
0'
0/
#809960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#809970000000
0!
0'
0/
#809980000000
1!
1'
1/
#809990000000
0!
0'
0/
#810000000000
1!
1'
1/
#810010000000
0!
0'
0/
#810020000000
1!
1'
1/
#810030000000
0!
0'
0/
#810040000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#810050000000
0!
0'
0/
#810060000000
1!
1'
1/
#810070000000
0!
0'
0/
#810080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#810090000000
0!
0'
0/
#810100000000
1!
1'
1/
#810110000000
0!
0'
0/
#810120000000
#810130000000
1!
1'
1/
#810140000000
0!
0'
0/
#810150000000
1!
1'
1/
#810160000000
0!
1"
0'
1(
0/
10
#810170000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#810180000000
0!
0'
0/
#810190000000
1!
1'
1/
#810200000000
0!
0'
0/
#810210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#810220000000
0!
0'
0/
#810230000000
1!
1'
1/
#810240000000
0!
1"
0'
1(
0/
10
#810250000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#810260000000
0!
1$
0'
1+
0/
#810270000000
1!
1'
1/
#810280000000
0!
0'
0/
#810290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#810300000000
0!
0'
0/
#810310000000
1!
1'
1/
#810320000000
0!
0'
0/
#810330000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#810340000000
0!
0'
0/
#810350000000
1!
1'
1/
#810360000000
0!
0'
0/
#810370000000
1!
1'
1/
#810380000000
0!
0'
0/
#810390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#810400000000
0!
0'
0/
#810410000000
1!
1'
1/
#810420000000
0!
0'
0/
#810430000000
1!
1'
1/
#810440000000
0!
0'
0/
#810450000000
1!
1'
1/
#810460000000
0!
0'
0/
#810470000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#810480000000
0!
0'
0/
#810490000000
1!
1'
1/
#810500000000
0!
0'
0/
#810510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#810520000000
0!
0'
0/
#810530000000
1!
1'
1/
#810540000000
0!
0'
0/
#810550000000
#810560000000
1!
1'
1/
#810570000000
0!
0'
0/
#810580000000
1!
1'
1/
#810590000000
0!
1"
0'
1(
0/
10
#810600000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#810610000000
0!
0'
0/
#810620000000
1!
1'
1/
#810630000000
0!
0'
0/
#810640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#810650000000
0!
0'
0/
#810660000000
1!
1'
1/
#810670000000
0!
1"
0'
1(
0/
10
#810680000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#810690000000
0!
1$
0'
1+
0/
#810700000000
1!
1'
1/
#810710000000
0!
0'
0/
#810720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#810730000000
0!
0'
0/
#810740000000
1!
1'
1/
#810750000000
0!
0'
0/
#810760000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#810770000000
0!
0'
0/
#810780000000
1!
1'
1/
#810790000000
0!
0'
0/
#810800000000
1!
1'
1/
#810810000000
0!
0'
0/
#810820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#810830000000
0!
0'
0/
#810840000000
1!
1'
1/
#810850000000
0!
0'
0/
#810860000000
1!
1'
1/
#810870000000
0!
0'
0/
#810880000000
1!
1'
1/
#810890000000
0!
0'
0/
#810900000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#810910000000
0!
0'
0/
#810920000000
1!
1'
1/
#810930000000
0!
0'
0/
#810940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#810950000000
0!
0'
0/
#810960000000
1!
1'
1/
#810970000000
0!
0'
0/
#810980000000
#810990000000
1!
1'
1/
#811000000000
0!
0'
0/
#811010000000
1!
1'
1/
#811020000000
0!
1"
0'
1(
0/
10
#811030000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#811040000000
0!
0'
0/
#811050000000
1!
1'
1/
#811060000000
0!
0'
0/
#811070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#811080000000
0!
0'
0/
#811090000000
1!
1'
1/
#811100000000
0!
1"
0'
1(
0/
10
#811110000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#811120000000
0!
1$
0'
1+
0/
#811130000000
1!
1'
1/
#811140000000
0!
0'
0/
#811150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#811160000000
0!
0'
0/
#811170000000
1!
1'
1/
#811180000000
0!
0'
0/
#811190000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#811200000000
0!
0'
0/
#811210000000
1!
1'
1/
#811220000000
0!
0'
0/
#811230000000
1!
1'
1/
#811240000000
0!
0'
0/
#811250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#811260000000
0!
0'
0/
#811270000000
1!
1'
1/
#811280000000
0!
0'
0/
#811290000000
1!
1'
1/
#811300000000
0!
0'
0/
#811310000000
1!
1'
1/
#811320000000
0!
0'
0/
#811330000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#811340000000
0!
0'
0/
#811350000000
1!
1'
1/
#811360000000
0!
0'
0/
#811370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#811380000000
0!
0'
0/
#811390000000
1!
1'
1/
#811400000000
0!
0'
0/
#811410000000
#811420000000
1!
1'
1/
#811430000000
0!
0'
0/
#811440000000
1!
1'
1/
#811450000000
0!
1"
0'
1(
0/
10
#811460000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#811470000000
0!
0'
0/
#811480000000
1!
1'
1/
#811490000000
0!
0'
0/
#811500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#811510000000
0!
0'
0/
#811520000000
1!
1'
1/
#811530000000
0!
1"
0'
1(
0/
10
#811540000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#811550000000
0!
1$
0'
1+
0/
#811560000000
1!
1'
1/
#811570000000
0!
0'
0/
#811580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#811590000000
0!
0'
0/
#811600000000
1!
1'
1/
#811610000000
0!
0'
0/
#811620000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#811630000000
0!
0'
0/
#811640000000
1!
1'
1/
#811650000000
0!
0'
0/
#811660000000
1!
1'
1/
#811670000000
0!
0'
0/
#811680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#811690000000
0!
0'
0/
#811700000000
1!
1'
1/
#811710000000
0!
0'
0/
#811720000000
1!
1'
1/
#811730000000
0!
0'
0/
#811740000000
1!
1'
1/
#811750000000
0!
0'
0/
#811760000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#811770000000
0!
0'
0/
#811780000000
1!
1'
1/
#811790000000
0!
0'
0/
#811800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#811810000000
0!
0'
0/
#811820000000
1!
1'
1/
#811830000000
0!
0'
0/
#811840000000
#811850000000
1!
1'
1/
#811860000000
0!
0'
0/
#811870000000
1!
1'
1/
#811880000000
0!
1"
0'
1(
0/
10
#811890000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#811900000000
0!
0'
0/
#811910000000
1!
1'
1/
#811920000000
0!
0'
0/
#811930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#811940000000
0!
0'
0/
#811950000000
1!
1'
1/
#811960000000
0!
1"
0'
1(
0/
10
#811970000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#811980000000
0!
1$
0'
1+
0/
#811990000000
1!
1'
1/
#812000000000
0!
0'
0/
#812010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#812020000000
0!
0'
0/
#812030000000
1!
1'
1/
#812040000000
0!
0'
0/
#812050000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#812060000000
0!
0'
0/
#812070000000
1!
1'
1/
#812080000000
0!
0'
0/
#812090000000
1!
1'
1/
#812100000000
0!
0'
0/
#812110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#812120000000
0!
0'
0/
#812130000000
1!
1'
1/
#812140000000
0!
0'
0/
#812150000000
1!
1'
1/
#812160000000
0!
0'
0/
#812170000000
1!
1'
1/
#812180000000
0!
0'
0/
#812190000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#812200000000
0!
0'
0/
#812210000000
1!
1'
1/
#812220000000
0!
0'
0/
#812230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#812240000000
0!
0'
0/
#812250000000
1!
1'
1/
#812260000000
0!
0'
0/
#812270000000
#812280000000
1!
1'
1/
#812290000000
0!
0'
0/
#812300000000
1!
1'
1/
#812310000000
0!
1"
0'
1(
0/
10
#812320000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#812330000000
0!
0'
0/
#812340000000
1!
1'
1/
#812350000000
0!
0'
0/
#812360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#812370000000
0!
0'
0/
#812380000000
1!
1'
1/
#812390000000
0!
1"
0'
1(
0/
10
#812400000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#812410000000
0!
1$
0'
1+
0/
#812420000000
1!
1'
1/
#812430000000
0!
0'
0/
#812440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#812450000000
0!
0'
0/
#812460000000
1!
1'
1/
#812470000000
0!
0'
0/
#812480000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#812490000000
0!
0'
0/
#812500000000
1!
1'
1/
#812510000000
0!
0'
0/
#812520000000
1!
1'
1/
#812530000000
0!
0'
0/
#812540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#812550000000
0!
0'
0/
#812560000000
1!
1'
1/
#812570000000
0!
0'
0/
#812580000000
1!
1'
1/
#812590000000
0!
0'
0/
#812600000000
1!
1'
1/
#812610000000
0!
0'
0/
#812620000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#812630000000
0!
0'
0/
#812640000000
1!
1'
1/
#812650000000
0!
0'
0/
#812660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#812670000000
0!
0'
0/
#812680000000
1!
1'
1/
#812690000000
0!
0'
0/
#812700000000
#812710000000
1!
1'
1/
#812720000000
0!
0'
0/
#812730000000
1!
1'
1/
#812740000000
0!
1"
0'
1(
0/
10
#812750000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#812760000000
0!
0'
0/
#812770000000
1!
1'
1/
#812780000000
0!
0'
0/
#812790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#812800000000
0!
0'
0/
#812810000000
1!
1'
1/
#812820000000
0!
1"
0'
1(
0/
10
#812830000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#812840000000
0!
1$
0'
1+
0/
#812850000000
1!
1'
1/
#812860000000
0!
0'
0/
#812870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#812880000000
0!
0'
0/
#812890000000
1!
1'
1/
#812900000000
0!
0'
0/
#812910000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#812920000000
0!
0'
0/
#812930000000
1!
1'
1/
#812940000000
0!
0'
0/
#812950000000
1!
1'
1/
#812960000000
0!
0'
0/
#812970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#812980000000
0!
0'
0/
#812990000000
1!
1'
1/
#813000000000
0!
0'
0/
#813010000000
1!
1'
1/
#813020000000
0!
0'
0/
#813030000000
1!
1'
1/
#813040000000
0!
0'
0/
#813050000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#813060000000
0!
0'
0/
#813070000000
1!
1'
1/
#813080000000
0!
0'
0/
#813090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#813100000000
0!
0'
0/
#813110000000
1!
1'
1/
#813120000000
0!
0'
0/
#813130000000
#813140000000
1!
1'
1/
#813150000000
0!
0'
0/
#813160000000
1!
1'
1/
#813170000000
0!
1"
0'
1(
0/
10
#813180000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#813190000000
0!
0'
0/
#813200000000
1!
1'
1/
#813210000000
0!
0'
0/
#813220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#813230000000
0!
0'
0/
#813240000000
1!
1'
1/
#813250000000
0!
1"
0'
1(
0/
10
#813260000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#813270000000
0!
1$
0'
1+
0/
#813280000000
1!
1'
1/
#813290000000
0!
0'
0/
#813300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#813310000000
0!
0'
0/
#813320000000
1!
1'
1/
#813330000000
0!
0'
0/
#813340000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#813350000000
0!
0'
0/
#813360000000
1!
1'
1/
#813370000000
0!
0'
0/
#813380000000
1!
1'
1/
#813390000000
0!
0'
0/
#813400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#813410000000
0!
0'
0/
#813420000000
1!
1'
1/
#813430000000
0!
0'
0/
#813440000000
1!
1'
1/
#813450000000
0!
0'
0/
#813460000000
1!
1'
1/
#813470000000
0!
0'
0/
#813480000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#813490000000
0!
0'
0/
#813500000000
1!
1'
1/
#813510000000
0!
0'
0/
#813520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#813530000000
0!
0'
0/
#813540000000
1!
1'
1/
#813550000000
0!
0'
0/
#813560000000
#813570000000
1!
1'
1/
#813580000000
0!
0'
0/
#813590000000
1!
1'
1/
#813600000000
0!
1"
0'
1(
0/
10
#813610000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#813620000000
0!
0'
0/
#813630000000
1!
1'
1/
#813640000000
0!
0'
0/
#813650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#813660000000
0!
0'
0/
#813670000000
1!
1'
1/
#813680000000
0!
1"
0'
1(
0/
10
#813690000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#813700000000
0!
1$
0'
1+
0/
#813710000000
1!
1'
1/
#813720000000
0!
0'
0/
#813730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#813740000000
0!
0'
0/
#813750000000
1!
1'
1/
#813760000000
0!
0'
0/
#813770000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#813780000000
0!
0'
0/
#813790000000
1!
1'
1/
#813800000000
0!
0'
0/
#813810000000
1!
1'
1/
#813820000000
0!
0'
0/
#813830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#813840000000
0!
0'
0/
#813850000000
1!
1'
1/
#813860000000
0!
0'
0/
#813870000000
1!
1'
1/
#813880000000
0!
0'
0/
#813890000000
1!
1'
1/
#813900000000
0!
0'
0/
#813910000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#813920000000
0!
0'
0/
#813930000000
1!
1'
1/
#813940000000
0!
0'
0/
#813950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#813960000000
0!
0'
0/
#813970000000
1!
1'
1/
#813980000000
0!
0'
0/
#813990000000
#814000000000
1!
1'
1/
#814010000000
0!
0'
0/
#814020000000
1!
1'
1/
#814030000000
0!
1"
0'
1(
0/
10
#814040000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#814050000000
0!
0'
0/
#814060000000
1!
1'
1/
#814070000000
0!
0'
0/
#814080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#814090000000
0!
0'
0/
#814100000000
1!
1'
1/
#814110000000
0!
1"
0'
1(
0/
10
#814120000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#814130000000
0!
1$
0'
1+
0/
#814140000000
1!
1'
1/
#814150000000
0!
0'
0/
#814160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#814170000000
0!
0'
0/
#814180000000
1!
1'
1/
#814190000000
0!
0'
0/
#814200000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#814210000000
0!
0'
0/
#814220000000
1!
1'
1/
#814230000000
0!
0'
0/
#814240000000
1!
1'
1/
#814250000000
0!
0'
0/
#814260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#814270000000
0!
0'
0/
#814280000000
1!
1'
1/
#814290000000
0!
0'
0/
#814300000000
1!
1'
1/
#814310000000
0!
0'
0/
#814320000000
1!
1'
1/
#814330000000
0!
0'
0/
#814340000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#814350000000
0!
0'
0/
#814360000000
1!
1'
1/
#814370000000
0!
0'
0/
#814380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#814390000000
0!
0'
0/
#814400000000
1!
1'
1/
#814410000000
0!
0'
0/
#814420000000
#814430000000
1!
1'
1/
#814440000000
0!
0'
0/
#814450000000
1!
1'
1/
#814460000000
0!
1"
0'
1(
0/
10
#814470000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#814480000000
0!
0'
0/
#814490000000
1!
1'
1/
#814500000000
0!
0'
0/
#814510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#814520000000
0!
0'
0/
#814530000000
1!
1'
1/
#814540000000
0!
1"
0'
1(
0/
10
#814550000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#814560000000
0!
1$
0'
1+
0/
#814570000000
1!
1'
1/
#814580000000
0!
0'
0/
#814590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#814600000000
0!
0'
0/
#814610000000
1!
1'
1/
#814620000000
0!
0'
0/
#814630000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#814640000000
0!
0'
0/
#814650000000
1!
1'
1/
#814660000000
0!
0'
0/
#814670000000
1!
1'
1/
#814680000000
0!
0'
0/
#814690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#814700000000
0!
0'
0/
#814710000000
1!
1'
1/
#814720000000
0!
0'
0/
#814730000000
1!
1'
1/
#814740000000
0!
0'
0/
#814750000000
1!
1'
1/
#814760000000
0!
0'
0/
#814770000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#814780000000
0!
0'
0/
#814790000000
1!
1'
1/
#814800000000
0!
0'
0/
#814810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#814820000000
0!
0'
0/
#814830000000
1!
1'
1/
#814840000000
0!
0'
0/
#814850000000
#814860000000
1!
1'
1/
#814870000000
0!
0'
0/
#814880000000
1!
1'
1/
#814890000000
0!
1"
0'
1(
0/
10
#814900000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#814910000000
0!
0'
0/
#814920000000
1!
1'
1/
#814930000000
0!
0'
0/
#814940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#814950000000
0!
0'
0/
#814960000000
1!
1'
1/
#814970000000
0!
1"
0'
1(
0/
10
#814980000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#814990000000
0!
1$
0'
1+
0/
#815000000000
1!
1'
1/
#815010000000
0!
0'
0/
#815020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#815030000000
0!
0'
0/
#815040000000
1!
1'
1/
#815050000000
0!
0'
0/
#815060000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#815070000000
0!
0'
0/
#815080000000
1!
1'
1/
#815090000000
0!
0'
0/
#815100000000
1!
1'
1/
#815110000000
0!
0'
0/
#815120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#815130000000
0!
0'
0/
#815140000000
1!
1'
1/
#815150000000
0!
0'
0/
#815160000000
1!
1'
1/
#815170000000
0!
0'
0/
#815180000000
1!
1'
1/
#815190000000
0!
0'
0/
#815200000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#815210000000
0!
0'
0/
#815220000000
1!
1'
1/
#815230000000
0!
0'
0/
#815240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#815250000000
0!
0'
0/
#815260000000
1!
1'
1/
#815270000000
0!
0'
0/
#815280000000
#815290000000
1!
1'
1/
#815300000000
0!
0'
0/
#815310000000
1!
1'
1/
#815320000000
0!
1"
0'
1(
0/
10
#815330000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#815340000000
0!
0'
0/
#815350000000
1!
1'
1/
#815360000000
0!
0'
0/
#815370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#815380000000
0!
0'
0/
#815390000000
1!
1'
1/
#815400000000
0!
1"
0'
1(
0/
10
#815410000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#815420000000
0!
1$
0'
1+
0/
#815430000000
1!
1'
1/
#815440000000
0!
0'
0/
#815450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#815460000000
0!
0'
0/
#815470000000
1!
1'
1/
#815480000000
0!
0'
0/
#815490000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#815500000000
0!
0'
0/
#815510000000
1!
1'
1/
#815520000000
0!
0'
0/
#815530000000
1!
1'
1/
#815540000000
0!
0'
0/
#815550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#815560000000
0!
0'
0/
#815570000000
1!
1'
1/
#815580000000
0!
0'
0/
#815590000000
1!
1'
1/
#815600000000
0!
0'
0/
#815610000000
1!
1'
1/
#815620000000
0!
0'
0/
#815630000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#815640000000
0!
0'
0/
#815650000000
1!
1'
1/
#815660000000
0!
0'
0/
#815670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#815680000000
0!
0'
0/
#815690000000
1!
1'
1/
#815700000000
0!
0'
0/
#815710000000
#815720000000
1!
1'
1/
#815730000000
0!
0'
0/
#815740000000
1!
1'
1/
#815750000000
0!
1"
0'
1(
0/
10
#815760000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#815770000000
0!
0'
0/
#815780000000
1!
1'
1/
#815790000000
0!
0'
0/
#815800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#815810000000
0!
0'
0/
#815820000000
1!
1'
1/
#815830000000
0!
1"
0'
1(
0/
10
#815840000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#815850000000
0!
1$
0'
1+
0/
#815860000000
1!
1'
1/
#815870000000
0!
0'
0/
#815880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#815890000000
0!
0'
0/
#815900000000
1!
1'
1/
#815910000000
0!
0'
0/
#815920000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#815930000000
0!
0'
0/
#815940000000
1!
1'
1/
#815950000000
0!
0'
0/
#815960000000
1!
1'
1/
#815970000000
0!
0'
0/
#815980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#815990000000
0!
0'
0/
#816000000000
1!
1'
1/
#816010000000
0!
0'
0/
#816020000000
1!
1'
1/
#816030000000
0!
0'
0/
#816040000000
1!
1'
1/
#816050000000
0!
0'
0/
#816060000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#816070000000
0!
0'
0/
#816080000000
1!
1'
1/
#816090000000
0!
0'
0/
#816100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#816110000000
0!
0'
0/
#816120000000
1!
1'
1/
#816130000000
0!
0'
0/
#816140000000
#816150000000
1!
1'
1/
#816160000000
0!
0'
0/
#816170000000
1!
1'
1/
#816180000000
0!
1"
0'
1(
0/
10
#816190000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#816200000000
0!
0'
0/
#816210000000
1!
1'
1/
#816220000000
0!
0'
0/
#816230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#816240000000
0!
0'
0/
#816250000000
1!
1'
1/
#816260000000
0!
1"
0'
1(
0/
10
#816270000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#816280000000
0!
1$
0'
1+
0/
#816290000000
1!
1'
1/
#816300000000
0!
0'
0/
#816310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#816320000000
0!
0'
0/
#816330000000
1!
1'
1/
#816340000000
0!
0'
0/
#816350000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#816360000000
0!
0'
0/
#816370000000
1!
1'
1/
#816380000000
0!
0'
0/
#816390000000
1!
1'
1/
#816400000000
0!
0'
0/
#816410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#816420000000
0!
0'
0/
#816430000000
1!
1'
1/
#816440000000
0!
0'
0/
#816450000000
1!
1'
1/
#816460000000
0!
0'
0/
#816470000000
1!
1'
1/
#816480000000
0!
0'
0/
#816490000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#816500000000
0!
0'
0/
#816510000000
1!
1'
1/
#816520000000
0!
0'
0/
#816530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#816540000000
0!
0'
0/
#816550000000
1!
1'
1/
#816560000000
0!
0'
0/
#816570000000
#816580000000
1!
1'
1/
#816590000000
0!
0'
0/
#816600000000
1!
1'
1/
#816610000000
0!
1"
0'
1(
0/
10
#816620000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#816630000000
0!
0'
0/
#816640000000
1!
1'
1/
#816650000000
0!
0'
0/
#816660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#816670000000
0!
0'
0/
#816680000000
1!
1'
1/
#816690000000
0!
1"
0'
1(
0/
10
#816700000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#816710000000
0!
1$
0'
1+
0/
#816720000000
1!
1'
1/
#816730000000
0!
0'
0/
#816740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#816750000000
0!
0'
0/
#816760000000
1!
1'
1/
#816770000000
0!
0'
0/
#816780000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#816790000000
0!
0'
0/
#816800000000
1!
1'
1/
#816810000000
0!
0'
0/
#816820000000
1!
1'
1/
#816830000000
0!
0'
0/
#816840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#816850000000
0!
0'
0/
#816860000000
1!
1'
1/
#816870000000
0!
0'
0/
#816880000000
1!
1'
1/
#816890000000
0!
0'
0/
#816900000000
1!
1'
1/
#816910000000
0!
0'
0/
#816920000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#816930000000
0!
0'
0/
#816940000000
1!
1'
1/
#816950000000
0!
0'
0/
#816960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#816970000000
0!
0'
0/
#816980000000
1!
1'
1/
#816990000000
0!
0'
0/
#817000000000
#817010000000
1!
1'
1/
#817020000000
0!
0'
0/
#817030000000
1!
1'
1/
#817040000000
0!
1"
0'
1(
0/
10
#817050000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#817060000000
0!
0'
0/
#817070000000
1!
1'
1/
#817080000000
0!
0'
0/
#817090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#817100000000
0!
0'
0/
#817110000000
1!
1'
1/
#817120000000
0!
1"
0'
1(
0/
10
#817130000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#817140000000
0!
1$
0'
1+
0/
#817150000000
1!
1'
1/
#817160000000
0!
0'
0/
#817170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#817180000000
0!
0'
0/
#817190000000
1!
1'
1/
#817200000000
0!
0'
0/
#817210000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#817220000000
0!
0'
0/
#817230000000
1!
1'
1/
#817240000000
0!
0'
0/
#817250000000
1!
1'
1/
#817260000000
0!
0'
0/
#817270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#817280000000
0!
0'
0/
#817290000000
1!
1'
1/
#817300000000
0!
0'
0/
#817310000000
1!
1'
1/
#817320000000
0!
0'
0/
#817330000000
1!
1'
1/
#817340000000
0!
0'
0/
#817350000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#817360000000
0!
0'
0/
#817370000000
1!
1'
1/
#817380000000
0!
0'
0/
#817390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#817400000000
0!
0'
0/
#817410000000
1!
1'
1/
#817420000000
0!
0'
0/
#817430000000
#817440000000
1!
1'
1/
#817450000000
0!
0'
0/
#817460000000
1!
1'
1/
#817470000000
0!
1"
0'
1(
0/
10
#817480000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#817490000000
0!
0'
0/
#817500000000
1!
1'
1/
#817510000000
0!
0'
0/
#817520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#817530000000
0!
0'
0/
#817540000000
1!
1'
1/
#817550000000
0!
1"
0'
1(
0/
10
#817560000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#817570000000
0!
1$
0'
1+
0/
#817580000000
1!
1'
1/
#817590000000
0!
0'
0/
#817600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#817610000000
0!
0'
0/
#817620000000
1!
1'
1/
#817630000000
0!
0'
0/
#817640000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#817650000000
0!
0'
0/
#817660000000
1!
1'
1/
#817670000000
0!
0'
0/
#817680000000
1!
1'
1/
#817690000000
0!
0'
0/
#817700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#817710000000
0!
0'
0/
#817720000000
1!
1'
1/
#817730000000
0!
0'
0/
#817740000000
1!
1'
1/
#817750000000
0!
0'
0/
#817760000000
1!
1'
1/
#817770000000
0!
0'
0/
#817780000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#817790000000
0!
0'
0/
#817800000000
1!
1'
1/
#817810000000
0!
0'
0/
#817820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#817830000000
0!
0'
0/
#817840000000
1!
1'
1/
#817850000000
0!
0'
0/
#817860000000
#817870000000
1!
1'
1/
#817880000000
0!
0'
0/
#817890000000
1!
1'
1/
#817900000000
0!
1"
0'
1(
0/
10
#817910000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#817920000000
0!
0'
0/
#817930000000
1!
1'
1/
#817940000000
0!
0'
0/
#817950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#817960000000
0!
0'
0/
#817970000000
1!
1'
1/
#817980000000
0!
1"
0'
1(
0/
10
#817990000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#818000000000
0!
1$
0'
1+
0/
#818010000000
1!
1'
1/
#818020000000
0!
0'
0/
#818030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#818040000000
0!
0'
0/
#818050000000
1!
1'
1/
#818060000000
0!
0'
0/
#818070000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#818080000000
0!
0'
0/
#818090000000
1!
1'
1/
#818100000000
0!
0'
0/
#818110000000
1!
1'
1/
#818120000000
0!
0'
0/
#818130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#818140000000
0!
0'
0/
#818150000000
1!
1'
1/
#818160000000
0!
0'
0/
#818170000000
1!
1'
1/
#818180000000
0!
0'
0/
#818190000000
1!
1'
1/
#818200000000
0!
0'
0/
#818210000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#818220000000
0!
0'
0/
#818230000000
1!
1'
1/
#818240000000
0!
0'
0/
#818250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#818260000000
0!
0'
0/
#818270000000
1!
1'
1/
#818280000000
0!
0'
0/
#818290000000
#818300000000
1!
1'
1/
#818310000000
0!
0'
0/
#818320000000
1!
1'
1/
#818330000000
0!
1"
0'
1(
0/
10
#818340000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#818350000000
0!
0'
0/
#818360000000
1!
1'
1/
#818370000000
0!
0'
0/
#818380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#818390000000
0!
0'
0/
#818400000000
1!
1'
1/
#818410000000
0!
1"
0'
1(
0/
10
#818420000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#818430000000
0!
1$
0'
1+
0/
#818440000000
1!
1'
1/
#818450000000
0!
0'
0/
#818460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#818470000000
0!
0'
0/
#818480000000
1!
1'
1/
#818490000000
0!
0'
0/
#818500000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#818510000000
0!
0'
0/
#818520000000
1!
1'
1/
#818530000000
0!
0'
0/
#818540000000
1!
1'
1/
#818550000000
0!
0'
0/
#818560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#818570000000
0!
0'
0/
#818580000000
1!
1'
1/
#818590000000
0!
0'
0/
#818600000000
1!
1'
1/
#818610000000
0!
0'
0/
#818620000000
1!
1'
1/
#818630000000
0!
0'
0/
#818640000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#818650000000
0!
0'
0/
#818660000000
1!
1'
1/
#818670000000
0!
0'
0/
#818680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#818690000000
0!
0'
0/
#818700000000
1!
1'
1/
#818710000000
0!
0'
0/
#818720000000
#818730000000
1!
1'
1/
#818740000000
0!
0'
0/
#818750000000
1!
1'
1/
#818760000000
0!
1"
0'
1(
0/
10
#818770000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#818780000000
0!
0'
0/
#818790000000
1!
1'
1/
#818800000000
0!
0'
0/
#818810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#818820000000
0!
0'
0/
#818830000000
1!
1'
1/
#818840000000
0!
1"
0'
1(
0/
10
#818850000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#818860000000
0!
1$
0'
1+
0/
#818870000000
1!
1'
1/
#818880000000
0!
0'
0/
#818890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#818900000000
0!
0'
0/
#818910000000
1!
1'
1/
#818920000000
0!
0'
0/
#818930000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#818940000000
0!
0'
0/
#818950000000
1!
1'
1/
#818960000000
0!
0'
0/
#818970000000
1!
1'
1/
#818980000000
0!
0'
0/
#818990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#819000000000
0!
0'
0/
#819010000000
1!
1'
1/
#819020000000
0!
0'
0/
#819030000000
1!
1'
1/
#819040000000
0!
0'
0/
#819050000000
1!
1'
1/
#819060000000
0!
0'
0/
#819070000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#819080000000
0!
0'
0/
#819090000000
1!
1'
1/
#819100000000
0!
0'
0/
#819110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#819120000000
0!
0'
0/
#819130000000
1!
1'
1/
#819140000000
0!
0'
0/
#819150000000
#819160000000
1!
1'
1/
#819170000000
0!
0'
0/
#819180000000
1!
1'
1/
#819190000000
0!
1"
0'
1(
0/
10
#819200000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#819210000000
0!
0'
0/
#819220000000
1!
1'
1/
#819230000000
0!
0'
0/
#819240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#819250000000
0!
0'
0/
#819260000000
1!
1'
1/
#819270000000
0!
1"
0'
1(
0/
10
#819280000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#819290000000
0!
1$
0'
1+
0/
#819300000000
1!
1'
1/
#819310000000
0!
0'
0/
#819320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#819330000000
0!
0'
0/
#819340000000
1!
1'
1/
#819350000000
0!
0'
0/
#819360000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#819370000000
0!
0'
0/
#819380000000
1!
1'
1/
#819390000000
0!
0'
0/
#819400000000
1!
1'
1/
#819410000000
0!
0'
0/
#819420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#819430000000
0!
0'
0/
#819440000000
1!
1'
1/
#819450000000
0!
0'
0/
#819460000000
1!
1'
1/
#819470000000
0!
0'
0/
#819480000000
1!
1'
1/
#819490000000
0!
0'
0/
#819500000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#819510000000
0!
0'
0/
#819520000000
1!
1'
1/
#819530000000
0!
0'
0/
#819540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#819550000000
0!
0'
0/
#819560000000
1!
1'
1/
#819570000000
0!
0'
0/
#819580000000
#819590000000
1!
1'
1/
#819600000000
0!
0'
0/
#819610000000
1!
1'
1/
#819620000000
0!
1"
0'
1(
0/
10
#819630000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#819640000000
0!
0'
0/
#819650000000
1!
1'
1/
#819660000000
0!
0'
0/
#819670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#819680000000
0!
0'
0/
#819690000000
1!
1'
1/
#819700000000
0!
1"
0'
1(
0/
10
#819710000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#819720000000
0!
1$
0'
1+
0/
#819730000000
1!
1'
1/
#819740000000
0!
0'
0/
#819750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#819760000000
0!
0'
0/
#819770000000
1!
1'
1/
#819780000000
0!
0'
0/
#819790000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#819800000000
0!
0'
0/
#819810000000
1!
1'
1/
#819820000000
0!
0'
0/
#819830000000
1!
1'
1/
#819840000000
0!
0'
0/
#819850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#819860000000
0!
0'
0/
#819870000000
1!
1'
1/
#819880000000
0!
0'
0/
#819890000000
1!
1'
1/
#819900000000
0!
0'
0/
#819910000000
1!
1'
1/
#819920000000
0!
0'
0/
#819930000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#819940000000
0!
0'
0/
#819950000000
1!
1'
1/
#819960000000
0!
0'
0/
#819970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#819980000000
0!
0'
0/
#819990000000
1!
1'
1/
#820000000000
0!
0'
0/
#820010000000
#820020000000
1!
1'
1/
#820030000000
0!
0'
0/
#820040000000
1!
1'
1/
#820050000000
0!
1"
0'
1(
0/
10
#820060000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#820070000000
0!
0'
0/
#820080000000
1!
1'
1/
#820090000000
0!
0'
0/
#820100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#820110000000
0!
0'
0/
#820120000000
1!
1'
1/
#820130000000
0!
1"
0'
1(
0/
10
#820140000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#820150000000
0!
1$
0'
1+
0/
#820160000000
1!
1'
1/
#820170000000
0!
0'
0/
#820180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#820190000000
0!
0'
0/
#820200000000
1!
1'
1/
#820210000000
0!
0'
0/
#820220000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#820230000000
0!
0'
0/
#820240000000
1!
1'
1/
#820250000000
0!
0'
0/
#820260000000
1!
1'
1/
#820270000000
0!
0'
0/
#820280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#820290000000
0!
0'
0/
#820300000000
1!
1'
1/
#820310000000
0!
0'
0/
#820320000000
1!
1'
1/
#820330000000
0!
0'
0/
#820340000000
1!
1'
1/
#820350000000
0!
0'
0/
#820360000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#820370000000
0!
0'
0/
#820380000000
1!
1'
1/
#820390000000
0!
0'
0/
#820400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#820410000000
0!
0'
0/
#820420000000
1!
1'
1/
#820430000000
0!
0'
0/
#820440000000
#820450000000
1!
1'
1/
#820460000000
0!
0'
0/
#820470000000
1!
1'
1/
#820480000000
0!
1"
0'
1(
0/
10
#820490000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#820500000000
0!
0'
0/
#820510000000
1!
1'
1/
#820520000000
0!
0'
0/
#820530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#820540000000
0!
0'
0/
#820550000000
1!
1'
1/
#820560000000
0!
1"
0'
1(
0/
10
#820570000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#820580000000
0!
1$
0'
1+
0/
#820590000000
1!
1'
1/
#820600000000
0!
0'
0/
#820610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#820620000000
0!
0'
0/
#820630000000
1!
1'
1/
#820640000000
0!
0'
0/
#820650000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#820660000000
0!
0'
0/
#820670000000
1!
1'
1/
#820680000000
0!
0'
0/
#820690000000
1!
1'
1/
#820700000000
0!
0'
0/
#820710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#820720000000
0!
0'
0/
#820730000000
1!
1'
1/
#820740000000
0!
0'
0/
#820750000000
1!
1'
1/
#820760000000
0!
0'
0/
#820770000000
1!
1'
1/
#820780000000
0!
0'
0/
#820790000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#820800000000
0!
0'
0/
#820810000000
1!
1'
1/
#820820000000
0!
0'
0/
#820830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#820840000000
0!
0'
0/
#820850000000
1!
1'
1/
#820860000000
0!
0'
0/
#820870000000
#820880000000
1!
1'
1/
#820890000000
0!
0'
0/
#820900000000
1!
1'
1/
#820910000000
0!
1"
0'
1(
0/
10
#820920000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#820930000000
0!
0'
0/
#820940000000
1!
1'
1/
#820950000000
0!
0'
0/
#820960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#820970000000
0!
0'
0/
#820980000000
1!
1'
1/
#820990000000
0!
1"
0'
1(
0/
10
#821000000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#821010000000
0!
1$
0'
1+
0/
#821020000000
1!
1'
1/
#821030000000
0!
0'
0/
#821040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#821050000000
0!
0'
0/
#821060000000
1!
1'
1/
#821070000000
0!
0'
0/
#821080000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#821090000000
0!
0'
0/
#821100000000
1!
1'
1/
#821110000000
0!
0'
0/
#821120000000
1!
1'
1/
#821130000000
0!
0'
0/
#821140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#821150000000
0!
0'
0/
#821160000000
1!
1'
1/
#821170000000
0!
0'
0/
#821180000000
1!
1'
1/
#821190000000
0!
0'
0/
#821200000000
1!
1'
1/
#821210000000
0!
0'
0/
#821220000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#821230000000
0!
0'
0/
#821240000000
1!
1'
1/
#821250000000
0!
0'
0/
#821260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#821270000000
0!
0'
0/
#821280000000
1!
1'
1/
#821290000000
0!
0'
0/
#821300000000
#821310000000
1!
1'
1/
#821320000000
0!
0'
0/
#821330000000
1!
1'
1/
#821340000000
0!
1"
0'
1(
0/
10
#821350000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#821360000000
0!
0'
0/
#821370000000
1!
1'
1/
#821380000000
0!
0'
0/
#821390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#821400000000
0!
0'
0/
#821410000000
1!
1'
1/
#821420000000
0!
1"
0'
1(
0/
10
#821430000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#821440000000
0!
1$
0'
1+
0/
#821450000000
1!
1'
1/
#821460000000
0!
0'
0/
#821470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#821480000000
0!
0'
0/
#821490000000
1!
1'
1/
#821500000000
0!
0'
0/
#821510000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#821520000000
0!
0'
0/
#821530000000
1!
1'
1/
#821540000000
0!
0'
0/
#821550000000
1!
1'
1/
#821560000000
0!
0'
0/
#821570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#821580000000
0!
0'
0/
#821590000000
1!
1'
1/
#821600000000
0!
0'
0/
#821610000000
1!
1'
1/
#821620000000
0!
0'
0/
#821630000000
1!
1'
1/
#821640000000
0!
0'
0/
#821650000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#821660000000
0!
0'
0/
#821670000000
1!
1'
1/
#821680000000
0!
0'
0/
#821690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#821700000000
0!
0'
0/
#821710000000
1!
1'
1/
#821720000000
0!
0'
0/
#821730000000
#821740000000
1!
1'
1/
#821750000000
0!
0'
0/
#821760000000
1!
1'
1/
#821770000000
0!
1"
0'
1(
0/
10
#821780000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#821790000000
0!
0'
0/
#821800000000
1!
1'
1/
#821810000000
0!
0'
0/
#821820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#821830000000
0!
0'
0/
#821840000000
1!
1'
1/
#821850000000
0!
1"
0'
1(
0/
10
#821860000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#821870000000
0!
1$
0'
1+
0/
#821880000000
1!
1'
1/
#821890000000
0!
0'
0/
#821900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#821910000000
0!
0'
0/
#821920000000
1!
1'
1/
#821930000000
0!
0'
0/
#821940000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#821950000000
0!
0'
0/
#821960000000
1!
1'
1/
#821970000000
0!
0'
0/
#821980000000
1!
1'
1/
#821990000000
0!
0'
0/
#822000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#822010000000
0!
0'
0/
#822020000000
1!
1'
1/
#822030000000
0!
0'
0/
#822040000000
1!
1'
1/
#822050000000
0!
0'
0/
#822060000000
1!
1'
1/
#822070000000
0!
0'
0/
#822080000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#822090000000
0!
0'
0/
#822100000000
1!
1'
1/
#822110000000
0!
0'
0/
#822120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#822130000000
0!
0'
0/
#822140000000
1!
1'
1/
#822150000000
0!
0'
0/
#822160000000
#822170000000
1!
1'
1/
#822180000000
0!
0'
0/
#822190000000
1!
1'
1/
#822200000000
0!
1"
0'
1(
0/
10
#822210000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#822220000000
0!
0'
0/
#822230000000
1!
1'
1/
#822240000000
0!
0'
0/
#822250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#822260000000
0!
0'
0/
#822270000000
1!
1'
1/
#822280000000
0!
1"
0'
1(
0/
10
#822290000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#822300000000
0!
1$
0'
1+
0/
#822310000000
1!
1'
1/
#822320000000
0!
0'
0/
#822330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#822340000000
0!
0'
0/
#822350000000
1!
1'
1/
#822360000000
0!
0'
0/
#822370000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#822380000000
0!
0'
0/
#822390000000
1!
1'
1/
#822400000000
0!
0'
0/
#822410000000
1!
1'
1/
#822420000000
0!
0'
0/
#822430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#822440000000
0!
0'
0/
#822450000000
1!
1'
1/
#822460000000
0!
0'
0/
#822470000000
1!
1'
1/
#822480000000
0!
0'
0/
#822490000000
1!
1'
1/
#822500000000
0!
0'
0/
#822510000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#822520000000
0!
0'
0/
#822530000000
1!
1'
1/
#822540000000
0!
0'
0/
#822550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#822560000000
0!
0'
0/
#822570000000
1!
1'
1/
#822580000000
0!
0'
0/
#822590000000
#822600000000
1!
1'
1/
#822610000000
0!
0'
0/
#822620000000
1!
1'
1/
#822630000000
0!
1"
0'
1(
0/
10
#822640000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#822650000000
0!
0'
0/
#822660000000
1!
1'
1/
#822670000000
0!
0'
0/
#822680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#822690000000
0!
0'
0/
#822700000000
1!
1'
1/
#822710000000
0!
1"
0'
1(
0/
10
#822720000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#822730000000
0!
1$
0'
1+
0/
#822740000000
1!
1'
1/
#822750000000
0!
0'
0/
#822760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#822770000000
0!
0'
0/
#822780000000
1!
1'
1/
#822790000000
0!
0'
0/
#822800000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#822810000000
0!
0'
0/
#822820000000
1!
1'
1/
#822830000000
0!
0'
0/
#822840000000
1!
1'
1/
#822850000000
0!
0'
0/
#822860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#822870000000
0!
0'
0/
#822880000000
1!
1'
1/
#822890000000
0!
0'
0/
#822900000000
1!
1'
1/
#822910000000
0!
0'
0/
#822920000000
1!
1'
1/
#822930000000
0!
0'
0/
#822940000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#822950000000
0!
0'
0/
#822960000000
1!
1'
1/
#822970000000
0!
0'
0/
#822980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#822990000000
0!
0'
0/
#823000000000
1!
1'
1/
#823010000000
0!
0'
0/
#823020000000
#823030000000
1!
1'
1/
#823040000000
0!
0'
0/
#823050000000
1!
1'
1/
#823060000000
0!
1"
0'
1(
0/
10
#823070000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#823080000000
0!
0'
0/
#823090000000
1!
1'
1/
#823100000000
0!
0'
0/
#823110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#823120000000
0!
0'
0/
#823130000000
1!
1'
1/
#823140000000
0!
1"
0'
1(
0/
10
#823150000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#823160000000
0!
1$
0'
1+
0/
#823170000000
1!
1'
1/
#823180000000
0!
0'
0/
#823190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#823200000000
0!
0'
0/
#823210000000
1!
1'
1/
#823220000000
0!
0'
0/
#823230000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#823240000000
0!
0'
0/
#823250000000
1!
1'
1/
#823260000000
0!
0'
0/
#823270000000
1!
1'
1/
#823280000000
0!
0'
0/
#823290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#823300000000
0!
0'
0/
#823310000000
1!
1'
1/
#823320000000
0!
0'
0/
#823330000000
1!
1'
1/
#823340000000
0!
0'
0/
#823350000000
1!
1'
1/
#823360000000
0!
0'
0/
#823370000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#823380000000
0!
0'
0/
#823390000000
1!
1'
1/
#823400000000
0!
0'
0/
#823410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#823420000000
0!
0'
0/
#823430000000
1!
1'
1/
#823440000000
0!
0'
0/
#823450000000
#823460000000
1!
1'
1/
#823470000000
0!
0'
0/
#823480000000
1!
1'
1/
#823490000000
0!
1"
0'
1(
0/
10
#823500000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#823510000000
0!
0'
0/
#823520000000
1!
1'
1/
#823530000000
0!
0'
0/
#823540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#823550000000
0!
0'
0/
#823560000000
1!
1'
1/
#823570000000
0!
1"
0'
1(
0/
10
#823580000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#823590000000
0!
1$
0'
1+
0/
#823600000000
1!
1'
1/
#823610000000
0!
0'
0/
#823620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#823630000000
0!
0'
0/
#823640000000
1!
1'
1/
#823650000000
0!
0'
0/
#823660000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#823670000000
0!
0'
0/
#823680000000
1!
1'
1/
#823690000000
0!
0'
0/
#823700000000
1!
1'
1/
#823710000000
0!
0'
0/
#823720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#823730000000
0!
0'
0/
#823740000000
1!
1'
1/
#823750000000
0!
0'
0/
#823760000000
1!
1'
1/
#823770000000
0!
0'
0/
#823780000000
1!
1'
1/
#823790000000
0!
0'
0/
#823800000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#823810000000
0!
0'
0/
#823820000000
1!
1'
1/
#823830000000
0!
0'
0/
#823840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#823850000000
0!
0'
0/
#823860000000
1!
1'
1/
#823870000000
0!
0'
0/
#823880000000
#823890000000
1!
1'
1/
#823900000000
0!
0'
0/
#823910000000
1!
1'
1/
#823920000000
0!
1"
0'
1(
0/
10
#823930000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#823940000000
0!
0'
0/
#823950000000
1!
1'
1/
#823960000000
0!
0'
0/
#823970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#823980000000
0!
0'
0/
#823990000000
1!
1'
1/
#824000000000
0!
1"
0'
1(
0/
10
#824010000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#824020000000
0!
1$
0'
1+
0/
#824030000000
1!
1'
1/
#824040000000
0!
0'
0/
#824050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#824060000000
0!
0'
0/
#824070000000
1!
1'
1/
#824080000000
0!
0'
0/
#824090000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#824100000000
0!
0'
0/
#824110000000
1!
1'
1/
#824120000000
0!
0'
0/
#824130000000
1!
1'
1/
#824140000000
0!
0'
0/
#824150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#824160000000
0!
0'
0/
#824170000000
1!
1'
1/
#824180000000
0!
0'
0/
#824190000000
1!
1'
1/
#824200000000
0!
0'
0/
#824210000000
1!
1'
1/
#824220000000
0!
0'
0/
#824230000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#824240000000
0!
0'
0/
#824250000000
1!
1'
1/
#824260000000
0!
0'
0/
#824270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#824280000000
0!
0'
0/
#824290000000
1!
1'
1/
#824300000000
0!
0'
0/
#824310000000
#824320000000
1!
1'
1/
#824330000000
0!
0'
0/
#824340000000
1!
1'
1/
#824350000000
0!
1"
0'
1(
0/
10
#824360000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#824370000000
0!
0'
0/
#824380000000
1!
1'
1/
#824390000000
0!
0'
0/
#824400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#824410000000
0!
0'
0/
#824420000000
1!
1'
1/
#824430000000
0!
1"
0'
1(
0/
10
#824440000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#824450000000
0!
1$
0'
1+
0/
#824460000000
1!
1'
1/
#824470000000
0!
0'
0/
#824480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#824490000000
0!
0'
0/
#824500000000
1!
1'
1/
#824510000000
0!
0'
0/
#824520000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#824530000000
0!
0'
0/
#824540000000
1!
1'
1/
#824550000000
0!
0'
0/
#824560000000
1!
1'
1/
#824570000000
0!
0'
0/
#824580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#824590000000
0!
0'
0/
#824600000000
1!
1'
1/
#824610000000
0!
0'
0/
#824620000000
1!
1'
1/
#824630000000
0!
0'
0/
#824640000000
1!
1'
1/
#824650000000
0!
0'
0/
#824660000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#824670000000
0!
0'
0/
#824680000000
1!
1'
1/
#824690000000
0!
0'
0/
#824700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#824710000000
0!
0'
0/
#824720000000
1!
1'
1/
#824730000000
0!
0'
0/
#824740000000
#824750000000
1!
1'
1/
#824760000000
0!
0'
0/
#824770000000
1!
1'
1/
#824780000000
0!
1"
0'
1(
0/
10
#824790000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#824800000000
0!
0'
0/
#824810000000
1!
1'
1/
#824820000000
0!
0'
0/
#824830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#824840000000
0!
0'
0/
#824850000000
1!
1'
1/
#824860000000
0!
1"
0'
1(
0/
10
#824870000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#824880000000
0!
1$
0'
1+
0/
#824890000000
1!
1'
1/
#824900000000
0!
0'
0/
#824910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#824920000000
0!
0'
0/
#824930000000
1!
1'
1/
#824940000000
0!
0'
0/
#824950000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#824960000000
0!
0'
0/
#824970000000
1!
1'
1/
#824980000000
0!
0'
0/
#824990000000
1!
1'
1/
#825000000000
0!
0'
0/
#825010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#825020000000
0!
0'
0/
#825030000000
1!
1'
1/
#825040000000
0!
0'
0/
#825050000000
1!
1'
1/
#825060000000
0!
0'
0/
#825070000000
1!
1'
1/
#825080000000
0!
0'
0/
#825090000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#825100000000
0!
0'
0/
#825110000000
1!
1'
1/
#825120000000
0!
0'
0/
#825130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#825140000000
0!
0'
0/
#825150000000
1!
1'
1/
#825160000000
0!
0'
0/
#825170000000
#825180000000
1!
1'
1/
#825190000000
0!
0'
0/
#825200000000
1!
1'
1/
#825210000000
0!
1"
0'
1(
0/
10
#825220000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#825230000000
0!
0'
0/
#825240000000
1!
1'
1/
#825250000000
0!
0'
0/
#825260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#825270000000
0!
0'
0/
#825280000000
1!
1'
1/
#825290000000
0!
1"
0'
1(
0/
10
#825300000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#825310000000
0!
1$
0'
1+
0/
#825320000000
1!
1'
1/
#825330000000
0!
0'
0/
#825340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#825350000000
0!
0'
0/
#825360000000
1!
1'
1/
#825370000000
0!
0'
0/
#825380000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#825390000000
0!
0'
0/
#825400000000
1!
1'
1/
#825410000000
0!
0'
0/
#825420000000
1!
1'
1/
#825430000000
0!
0'
0/
#825440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#825450000000
0!
0'
0/
#825460000000
1!
1'
1/
#825470000000
0!
0'
0/
#825480000000
1!
1'
1/
#825490000000
0!
0'
0/
#825500000000
1!
1'
1/
#825510000000
0!
0'
0/
#825520000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#825530000000
0!
0'
0/
#825540000000
1!
1'
1/
#825550000000
0!
0'
0/
#825560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#825570000000
0!
0'
0/
#825580000000
1!
1'
1/
#825590000000
0!
0'
0/
#825600000000
#825610000000
1!
1'
1/
#825620000000
0!
0'
0/
#825630000000
1!
1'
1/
#825640000000
0!
1"
0'
1(
0/
10
#825650000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#825660000000
0!
0'
0/
#825670000000
1!
1'
1/
#825680000000
0!
0'
0/
#825690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#825700000000
0!
0'
0/
#825710000000
1!
1'
1/
#825720000000
0!
1"
0'
1(
0/
10
#825730000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#825740000000
0!
1$
0'
1+
0/
#825750000000
1!
1'
1/
#825760000000
0!
0'
0/
#825770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#825780000000
0!
0'
0/
#825790000000
1!
1'
1/
#825800000000
0!
0'
0/
#825810000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#825820000000
0!
0'
0/
#825830000000
1!
1'
1/
#825840000000
0!
0'
0/
#825850000000
1!
1'
1/
#825860000000
0!
0'
0/
#825870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#825880000000
0!
0'
0/
#825890000000
1!
1'
1/
#825900000000
0!
0'
0/
#825910000000
1!
1'
1/
#825920000000
0!
0'
0/
#825930000000
1!
1'
1/
#825940000000
0!
0'
0/
#825950000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#825960000000
0!
0'
0/
#825970000000
1!
1'
1/
#825980000000
0!
0'
0/
#825990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#826000000000
0!
0'
0/
#826010000000
1!
1'
1/
#826020000000
0!
0'
0/
#826030000000
#826040000000
1!
1'
1/
#826050000000
0!
0'
0/
#826060000000
1!
1'
1/
#826070000000
0!
1"
0'
1(
0/
10
#826080000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#826090000000
0!
0'
0/
#826100000000
1!
1'
1/
#826110000000
0!
0'
0/
#826120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#826130000000
0!
0'
0/
#826140000000
1!
1'
1/
#826150000000
0!
1"
0'
1(
0/
10
#826160000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#826170000000
0!
1$
0'
1+
0/
#826180000000
1!
1'
1/
#826190000000
0!
0'
0/
#826200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#826210000000
0!
0'
0/
#826220000000
1!
1'
1/
#826230000000
0!
0'
0/
#826240000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#826250000000
0!
0'
0/
#826260000000
1!
1'
1/
#826270000000
0!
0'
0/
#826280000000
1!
1'
1/
#826290000000
0!
0'
0/
#826300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#826310000000
0!
0'
0/
#826320000000
1!
1'
1/
#826330000000
0!
0'
0/
#826340000000
1!
1'
1/
#826350000000
0!
0'
0/
#826360000000
1!
1'
1/
#826370000000
0!
0'
0/
#826380000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#826390000000
0!
0'
0/
#826400000000
1!
1'
1/
#826410000000
0!
0'
0/
#826420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#826430000000
0!
0'
0/
#826440000000
1!
1'
1/
#826450000000
0!
0'
0/
#826460000000
#826470000000
1!
1'
1/
#826480000000
0!
0'
0/
#826490000000
1!
1'
1/
#826500000000
0!
1"
0'
1(
0/
10
#826510000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#826520000000
0!
0'
0/
#826530000000
1!
1'
1/
#826540000000
0!
0'
0/
#826550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#826560000000
0!
0'
0/
#826570000000
1!
1'
1/
#826580000000
0!
1"
0'
1(
0/
10
#826590000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#826600000000
0!
1$
0'
1+
0/
#826610000000
1!
1'
1/
#826620000000
0!
0'
0/
#826630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#826640000000
0!
0'
0/
#826650000000
1!
1'
1/
#826660000000
0!
0'
0/
#826670000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#826680000000
0!
0'
0/
#826690000000
1!
1'
1/
#826700000000
0!
0'
0/
#826710000000
1!
1'
1/
#826720000000
0!
0'
0/
#826730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#826740000000
0!
0'
0/
#826750000000
1!
1'
1/
#826760000000
0!
0'
0/
#826770000000
1!
1'
1/
#826780000000
0!
0'
0/
#826790000000
1!
1'
1/
#826800000000
0!
0'
0/
#826810000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#826820000000
0!
0'
0/
#826830000000
1!
1'
1/
#826840000000
0!
0'
0/
#826850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#826860000000
0!
0'
0/
#826870000000
1!
1'
1/
#826880000000
0!
0'
0/
#826890000000
#826900000000
1!
1'
1/
#826910000000
0!
0'
0/
#826920000000
1!
1'
1/
#826930000000
0!
1"
0'
1(
0/
10
#826940000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#826950000000
0!
0'
0/
#826960000000
1!
1'
1/
#826970000000
0!
0'
0/
#826980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#826990000000
0!
0'
0/
#827000000000
1!
1'
1/
#827010000000
0!
1"
0'
1(
0/
10
#827020000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#827030000000
0!
1$
0'
1+
0/
#827040000000
1!
1'
1/
#827050000000
0!
0'
0/
#827060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#827070000000
0!
0'
0/
#827080000000
1!
1'
1/
#827090000000
0!
0'
0/
#827100000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#827110000000
0!
0'
0/
#827120000000
1!
1'
1/
#827130000000
0!
0'
0/
#827140000000
1!
1'
1/
#827150000000
0!
0'
0/
#827160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#827170000000
0!
0'
0/
#827180000000
1!
1'
1/
#827190000000
0!
0'
0/
#827200000000
1!
1'
1/
#827210000000
0!
0'
0/
#827220000000
1!
1'
1/
#827230000000
0!
0'
0/
#827240000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#827250000000
0!
0'
0/
#827260000000
1!
1'
1/
#827270000000
0!
0'
0/
#827280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#827290000000
0!
0'
0/
#827300000000
1!
1'
1/
#827310000000
0!
0'
0/
#827320000000
#827330000000
1!
1'
1/
#827340000000
0!
0'
0/
#827350000000
1!
1'
1/
#827360000000
0!
1"
0'
1(
0/
10
#827370000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#827380000000
0!
0'
0/
#827390000000
1!
1'
1/
#827400000000
0!
0'
0/
#827410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#827420000000
0!
0'
0/
#827430000000
1!
1'
1/
#827440000000
0!
1"
0'
1(
0/
10
#827450000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#827460000000
0!
1$
0'
1+
0/
#827470000000
1!
1'
1/
#827480000000
0!
0'
0/
#827490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#827500000000
0!
0'
0/
#827510000000
1!
1'
1/
#827520000000
0!
0'
0/
#827530000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#827540000000
0!
0'
0/
#827550000000
1!
1'
1/
#827560000000
0!
0'
0/
#827570000000
1!
1'
1/
#827580000000
0!
0'
0/
#827590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#827600000000
0!
0'
0/
#827610000000
1!
1'
1/
#827620000000
0!
0'
0/
#827630000000
1!
1'
1/
#827640000000
0!
0'
0/
#827650000000
1!
1'
1/
#827660000000
0!
0'
0/
#827670000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#827680000000
0!
0'
0/
#827690000000
1!
1'
1/
#827700000000
0!
0'
0/
#827710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#827720000000
0!
0'
0/
#827730000000
1!
1'
1/
#827740000000
0!
0'
0/
#827750000000
#827760000000
1!
1'
1/
#827770000000
0!
0'
0/
#827780000000
1!
1'
1/
#827790000000
0!
1"
0'
1(
0/
10
#827800000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#827810000000
0!
0'
0/
#827820000000
1!
1'
1/
#827830000000
0!
0'
0/
#827840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#827850000000
0!
0'
0/
#827860000000
1!
1'
1/
#827870000000
0!
1"
0'
1(
0/
10
#827880000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#827890000000
0!
1$
0'
1+
0/
#827900000000
1!
1'
1/
#827910000000
0!
0'
0/
#827920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#827930000000
0!
0'
0/
#827940000000
1!
1'
1/
#827950000000
0!
0'
0/
#827960000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#827970000000
0!
0'
0/
#827980000000
1!
1'
1/
#827990000000
0!
0'
0/
#828000000000
1!
1'
1/
#828010000000
0!
0'
0/
#828020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#828030000000
0!
0'
0/
#828040000000
1!
1'
1/
#828050000000
0!
0'
0/
#828060000000
1!
1'
1/
#828070000000
0!
0'
0/
#828080000000
1!
1'
1/
#828090000000
0!
0'
0/
#828100000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#828110000000
0!
0'
0/
#828120000000
1!
1'
1/
#828130000000
0!
0'
0/
#828140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#828150000000
0!
0'
0/
#828160000000
1!
1'
1/
#828170000000
0!
0'
0/
#828180000000
#828190000000
1!
1'
1/
#828200000000
0!
0'
0/
#828210000000
1!
1'
1/
#828220000000
0!
1"
0'
1(
0/
10
#828230000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#828240000000
0!
0'
0/
#828250000000
1!
1'
1/
#828260000000
0!
0'
0/
#828270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#828280000000
0!
0'
0/
#828290000000
1!
1'
1/
#828300000000
0!
1"
0'
1(
0/
10
#828310000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#828320000000
0!
1$
0'
1+
0/
#828330000000
1!
1'
1/
#828340000000
0!
0'
0/
#828350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#828360000000
0!
0'
0/
#828370000000
1!
1'
1/
#828380000000
0!
0'
0/
#828390000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#828400000000
0!
0'
0/
#828410000000
1!
1'
1/
#828420000000
0!
0'
0/
#828430000000
1!
1'
1/
#828440000000
0!
0'
0/
#828450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#828460000000
0!
0'
0/
#828470000000
1!
1'
1/
#828480000000
0!
0'
0/
#828490000000
1!
1'
1/
#828500000000
0!
0'
0/
#828510000000
1!
1'
1/
#828520000000
0!
0'
0/
#828530000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#828540000000
0!
0'
0/
#828550000000
1!
1'
1/
#828560000000
0!
0'
0/
#828570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#828580000000
0!
0'
0/
#828590000000
1!
1'
1/
#828600000000
0!
0'
0/
#828610000000
#828620000000
1!
1'
1/
#828630000000
0!
0'
0/
#828640000000
1!
1'
1/
#828650000000
0!
1"
0'
1(
0/
10
#828660000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#828670000000
0!
0'
0/
#828680000000
1!
1'
1/
#828690000000
0!
0'
0/
#828700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#828710000000
0!
0'
0/
#828720000000
1!
1'
1/
#828730000000
0!
1"
0'
1(
0/
10
#828740000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#828750000000
0!
1$
0'
1+
0/
#828760000000
1!
1'
1/
#828770000000
0!
0'
0/
#828780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#828790000000
0!
0'
0/
#828800000000
1!
1'
1/
#828810000000
0!
0'
0/
#828820000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#828830000000
0!
0'
0/
#828840000000
1!
1'
1/
#828850000000
0!
0'
0/
#828860000000
1!
1'
1/
#828870000000
0!
0'
0/
#828880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#828890000000
0!
0'
0/
#828900000000
1!
1'
1/
#828910000000
0!
0'
0/
#828920000000
1!
1'
1/
#828930000000
0!
0'
0/
#828940000000
1!
1'
1/
#828950000000
0!
0'
0/
#828960000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#828970000000
0!
0'
0/
#828980000000
1!
1'
1/
#828990000000
0!
0'
0/
#829000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#829010000000
0!
0'
0/
#829020000000
1!
1'
1/
#829030000000
0!
0'
0/
#829040000000
#829050000000
1!
1'
1/
#829060000000
0!
0'
0/
#829070000000
1!
1'
1/
#829080000000
0!
1"
0'
1(
0/
10
#829090000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#829100000000
0!
0'
0/
#829110000000
1!
1'
1/
#829120000000
0!
0'
0/
#829130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#829140000000
0!
0'
0/
#829150000000
1!
1'
1/
#829160000000
0!
1"
0'
1(
0/
10
#829170000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#829180000000
0!
1$
0'
1+
0/
#829190000000
1!
1'
1/
#829200000000
0!
0'
0/
#829210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#829220000000
0!
0'
0/
#829230000000
1!
1'
1/
#829240000000
0!
0'
0/
#829250000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#829260000000
0!
0'
0/
#829270000000
1!
1'
1/
#829280000000
0!
0'
0/
#829290000000
1!
1'
1/
#829300000000
0!
0'
0/
#829310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#829320000000
0!
0'
0/
#829330000000
1!
1'
1/
#829340000000
0!
0'
0/
#829350000000
1!
1'
1/
#829360000000
0!
0'
0/
#829370000000
1!
1'
1/
#829380000000
0!
0'
0/
#829390000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#829400000000
0!
0'
0/
#829410000000
1!
1'
1/
#829420000000
0!
0'
0/
#829430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#829440000000
0!
0'
0/
#829450000000
1!
1'
1/
#829460000000
0!
0'
0/
#829470000000
#829480000000
1!
1'
1/
#829490000000
0!
0'
0/
#829500000000
1!
1'
1/
#829510000000
0!
1"
0'
1(
0/
10
#829520000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#829530000000
0!
0'
0/
#829540000000
1!
1'
1/
#829550000000
0!
0'
0/
#829560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#829570000000
0!
0'
0/
#829580000000
1!
1'
1/
#829590000000
0!
1"
0'
1(
0/
10
#829600000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#829610000000
0!
1$
0'
1+
0/
#829620000000
1!
1'
1/
#829630000000
0!
0'
0/
#829640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#829650000000
0!
0'
0/
#829660000000
1!
1'
1/
#829670000000
0!
0'
0/
#829680000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#829690000000
0!
0'
0/
#829700000000
1!
1'
1/
#829710000000
0!
0'
0/
#829720000000
1!
1'
1/
#829730000000
0!
0'
0/
#829740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#829750000000
0!
0'
0/
#829760000000
1!
1'
1/
#829770000000
0!
0'
0/
#829780000000
1!
1'
1/
#829790000000
0!
0'
0/
#829800000000
1!
1'
1/
#829810000000
0!
0'
0/
#829820000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#829830000000
0!
0'
0/
#829840000000
1!
1'
1/
#829850000000
0!
0'
0/
#829860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#829870000000
0!
0'
0/
#829880000000
1!
1'
1/
#829890000000
0!
0'
0/
#829900000000
#829910000000
1!
1'
1/
#829920000000
0!
0'
0/
#829930000000
1!
1'
1/
#829940000000
0!
1"
0'
1(
0/
10
#829950000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#829960000000
0!
0'
0/
#829970000000
1!
1'
1/
#829980000000
0!
0'
0/
#829990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#830000000000
0!
0'
0/
#830010000000
1!
1'
1/
#830020000000
0!
1"
0'
1(
0/
10
#830030000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#830040000000
0!
1$
0'
1+
0/
#830050000000
1!
1'
1/
#830060000000
0!
0'
0/
#830070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#830080000000
0!
0'
0/
#830090000000
1!
1'
1/
#830100000000
0!
0'
0/
#830110000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#830120000000
0!
0'
0/
#830130000000
1!
1'
1/
#830140000000
0!
0'
0/
#830150000000
1!
1'
1/
#830160000000
0!
0'
0/
#830170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#830180000000
0!
0'
0/
#830190000000
1!
1'
1/
#830200000000
0!
0'
0/
#830210000000
1!
1'
1/
#830220000000
0!
0'
0/
#830230000000
1!
1'
1/
#830240000000
0!
0'
0/
#830250000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#830260000000
0!
0'
0/
#830270000000
1!
1'
1/
#830280000000
0!
0'
0/
#830290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#830300000000
0!
0'
0/
#830310000000
1!
1'
1/
#830320000000
0!
0'
0/
#830330000000
#830340000000
1!
1'
1/
#830350000000
0!
0'
0/
#830360000000
1!
1'
1/
#830370000000
0!
1"
0'
1(
0/
10
#830380000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#830390000000
0!
0'
0/
#830400000000
1!
1'
1/
#830410000000
0!
0'
0/
#830420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#830430000000
0!
0'
0/
#830440000000
1!
1'
1/
#830450000000
0!
1"
0'
1(
0/
10
#830460000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#830470000000
0!
1$
0'
1+
0/
#830480000000
1!
1'
1/
#830490000000
0!
0'
0/
#830500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#830510000000
0!
0'
0/
#830520000000
1!
1'
1/
#830530000000
0!
0'
0/
#830540000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#830550000000
0!
0'
0/
#830560000000
1!
1'
1/
#830570000000
0!
0'
0/
#830580000000
1!
1'
1/
#830590000000
0!
0'
0/
#830600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#830610000000
0!
0'
0/
#830620000000
1!
1'
1/
#830630000000
0!
0'
0/
#830640000000
1!
1'
1/
#830650000000
0!
0'
0/
#830660000000
1!
1'
1/
#830670000000
0!
0'
0/
#830680000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#830690000000
0!
0'
0/
#830700000000
1!
1'
1/
#830710000000
0!
0'
0/
#830720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#830730000000
0!
0'
0/
#830740000000
1!
1'
1/
#830750000000
0!
0'
0/
#830760000000
#830770000000
1!
1'
1/
#830780000000
0!
0'
0/
#830790000000
1!
1'
1/
#830800000000
0!
1"
0'
1(
0/
10
#830810000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#830820000000
0!
0'
0/
#830830000000
1!
1'
1/
#830840000000
0!
0'
0/
#830850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#830860000000
0!
0'
0/
#830870000000
1!
1'
1/
#830880000000
0!
1"
0'
1(
0/
10
#830890000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#830900000000
0!
1$
0'
1+
0/
#830910000000
1!
1'
1/
#830920000000
0!
0'
0/
#830930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#830940000000
0!
0'
0/
#830950000000
1!
1'
1/
#830960000000
0!
0'
0/
#830970000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#830980000000
0!
0'
0/
#830990000000
1!
1'
1/
#831000000000
0!
0'
0/
#831010000000
1!
1'
1/
#831020000000
0!
0'
0/
#831030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#831040000000
0!
0'
0/
#831050000000
1!
1'
1/
#831060000000
0!
0'
0/
#831070000000
1!
1'
1/
#831080000000
0!
0'
0/
#831090000000
1!
1'
1/
#831100000000
0!
0'
0/
#831110000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#831120000000
0!
0'
0/
#831130000000
1!
1'
1/
#831140000000
0!
0'
0/
#831150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#831160000000
0!
0'
0/
#831170000000
1!
1'
1/
#831180000000
0!
0'
0/
#831190000000
#831200000000
1!
1'
1/
#831210000000
0!
0'
0/
#831220000000
1!
1'
1/
#831230000000
0!
1"
0'
1(
0/
10
#831240000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#831250000000
0!
0'
0/
#831260000000
1!
1'
1/
#831270000000
0!
0'
0/
#831280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#831290000000
0!
0'
0/
#831300000000
1!
1'
1/
#831310000000
0!
1"
0'
1(
0/
10
#831320000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#831330000000
0!
1$
0'
1+
0/
#831340000000
1!
1'
1/
#831350000000
0!
0'
0/
#831360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#831370000000
0!
0'
0/
#831380000000
1!
1'
1/
#831390000000
0!
0'
0/
#831400000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#831410000000
0!
0'
0/
#831420000000
1!
1'
1/
#831430000000
0!
0'
0/
#831440000000
1!
1'
1/
#831450000000
0!
0'
0/
#831460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#831470000000
0!
0'
0/
#831480000000
1!
1'
1/
#831490000000
0!
0'
0/
#831500000000
1!
1'
1/
#831510000000
0!
0'
0/
#831520000000
1!
1'
1/
#831530000000
0!
0'
0/
#831540000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#831550000000
0!
0'
0/
#831560000000
1!
1'
1/
#831570000000
0!
0'
0/
#831580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#831590000000
0!
0'
0/
#831600000000
1!
1'
1/
#831610000000
0!
0'
0/
#831620000000
#831630000000
1!
1'
1/
#831640000000
0!
0'
0/
#831650000000
1!
1'
1/
#831660000000
0!
1"
0'
1(
0/
10
#831670000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#831680000000
0!
0'
0/
#831690000000
1!
1'
1/
#831700000000
0!
0'
0/
#831710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#831720000000
0!
0'
0/
#831730000000
1!
1'
1/
#831740000000
0!
1"
0'
1(
0/
10
#831750000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#831760000000
0!
1$
0'
1+
0/
#831770000000
1!
1'
1/
#831780000000
0!
0'
0/
#831790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#831800000000
0!
0'
0/
#831810000000
1!
1'
1/
#831820000000
0!
0'
0/
#831830000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#831840000000
0!
0'
0/
#831850000000
1!
1'
1/
#831860000000
0!
0'
0/
#831870000000
1!
1'
1/
#831880000000
0!
0'
0/
#831890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#831900000000
0!
0'
0/
#831910000000
1!
1'
1/
#831920000000
0!
0'
0/
#831930000000
1!
1'
1/
#831940000000
0!
0'
0/
#831950000000
1!
1'
1/
#831960000000
0!
0'
0/
#831970000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#831980000000
0!
0'
0/
#831990000000
1!
1'
1/
#832000000000
0!
0'
0/
#832010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#832020000000
0!
0'
0/
#832030000000
1!
1'
1/
#832040000000
0!
0'
0/
#832050000000
#832060000000
1!
1'
1/
#832070000000
0!
0'
0/
#832080000000
1!
1'
1/
#832090000000
0!
1"
0'
1(
0/
10
#832100000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#832110000000
0!
0'
0/
#832120000000
1!
1'
1/
#832130000000
0!
0'
0/
#832140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#832150000000
0!
0'
0/
#832160000000
1!
1'
1/
#832170000000
0!
1"
0'
1(
0/
10
#832180000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#832190000000
0!
1$
0'
1+
0/
#832200000000
1!
1'
1/
#832210000000
0!
0'
0/
#832220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#832230000000
0!
0'
0/
#832240000000
1!
1'
1/
#832250000000
0!
0'
0/
#832260000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#832270000000
0!
0'
0/
#832280000000
1!
1'
1/
#832290000000
0!
0'
0/
#832300000000
1!
1'
1/
#832310000000
0!
0'
0/
#832320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#832330000000
0!
0'
0/
#832340000000
1!
1'
1/
#832350000000
0!
0'
0/
#832360000000
1!
1'
1/
#832370000000
0!
0'
0/
#832380000000
1!
1'
1/
#832390000000
0!
0'
0/
#832400000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#832410000000
0!
0'
0/
#832420000000
1!
1'
1/
#832430000000
0!
0'
0/
#832440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#832450000000
0!
0'
0/
#832460000000
1!
1'
1/
#832470000000
0!
0'
0/
#832480000000
#832490000000
1!
1'
1/
#832500000000
0!
0'
0/
#832510000000
1!
1'
1/
#832520000000
0!
1"
0'
1(
0/
10
#832530000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#832540000000
0!
0'
0/
#832550000000
1!
1'
1/
#832560000000
0!
0'
0/
#832570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#832580000000
0!
0'
0/
#832590000000
1!
1'
1/
#832600000000
0!
1"
0'
1(
0/
10
#832610000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#832620000000
0!
1$
0'
1+
0/
#832630000000
1!
1'
1/
#832640000000
0!
0'
0/
#832650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#832660000000
0!
0'
0/
#832670000000
1!
1'
1/
#832680000000
0!
0'
0/
#832690000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#832700000000
0!
0'
0/
#832710000000
1!
1'
1/
#832720000000
0!
0'
0/
#832730000000
1!
1'
1/
#832740000000
0!
0'
0/
#832750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#832760000000
0!
0'
0/
#832770000000
1!
1'
1/
#832780000000
0!
0'
0/
#832790000000
1!
1'
1/
#832800000000
0!
0'
0/
#832810000000
1!
1'
1/
#832820000000
0!
0'
0/
#832830000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#832840000000
0!
0'
0/
#832850000000
1!
1'
1/
#832860000000
0!
0'
0/
#832870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#832880000000
0!
0'
0/
#832890000000
1!
1'
1/
#832900000000
0!
0'
0/
#832910000000
#832920000000
1!
1'
1/
#832930000000
0!
0'
0/
#832940000000
1!
1'
1/
#832950000000
0!
1"
0'
1(
0/
10
#832960000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#832970000000
0!
0'
0/
#832980000000
1!
1'
1/
#832990000000
0!
0'
0/
#833000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#833010000000
0!
0'
0/
#833020000000
1!
1'
1/
#833030000000
0!
1"
0'
1(
0/
10
#833040000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#833050000000
0!
1$
0'
1+
0/
#833060000000
1!
1'
1/
#833070000000
0!
0'
0/
#833080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#833090000000
0!
0'
0/
#833100000000
1!
1'
1/
#833110000000
0!
0'
0/
#833120000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#833130000000
0!
0'
0/
#833140000000
1!
1'
1/
#833150000000
0!
0'
0/
#833160000000
1!
1'
1/
#833170000000
0!
0'
0/
#833180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#833190000000
0!
0'
0/
#833200000000
1!
1'
1/
#833210000000
0!
0'
0/
#833220000000
1!
1'
1/
#833230000000
0!
0'
0/
#833240000000
1!
1'
1/
#833250000000
0!
0'
0/
#833260000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#833270000000
0!
0'
0/
#833280000000
1!
1'
1/
#833290000000
0!
0'
0/
#833300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#833310000000
0!
0'
0/
#833320000000
1!
1'
1/
#833330000000
0!
0'
0/
#833340000000
#833350000000
1!
1'
1/
#833360000000
0!
0'
0/
#833370000000
1!
1'
1/
#833380000000
0!
1"
0'
1(
0/
10
#833390000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#833400000000
0!
0'
0/
#833410000000
1!
1'
1/
#833420000000
0!
0'
0/
#833430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#833440000000
0!
0'
0/
#833450000000
1!
1'
1/
#833460000000
0!
1"
0'
1(
0/
10
#833470000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#833480000000
0!
1$
0'
1+
0/
#833490000000
1!
1'
1/
#833500000000
0!
0'
0/
#833510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#833520000000
0!
0'
0/
#833530000000
1!
1'
1/
#833540000000
0!
0'
0/
#833550000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#833560000000
0!
0'
0/
#833570000000
1!
1'
1/
#833580000000
0!
0'
0/
#833590000000
1!
1'
1/
#833600000000
0!
0'
0/
#833610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#833620000000
0!
0'
0/
#833630000000
1!
1'
1/
#833640000000
0!
0'
0/
#833650000000
1!
1'
1/
#833660000000
0!
0'
0/
#833670000000
1!
1'
1/
#833680000000
0!
0'
0/
#833690000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#833700000000
0!
0'
0/
#833710000000
1!
1'
1/
#833720000000
0!
0'
0/
#833730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#833740000000
0!
0'
0/
#833750000000
1!
1'
1/
#833760000000
0!
0'
0/
#833770000000
#833780000000
1!
1'
1/
#833790000000
0!
0'
0/
#833800000000
1!
1'
1/
#833810000000
0!
1"
0'
1(
0/
10
#833820000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#833830000000
0!
0'
0/
#833840000000
1!
1'
1/
#833850000000
0!
0'
0/
#833860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#833870000000
0!
0'
0/
#833880000000
1!
1'
1/
#833890000000
0!
1"
0'
1(
0/
10
#833900000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#833910000000
0!
1$
0'
1+
0/
#833920000000
1!
1'
1/
#833930000000
0!
0'
0/
#833940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#833950000000
0!
0'
0/
#833960000000
1!
1'
1/
#833970000000
0!
0'
0/
#833980000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#833990000000
0!
0'
0/
#834000000000
1!
1'
1/
#834010000000
0!
0'
0/
#834020000000
1!
1'
1/
#834030000000
0!
0'
0/
#834040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#834050000000
0!
0'
0/
#834060000000
1!
1'
1/
#834070000000
0!
0'
0/
#834080000000
1!
1'
1/
#834090000000
0!
0'
0/
#834100000000
1!
1'
1/
#834110000000
0!
0'
0/
#834120000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#834130000000
0!
0'
0/
#834140000000
1!
1'
1/
#834150000000
0!
0'
0/
#834160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#834170000000
0!
0'
0/
#834180000000
1!
1'
1/
#834190000000
0!
0'
0/
#834200000000
#834210000000
1!
1'
1/
#834220000000
0!
0'
0/
#834230000000
1!
1'
1/
#834240000000
0!
1"
0'
1(
0/
10
#834250000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#834260000000
0!
0'
0/
#834270000000
1!
1'
1/
#834280000000
0!
0'
0/
#834290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#834300000000
0!
0'
0/
#834310000000
1!
1'
1/
#834320000000
0!
1"
0'
1(
0/
10
#834330000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#834340000000
0!
1$
0'
1+
0/
#834350000000
1!
1'
1/
#834360000000
0!
0'
0/
#834370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#834380000000
0!
0'
0/
#834390000000
1!
1'
1/
#834400000000
0!
0'
0/
#834410000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#834420000000
0!
0'
0/
#834430000000
1!
1'
1/
#834440000000
0!
0'
0/
#834450000000
1!
1'
1/
#834460000000
0!
0'
0/
#834470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#834480000000
0!
0'
0/
#834490000000
1!
1'
1/
#834500000000
0!
0'
0/
#834510000000
1!
1'
1/
#834520000000
0!
0'
0/
#834530000000
1!
1'
1/
#834540000000
0!
0'
0/
#834550000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#834560000000
0!
0'
0/
#834570000000
1!
1'
1/
#834580000000
0!
0'
0/
#834590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#834600000000
0!
0'
0/
#834610000000
1!
1'
1/
#834620000000
0!
0'
0/
#834630000000
#834640000000
1!
1'
1/
#834650000000
0!
0'
0/
#834660000000
1!
1'
1/
#834670000000
0!
1"
0'
1(
0/
10
#834680000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#834690000000
0!
0'
0/
#834700000000
1!
1'
1/
#834710000000
0!
0'
0/
#834720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#834730000000
0!
0'
0/
#834740000000
1!
1'
1/
#834750000000
0!
1"
0'
1(
0/
10
#834760000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#834770000000
0!
1$
0'
1+
0/
#834780000000
1!
1'
1/
#834790000000
0!
0'
0/
#834800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#834810000000
0!
0'
0/
#834820000000
1!
1'
1/
#834830000000
0!
0'
0/
#834840000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#834850000000
0!
0'
0/
#834860000000
1!
1'
1/
#834870000000
0!
0'
0/
#834880000000
1!
1'
1/
#834890000000
0!
0'
0/
#834900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#834910000000
0!
0'
0/
#834920000000
1!
1'
1/
#834930000000
0!
0'
0/
#834940000000
1!
1'
1/
#834950000000
0!
0'
0/
#834960000000
1!
1'
1/
#834970000000
0!
0'
0/
#834980000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#834990000000
0!
0'
0/
#835000000000
1!
1'
1/
#835010000000
0!
0'
0/
#835020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#835030000000
0!
0'
0/
#835040000000
1!
1'
1/
#835050000000
0!
0'
0/
#835060000000
#835070000000
1!
1'
1/
#835080000000
0!
0'
0/
#835090000000
1!
1'
1/
#835100000000
0!
1"
0'
1(
0/
10
#835110000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#835120000000
0!
0'
0/
#835130000000
1!
1'
1/
#835140000000
0!
0'
0/
#835150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#835160000000
0!
0'
0/
#835170000000
1!
1'
1/
#835180000000
0!
1"
0'
1(
0/
10
#835190000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#835200000000
0!
1$
0'
1+
0/
#835210000000
1!
1'
1/
#835220000000
0!
0'
0/
#835230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#835240000000
0!
0'
0/
#835250000000
1!
1'
1/
#835260000000
0!
0'
0/
#835270000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#835280000000
0!
0'
0/
#835290000000
1!
1'
1/
#835300000000
0!
0'
0/
#835310000000
1!
1'
1/
#835320000000
0!
0'
0/
#835330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#835340000000
0!
0'
0/
#835350000000
1!
1'
1/
#835360000000
0!
0'
0/
#835370000000
1!
1'
1/
#835380000000
0!
0'
0/
#835390000000
1!
1'
1/
#835400000000
0!
0'
0/
#835410000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#835420000000
0!
0'
0/
#835430000000
1!
1'
1/
#835440000000
0!
0'
0/
#835450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#835460000000
0!
0'
0/
#835470000000
1!
1'
1/
#835480000000
0!
0'
0/
#835490000000
#835500000000
1!
1'
1/
#835510000000
0!
0'
0/
#835520000000
1!
1'
1/
#835530000000
0!
1"
0'
1(
0/
10
#835540000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#835550000000
0!
0'
0/
#835560000000
1!
1'
1/
#835570000000
0!
0'
0/
#835580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#835590000000
0!
0'
0/
#835600000000
1!
1'
1/
#835610000000
0!
1"
0'
1(
0/
10
#835620000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#835630000000
0!
1$
0'
1+
0/
#835640000000
1!
1'
1/
#835650000000
0!
0'
0/
#835660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#835670000000
0!
0'
0/
#835680000000
1!
1'
1/
#835690000000
0!
0'
0/
#835700000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#835710000000
0!
0'
0/
#835720000000
1!
1'
1/
#835730000000
0!
0'
0/
#835740000000
1!
1'
1/
#835750000000
0!
0'
0/
#835760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#835770000000
0!
0'
0/
#835780000000
1!
1'
1/
#835790000000
0!
0'
0/
#835800000000
1!
1'
1/
#835810000000
0!
0'
0/
#835820000000
1!
1'
1/
#835830000000
0!
0'
0/
#835840000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#835850000000
0!
0'
0/
#835860000000
1!
1'
1/
#835870000000
0!
0'
0/
#835880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#835890000000
0!
0'
0/
#835900000000
1!
1'
1/
#835910000000
0!
0'
0/
#835920000000
#835930000000
1!
1'
1/
#835940000000
0!
0'
0/
#835950000000
1!
1'
1/
#835960000000
0!
1"
0'
1(
0/
10
#835970000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#835980000000
0!
0'
0/
#835990000000
1!
1'
1/
#836000000000
0!
0'
0/
#836010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#836020000000
0!
0'
0/
#836030000000
1!
1'
1/
#836040000000
0!
1"
0'
1(
0/
10
#836050000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#836060000000
0!
1$
0'
1+
0/
#836070000000
1!
1'
1/
#836080000000
0!
0'
0/
#836090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#836100000000
0!
0'
0/
#836110000000
1!
1'
1/
#836120000000
0!
0'
0/
#836130000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#836140000000
0!
0'
0/
#836150000000
1!
1'
1/
#836160000000
0!
0'
0/
#836170000000
1!
1'
1/
#836180000000
0!
0'
0/
#836190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#836200000000
0!
0'
0/
#836210000000
1!
1'
1/
#836220000000
0!
0'
0/
#836230000000
1!
1'
1/
#836240000000
0!
0'
0/
#836250000000
1!
1'
1/
#836260000000
0!
0'
0/
#836270000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#836280000000
0!
0'
0/
#836290000000
1!
1'
1/
#836300000000
0!
0'
0/
#836310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#836320000000
0!
0'
0/
#836330000000
1!
1'
1/
#836340000000
0!
0'
0/
#836350000000
#836360000000
1!
1'
1/
#836370000000
0!
0'
0/
#836380000000
1!
1'
1/
#836390000000
0!
1"
0'
1(
0/
10
#836400000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#836410000000
0!
0'
0/
#836420000000
1!
1'
1/
#836430000000
0!
0'
0/
#836440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#836450000000
0!
0'
0/
#836460000000
1!
1'
1/
#836470000000
0!
1"
0'
1(
0/
10
#836480000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#836490000000
0!
1$
0'
1+
0/
#836500000000
1!
1'
1/
#836510000000
0!
0'
0/
#836520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#836530000000
0!
0'
0/
#836540000000
1!
1'
1/
#836550000000
0!
0'
0/
#836560000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#836570000000
0!
0'
0/
#836580000000
1!
1'
1/
#836590000000
0!
0'
0/
#836600000000
1!
1'
1/
#836610000000
0!
0'
0/
#836620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#836630000000
0!
0'
0/
#836640000000
1!
1'
1/
#836650000000
0!
0'
0/
#836660000000
1!
1'
1/
#836670000000
0!
0'
0/
#836680000000
1!
1'
1/
#836690000000
0!
0'
0/
#836700000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#836710000000
0!
0'
0/
#836720000000
1!
1'
1/
#836730000000
0!
0'
0/
#836740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#836750000000
0!
0'
0/
#836760000000
1!
1'
1/
#836770000000
0!
0'
0/
#836780000000
#836790000000
1!
1'
1/
#836800000000
0!
0'
0/
#836810000000
1!
1'
1/
#836820000000
0!
1"
0'
1(
0/
10
#836830000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#836840000000
0!
0'
0/
#836850000000
1!
1'
1/
#836860000000
0!
0'
0/
#836870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#836880000000
0!
0'
0/
#836890000000
1!
1'
1/
#836900000000
0!
1"
0'
1(
0/
10
#836910000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#836920000000
0!
1$
0'
1+
0/
#836930000000
1!
1'
1/
#836940000000
0!
0'
0/
#836950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#836960000000
0!
0'
0/
#836970000000
1!
1'
1/
#836980000000
0!
0'
0/
#836990000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#837000000000
0!
0'
0/
#837010000000
1!
1'
1/
#837020000000
0!
0'
0/
#837030000000
1!
1'
1/
#837040000000
0!
0'
0/
#837050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#837060000000
0!
0'
0/
#837070000000
1!
1'
1/
#837080000000
0!
0'
0/
#837090000000
1!
1'
1/
#837100000000
0!
0'
0/
#837110000000
1!
1'
1/
#837120000000
0!
0'
0/
#837130000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#837140000000
0!
0'
0/
#837150000000
1!
1'
1/
#837160000000
0!
0'
0/
#837170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#837180000000
0!
0'
0/
#837190000000
1!
1'
1/
#837200000000
0!
0'
0/
#837210000000
#837220000000
1!
1'
1/
#837230000000
0!
0'
0/
#837240000000
1!
1'
1/
#837250000000
0!
1"
0'
1(
0/
10
#837260000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#837270000000
0!
0'
0/
#837280000000
1!
1'
1/
#837290000000
0!
0'
0/
#837300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#837310000000
0!
0'
0/
#837320000000
1!
1'
1/
#837330000000
0!
1"
0'
1(
0/
10
#837340000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#837350000000
0!
1$
0'
1+
0/
#837360000000
1!
1'
1/
#837370000000
0!
0'
0/
#837380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#837390000000
0!
0'
0/
#837400000000
1!
1'
1/
#837410000000
0!
0'
0/
#837420000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#837430000000
0!
0'
0/
#837440000000
1!
1'
1/
#837450000000
0!
0'
0/
#837460000000
1!
1'
1/
#837470000000
0!
0'
0/
#837480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#837490000000
0!
0'
0/
#837500000000
1!
1'
1/
#837510000000
0!
0'
0/
#837520000000
1!
1'
1/
#837530000000
0!
0'
0/
#837540000000
1!
1'
1/
#837550000000
0!
0'
0/
#837560000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#837570000000
0!
0'
0/
#837580000000
1!
1'
1/
#837590000000
0!
0'
0/
#837600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#837610000000
0!
0'
0/
#837620000000
1!
1'
1/
#837630000000
0!
0'
0/
#837640000000
#837650000000
1!
1'
1/
#837660000000
0!
0'
0/
#837670000000
1!
1'
1/
#837680000000
0!
1"
0'
1(
0/
10
#837690000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#837700000000
0!
0'
0/
#837710000000
1!
1'
1/
#837720000000
0!
0'
0/
#837730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#837740000000
0!
0'
0/
#837750000000
1!
1'
1/
#837760000000
0!
1"
0'
1(
0/
10
#837770000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#837780000000
0!
1$
0'
1+
0/
#837790000000
1!
1'
1/
#837800000000
0!
0'
0/
#837810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#837820000000
0!
0'
0/
#837830000000
1!
1'
1/
#837840000000
0!
0'
0/
#837850000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#837860000000
0!
0'
0/
#837870000000
1!
1'
1/
#837880000000
0!
0'
0/
#837890000000
1!
1'
1/
#837900000000
0!
0'
0/
#837910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#837920000000
0!
0'
0/
#837930000000
1!
1'
1/
#837940000000
0!
0'
0/
#837950000000
1!
1'
1/
#837960000000
0!
0'
0/
#837970000000
1!
1'
1/
#837980000000
0!
0'
0/
#837990000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#838000000000
0!
0'
0/
#838010000000
1!
1'
1/
#838020000000
0!
0'
0/
#838030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#838040000000
0!
0'
0/
#838050000000
1!
1'
1/
#838060000000
0!
0'
0/
#838070000000
#838080000000
1!
1'
1/
#838090000000
0!
0'
0/
#838100000000
1!
1'
1/
#838110000000
0!
1"
0'
1(
0/
10
#838120000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#838130000000
0!
0'
0/
#838140000000
1!
1'
1/
#838150000000
0!
0'
0/
#838160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#838170000000
0!
0'
0/
#838180000000
1!
1'
1/
#838190000000
0!
1"
0'
1(
0/
10
#838200000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#838210000000
0!
1$
0'
1+
0/
#838220000000
1!
1'
1/
#838230000000
0!
0'
0/
#838240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#838250000000
0!
0'
0/
#838260000000
1!
1'
1/
#838270000000
0!
0'
0/
#838280000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#838290000000
0!
0'
0/
#838300000000
1!
1'
1/
#838310000000
0!
0'
0/
#838320000000
1!
1'
1/
#838330000000
0!
0'
0/
#838340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#838350000000
0!
0'
0/
#838360000000
1!
1'
1/
#838370000000
0!
0'
0/
#838380000000
1!
1'
1/
#838390000000
0!
0'
0/
#838400000000
1!
1'
1/
#838410000000
0!
0'
0/
#838420000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#838430000000
0!
0'
0/
#838440000000
1!
1'
1/
#838450000000
0!
0'
0/
#838460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#838470000000
0!
0'
0/
#838480000000
1!
1'
1/
#838490000000
0!
0'
0/
#838500000000
#838510000000
1!
1'
1/
#838520000000
0!
0'
0/
#838530000000
1!
1'
1/
#838540000000
0!
1"
0'
1(
0/
10
#838550000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#838560000000
0!
0'
0/
#838570000000
1!
1'
1/
#838580000000
0!
0'
0/
#838590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#838600000000
0!
0'
0/
#838610000000
1!
1'
1/
#838620000000
0!
1"
0'
1(
0/
10
#838630000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#838640000000
0!
1$
0'
1+
0/
#838650000000
1!
1'
1/
#838660000000
0!
0'
0/
#838670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#838680000000
0!
0'
0/
#838690000000
1!
1'
1/
#838700000000
0!
0'
0/
#838710000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#838720000000
0!
0'
0/
#838730000000
1!
1'
1/
#838740000000
0!
0'
0/
#838750000000
1!
1'
1/
#838760000000
0!
0'
0/
#838770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#838780000000
0!
0'
0/
#838790000000
1!
1'
1/
#838800000000
0!
0'
0/
#838810000000
1!
1'
1/
#838820000000
0!
0'
0/
#838830000000
1!
1'
1/
#838840000000
0!
0'
0/
#838850000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#838860000000
0!
0'
0/
#838870000000
1!
1'
1/
#838880000000
0!
0'
0/
#838890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#838900000000
0!
0'
0/
#838910000000
1!
1'
1/
#838920000000
0!
0'
0/
#838930000000
#838940000000
1!
1'
1/
#838950000000
0!
0'
0/
#838960000000
1!
1'
1/
#838970000000
0!
1"
0'
1(
0/
10
#838980000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#838990000000
0!
0'
0/
#839000000000
1!
1'
1/
#839010000000
0!
0'
0/
#839020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#839030000000
0!
0'
0/
#839040000000
1!
1'
1/
#839050000000
0!
1"
0'
1(
0/
10
#839060000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#839070000000
0!
1$
0'
1+
0/
#839080000000
1!
1'
1/
#839090000000
0!
0'
0/
#839100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#839110000000
0!
0'
0/
#839120000000
1!
1'
1/
#839130000000
0!
0'
0/
#839140000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#839150000000
0!
0'
0/
#839160000000
1!
1'
1/
#839170000000
0!
0'
0/
#839180000000
1!
1'
1/
#839190000000
0!
0'
0/
#839200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#839210000000
0!
0'
0/
#839220000000
1!
1'
1/
#839230000000
0!
0'
0/
#839240000000
1!
1'
1/
#839250000000
0!
0'
0/
#839260000000
1!
1'
1/
#839270000000
0!
0'
0/
#839280000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#839290000000
0!
0'
0/
#839300000000
1!
1'
1/
#839310000000
0!
0'
0/
#839320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#839330000000
0!
0'
0/
#839340000000
1!
1'
1/
#839350000000
0!
0'
0/
#839360000000
#839370000000
1!
1'
1/
#839380000000
0!
0'
0/
#839390000000
1!
1'
1/
#839400000000
0!
1"
0'
1(
0/
10
#839410000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#839420000000
0!
0'
0/
#839430000000
1!
1'
1/
#839440000000
0!
0'
0/
#839450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#839460000000
0!
0'
0/
#839470000000
1!
1'
1/
#839480000000
0!
1"
0'
1(
0/
10
#839490000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#839500000000
0!
1$
0'
1+
0/
#839510000000
1!
1'
1/
#839520000000
0!
0'
0/
#839530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#839540000000
0!
0'
0/
#839550000000
1!
1'
1/
#839560000000
0!
0'
0/
#839570000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#839580000000
0!
0'
0/
#839590000000
1!
1'
1/
#839600000000
0!
0'
0/
#839610000000
1!
1'
1/
#839620000000
0!
0'
0/
#839630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#839640000000
0!
0'
0/
#839650000000
1!
1'
1/
#839660000000
0!
0'
0/
#839670000000
1!
1'
1/
#839680000000
0!
0'
0/
#839690000000
1!
1'
1/
#839700000000
0!
0'
0/
#839710000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#839720000000
0!
0'
0/
#839730000000
1!
1'
1/
#839740000000
0!
0'
0/
#839750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#839760000000
0!
0'
0/
#839770000000
1!
1'
1/
#839780000000
0!
0'
0/
#839790000000
#839800000000
1!
1'
1/
#839810000000
0!
0'
0/
#839820000000
1!
1'
1/
#839830000000
0!
1"
0'
1(
0/
10
#839840000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#839850000000
0!
0'
0/
#839860000000
1!
1'
1/
#839870000000
0!
0'
0/
#839880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#839890000000
0!
0'
0/
#839900000000
1!
1'
1/
#839910000000
0!
1"
0'
1(
0/
10
#839920000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#839930000000
0!
1$
0'
1+
0/
#839940000000
1!
1'
1/
#839950000000
0!
0'
0/
#839960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#839970000000
0!
0'
0/
#839980000000
1!
1'
1/
#839990000000
0!
0'
0/
#840000000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#840010000000
0!
0'
0/
#840020000000
1!
1'
1/
#840030000000
0!
0'
0/
#840040000000
1!
1'
1/
#840050000000
0!
0'
0/
#840060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#840070000000
0!
0'
0/
#840080000000
1!
1'
1/
#840090000000
0!
0'
0/
#840100000000
1!
1'
1/
#840110000000
0!
0'
0/
#840120000000
1!
1'
1/
#840130000000
0!
0'
0/
#840140000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#840150000000
0!
0'
0/
#840160000000
1!
1'
1/
#840170000000
0!
0'
0/
#840180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#840190000000
0!
0'
0/
#840200000000
1!
1'
1/
#840210000000
0!
0'
0/
#840220000000
#840230000000
1!
1'
1/
#840240000000
0!
0'
0/
#840250000000
1!
1'
1/
#840260000000
0!
1"
0'
1(
0/
10
#840270000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#840280000000
0!
0'
0/
#840290000000
1!
1'
1/
#840300000000
0!
0'
0/
#840310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#840320000000
0!
0'
0/
#840330000000
1!
1'
1/
#840340000000
0!
1"
0'
1(
0/
10
#840350000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#840360000000
0!
1$
0'
1+
0/
#840370000000
1!
1'
1/
#840380000000
0!
0'
0/
#840390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#840400000000
0!
0'
0/
#840410000000
1!
1'
1/
#840420000000
0!
0'
0/
#840430000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#840440000000
0!
0'
0/
#840450000000
1!
1'
1/
#840460000000
0!
0'
0/
#840470000000
1!
1'
1/
#840480000000
0!
0'
0/
#840490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#840500000000
0!
0'
0/
#840510000000
1!
1'
1/
#840520000000
0!
0'
0/
#840530000000
1!
1'
1/
#840540000000
0!
0'
0/
#840550000000
1!
1'
1/
#840560000000
0!
0'
0/
#840570000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#840580000000
0!
0'
0/
#840590000000
1!
1'
1/
#840600000000
0!
0'
0/
#840610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#840620000000
0!
0'
0/
#840630000000
1!
1'
1/
#840640000000
0!
0'
0/
#840650000000
#840660000000
1!
1'
1/
#840670000000
0!
0'
0/
#840680000000
1!
1'
1/
#840690000000
0!
1"
0'
1(
0/
10
#840700000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#840710000000
0!
0'
0/
#840720000000
1!
1'
1/
#840730000000
0!
0'
0/
#840740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#840750000000
0!
0'
0/
#840760000000
1!
1'
1/
#840770000000
0!
1"
0'
1(
0/
10
#840780000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#840790000000
0!
1$
0'
1+
0/
#840800000000
1!
1'
1/
#840810000000
0!
0'
0/
#840820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#840830000000
0!
0'
0/
#840840000000
1!
1'
1/
#840850000000
0!
0'
0/
#840860000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#840870000000
0!
0'
0/
#840880000000
1!
1'
1/
#840890000000
0!
0'
0/
#840900000000
1!
1'
1/
#840910000000
0!
0'
0/
#840920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#840930000000
0!
0'
0/
#840940000000
1!
1'
1/
#840950000000
0!
0'
0/
#840960000000
1!
1'
1/
#840970000000
0!
0'
0/
#840980000000
1!
1'
1/
#840990000000
0!
0'
0/
#841000000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#841010000000
0!
0'
0/
#841020000000
1!
1'
1/
#841030000000
0!
0'
0/
#841040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#841050000000
0!
0'
0/
#841060000000
1!
1'
1/
#841070000000
0!
0'
0/
#841080000000
#841090000000
1!
1'
1/
#841100000000
0!
0'
0/
#841110000000
1!
1'
1/
#841120000000
0!
1"
0'
1(
0/
10
#841130000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#841140000000
0!
0'
0/
#841150000000
1!
1'
1/
#841160000000
0!
0'
0/
#841170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#841180000000
0!
0'
0/
#841190000000
1!
1'
1/
#841200000000
0!
1"
0'
1(
0/
10
#841210000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#841220000000
0!
1$
0'
1+
0/
#841230000000
1!
1'
1/
#841240000000
0!
0'
0/
#841250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#841260000000
0!
0'
0/
#841270000000
1!
1'
1/
#841280000000
0!
0'
0/
#841290000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#841300000000
0!
0'
0/
#841310000000
1!
1'
1/
#841320000000
0!
0'
0/
#841330000000
1!
1'
1/
#841340000000
0!
0'
0/
#841350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#841360000000
0!
0'
0/
#841370000000
1!
1'
1/
#841380000000
0!
0'
0/
#841390000000
1!
1'
1/
#841400000000
0!
0'
0/
#841410000000
1!
1'
1/
#841420000000
0!
0'
0/
#841430000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#841440000000
0!
0'
0/
#841450000000
1!
1'
1/
#841460000000
0!
0'
0/
#841470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#841480000000
0!
0'
0/
#841490000000
1!
1'
1/
#841500000000
0!
0'
0/
#841510000000
#841520000000
1!
1'
1/
#841530000000
0!
0'
0/
#841540000000
1!
1'
1/
#841550000000
0!
1"
0'
1(
0/
10
#841560000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#841570000000
0!
0'
0/
#841580000000
1!
1'
1/
#841590000000
0!
0'
0/
#841600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#841610000000
0!
0'
0/
#841620000000
1!
1'
1/
#841630000000
0!
1"
0'
1(
0/
10
#841640000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#841650000000
0!
1$
0'
1+
0/
#841660000000
1!
1'
1/
#841670000000
0!
0'
0/
#841680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#841690000000
0!
0'
0/
#841700000000
1!
1'
1/
#841710000000
0!
0'
0/
#841720000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#841730000000
0!
0'
0/
#841740000000
1!
1'
1/
#841750000000
0!
0'
0/
#841760000000
1!
1'
1/
#841770000000
0!
0'
0/
#841780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#841790000000
0!
0'
0/
#841800000000
1!
1'
1/
#841810000000
0!
0'
0/
#841820000000
1!
1'
1/
#841830000000
0!
0'
0/
#841840000000
1!
1'
1/
#841850000000
0!
0'
0/
#841860000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#841870000000
0!
0'
0/
#841880000000
1!
1'
1/
#841890000000
0!
0'
0/
#841900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#841910000000
0!
0'
0/
#841920000000
1!
1'
1/
#841930000000
0!
0'
0/
#841940000000
#841950000000
1!
1'
1/
#841960000000
0!
0'
0/
#841970000000
1!
1'
1/
#841980000000
0!
1"
0'
1(
0/
10
#841990000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#842000000000
0!
0'
0/
#842010000000
1!
1'
1/
#842020000000
0!
0'
0/
#842030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#842040000000
0!
0'
0/
#842050000000
1!
1'
1/
#842060000000
0!
1"
0'
1(
0/
10
#842070000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#842080000000
0!
1$
0'
1+
0/
#842090000000
1!
1'
1/
#842100000000
0!
0'
0/
#842110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#842120000000
0!
0'
0/
#842130000000
1!
1'
1/
#842140000000
0!
0'
0/
#842150000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#842160000000
0!
0'
0/
#842170000000
1!
1'
1/
#842180000000
0!
0'
0/
#842190000000
1!
1'
1/
#842200000000
0!
0'
0/
#842210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#842220000000
0!
0'
0/
#842230000000
1!
1'
1/
#842240000000
0!
0'
0/
#842250000000
1!
1'
1/
#842260000000
0!
0'
0/
#842270000000
1!
1'
1/
#842280000000
0!
0'
0/
#842290000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#842300000000
0!
0'
0/
#842310000000
1!
1'
1/
#842320000000
0!
0'
0/
#842330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#842340000000
0!
0'
0/
#842350000000
1!
1'
1/
#842360000000
0!
0'
0/
#842370000000
#842380000000
1!
1'
1/
#842390000000
0!
0'
0/
#842400000000
1!
1'
1/
#842410000000
0!
1"
0'
1(
0/
10
#842420000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#842430000000
0!
0'
0/
#842440000000
1!
1'
1/
#842450000000
0!
0'
0/
#842460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#842470000000
0!
0'
0/
#842480000000
1!
1'
1/
#842490000000
0!
1"
0'
1(
0/
10
#842500000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#842510000000
0!
1$
0'
1+
0/
#842520000000
1!
1'
1/
#842530000000
0!
0'
0/
#842540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#842550000000
0!
0'
0/
#842560000000
1!
1'
1/
#842570000000
0!
0'
0/
#842580000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#842590000000
0!
0'
0/
#842600000000
1!
1'
1/
#842610000000
0!
0'
0/
#842620000000
1!
1'
1/
#842630000000
0!
0'
0/
#842640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#842650000000
0!
0'
0/
#842660000000
1!
1'
1/
#842670000000
0!
0'
0/
#842680000000
1!
1'
1/
#842690000000
0!
0'
0/
#842700000000
1!
1'
1/
#842710000000
0!
0'
0/
#842720000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#842730000000
0!
0'
0/
#842740000000
1!
1'
1/
#842750000000
0!
0'
0/
#842760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#842770000000
0!
0'
0/
#842780000000
1!
1'
1/
#842790000000
0!
0'
0/
#842800000000
#842810000000
1!
1'
1/
#842820000000
0!
0'
0/
#842830000000
1!
1'
1/
#842840000000
0!
1"
0'
1(
0/
10
#842850000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#842860000000
0!
0'
0/
#842870000000
1!
1'
1/
#842880000000
0!
0'
0/
#842890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#842900000000
0!
0'
0/
#842910000000
1!
1'
1/
#842920000000
0!
1"
0'
1(
0/
10
#842930000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#842940000000
0!
1$
0'
1+
0/
#842950000000
1!
1'
1/
#842960000000
0!
0'
0/
#842970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#842980000000
0!
0'
0/
#842990000000
1!
1'
1/
#843000000000
0!
0'
0/
#843010000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#843020000000
0!
0'
0/
#843030000000
1!
1'
1/
#843040000000
0!
0'
0/
#843050000000
1!
1'
1/
#843060000000
0!
0'
0/
#843070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#843080000000
0!
0'
0/
#843090000000
1!
1'
1/
#843100000000
0!
0'
0/
#843110000000
1!
1'
1/
#843120000000
0!
0'
0/
#843130000000
1!
1'
1/
#843140000000
0!
0'
0/
#843150000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#843160000000
0!
0'
0/
#843170000000
1!
1'
1/
#843180000000
0!
0'
0/
#843190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#843200000000
0!
0'
0/
#843210000000
1!
1'
1/
#843220000000
0!
0'
0/
#843230000000
#843240000000
1!
1'
1/
#843250000000
0!
0'
0/
#843260000000
1!
1'
1/
#843270000000
0!
1"
0'
1(
0/
10
#843280000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#843290000000
0!
0'
0/
#843300000000
1!
1'
1/
#843310000000
0!
0'
0/
#843320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#843330000000
0!
0'
0/
#843340000000
1!
1'
1/
#843350000000
0!
1"
0'
1(
0/
10
#843360000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#843370000000
0!
1$
0'
1+
0/
#843380000000
1!
1'
1/
#843390000000
0!
0'
0/
#843400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#843410000000
0!
0'
0/
#843420000000
1!
1'
1/
#843430000000
0!
0'
0/
#843440000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#843450000000
0!
0'
0/
#843460000000
1!
1'
1/
#843470000000
0!
0'
0/
#843480000000
1!
1'
1/
#843490000000
0!
0'
0/
#843500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#843510000000
0!
0'
0/
#843520000000
1!
1'
1/
#843530000000
0!
0'
0/
#843540000000
1!
1'
1/
#843550000000
0!
0'
0/
#843560000000
1!
1'
1/
#843570000000
0!
0'
0/
#843580000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#843590000000
0!
0'
0/
#843600000000
1!
1'
1/
#843610000000
0!
0'
0/
#843620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#843630000000
0!
0'
0/
#843640000000
1!
1'
1/
#843650000000
0!
0'
0/
#843660000000
#843670000000
1!
1'
1/
#843680000000
0!
0'
0/
#843690000000
1!
1'
1/
#843700000000
0!
1"
0'
1(
0/
10
#843710000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#843720000000
0!
0'
0/
#843730000000
1!
1'
1/
#843740000000
0!
0'
0/
#843750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#843760000000
0!
0'
0/
#843770000000
1!
1'
1/
#843780000000
0!
1"
0'
1(
0/
10
#843790000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#843800000000
0!
1$
0'
1+
0/
#843810000000
1!
1'
1/
#843820000000
0!
0'
0/
#843830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#843840000000
0!
0'
0/
#843850000000
1!
1'
1/
#843860000000
0!
0'
0/
#843870000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#843880000000
0!
0'
0/
#843890000000
1!
1'
1/
#843900000000
0!
0'
0/
#843910000000
1!
1'
1/
#843920000000
0!
0'
0/
#843930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#843940000000
0!
0'
0/
#843950000000
1!
1'
1/
#843960000000
0!
0'
0/
#843970000000
1!
1'
1/
#843980000000
0!
0'
0/
#843990000000
1!
1'
1/
#844000000000
0!
0'
0/
#844010000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#844020000000
0!
0'
0/
#844030000000
1!
1'
1/
#844040000000
0!
0'
0/
#844050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#844060000000
0!
0'
0/
#844070000000
1!
1'
1/
#844080000000
0!
0'
0/
#844090000000
#844100000000
1!
1'
1/
#844110000000
0!
0'
0/
#844120000000
1!
1'
1/
#844130000000
0!
1"
0'
1(
0/
10
#844140000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#844150000000
0!
0'
0/
#844160000000
1!
1'
1/
#844170000000
0!
0'
0/
#844180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#844190000000
0!
0'
0/
#844200000000
1!
1'
1/
#844210000000
0!
1"
0'
1(
0/
10
#844220000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#844230000000
0!
1$
0'
1+
0/
#844240000000
1!
1'
1/
#844250000000
0!
0'
0/
#844260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#844270000000
0!
0'
0/
#844280000000
1!
1'
1/
#844290000000
0!
0'
0/
#844300000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#844310000000
0!
0'
0/
#844320000000
1!
1'
1/
#844330000000
0!
0'
0/
#844340000000
1!
1'
1/
#844350000000
0!
0'
0/
#844360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#844370000000
0!
0'
0/
#844380000000
1!
1'
1/
#844390000000
0!
0'
0/
#844400000000
1!
1'
1/
#844410000000
0!
0'
0/
#844420000000
1!
1'
1/
#844430000000
0!
0'
0/
#844440000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#844450000000
0!
0'
0/
#844460000000
1!
1'
1/
#844470000000
0!
0'
0/
#844480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#844490000000
0!
0'
0/
#844500000000
1!
1'
1/
#844510000000
0!
0'
0/
#844520000000
#844530000000
1!
1'
1/
#844540000000
0!
0'
0/
#844550000000
1!
1'
1/
#844560000000
0!
1"
0'
1(
0/
10
#844570000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#844580000000
0!
0'
0/
#844590000000
1!
1'
1/
#844600000000
0!
0'
0/
#844610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#844620000000
0!
0'
0/
#844630000000
1!
1'
1/
#844640000000
0!
1"
0'
1(
0/
10
#844650000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#844660000000
0!
1$
0'
1+
0/
#844670000000
1!
1'
1/
#844680000000
0!
0'
0/
#844690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#844700000000
0!
0'
0/
#844710000000
1!
1'
1/
#844720000000
0!
0'
0/
#844730000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#844740000000
0!
0'
0/
#844750000000
1!
1'
1/
#844760000000
0!
0'
0/
#844770000000
1!
1'
1/
#844780000000
0!
0'
0/
#844790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#844800000000
0!
0'
0/
#844810000000
1!
1'
1/
#844820000000
0!
0'
0/
#844830000000
1!
1'
1/
#844840000000
0!
0'
0/
#844850000000
1!
1'
1/
#844860000000
0!
0'
0/
#844870000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#844880000000
0!
0'
0/
#844890000000
1!
1'
1/
#844900000000
0!
0'
0/
#844910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#844920000000
0!
0'
0/
#844930000000
1!
1'
1/
#844940000000
0!
0'
0/
#844950000000
#844960000000
1!
1'
1/
#844970000000
0!
0'
0/
#844980000000
1!
1'
1/
#844990000000
0!
1"
0'
1(
0/
10
#845000000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#845010000000
0!
0'
0/
#845020000000
1!
1'
1/
#845030000000
0!
0'
0/
#845040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#845050000000
0!
0'
0/
#845060000000
1!
1'
1/
#845070000000
0!
1"
0'
1(
0/
10
#845080000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#845090000000
0!
1$
0'
1+
0/
#845100000000
1!
1'
1/
#845110000000
0!
0'
0/
#845120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#845130000000
0!
0'
0/
#845140000000
1!
1'
1/
#845150000000
0!
0'
0/
#845160000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#845170000000
0!
0'
0/
#845180000000
1!
1'
1/
#845190000000
0!
0'
0/
#845200000000
1!
1'
1/
#845210000000
0!
0'
0/
#845220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#845230000000
0!
0'
0/
#845240000000
1!
1'
1/
#845250000000
0!
0'
0/
#845260000000
1!
1'
1/
#845270000000
0!
0'
0/
#845280000000
1!
1'
1/
#845290000000
0!
0'
0/
#845300000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#845310000000
0!
0'
0/
#845320000000
1!
1'
1/
#845330000000
0!
0'
0/
#845340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#845350000000
0!
0'
0/
#845360000000
1!
1'
1/
#845370000000
0!
0'
0/
#845380000000
#845390000000
1!
1'
1/
#845400000000
0!
0'
0/
#845410000000
1!
1'
1/
#845420000000
0!
1"
0'
1(
0/
10
#845430000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#845440000000
0!
0'
0/
#845450000000
1!
1'
1/
#845460000000
0!
0'
0/
#845470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#845480000000
0!
0'
0/
#845490000000
1!
1'
1/
#845500000000
0!
1"
0'
1(
0/
10
#845510000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#845520000000
0!
1$
0'
1+
0/
#845530000000
1!
1'
1/
#845540000000
0!
0'
0/
#845550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#845560000000
0!
0'
0/
#845570000000
1!
1'
1/
#845580000000
0!
0'
0/
#845590000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#845600000000
0!
0'
0/
#845610000000
1!
1'
1/
#845620000000
0!
0'
0/
#845630000000
1!
1'
1/
#845640000000
0!
0'
0/
#845650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#845660000000
0!
0'
0/
#845670000000
1!
1'
1/
#845680000000
0!
0'
0/
#845690000000
1!
1'
1/
#845700000000
0!
0'
0/
#845710000000
1!
1'
1/
#845720000000
0!
0'
0/
#845730000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#845740000000
0!
0'
0/
#845750000000
1!
1'
1/
#845760000000
0!
0'
0/
#845770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#845780000000
0!
0'
0/
#845790000000
1!
1'
1/
#845800000000
0!
0'
0/
#845810000000
#845820000000
1!
1'
1/
#845830000000
0!
0'
0/
#845840000000
1!
1'
1/
#845850000000
0!
1"
0'
1(
0/
10
#845860000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#845870000000
0!
0'
0/
#845880000000
1!
1'
1/
#845890000000
0!
0'
0/
#845900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#845910000000
0!
0'
0/
#845920000000
1!
1'
1/
#845930000000
0!
1"
0'
1(
0/
10
#845940000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#845950000000
0!
1$
0'
1+
0/
#845960000000
1!
1'
1/
#845970000000
0!
0'
0/
#845980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#845990000000
0!
0'
0/
#846000000000
1!
1'
1/
#846010000000
0!
0'
0/
#846020000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#846030000000
0!
0'
0/
#846040000000
1!
1'
1/
#846050000000
0!
0'
0/
#846060000000
1!
1'
1/
#846070000000
0!
0'
0/
#846080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#846090000000
0!
0'
0/
#846100000000
1!
1'
1/
#846110000000
0!
0'
0/
#846120000000
1!
1'
1/
#846130000000
0!
0'
0/
#846140000000
1!
1'
1/
#846150000000
0!
0'
0/
#846160000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#846170000000
0!
0'
0/
#846180000000
1!
1'
1/
#846190000000
0!
0'
0/
#846200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#846210000000
0!
0'
0/
#846220000000
1!
1'
1/
#846230000000
0!
0'
0/
#846240000000
#846250000000
1!
1'
1/
#846260000000
0!
0'
0/
#846270000000
1!
1'
1/
#846280000000
0!
1"
0'
1(
0/
10
#846290000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#846300000000
0!
0'
0/
#846310000000
1!
1'
1/
#846320000000
0!
0'
0/
#846330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#846340000000
0!
0'
0/
#846350000000
1!
1'
1/
#846360000000
0!
1"
0'
1(
0/
10
#846370000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#846380000000
0!
1$
0'
1+
0/
#846390000000
1!
1'
1/
#846400000000
0!
0'
0/
#846410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#846420000000
0!
0'
0/
#846430000000
1!
1'
1/
#846440000000
0!
0'
0/
#846450000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#846460000000
0!
0'
0/
#846470000000
1!
1'
1/
#846480000000
0!
0'
0/
#846490000000
1!
1'
1/
#846500000000
0!
0'
0/
#846510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#846520000000
0!
0'
0/
#846530000000
1!
1'
1/
#846540000000
0!
0'
0/
#846550000000
1!
1'
1/
#846560000000
0!
0'
0/
#846570000000
1!
1'
1/
#846580000000
0!
0'
0/
#846590000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#846600000000
0!
0'
0/
#846610000000
1!
1'
1/
#846620000000
0!
0'
0/
#846630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#846640000000
0!
0'
0/
#846650000000
1!
1'
1/
#846660000000
0!
0'
0/
#846670000000
#846680000000
1!
1'
1/
#846690000000
0!
0'
0/
#846700000000
1!
1'
1/
#846710000000
0!
1"
0'
1(
0/
10
#846720000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#846730000000
0!
0'
0/
#846740000000
1!
1'
1/
#846750000000
0!
0'
0/
#846760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#846770000000
0!
0'
0/
#846780000000
1!
1'
1/
#846790000000
0!
1"
0'
1(
0/
10
#846800000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#846810000000
0!
1$
0'
1+
0/
#846820000000
1!
1'
1/
#846830000000
0!
0'
0/
#846840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#846850000000
0!
0'
0/
#846860000000
1!
1'
1/
#846870000000
0!
0'
0/
#846880000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#846890000000
0!
0'
0/
#846900000000
1!
1'
1/
#846910000000
0!
0'
0/
#846920000000
1!
1'
1/
#846930000000
0!
0'
0/
#846940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#846950000000
0!
0'
0/
#846960000000
1!
1'
1/
#846970000000
0!
0'
0/
#846980000000
1!
1'
1/
#846990000000
0!
0'
0/
#847000000000
1!
1'
1/
#847010000000
0!
0'
0/
#847020000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#847030000000
0!
0'
0/
#847040000000
1!
1'
1/
#847050000000
0!
0'
0/
#847060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#847070000000
0!
0'
0/
#847080000000
1!
1'
1/
#847090000000
0!
0'
0/
#847100000000
#847110000000
1!
1'
1/
#847120000000
0!
0'
0/
#847130000000
1!
1'
1/
#847140000000
0!
1"
0'
1(
0/
10
#847150000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#847160000000
0!
0'
0/
#847170000000
1!
1'
1/
#847180000000
0!
0'
0/
#847190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#847200000000
0!
0'
0/
#847210000000
1!
1'
1/
#847220000000
0!
1"
0'
1(
0/
10
#847230000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#847240000000
0!
1$
0'
1+
0/
#847250000000
1!
1'
1/
#847260000000
0!
0'
0/
#847270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#847280000000
0!
0'
0/
#847290000000
1!
1'
1/
#847300000000
0!
0'
0/
#847310000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#847320000000
0!
0'
0/
#847330000000
1!
1'
1/
#847340000000
0!
0'
0/
#847350000000
1!
1'
1/
#847360000000
0!
0'
0/
#847370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#847380000000
0!
0'
0/
#847390000000
1!
1'
1/
#847400000000
0!
0'
0/
#847410000000
1!
1'
1/
#847420000000
0!
0'
0/
#847430000000
1!
1'
1/
#847440000000
0!
0'
0/
#847450000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#847460000000
0!
0'
0/
#847470000000
1!
1'
1/
#847480000000
0!
0'
0/
#847490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#847500000000
0!
0'
0/
#847510000000
1!
1'
1/
#847520000000
0!
0'
0/
#847530000000
#847540000000
1!
1'
1/
#847550000000
0!
0'
0/
#847560000000
1!
1'
1/
#847570000000
0!
1"
0'
1(
0/
10
#847580000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#847590000000
0!
0'
0/
#847600000000
1!
1'
1/
#847610000000
0!
0'
0/
#847620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#847630000000
0!
0'
0/
#847640000000
1!
1'
1/
#847650000000
0!
1"
0'
1(
0/
10
#847660000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#847670000000
0!
1$
0'
1+
0/
#847680000000
1!
1'
1/
#847690000000
0!
0'
0/
#847700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#847710000000
0!
0'
0/
#847720000000
1!
1'
1/
#847730000000
0!
0'
0/
#847740000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#847750000000
0!
0'
0/
#847760000000
1!
1'
1/
#847770000000
0!
0'
0/
#847780000000
1!
1'
1/
#847790000000
0!
0'
0/
#847800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#847810000000
0!
0'
0/
#847820000000
1!
1'
1/
#847830000000
0!
0'
0/
#847840000000
1!
1'
1/
#847850000000
0!
0'
0/
#847860000000
1!
1'
1/
#847870000000
0!
0'
0/
#847880000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#847890000000
0!
0'
0/
#847900000000
1!
1'
1/
#847910000000
0!
0'
0/
#847920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#847930000000
0!
0'
0/
#847940000000
1!
1'
1/
#847950000000
0!
0'
0/
#847960000000
#847970000000
1!
1'
1/
#847980000000
0!
0'
0/
#847990000000
1!
1'
1/
#848000000000
0!
1"
0'
1(
0/
10
#848010000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#848020000000
0!
0'
0/
#848030000000
1!
1'
1/
#848040000000
0!
0'
0/
#848050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#848060000000
0!
0'
0/
#848070000000
1!
1'
1/
#848080000000
0!
1"
0'
1(
0/
10
#848090000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#848100000000
0!
1$
0'
1+
0/
#848110000000
1!
1'
1/
#848120000000
0!
0'
0/
#848130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#848140000000
0!
0'
0/
#848150000000
1!
1'
1/
#848160000000
0!
0'
0/
#848170000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#848180000000
0!
0'
0/
#848190000000
1!
1'
1/
#848200000000
0!
0'
0/
#848210000000
1!
1'
1/
#848220000000
0!
0'
0/
#848230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#848240000000
0!
0'
0/
#848250000000
1!
1'
1/
#848260000000
0!
0'
0/
#848270000000
1!
1'
1/
#848280000000
0!
0'
0/
#848290000000
1!
1'
1/
#848300000000
0!
0'
0/
#848310000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#848320000000
0!
0'
0/
#848330000000
1!
1'
1/
#848340000000
0!
0'
0/
#848350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#848360000000
0!
0'
0/
#848370000000
1!
1'
1/
#848380000000
0!
0'
0/
#848390000000
#848400000000
1!
1'
1/
#848410000000
0!
0'
0/
#848420000000
1!
1'
1/
#848430000000
0!
1"
0'
1(
0/
10
#848440000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#848450000000
0!
0'
0/
#848460000000
1!
1'
1/
#848470000000
0!
0'
0/
#848480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#848490000000
0!
0'
0/
#848500000000
1!
1'
1/
#848510000000
0!
1"
0'
1(
0/
10
#848520000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#848530000000
0!
1$
0'
1+
0/
#848540000000
1!
1'
1/
#848550000000
0!
0'
0/
#848560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#848570000000
0!
0'
0/
#848580000000
1!
1'
1/
#848590000000
0!
0'
0/
#848600000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#848610000000
0!
0'
0/
#848620000000
1!
1'
1/
#848630000000
0!
0'
0/
#848640000000
1!
1'
1/
#848650000000
0!
0'
0/
#848660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#848670000000
0!
0'
0/
#848680000000
1!
1'
1/
#848690000000
0!
0'
0/
#848700000000
1!
1'
1/
#848710000000
0!
0'
0/
#848720000000
1!
1'
1/
#848730000000
0!
0'
0/
#848740000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#848750000000
0!
0'
0/
#848760000000
1!
1'
1/
#848770000000
0!
0'
0/
#848780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#848790000000
0!
0'
0/
#848800000000
1!
1'
1/
#848810000000
0!
0'
0/
#848820000000
#848830000000
1!
1'
1/
#848840000000
0!
0'
0/
#848850000000
1!
1'
1/
#848860000000
0!
1"
0'
1(
0/
10
#848870000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#848880000000
0!
0'
0/
#848890000000
1!
1'
1/
#848900000000
0!
0'
0/
#848910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#848920000000
0!
0'
0/
#848930000000
1!
1'
1/
#848940000000
0!
1"
0'
1(
0/
10
#848950000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#848960000000
0!
1$
0'
1+
0/
#848970000000
1!
1'
1/
#848980000000
0!
0'
0/
#848990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#849000000000
0!
0'
0/
#849010000000
1!
1'
1/
#849020000000
0!
0'
0/
#849030000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#849040000000
0!
0'
0/
#849050000000
1!
1'
1/
#849060000000
0!
0'
0/
#849070000000
1!
1'
1/
#849080000000
0!
0'
0/
#849090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#849100000000
0!
0'
0/
#849110000000
1!
1'
1/
#849120000000
0!
0'
0/
#849130000000
1!
1'
1/
#849140000000
0!
0'
0/
#849150000000
1!
1'
1/
#849160000000
0!
0'
0/
#849170000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#849180000000
0!
0'
0/
#849190000000
1!
1'
1/
#849200000000
0!
0'
0/
#849210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#849220000000
0!
0'
0/
#849230000000
1!
1'
1/
#849240000000
0!
0'
0/
#849250000000
#849260000000
1!
1'
1/
#849270000000
0!
0'
0/
#849280000000
1!
1'
1/
#849290000000
0!
1"
0'
1(
0/
10
#849300000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#849310000000
0!
0'
0/
#849320000000
1!
1'
1/
#849330000000
0!
0'
0/
#849340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#849350000000
0!
0'
0/
#849360000000
1!
1'
1/
#849370000000
0!
1"
0'
1(
0/
10
#849380000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#849390000000
0!
1$
0'
1+
0/
#849400000000
1!
1'
1/
#849410000000
0!
0'
0/
#849420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#849430000000
0!
0'
0/
#849440000000
1!
1'
1/
#849450000000
0!
0'
0/
#849460000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#849470000000
0!
0'
0/
#849480000000
1!
1'
1/
#849490000000
0!
0'
0/
#849500000000
1!
1'
1/
#849510000000
0!
0'
0/
#849520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#849530000000
0!
0'
0/
#849540000000
1!
1'
1/
#849550000000
0!
0'
0/
#849560000000
1!
1'
1/
#849570000000
0!
0'
0/
#849580000000
1!
1'
1/
#849590000000
0!
0'
0/
#849600000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#849610000000
0!
0'
0/
#849620000000
1!
1'
1/
#849630000000
0!
0'
0/
#849640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#849650000000
0!
0'
0/
#849660000000
1!
1'
1/
#849670000000
0!
0'
0/
#849680000000
#849690000000
1!
1'
1/
#849700000000
0!
0'
0/
#849710000000
1!
1'
1/
#849720000000
0!
1"
0'
1(
0/
10
#849730000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#849740000000
0!
0'
0/
#849750000000
1!
1'
1/
#849760000000
0!
0'
0/
#849770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#849780000000
0!
0'
0/
#849790000000
1!
1'
1/
#849800000000
0!
1"
0'
1(
0/
10
#849810000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#849820000000
0!
1$
0'
1+
0/
#849830000000
1!
1'
1/
#849840000000
0!
0'
0/
#849850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#849860000000
0!
0'
0/
#849870000000
1!
1'
1/
#849880000000
0!
0'
0/
#849890000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#849900000000
0!
0'
0/
#849910000000
1!
1'
1/
#849920000000
0!
0'
0/
#849930000000
1!
1'
1/
#849940000000
0!
0'
0/
#849950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#849960000000
0!
0'
0/
#849970000000
1!
1'
1/
#849980000000
0!
0'
0/
#849990000000
1!
1'
1/
#850000000000
0!
0'
0/
#850010000000
1!
1'
1/
#850020000000
0!
0'
0/
#850030000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#850040000000
0!
0'
0/
#850050000000
1!
1'
1/
#850060000000
0!
0'
0/
#850070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#850080000000
0!
0'
0/
#850090000000
1!
1'
1/
#850100000000
0!
0'
0/
#850110000000
#850120000000
1!
1'
1/
#850130000000
0!
0'
0/
#850140000000
1!
1'
1/
#850150000000
0!
1"
0'
1(
0/
10
#850160000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#850170000000
0!
0'
0/
#850180000000
1!
1'
1/
#850190000000
0!
0'
0/
#850200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#850210000000
0!
0'
0/
#850220000000
1!
1'
1/
#850230000000
0!
1"
0'
1(
0/
10
#850240000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#850250000000
0!
1$
0'
1+
0/
#850260000000
1!
1'
1/
#850270000000
0!
0'
0/
#850280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#850290000000
0!
0'
0/
#850300000000
1!
1'
1/
#850310000000
0!
0'
0/
#850320000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#850330000000
0!
0'
0/
#850340000000
1!
1'
1/
#850350000000
0!
0'
0/
#850360000000
1!
1'
1/
#850370000000
0!
0'
0/
#850380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#850390000000
0!
0'
0/
#850400000000
1!
1'
1/
#850410000000
0!
0'
0/
#850420000000
1!
1'
1/
#850430000000
0!
0'
0/
#850440000000
1!
1'
1/
#850450000000
0!
0'
0/
#850460000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#850470000000
0!
0'
0/
#850480000000
1!
1'
1/
#850490000000
0!
0'
0/
#850500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#850510000000
0!
0'
0/
#850520000000
1!
1'
1/
#850530000000
0!
0'
0/
#850540000000
#850550000000
1!
1'
1/
#850560000000
0!
0'
0/
#850570000000
1!
1'
1/
#850580000000
0!
1"
0'
1(
0/
10
#850590000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#850600000000
0!
0'
0/
#850610000000
1!
1'
1/
#850620000000
0!
0'
0/
#850630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#850640000000
0!
0'
0/
#850650000000
1!
1'
1/
#850660000000
0!
1"
0'
1(
0/
10
#850670000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#850680000000
0!
1$
0'
1+
0/
#850690000000
1!
1'
1/
#850700000000
0!
0'
0/
#850710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#850720000000
0!
0'
0/
#850730000000
1!
1'
1/
#850740000000
0!
0'
0/
#850750000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#850760000000
0!
0'
0/
#850770000000
1!
1'
1/
#850780000000
0!
0'
0/
#850790000000
1!
1'
1/
#850800000000
0!
0'
0/
#850810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#850820000000
0!
0'
0/
#850830000000
1!
1'
1/
#850840000000
0!
0'
0/
#850850000000
1!
1'
1/
#850860000000
0!
0'
0/
#850870000000
1!
1'
1/
#850880000000
0!
0'
0/
#850890000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#850900000000
0!
0'
0/
#850910000000
1!
1'
1/
#850920000000
0!
0'
0/
#850930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#850940000000
0!
0'
0/
#850950000000
1!
1'
1/
#850960000000
0!
0'
0/
#850970000000
#850980000000
1!
1'
1/
#850990000000
0!
0'
0/
#851000000000
1!
1'
1/
#851010000000
0!
1"
0'
1(
0/
10
#851020000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#851030000000
0!
0'
0/
#851040000000
1!
1'
1/
#851050000000
0!
0'
0/
#851060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#851070000000
0!
0'
0/
#851080000000
1!
1'
1/
#851090000000
0!
1"
0'
1(
0/
10
#851100000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#851110000000
0!
1$
0'
1+
0/
#851120000000
1!
1'
1/
#851130000000
0!
0'
0/
#851140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#851150000000
0!
0'
0/
#851160000000
1!
1'
1/
#851170000000
0!
0'
0/
#851180000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#851190000000
0!
0'
0/
#851200000000
1!
1'
1/
#851210000000
0!
0'
0/
#851220000000
1!
1'
1/
#851230000000
0!
0'
0/
#851240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#851250000000
0!
0'
0/
#851260000000
1!
1'
1/
#851270000000
0!
0'
0/
#851280000000
1!
1'
1/
#851290000000
0!
0'
0/
#851300000000
1!
1'
1/
#851310000000
0!
0'
0/
#851320000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#851330000000
0!
0'
0/
#851340000000
1!
1'
1/
#851350000000
0!
0'
0/
#851360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#851370000000
0!
0'
0/
#851380000000
1!
1'
1/
#851390000000
0!
0'
0/
#851400000000
#851410000000
1!
1'
1/
#851420000000
0!
0'
0/
#851430000000
1!
1'
1/
#851440000000
0!
1"
0'
1(
0/
10
#851450000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#851460000000
0!
0'
0/
#851470000000
1!
1'
1/
#851480000000
0!
0'
0/
#851490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#851500000000
0!
0'
0/
#851510000000
1!
1'
1/
#851520000000
0!
1"
0'
1(
0/
10
#851530000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#851540000000
0!
1$
0'
1+
0/
#851550000000
1!
1'
1/
#851560000000
0!
0'
0/
#851570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#851580000000
0!
0'
0/
#851590000000
1!
1'
1/
#851600000000
0!
0'
0/
#851610000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#851620000000
0!
0'
0/
#851630000000
1!
1'
1/
#851640000000
0!
0'
0/
#851650000000
1!
1'
1/
#851660000000
0!
0'
0/
#851670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#851680000000
0!
0'
0/
#851690000000
1!
1'
1/
#851700000000
0!
0'
0/
#851710000000
1!
1'
1/
#851720000000
0!
0'
0/
#851730000000
1!
1'
1/
#851740000000
0!
0'
0/
#851750000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#851760000000
0!
0'
0/
#851770000000
1!
1'
1/
#851780000000
0!
0'
0/
#851790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#851800000000
0!
0'
0/
#851810000000
1!
1'
1/
#851820000000
0!
0'
0/
#851830000000
#851840000000
1!
1'
1/
#851850000000
0!
0'
0/
#851860000000
1!
1'
1/
#851870000000
0!
1"
0'
1(
0/
10
#851880000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#851890000000
0!
0'
0/
#851900000000
1!
1'
1/
#851910000000
0!
0'
0/
#851920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#851930000000
0!
0'
0/
#851940000000
1!
1'
1/
#851950000000
0!
1"
0'
1(
0/
10
#851960000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#851970000000
0!
1$
0'
1+
0/
#851980000000
1!
1'
1/
#851990000000
0!
0'
0/
#852000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#852010000000
0!
0'
0/
#852020000000
1!
1'
1/
#852030000000
0!
0'
0/
#852040000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#852050000000
0!
0'
0/
#852060000000
1!
1'
1/
#852070000000
0!
0'
0/
#852080000000
1!
1'
1/
#852090000000
0!
0'
0/
#852100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#852110000000
0!
0'
0/
#852120000000
1!
1'
1/
#852130000000
0!
0'
0/
#852140000000
1!
1'
1/
#852150000000
0!
0'
0/
#852160000000
1!
1'
1/
#852170000000
0!
0'
0/
#852180000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#852190000000
0!
0'
0/
#852200000000
1!
1'
1/
#852210000000
0!
0'
0/
#852220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#852230000000
0!
0'
0/
#852240000000
1!
1'
1/
#852250000000
0!
0'
0/
#852260000000
#852270000000
1!
1'
1/
#852280000000
0!
0'
0/
#852290000000
1!
1'
1/
#852300000000
0!
1"
0'
1(
0/
10
#852310000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#852320000000
0!
0'
0/
#852330000000
1!
1'
1/
#852340000000
0!
0'
0/
#852350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#852360000000
0!
0'
0/
#852370000000
1!
1'
1/
#852380000000
0!
1"
0'
1(
0/
10
#852390000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#852400000000
0!
1$
0'
1+
0/
#852410000000
1!
1'
1/
#852420000000
0!
0'
0/
#852430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#852440000000
0!
0'
0/
#852450000000
1!
1'
1/
#852460000000
0!
0'
0/
#852470000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#852480000000
0!
0'
0/
#852490000000
1!
1'
1/
#852500000000
0!
0'
0/
#852510000000
1!
1'
1/
#852520000000
0!
0'
0/
#852530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#852540000000
0!
0'
0/
#852550000000
1!
1'
1/
#852560000000
0!
0'
0/
#852570000000
1!
1'
1/
#852580000000
0!
0'
0/
#852590000000
1!
1'
1/
#852600000000
0!
0'
0/
#852610000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#852620000000
0!
0'
0/
#852630000000
1!
1'
1/
#852640000000
0!
0'
0/
#852650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#852660000000
0!
0'
0/
#852670000000
1!
1'
1/
#852680000000
0!
0'
0/
#852690000000
#852700000000
1!
1'
1/
#852710000000
0!
0'
0/
#852720000000
1!
1'
1/
#852730000000
0!
1"
0'
1(
0/
10
#852740000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#852750000000
0!
0'
0/
#852760000000
1!
1'
1/
#852770000000
0!
0'
0/
#852780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#852790000000
0!
0'
0/
#852800000000
1!
1'
1/
#852810000000
0!
1"
0'
1(
0/
10
#852820000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#852830000000
0!
1$
0'
1+
0/
#852840000000
1!
1'
1/
#852850000000
0!
0'
0/
#852860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#852870000000
0!
0'
0/
#852880000000
1!
1'
1/
#852890000000
0!
0'
0/
#852900000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#852910000000
0!
0'
0/
#852920000000
1!
1'
1/
#852930000000
0!
0'
0/
#852940000000
1!
1'
1/
#852950000000
0!
0'
0/
#852960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#852970000000
0!
0'
0/
#852980000000
1!
1'
1/
#852990000000
0!
0'
0/
#853000000000
1!
1'
1/
#853010000000
0!
0'
0/
#853020000000
1!
1'
1/
#853030000000
0!
0'
0/
#853040000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#853050000000
0!
0'
0/
#853060000000
1!
1'
1/
#853070000000
0!
0'
0/
#853080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#853090000000
0!
0'
0/
#853100000000
1!
1'
1/
#853110000000
0!
0'
0/
#853120000000
#853130000000
1!
1'
1/
#853140000000
0!
0'
0/
#853150000000
1!
1'
1/
#853160000000
0!
1"
0'
1(
0/
10
#853170000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#853180000000
0!
0'
0/
#853190000000
1!
1'
1/
#853200000000
0!
0'
0/
#853210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#853220000000
0!
0'
0/
#853230000000
1!
1'
1/
#853240000000
0!
1"
0'
1(
0/
10
#853250000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#853260000000
0!
1$
0'
1+
0/
#853270000000
1!
1'
1/
#853280000000
0!
0'
0/
#853290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#853300000000
0!
0'
0/
#853310000000
1!
1'
1/
#853320000000
0!
0'
0/
#853330000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#853340000000
0!
0'
0/
#853350000000
1!
1'
1/
#853360000000
0!
0'
0/
#853370000000
1!
1'
1/
#853380000000
0!
0'
0/
#853390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#853400000000
0!
0'
0/
#853410000000
1!
1'
1/
#853420000000
0!
0'
0/
#853430000000
1!
1'
1/
#853440000000
0!
0'
0/
#853450000000
1!
1'
1/
#853460000000
0!
0'
0/
#853470000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#853480000000
0!
0'
0/
#853490000000
1!
1'
1/
#853500000000
0!
0'
0/
#853510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#853520000000
0!
0'
0/
#853530000000
1!
1'
1/
#853540000000
0!
0'
0/
#853550000000
#853560000000
1!
1'
1/
#853570000000
0!
0'
0/
#853580000000
1!
1'
1/
#853590000000
0!
1"
0'
1(
0/
10
#853600000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#853610000000
0!
0'
0/
#853620000000
1!
1'
1/
#853630000000
0!
0'
0/
#853640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#853650000000
0!
0'
0/
#853660000000
1!
1'
1/
#853670000000
0!
1"
0'
1(
0/
10
#853680000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#853690000000
0!
1$
0'
1+
0/
#853700000000
1!
1'
1/
#853710000000
0!
0'
0/
#853720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#853730000000
0!
0'
0/
#853740000000
1!
1'
1/
#853750000000
0!
0'
0/
#853760000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#853770000000
0!
0'
0/
#853780000000
1!
1'
1/
#853790000000
0!
0'
0/
#853800000000
1!
1'
1/
#853810000000
0!
0'
0/
#853820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#853830000000
0!
0'
0/
#853840000000
1!
1'
1/
#853850000000
0!
0'
0/
#853860000000
1!
1'
1/
#853870000000
0!
0'
0/
#853880000000
1!
1'
1/
#853890000000
0!
0'
0/
#853900000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#853910000000
0!
0'
0/
#853920000000
1!
1'
1/
#853930000000
0!
0'
0/
#853940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#853950000000
0!
0'
0/
#853960000000
1!
1'
1/
#853970000000
0!
0'
0/
#853980000000
#853990000000
1!
1'
1/
#854000000000
0!
0'
0/
#854010000000
1!
1'
1/
#854020000000
0!
1"
0'
1(
0/
10
#854030000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#854040000000
0!
0'
0/
#854050000000
1!
1'
1/
#854060000000
0!
0'
0/
#854070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#854080000000
0!
0'
0/
#854090000000
1!
1'
1/
#854100000000
0!
1"
0'
1(
0/
10
#854110000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#854120000000
0!
1$
0'
1+
0/
#854130000000
1!
1'
1/
#854140000000
0!
0'
0/
#854150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#854160000000
0!
0'
0/
#854170000000
1!
1'
1/
#854180000000
0!
0'
0/
#854190000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#854200000000
0!
0'
0/
#854210000000
1!
1'
1/
#854220000000
0!
0'
0/
#854230000000
1!
1'
1/
#854240000000
0!
0'
0/
#854250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#854260000000
0!
0'
0/
#854270000000
1!
1'
1/
#854280000000
0!
0'
0/
#854290000000
1!
1'
1/
#854300000000
0!
0'
0/
#854310000000
1!
1'
1/
#854320000000
0!
0'
0/
#854330000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#854340000000
0!
0'
0/
#854350000000
1!
1'
1/
#854360000000
0!
0'
0/
#854370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#854380000000
0!
0'
0/
#854390000000
1!
1'
1/
#854400000000
0!
0'
0/
#854410000000
#854420000000
1!
1'
1/
#854430000000
0!
0'
0/
#854440000000
1!
1'
1/
#854450000000
0!
1"
0'
1(
0/
10
#854460000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#854470000000
0!
0'
0/
#854480000000
1!
1'
1/
#854490000000
0!
0'
0/
#854500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#854510000000
0!
0'
0/
#854520000000
1!
1'
1/
#854530000000
0!
1"
0'
1(
0/
10
#854540000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#854550000000
0!
1$
0'
1+
0/
#854560000000
1!
1'
1/
#854570000000
0!
0'
0/
#854580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#854590000000
0!
0'
0/
#854600000000
1!
1'
1/
#854610000000
0!
0'
0/
#854620000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#854630000000
0!
0'
0/
#854640000000
1!
1'
1/
#854650000000
0!
0'
0/
#854660000000
1!
1'
1/
#854670000000
0!
0'
0/
#854680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#854690000000
0!
0'
0/
#854700000000
1!
1'
1/
#854710000000
0!
0'
0/
#854720000000
1!
1'
1/
#854730000000
0!
0'
0/
#854740000000
1!
1'
1/
#854750000000
0!
0'
0/
#854760000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#854770000000
0!
0'
0/
#854780000000
1!
1'
1/
#854790000000
0!
0'
0/
#854800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#854810000000
0!
0'
0/
#854820000000
1!
1'
1/
#854830000000
0!
0'
0/
#854840000000
#854850000000
1!
1'
1/
#854860000000
0!
0'
0/
#854870000000
1!
1'
1/
#854880000000
0!
1"
0'
1(
0/
10
#854890000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#854900000000
0!
0'
0/
#854910000000
1!
1'
1/
#854920000000
0!
0'
0/
#854930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#854940000000
0!
0'
0/
#854950000000
1!
1'
1/
#854960000000
0!
1"
0'
1(
0/
10
#854970000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#854980000000
0!
1$
0'
1+
0/
#854990000000
1!
1'
1/
#855000000000
0!
0'
0/
#855010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#855020000000
0!
0'
0/
#855030000000
1!
1'
1/
#855040000000
0!
0'
0/
#855050000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#855060000000
0!
0'
0/
#855070000000
1!
1'
1/
#855080000000
0!
0'
0/
#855090000000
1!
1'
1/
#855100000000
0!
0'
0/
#855110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#855120000000
0!
0'
0/
#855130000000
1!
1'
1/
#855140000000
0!
0'
0/
#855150000000
1!
1'
1/
#855160000000
0!
0'
0/
#855170000000
1!
1'
1/
#855180000000
0!
0'
0/
#855190000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#855200000000
0!
0'
0/
#855210000000
1!
1'
1/
#855220000000
0!
0'
0/
#855230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#855240000000
0!
0'
0/
#855250000000
1!
1'
1/
#855260000000
0!
0'
0/
#855270000000
#855280000000
1!
1'
1/
#855290000000
0!
0'
0/
#855300000000
1!
1'
1/
#855310000000
0!
1"
0'
1(
0/
10
#855320000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#855330000000
0!
0'
0/
#855340000000
1!
1'
1/
#855350000000
0!
0'
0/
#855360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#855370000000
0!
0'
0/
#855380000000
1!
1'
1/
#855390000000
0!
1"
0'
1(
0/
10
#855400000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#855410000000
0!
1$
0'
1+
0/
#855420000000
1!
1'
1/
#855430000000
0!
0'
0/
#855440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#855450000000
0!
0'
0/
#855460000000
1!
1'
1/
#855470000000
0!
0'
0/
#855480000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#855490000000
0!
0'
0/
#855500000000
1!
1'
1/
#855510000000
0!
0'
0/
#855520000000
1!
1'
1/
#855530000000
0!
0'
0/
#855540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#855550000000
0!
0'
0/
#855560000000
1!
1'
1/
#855570000000
0!
0'
0/
#855580000000
1!
1'
1/
#855590000000
0!
0'
0/
#855600000000
1!
1'
1/
#855610000000
0!
0'
0/
#855620000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#855630000000
0!
0'
0/
#855640000000
1!
1'
1/
#855650000000
0!
0'
0/
#855660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#855670000000
0!
0'
0/
#855680000000
1!
1'
1/
#855690000000
0!
0'
0/
#855700000000
#855710000000
1!
1'
1/
#855720000000
0!
0'
0/
#855730000000
1!
1'
1/
#855740000000
0!
1"
0'
1(
0/
10
#855750000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#855760000000
0!
0'
0/
#855770000000
1!
1'
1/
#855780000000
0!
0'
0/
#855790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#855800000000
0!
0'
0/
#855810000000
1!
1'
1/
#855820000000
0!
1"
0'
1(
0/
10
#855830000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#855840000000
0!
1$
0'
1+
0/
#855850000000
1!
1'
1/
#855860000000
0!
0'
0/
#855870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#855880000000
0!
0'
0/
#855890000000
1!
1'
1/
#855900000000
0!
0'
0/
#855910000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#855920000000
0!
0'
0/
#855930000000
1!
1'
1/
#855940000000
0!
0'
0/
#855950000000
1!
1'
1/
#855960000000
0!
0'
0/
#855970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#855980000000
0!
0'
0/
#855990000000
1!
1'
1/
#856000000000
0!
0'
0/
#856010000000
1!
1'
1/
#856020000000
0!
0'
0/
#856030000000
1!
1'
1/
#856040000000
0!
0'
0/
#856050000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#856060000000
0!
0'
0/
#856070000000
1!
1'
1/
#856080000000
0!
0'
0/
#856090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#856100000000
0!
0'
0/
#856110000000
1!
1'
1/
#856120000000
0!
0'
0/
#856130000000
#856140000000
1!
1'
1/
#856150000000
0!
0'
0/
#856160000000
1!
1'
1/
#856170000000
0!
1"
0'
1(
0/
10
#856180000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#856190000000
0!
0'
0/
#856200000000
1!
1'
1/
#856210000000
0!
0'
0/
#856220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#856230000000
0!
0'
0/
#856240000000
1!
1'
1/
#856250000000
0!
1"
0'
1(
0/
10
#856260000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#856270000000
0!
1$
0'
1+
0/
#856280000000
1!
1'
1/
#856290000000
0!
0'
0/
#856300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#856310000000
0!
0'
0/
#856320000000
1!
1'
1/
#856330000000
0!
0'
0/
#856340000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#856350000000
0!
0'
0/
#856360000000
1!
1'
1/
#856370000000
0!
0'
0/
#856380000000
1!
1'
1/
#856390000000
0!
0'
0/
#856400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#856410000000
0!
0'
0/
#856420000000
1!
1'
1/
#856430000000
0!
0'
0/
#856440000000
1!
1'
1/
#856450000000
0!
0'
0/
#856460000000
1!
1'
1/
#856470000000
0!
0'
0/
#856480000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#856490000000
0!
0'
0/
#856500000000
1!
1'
1/
#856510000000
0!
0'
0/
#856520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#856530000000
0!
0'
0/
#856540000000
1!
1'
1/
#856550000000
0!
0'
0/
#856560000000
#856570000000
1!
1'
1/
#856580000000
0!
0'
0/
#856590000000
1!
1'
1/
#856600000000
0!
1"
0'
1(
0/
10
#856610000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#856620000000
0!
0'
0/
#856630000000
1!
1'
1/
#856640000000
0!
0'
0/
#856650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#856660000000
0!
0'
0/
#856670000000
1!
1'
1/
#856680000000
0!
1"
0'
1(
0/
10
#856690000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#856700000000
0!
1$
0'
1+
0/
#856710000000
1!
1'
1/
#856720000000
0!
0'
0/
#856730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#856740000000
0!
0'
0/
#856750000000
1!
1'
1/
#856760000000
0!
0'
0/
#856770000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#856780000000
0!
0'
0/
#856790000000
1!
1'
1/
#856800000000
0!
0'
0/
#856810000000
1!
1'
1/
#856820000000
0!
0'
0/
#856830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#856840000000
0!
0'
0/
#856850000000
1!
1'
1/
#856860000000
0!
0'
0/
#856870000000
1!
1'
1/
#856880000000
0!
0'
0/
#856890000000
1!
1'
1/
#856900000000
0!
0'
0/
#856910000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#856920000000
0!
0'
0/
#856930000000
1!
1'
1/
#856940000000
0!
0'
0/
#856950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#856960000000
0!
0'
0/
#856970000000
1!
1'
1/
#856980000000
0!
0'
0/
#856990000000
#857000000000
1!
1'
1/
#857010000000
0!
0'
0/
#857020000000
1!
1'
1/
#857030000000
0!
1"
0'
1(
0/
10
#857040000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#857050000000
0!
0'
0/
#857060000000
1!
1'
1/
#857070000000
0!
0'
0/
#857080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#857090000000
0!
0'
0/
#857100000000
1!
1'
1/
#857110000000
0!
1"
0'
1(
0/
10
#857120000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#857130000000
0!
1$
0'
1+
0/
#857140000000
1!
1'
1/
#857150000000
0!
0'
0/
#857160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#857170000000
0!
0'
0/
#857180000000
1!
1'
1/
#857190000000
0!
0'
0/
#857200000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#857210000000
0!
0'
0/
#857220000000
1!
1'
1/
#857230000000
0!
0'
0/
#857240000000
1!
1'
1/
#857250000000
0!
0'
0/
#857260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#857270000000
0!
0'
0/
#857280000000
1!
1'
1/
#857290000000
0!
0'
0/
#857300000000
1!
1'
1/
#857310000000
0!
0'
0/
#857320000000
1!
1'
1/
#857330000000
0!
0'
0/
#857340000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#857350000000
0!
0'
0/
#857360000000
1!
1'
1/
#857370000000
0!
0'
0/
#857380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#857390000000
0!
0'
0/
#857400000000
1!
1'
1/
#857410000000
0!
0'
0/
#857420000000
#857430000000
1!
1'
1/
#857440000000
0!
0'
0/
#857450000000
1!
1'
1/
#857460000000
0!
1"
0'
1(
0/
10
#857470000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#857480000000
0!
0'
0/
#857490000000
1!
1'
1/
#857500000000
0!
0'
0/
#857510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#857520000000
0!
0'
0/
#857530000000
1!
1'
1/
#857540000000
0!
1"
0'
1(
0/
10
#857550000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#857560000000
0!
1$
0'
1+
0/
#857570000000
1!
1'
1/
#857580000000
0!
0'
0/
#857590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#857600000000
0!
0'
0/
#857610000000
1!
1'
1/
#857620000000
0!
0'
0/
#857630000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#857640000000
0!
0'
0/
#857650000000
1!
1'
1/
#857660000000
0!
0'
0/
#857670000000
1!
1'
1/
#857680000000
0!
0'
0/
#857690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#857700000000
0!
0'
0/
#857710000000
1!
1'
1/
#857720000000
0!
0'
0/
#857730000000
1!
1'
1/
#857740000000
0!
0'
0/
#857750000000
1!
1'
1/
#857760000000
0!
0'
0/
#857770000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#857780000000
0!
0'
0/
#857790000000
1!
1'
1/
#857800000000
0!
0'
0/
#857810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#857820000000
0!
0'
0/
#857830000000
1!
1'
1/
#857840000000
0!
0'
0/
#857850000000
#857860000000
1!
1'
1/
#857870000000
0!
0'
0/
#857880000000
1!
1'
1/
#857890000000
0!
1"
0'
1(
0/
10
#857900000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#857910000000
0!
0'
0/
#857920000000
1!
1'
1/
#857930000000
0!
0'
0/
#857940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#857950000000
0!
0'
0/
#857960000000
1!
1'
1/
#857970000000
0!
1"
0'
1(
0/
10
#857980000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#857990000000
0!
1$
0'
1+
0/
#858000000000
1!
1'
1/
#858010000000
0!
0'
0/
#858020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#858030000000
0!
0'
0/
#858040000000
1!
1'
1/
#858050000000
0!
0'
0/
#858060000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#858070000000
0!
0'
0/
#858080000000
1!
1'
1/
#858090000000
0!
0'
0/
#858100000000
1!
1'
1/
#858110000000
0!
0'
0/
#858120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#858130000000
0!
0'
0/
#858140000000
1!
1'
1/
#858150000000
0!
0'
0/
#858160000000
1!
1'
1/
#858170000000
0!
0'
0/
#858180000000
1!
1'
1/
#858190000000
0!
0'
0/
#858200000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#858210000000
0!
0'
0/
#858220000000
1!
1'
1/
#858230000000
0!
0'
0/
#858240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#858250000000
0!
0'
0/
#858260000000
1!
1'
1/
#858270000000
0!
0'
0/
#858280000000
#858290000000
1!
1'
1/
#858300000000
0!
0'
0/
#858310000000
1!
1'
1/
#858320000000
0!
1"
0'
1(
0/
10
#858330000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#858340000000
0!
0'
0/
#858350000000
1!
1'
1/
#858360000000
0!
0'
0/
#858370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#858380000000
0!
0'
0/
#858390000000
1!
1'
1/
#858400000000
0!
1"
0'
1(
0/
10
#858410000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#858420000000
0!
1$
0'
1+
0/
#858430000000
1!
1'
1/
#858440000000
0!
0'
0/
#858450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#858460000000
0!
0'
0/
#858470000000
1!
1'
1/
#858480000000
0!
0'
0/
#858490000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#858500000000
0!
0'
0/
#858510000000
1!
1'
1/
#858520000000
0!
0'
0/
#858530000000
1!
1'
1/
#858540000000
0!
0'
0/
#858550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#858560000000
0!
0'
0/
#858570000000
1!
1'
1/
#858580000000
0!
0'
0/
#858590000000
1!
1'
1/
#858600000000
0!
0'
0/
#858610000000
1!
1'
1/
#858620000000
0!
0'
0/
#858630000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#858640000000
0!
0'
0/
#858650000000
1!
1'
1/
#858660000000
0!
0'
0/
#858670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#858680000000
0!
0'
0/
#858690000000
1!
1'
1/
#858700000000
0!
0'
0/
#858710000000
#858720000000
1!
1'
1/
#858730000000
0!
0'
0/
#858740000000
1!
1'
1/
#858750000000
0!
1"
0'
1(
0/
10
#858760000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#858770000000
0!
0'
0/
#858780000000
1!
1'
1/
#858790000000
0!
0'
0/
#858800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#858810000000
0!
0'
0/
#858820000000
1!
1'
1/
#858830000000
0!
1"
0'
1(
0/
10
#858840000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#858850000000
0!
1$
0'
1+
0/
#858860000000
1!
1'
1/
#858870000000
0!
0'
0/
#858880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#858890000000
0!
0'
0/
#858900000000
1!
1'
1/
#858910000000
0!
0'
0/
#858920000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#858930000000
0!
0'
0/
#858940000000
1!
1'
1/
#858950000000
0!
0'
0/
#858960000000
1!
1'
1/
#858970000000
0!
0'
0/
#858980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#858990000000
0!
0'
0/
#859000000000
1!
1'
1/
#859010000000
0!
0'
0/
#859020000000
1!
1'
1/
#859030000000
0!
0'
0/
#859040000000
1!
1'
1/
#859050000000
0!
0'
0/
#859060000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#859070000000
0!
0'
0/
#859080000000
1!
1'
1/
#859090000000
0!
0'
0/
#859100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#859110000000
0!
0'
0/
#859120000000
1!
1'
1/
#859130000000
0!
0'
0/
#859140000000
#859150000000
1!
1'
1/
#859160000000
0!
0'
0/
#859170000000
1!
1'
1/
#859180000000
0!
1"
0'
1(
0/
10
#859190000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#859200000000
0!
0'
0/
#859210000000
1!
1'
1/
#859220000000
0!
0'
0/
#859230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#859240000000
0!
0'
0/
#859250000000
1!
1'
1/
#859260000000
0!
1"
0'
1(
0/
10
#859270000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#859280000000
0!
1$
0'
1+
0/
#859290000000
1!
1'
1/
#859300000000
0!
0'
0/
#859310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#859320000000
0!
0'
0/
#859330000000
1!
1'
1/
#859340000000
0!
0'
0/
#859350000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#859360000000
0!
0'
0/
#859370000000
1!
1'
1/
#859380000000
0!
0'
0/
#859390000000
1!
1'
1/
#859400000000
0!
0'
0/
#859410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#859420000000
0!
0'
0/
#859430000000
1!
1'
1/
#859440000000
0!
0'
0/
#859450000000
1!
1'
1/
#859460000000
0!
0'
0/
#859470000000
1!
1'
1/
#859480000000
0!
0'
0/
#859490000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#859500000000
0!
0'
0/
#859510000000
1!
1'
1/
#859520000000
0!
0'
0/
#859530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#859540000000
0!
0'
0/
#859550000000
1!
1'
1/
#859560000000
0!
0'
0/
#859570000000
#859580000000
1!
1'
1/
#859590000000
0!
0'
0/
#859600000000
1!
1'
1/
#859610000000
0!
1"
0'
1(
0/
10
#859620000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#859630000000
0!
0'
0/
#859640000000
1!
1'
1/
#859650000000
0!
0'
0/
#859660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#859670000000
0!
0'
0/
#859680000000
1!
1'
1/
#859690000000
0!
1"
0'
1(
0/
10
#859700000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#859710000000
0!
1$
0'
1+
0/
#859720000000
1!
1'
1/
#859730000000
0!
0'
0/
#859740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#859750000000
0!
0'
0/
#859760000000
1!
1'
1/
#859770000000
0!
0'
0/
#859780000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#859790000000
0!
0'
0/
#859800000000
1!
1'
1/
#859810000000
0!
0'
0/
#859820000000
1!
1'
1/
#859830000000
0!
0'
0/
#859840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#859850000000
0!
0'
0/
#859860000000
1!
1'
1/
#859870000000
0!
0'
0/
#859880000000
1!
1'
1/
#859890000000
0!
0'
0/
#859900000000
1!
1'
1/
#859910000000
0!
0'
0/
#859920000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#859930000000
0!
0'
0/
#859940000000
1!
1'
1/
#859950000000
0!
0'
0/
#859960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#859970000000
0!
0'
0/
#859980000000
1!
1'
1/
#859990000000
0!
0'
0/
#860000000000
#860010000000
1!
1'
1/
#860020000000
0!
0'
0/
#860030000000
1!
1'
1/
#860040000000
0!
1"
0'
1(
0/
10
#860050000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#860060000000
0!
0'
0/
#860070000000
1!
1'
1/
#860080000000
0!
0'
0/
#860090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#860100000000
0!
0'
0/
#860110000000
1!
1'
1/
#860120000000
0!
1"
0'
1(
0/
10
#860130000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#860140000000
0!
1$
0'
1+
0/
#860150000000
1!
1'
1/
#860160000000
0!
0'
0/
#860170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#860180000000
0!
0'
0/
#860190000000
1!
1'
1/
#860200000000
0!
0'
0/
#860210000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#860220000000
0!
0'
0/
#860230000000
1!
1'
1/
#860240000000
0!
0'
0/
#860250000000
1!
1'
1/
#860260000000
0!
0'
0/
#860270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#860280000000
0!
0'
0/
#860290000000
1!
1'
1/
#860300000000
0!
0'
0/
#860310000000
1!
1'
1/
#860320000000
0!
0'
0/
#860330000000
1!
1'
1/
#860340000000
0!
0'
0/
#860350000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#860360000000
0!
0'
0/
#860370000000
1!
1'
1/
#860380000000
0!
0'
0/
#860390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#860400000000
0!
0'
0/
#860410000000
1!
1'
1/
#860420000000
0!
0'
0/
#860430000000
#860440000000
1!
1'
1/
#860450000000
0!
0'
0/
#860460000000
1!
1'
1/
#860470000000
0!
1"
0'
1(
0/
10
#860480000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#860490000000
0!
0'
0/
#860500000000
1!
1'
1/
#860510000000
0!
0'
0/
#860520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#860530000000
0!
0'
0/
#860540000000
1!
1'
1/
#860550000000
0!
1"
0'
1(
0/
10
#860560000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#860570000000
0!
1$
0'
1+
0/
#860580000000
1!
1'
1/
#860590000000
0!
0'
0/
#860600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#860610000000
0!
0'
0/
#860620000000
1!
1'
1/
#860630000000
0!
0'
0/
#860640000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#860650000000
0!
0'
0/
#860660000000
1!
1'
1/
#860670000000
0!
0'
0/
#860680000000
1!
1'
1/
#860690000000
0!
0'
0/
#860700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#860710000000
0!
0'
0/
#860720000000
1!
1'
1/
#860730000000
0!
0'
0/
#860740000000
1!
1'
1/
#860750000000
0!
0'
0/
#860760000000
1!
1'
1/
#860770000000
0!
0'
0/
#860780000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#860790000000
0!
0'
0/
#860800000000
1!
1'
1/
#860810000000
0!
0'
0/
#860820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#860830000000
0!
0'
0/
#860840000000
1!
1'
1/
#860850000000
0!
0'
0/
#860860000000
#860870000000
1!
1'
1/
#860880000000
0!
0'
0/
#860890000000
1!
1'
1/
#860900000000
0!
1"
0'
1(
0/
10
#860910000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#860920000000
0!
0'
0/
#860930000000
1!
1'
1/
#860940000000
0!
0'
0/
#860950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#860960000000
0!
0'
0/
#860970000000
1!
1'
1/
#860980000000
0!
1"
0'
1(
0/
10
#860990000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#861000000000
0!
1$
0'
1+
0/
#861010000000
1!
1'
1/
#861020000000
0!
0'
0/
#861030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#861040000000
0!
0'
0/
#861050000000
1!
1'
1/
#861060000000
0!
0'
0/
#861070000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#861080000000
0!
0'
0/
#861090000000
1!
1'
1/
#861100000000
0!
0'
0/
#861110000000
1!
1'
1/
#861120000000
0!
0'
0/
#861130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#861140000000
0!
0'
0/
#861150000000
1!
1'
1/
#861160000000
0!
0'
0/
#861170000000
1!
1'
1/
#861180000000
0!
0'
0/
#861190000000
1!
1'
1/
#861200000000
0!
0'
0/
#861210000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#861220000000
0!
0'
0/
#861230000000
1!
1'
1/
#861240000000
0!
0'
0/
#861250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#861260000000
0!
0'
0/
#861270000000
1!
1'
1/
#861280000000
0!
0'
0/
#861290000000
#861300000000
1!
1'
1/
#861310000000
0!
0'
0/
#861320000000
1!
1'
1/
#861330000000
0!
1"
0'
1(
0/
10
#861340000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#861350000000
0!
0'
0/
#861360000000
1!
1'
1/
#861370000000
0!
0'
0/
#861380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#861390000000
0!
0'
0/
#861400000000
1!
1'
1/
#861410000000
0!
1"
0'
1(
0/
10
#861420000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#861430000000
0!
1$
0'
1+
0/
#861440000000
1!
1'
1/
#861450000000
0!
0'
0/
#861460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#861470000000
0!
0'
0/
#861480000000
1!
1'
1/
#861490000000
0!
0'
0/
#861500000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#861510000000
0!
0'
0/
#861520000000
1!
1'
1/
#861530000000
0!
0'
0/
#861540000000
1!
1'
1/
#861550000000
0!
0'
0/
#861560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#861570000000
0!
0'
0/
#861580000000
1!
1'
1/
#861590000000
0!
0'
0/
#861600000000
1!
1'
1/
#861610000000
0!
0'
0/
#861620000000
1!
1'
1/
#861630000000
0!
0'
0/
#861640000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#861650000000
0!
0'
0/
#861660000000
1!
1'
1/
#861670000000
0!
0'
0/
#861680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#861690000000
0!
0'
0/
#861700000000
1!
1'
1/
#861710000000
0!
0'
0/
#861720000000
#861730000000
1!
1'
1/
#861740000000
0!
0'
0/
#861750000000
1!
1'
1/
#861760000000
0!
1"
0'
1(
0/
10
#861770000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#861780000000
0!
0'
0/
#861790000000
1!
1'
1/
#861800000000
0!
0'
0/
#861810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#861820000000
0!
0'
0/
#861830000000
1!
1'
1/
#861840000000
0!
1"
0'
1(
0/
10
#861850000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#861860000000
0!
1$
0'
1+
0/
#861870000000
1!
1'
1/
#861880000000
0!
0'
0/
#861890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#861900000000
0!
0'
0/
#861910000000
1!
1'
1/
#861920000000
0!
0'
0/
#861930000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#861940000000
0!
0'
0/
#861950000000
1!
1'
1/
#861960000000
0!
0'
0/
#861970000000
1!
1'
1/
#861980000000
0!
0'
0/
#861990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#862000000000
0!
0'
0/
#862010000000
1!
1'
1/
#862020000000
0!
0'
0/
#862030000000
1!
1'
1/
#862040000000
0!
0'
0/
#862050000000
1!
1'
1/
#862060000000
0!
0'
0/
#862070000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#862080000000
0!
0'
0/
#862090000000
1!
1'
1/
#862100000000
0!
0'
0/
#862110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#862120000000
0!
0'
0/
#862130000000
1!
1'
1/
#862140000000
0!
0'
0/
#862150000000
#862160000000
1!
1'
1/
#862170000000
0!
0'
0/
#862180000000
1!
1'
1/
#862190000000
0!
1"
0'
1(
0/
10
#862200000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#862210000000
0!
0'
0/
#862220000000
1!
1'
1/
#862230000000
0!
0'
0/
#862240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#862250000000
0!
0'
0/
#862260000000
1!
1'
1/
#862270000000
0!
1"
0'
1(
0/
10
#862280000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#862290000000
0!
1$
0'
1+
0/
#862300000000
1!
1'
1/
#862310000000
0!
0'
0/
#862320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#862330000000
0!
0'
0/
#862340000000
1!
1'
1/
#862350000000
0!
0'
0/
#862360000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#862370000000
0!
0'
0/
#862380000000
1!
1'
1/
#862390000000
0!
0'
0/
#862400000000
1!
1'
1/
#862410000000
0!
0'
0/
#862420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#862430000000
0!
0'
0/
#862440000000
1!
1'
1/
#862450000000
0!
0'
0/
#862460000000
1!
1'
1/
#862470000000
0!
0'
0/
#862480000000
1!
1'
1/
#862490000000
0!
0'
0/
#862500000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#862510000000
0!
0'
0/
#862520000000
1!
1'
1/
#862530000000
0!
0'
0/
#862540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#862550000000
0!
0'
0/
#862560000000
1!
1'
1/
#862570000000
0!
0'
0/
#862580000000
#862590000000
1!
1'
1/
#862600000000
0!
0'
0/
#862610000000
1!
1'
1/
#862620000000
0!
1"
0'
1(
0/
10
#862630000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#862640000000
0!
0'
0/
#862650000000
1!
1'
1/
#862660000000
0!
0'
0/
#862670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#862680000000
0!
0'
0/
#862690000000
1!
1'
1/
#862700000000
0!
1"
0'
1(
0/
10
#862710000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#862720000000
0!
1$
0'
1+
0/
#862730000000
1!
1'
1/
#862740000000
0!
0'
0/
#862750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#862760000000
0!
0'
0/
#862770000000
1!
1'
1/
#862780000000
0!
0'
0/
#862790000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#862800000000
0!
0'
0/
#862810000000
1!
1'
1/
#862820000000
0!
0'
0/
#862830000000
1!
1'
1/
#862840000000
0!
0'
0/
#862850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#862860000000
0!
0'
0/
#862870000000
1!
1'
1/
#862880000000
0!
0'
0/
#862890000000
1!
1'
1/
#862900000000
0!
0'
0/
#862910000000
1!
1'
1/
#862920000000
0!
0'
0/
#862930000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#862940000000
0!
0'
0/
#862950000000
1!
1'
1/
#862960000000
0!
0'
0/
#862970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#862980000000
0!
0'
0/
#862990000000
1!
1'
1/
#863000000000
0!
0'
0/
#863010000000
#863020000000
1!
1'
1/
#863030000000
0!
0'
0/
#863040000000
1!
1'
1/
#863050000000
0!
1"
0'
1(
0/
10
#863060000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#863070000000
0!
0'
0/
#863080000000
1!
1'
1/
#863090000000
0!
0'
0/
#863100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#863110000000
0!
0'
0/
#863120000000
1!
1'
1/
#863130000000
0!
1"
0'
1(
0/
10
#863140000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#863150000000
0!
1$
0'
1+
0/
#863160000000
1!
1'
1/
#863170000000
0!
0'
0/
#863180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#863190000000
0!
0'
0/
#863200000000
1!
1'
1/
#863210000000
0!
0'
0/
#863220000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#863230000000
0!
0'
0/
#863240000000
1!
1'
1/
#863250000000
0!
0'
0/
#863260000000
1!
1'
1/
#863270000000
0!
0'
0/
#863280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#863290000000
0!
0'
0/
#863300000000
1!
1'
1/
#863310000000
0!
0'
0/
#863320000000
1!
1'
1/
#863330000000
0!
0'
0/
#863340000000
1!
1'
1/
#863350000000
0!
0'
0/
#863360000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#863370000000
0!
0'
0/
#863380000000
1!
1'
1/
#863390000000
0!
0'
0/
#863400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#863410000000
0!
0'
0/
#863420000000
1!
1'
1/
#863430000000
0!
0'
0/
#863440000000
#863450000000
1!
1'
1/
#863460000000
0!
0'
0/
#863470000000
1!
1'
1/
#863480000000
0!
1"
0'
1(
0/
10
#863490000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#863500000000
0!
0'
0/
#863510000000
1!
1'
1/
#863520000000
0!
0'
0/
#863530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#863540000000
0!
0'
0/
#863550000000
1!
1'
1/
#863560000000
0!
1"
0'
1(
0/
10
#863570000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#863580000000
0!
1$
0'
1+
0/
#863590000000
1!
1'
1/
#863600000000
0!
0'
0/
#863610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#863620000000
0!
0'
0/
#863630000000
1!
1'
1/
#863640000000
0!
0'
0/
#863650000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#863660000000
0!
0'
0/
#863670000000
1!
1'
1/
#863680000000
0!
0'
0/
#863690000000
1!
1'
1/
#863700000000
0!
0'
0/
#863710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#863720000000
0!
0'
0/
#863730000000
1!
1'
1/
#863740000000
0!
0'
0/
#863750000000
1!
1'
1/
#863760000000
0!
0'
0/
#863770000000
1!
1'
1/
#863780000000
0!
0'
0/
#863790000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#863800000000
0!
0'
0/
#863810000000
1!
1'
1/
#863820000000
0!
0'
0/
#863830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#863840000000
0!
0'
0/
#863850000000
1!
1'
1/
#863860000000
0!
0'
0/
#863870000000
#863880000000
1!
1'
1/
#863890000000
0!
0'
0/
#863900000000
1!
1'
1/
#863910000000
0!
1"
0'
1(
0/
10
#863920000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#863930000000
0!
0'
0/
#863940000000
1!
1'
1/
#863950000000
0!
0'
0/
#863960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#863970000000
0!
0'
0/
#863980000000
1!
1'
1/
#863990000000
0!
1"
0'
1(
0/
10
#864000000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#864010000000
0!
1$
0'
1+
0/
#864020000000
1!
1'
1/
#864030000000
0!
0'
0/
#864040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#864050000000
0!
0'
0/
#864060000000
1!
1'
1/
#864070000000
0!
0'
0/
#864080000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#864090000000
0!
0'
0/
#864100000000
1!
1'
1/
#864110000000
0!
0'
0/
#864120000000
1!
1'
1/
#864130000000
0!
0'
0/
#864140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#864150000000
0!
0'
0/
#864160000000
1!
1'
1/
#864170000000
0!
0'
0/
#864180000000
1!
1'
1/
#864190000000
0!
0'
0/
#864200000000
1!
1'
1/
#864210000000
0!
0'
0/
#864220000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#864230000000
0!
0'
0/
#864240000000
1!
1'
1/
#864250000000
0!
0'
0/
#864260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#864270000000
0!
0'
0/
#864280000000
1!
1'
1/
#864290000000
0!
0'
0/
#864300000000
#864310000000
1!
1'
1/
#864320000000
0!
0'
0/
#864330000000
1!
1'
1/
#864340000000
0!
1"
0'
1(
0/
10
#864350000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#864360000000
0!
0'
0/
#864370000000
1!
1'
1/
#864380000000
0!
0'
0/
#864390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#864400000000
0!
0'
0/
#864410000000
1!
1'
1/
#864420000000
0!
1"
0'
1(
0/
10
#864430000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#864440000000
0!
1$
0'
1+
0/
#864450000000
1!
1'
1/
#864460000000
0!
0'
0/
#864470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#864480000000
0!
0'
0/
#864490000000
1!
1'
1/
#864500000000
0!
0'
0/
#864510000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#864520000000
0!
0'
0/
#864530000000
1!
1'
1/
#864540000000
0!
0'
0/
#864550000000
1!
1'
1/
#864560000000
0!
0'
0/
#864570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#864580000000
0!
0'
0/
#864590000000
1!
1'
1/
#864600000000
0!
0'
0/
#864610000000
1!
1'
1/
#864620000000
0!
0'
0/
#864630000000
1!
1'
1/
#864640000000
0!
0'
0/
#864650000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#864660000000
0!
0'
0/
#864670000000
1!
1'
1/
#864680000000
0!
0'
0/
#864690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#864700000000
0!
0'
0/
#864710000000
1!
1'
1/
#864720000000
0!
0'
0/
#864730000000
#864740000000
1!
1'
1/
#864750000000
0!
0'
0/
#864760000000
1!
1'
1/
#864770000000
0!
1"
0'
1(
0/
10
#864780000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#864790000000
0!
0'
0/
#864800000000
1!
1'
1/
#864810000000
0!
0'
0/
#864820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#864830000000
0!
0'
0/
#864840000000
1!
1'
1/
#864850000000
0!
1"
0'
1(
0/
10
#864860000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#864870000000
0!
1$
0'
1+
0/
#864880000000
1!
1'
1/
#864890000000
0!
0'
0/
#864900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#864910000000
0!
0'
0/
#864920000000
1!
1'
1/
#864930000000
0!
0'
0/
#864940000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#864950000000
0!
0'
0/
#864960000000
1!
1'
1/
#864970000000
0!
0'
0/
#864980000000
1!
1'
1/
#864990000000
0!
0'
0/
#865000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#865010000000
0!
0'
0/
#865020000000
1!
1'
1/
#865030000000
0!
0'
0/
#865040000000
1!
1'
1/
#865050000000
0!
0'
0/
#865060000000
1!
1'
1/
#865070000000
0!
0'
0/
#865080000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#865090000000
0!
0'
0/
#865100000000
1!
1'
1/
#865110000000
0!
0'
0/
#865120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#865130000000
0!
0'
0/
#865140000000
1!
1'
1/
#865150000000
0!
0'
0/
#865160000000
#865170000000
1!
1'
1/
#865180000000
0!
0'
0/
#865190000000
1!
1'
1/
#865200000000
0!
1"
0'
1(
0/
10
#865210000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#865220000000
0!
0'
0/
#865230000000
1!
1'
1/
#865240000000
0!
0'
0/
#865250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#865260000000
0!
0'
0/
#865270000000
1!
1'
1/
#865280000000
0!
1"
0'
1(
0/
10
#865290000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#865300000000
0!
1$
0'
1+
0/
#865310000000
1!
1'
1/
#865320000000
0!
0'
0/
#865330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#865340000000
0!
0'
0/
#865350000000
1!
1'
1/
#865360000000
0!
0'
0/
#865370000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#865380000000
0!
0'
0/
#865390000000
1!
1'
1/
#865400000000
0!
0'
0/
#865410000000
1!
1'
1/
#865420000000
0!
0'
0/
#865430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#865440000000
0!
0'
0/
#865450000000
1!
1'
1/
#865460000000
0!
0'
0/
#865470000000
1!
1'
1/
#865480000000
0!
0'
0/
#865490000000
1!
1'
1/
#865500000000
0!
0'
0/
#865510000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#865520000000
0!
0'
0/
#865530000000
1!
1'
1/
#865540000000
0!
0'
0/
#865550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#865560000000
0!
0'
0/
#865570000000
1!
1'
1/
#865580000000
0!
0'
0/
#865590000000
#865600000000
1!
1'
1/
#865610000000
0!
0'
0/
#865620000000
1!
1'
1/
#865630000000
0!
1"
0'
1(
0/
10
#865640000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#865650000000
0!
0'
0/
#865660000000
1!
1'
1/
#865670000000
0!
0'
0/
#865680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#865690000000
0!
0'
0/
#865700000000
1!
1'
1/
#865710000000
0!
1"
0'
1(
0/
10
#865720000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#865730000000
0!
1$
0'
1+
0/
#865740000000
1!
1'
1/
#865750000000
0!
0'
0/
#865760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#865770000000
0!
0'
0/
#865780000000
1!
1'
1/
#865790000000
0!
0'
0/
#865800000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#865810000000
0!
0'
0/
#865820000000
1!
1'
1/
#865830000000
0!
0'
0/
#865840000000
1!
1'
1/
#865850000000
0!
0'
0/
#865860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#865870000000
0!
0'
0/
#865880000000
1!
1'
1/
#865890000000
0!
0'
0/
#865900000000
1!
1'
1/
#865910000000
0!
0'
0/
#865920000000
1!
1'
1/
#865930000000
0!
0'
0/
#865940000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#865950000000
0!
0'
0/
#865960000000
1!
1'
1/
#865970000000
0!
0'
0/
#865980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#865990000000
0!
0'
0/
#866000000000
1!
1'
1/
#866010000000
0!
0'
0/
#866020000000
#866030000000
1!
1'
1/
#866040000000
0!
0'
0/
#866050000000
1!
1'
1/
#866060000000
0!
1"
0'
1(
0/
10
#866070000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#866080000000
0!
0'
0/
#866090000000
1!
1'
1/
#866100000000
0!
0'
0/
#866110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#866120000000
0!
0'
0/
#866130000000
1!
1'
1/
#866140000000
0!
1"
0'
1(
0/
10
#866150000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#866160000000
0!
1$
0'
1+
0/
#866170000000
1!
1'
1/
#866180000000
0!
0'
0/
#866190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#866200000000
0!
0'
0/
#866210000000
1!
1'
1/
#866220000000
0!
0'
0/
#866230000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#866240000000
0!
0'
0/
#866250000000
1!
1'
1/
#866260000000
0!
0'
0/
#866270000000
1!
1'
1/
#866280000000
0!
0'
0/
#866290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#866300000000
0!
0'
0/
#866310000000
1!
1'
1/
#866320000000
0!
0'
0/
#866330000000
1!
1'
1/
#866340000000
0!
0'
0/
#866350000000
1!
1'
1/
#866360000000
0!
0'
0/
#866370000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#866380000000
0!
0'
0/
#866390000000
1!
1'
1/
#866400000000
0!
0'
0/
#866410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#866420000000
0!
0'
0/
#866430000000
1!
1'
1/
#866440000000
0!
0'
0/
#866450000000
#866460000000
1!
1'
1/
#866470000000
0!
0'
0/
#866480000000
1!
1'
1/
#866490000000
0!
1"
0'
1(
0/
10
#866500000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#866510000000
0!
0'
0/
#866520000000
1!
1'
1/
#866530000000
0!
0'
0/
#866540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#866550000000
0!
0'
0/
#866560000000
1!
1'
1/
#866570000000
0!
1"
0'
1(
0/
10
#866580000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#866590000000
0!
1$
0'
1+
0/
#866600000000
1!
1'
1/
#866610000000
0!
0'
0/
#866620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#866630000000
0!
0'
0/
#866640000000
1!
1'
1/
#866650000000
0!
0'
0/
#866660000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#866670000000
0!
0'
0/
#866680000000
1!
1'
1/
#866690000000
0!
0'
0/
#866700000000
1!
1'
1/
#866710000000
0!
0'
0/
#866720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#866730000000
0!
0'
0/
#866740000000
1!
1'
1/
#866750000000
0!
0'
0/
#866760000000
1!
1'
1/
#866770000000
0!
0'
0/
#866780000000
1!
1'
1/
#866790000000
0!
0'
0/
#866800000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#866810000000
0!
0'
0/
#866820000000
1!
1'
1/
#866830000000
0!
0'
0/
#866840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#866850000000
0!
0'
0/
#866860000000
1!
1'
1/
#866870000000
0!
0'
0/
#866880000000
#866890000000
1!
1'
1/
#866900000000
0!
0'
0/
#866910000000
1!
1'
1/
#866920000000
0!
1"
0'
1(
0/
10
#866930000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#866940000000
0!
0'
0/
#866950000000
1!
1'
1/
#866960000000
0!
0'
0/
#866970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#866980000000
0!
0'
0/
#866990000000
1!
1'
1/
#867000000000
0!
1"
0'
1(
0/
10
#867010000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#867020000000
0!
1$
0'
1+
0/
#867030000000
1!
1'
1/
#867040000000
0!
0'
0/
#867050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#867060000000
0!
0'
0/
#867070000000
1!
1'
1/
#867080000000
0!
0'
0/
#867090000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#867100000000
0!
0'
0/
#867110000000
1!
1'
1/
#867120000000
0!
0'
0/
#867130000000
1!
1'
1/
#867140000000
0!
0'
0/
#867150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#867160000000
0!
0'
0/
#867170000000
1!
1'
1/
#867180000000
0!
0'
0/
#867190000000
1!
1'
1/
#867200000000
0!
0'
0/
#867210000000
1!
1'
1/
#867220000000
0!
0'
0/
#867230000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#867240000000
0!
0'
0/
#867250000000
1!
1'
1/
#867260000000
0!
0'
0/
#867270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#867280000000
0!
0'
0/
#867290000000
1!
1'
1/
#867300000000
0!
0'
0/
#867310000000
#867320000000
1!
1'
1/
#867330000000
0!
0'
0/
#867340000000
1!
1'
1/
#867350000000
0!
1"
0'
1(
0/
10
#867360000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#867370000000
0!
0'
0/
#867380000000
1!
1'
1/
#867390000000
0!
0'
0/
#867400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#867410000000
0!
0'
0/
#867420000000
1!
1'
1/
#867430000000
0!
1"
0'
1(
0/
10
#867440000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#867450000000
0!
1$
0'
1+
0/
#867460000000
1!
1'
1/
#867470000000
0!
0'
0/
#867480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#867490000000
0!
0'
0/
#867500000000
1!
1'
1/
#867510000000
0!
0'
0/
#867520000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#867530000000
0!
0'
0/
#867540000000
1!
1'
1/
#867550000000
0!
0'
0/
#867560000000
1!
1'
1/
#867570000000
0!
0'
0/
#867580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#867590000000
0!
0'
0/
#867600000000
1!
1'
1/
#867610000000
0!
0'
0/
#867620000000
1!
1'
1/
#867630000000
0!
0'
0/
#867640000000
1!
1'
1/
#867650000000
0!
0'
0/
#867660000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#867670000000
0!
0'
0/
#867680000000
1!
1'
1/
#867690000000
0!
0'
0/
#867700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#867710000000
0!
0'
0/
#867720000000
1!
1'
1/
#867730000000
0!
0'
0/
#867740000000
#867750000000
1!
1'
1/
#867760000000
0!
0'
0/
#867770000000
1!
1'
1/
#867780000000
0!
1"
0'
1(
0/
10
#867790000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#867800000000
0!
0'
0/
#867810000000
1!
1'
1/
#867820000000
0!
0'
0/
#867830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#867840000000
0!
0'
0/
#867850000000
1!
1'
1/
#867860000000
0!
1"
0'
1(
0/
10
#867870000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#867880000000
0!
1$
0'
1+
0/
#867890000000
1!
1'
1/
#867900000000
0!
0'
0/
#867910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#867920000000
0!
0'
0/
#867930000000
1!
1'
1/
#867940000000
0!
0'
0/
#867950000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#867960000000
0!
0'
0/
#867970000000
1!
1'
1/
#867980000000
0!
0'
0/
#867990000000
1!
1'
1/
#868000000000
0!
0'
0/
#868010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#868020000000
0!
0'
0/
#868030000000
1!
1'
1/
#868040000000
0!
0'
0/
#868050000000
1!
1'
1/
#868060000000
0!
0'
0/
#868070000000
1!
1'
1/
#868080000000
0!
0'
0/
#868090000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#868100000000
0!
0'
0/
#868110000000
1!
1'
1/
#868120000000
0!
0'
0/
#868130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#868140000000
0!
0'
0/
#868150000000
1!
1'
1/
#868160000000
0!
0'
0/
#868170000000
#868180000000
1!
1'
1/
#868190000000
0!
0'
0/
#868200000000
1!
1'
1/
#868210000000
0!
1"
0'
1(
0/
10
#868220000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#868230000000
0!
0'
0/
#868240000000
1!
1'
1/
#868250000000
0!
0'
0/
#868260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#868270000000
0!
0'
0/
#868280000000
1!
1'
1/
#868290000000
0!
1"
0'
1(
0/
10
#868300000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#868310000000
0!
1$
0'
1+
0/
#868320000000
1!
1'
1/
#868330000000
0!
0'
0/
#868340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#868350000000
0!
0'
0/
#868360000000
1!
1'
1/
#868370000000
0!
0'
0/
#868380000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#868390000000
0!
0'
0/
#868400000000
1!
1'
1/
#868410000000
0!
0'
0/
#868420000000
1!
1'
1/
#868430000000
0!
0'
0/
#868440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#868450000000
0!
0'
0/
#868460000000
1!
1'
1/
#868470000000
0!
0'
0/
#868480000000
1!
1'
1/
#868490000000
0!
0'
0/
#868500000000
1!
1'
1/
#868510000000
0!
0'
0/
#868520000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#868530000000
0!
0'
0/
#868540000000
1!
1'
1/
#868550000000
0!
0'
0/
#868560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#868570000000
0!
0'
0/
#868580000000
1!
1'
1/
#868590000000
0!
0'
0/
#868600000000
#868610000000
1!
1'
1/
#868620000000
0!
0'
0/
#868630000000
1!
1'
1/
#868640000000
0!
1"
0'
1(
0/
10
#868650000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#868660000000
0!
0'
0/
#868670000000
1!
1'
1/
#868680000000
0!
0'
0/
#868690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#868700000000
0!
0'
0/
#868710000000
1!
1'
1/
#868720000000
0!
1"
0'
1(
0/
10
#868730000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#868740000000
0!
1$
0'
1+
0/
#868750000000
1!
1'
1/
#868760000000
0!
0'
0/
#868770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#868780000000
0!
0'
0/
#868790000000
1!
1'
1/
#868800000000
0!
0'
0/
#868810000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#868820000000
0!
0'
0/
#868830000000
1!
1'
1/
#868840000000
0!
0'
0/
#868850000000
1!
1'
1/
#868860000000
0!
0'
0/
#868870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#868880000000
0!
0'
0/
#868890000000
1!
1'
1/
#868900000000
0!
0'
0/
#868910000000
1!
1'
1/
#868920000000
0!
0'
0/
#868930000000
1!
1'
1/
#868940000000
0!
0'
0/
#868950000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#868960000000
0!
0'
0/
#868970000000
1!
1'
1/
#868980000000
0!
0'
0/
#868990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#869000000000
0!
0'
0/
#869010000000
1!
1'
1/
#869020000000
0!
0'
0/
#869030000000
#869040000000
1!
1'
1/
#869050000000
0!
0'
0/
#869060000000
1!
1'
1/
#869070000000
0!
1"
0'
1(
0/
10
#869080000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#869090000000
0!
0'
0/
#869100000000
1!
1'
1/
#869110000000
0!
0'
0/
#869120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#869130000000
0!
0'
0/
#869140000000
1!
1'
1/
#869150000000
0!
1"
0'
1(
0/
10
#869160000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#869170000000
0!
1$
0'
1+
0/
#869180000000
1!
1'
1/
#869190000000
0!
0'
0/
#869200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#869210000000
0!
0'
0/
#869220000000
1!
1'
1/
#869230000000
0!
0'
0/
#869240000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#869250000000
0!
0'
0/
#869260000000
1!
1'
1/
#869270000000
0!
0'
0/
#869280000000
1!
1'
1/
#869290000000
0!
0'
0/
#869300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#869310000000
0!
0'
0/
#869320000000
1!
1'
1/
#869330000000
0!
0'
0/
#869340000000
1!
1'
1/
#869350000000
0!
0'
0/
#869360000000
1!
1'
1/
#869370000000
0!
0'
0/
#869380000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#869390000000
0!
0'
0/
#869400000000
1!
1'
1/
#869410000000
0!
0'
0/
#869420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#869430000000
0!
0'
0/
#869440000000
1!
1'
1/
#869450000000
0!
0'
0/
#869460000000
#869470000000
1!
1'
1/
#869480000000
0!
0'
0/
#869490000000
1!
1'
1/
#869500000000
0!
1"
0'
1(
0/
10
#869510000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#869520000000
0!
0'
0/
#869530000000
1!
1'
1/
#869540000000
0!
0'
0/
#869550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#869560000000
0!
0'
0/
#869570000000
1!
1'
1/
#869580000000
0!
1"
0'
1(
0/
10
#869590000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#869600000000
0!
1$
0'
1+
0/
#869610000000
1!
1'
1/
#869620000000
0!
0'
0/
#869630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#869640000000
0!
0'
0/
#869650000000
1!
1'
1/
#869660000000
0!
0'
0/
#869670000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#869680000000
0!
0'
0/
#869690000000
1!
1'
1/
#869700000000
0!
0'
0/
#869710000000
1!
1'
1/
#869720000000
0!
0'
0/
#869730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#869740000000
0!
0'
0/
#869750000000
1!
1'
1/
#869760000000
0!
0'
0/
#869770000000
1!
1'
1/
#869780000000
0!
0'
0/
#869790000000
1!
1'
1/
#869800000000
0!
0'
0/
#869810000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#869820000000
0!
0'
0/
#869830000000
1!
1'
1/
#869840000000
0!
0'
0/
#869850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#869860000000
0!
0'
0/
#869870000000
1!
1'
1/
#869880000000
0!
0'
0/
#869890000000
#869900000000
1!
1'
1/
#869910000000
0!
0'
0/
#869920000000
1!
1'
1/
#869930000000
0!
1"
0'
1(
0/
10
#869940000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#869950000000
0!
0'
0/
#869960000000
1!
1'
1/
#869970000000
0!
0'
0/
#869980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#869990000000
0!
0'
0/
#870000000000
1!
1'
1/
#870010000000
0!
1"
0'
1(
0/
10
#870020000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#870030000000
0!
1$
0'
1+
0/
#870040000000
1!
1'
1/
#870050000000
0!
0'
0/
#870060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#870070000000
0!
0'
0/
#870080000000
1!
1'
1/
#870090000000
0!
0'
0/
#870100000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#870110000000
0!
0'
0/
#870120000000
1!
1'
1/
#870130000000
0!
0'
0/
#870140000000
1!
1'
1/
#870150000000
0!
0'
0/
#870160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#870170000000
0!
0'
0/
#870180000000
1!
1'
1/
#870190000000
0!
0'
0/
#870200000000
1!
1'
1/
#870210000000
0!
0'
0/
#870220000000
1!
1'
1/
#870230000000
0!
0'
0/
#870240000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#870250000000
0!
0'
0/
#870260000000
1!
1'
1/
#870270000000
0!
0'
0/
#870280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#870290000000
0!
0'
0/
#870300000000
1!
1'
1/
#870310000000
0!
0'
0/
#870320000000
#870330000000
1!
1'
1/
#870340000000
0!
0'
0/
#870350000000
1!
1'
1/
#870360000000
0!
1"
0'
1(
0/
10
#870370000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#870380000000
0!
0'
0/
#870390000000
1!
1'
1/
#870400000000
0!
0'
0/
#870410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#870420000000
0!
0'
0/
#870430000000
1!
1'
1/
#870440000000
0!
1"
0'
1(
0/
10
#870450000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#870460000000
0!
1$
0'
1+
0/
#870470000000
1!
1'
1/
#870480000000
0!
0'
0/
#870490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#870500000000
0!
0'
0/
#870510000000
1!
1'
1/
#870520000000
0!
0'
0/
#870530000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#870540000000
0!
0'
0/
#870550000000
1!
1'
1/
#870560000000
0!
0'
0/
#870570000000
1!
1'
1/
#870580000000
0!
0'
0/
#870590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#870600000000
0!
0'
0/
#870610000000
1!
1'
1/
#870620000000
0!
0'
0/
#870630000000
1!
1'
1/
#870640000000
0!
0'
0/
#870650000000
1!
1'
1/
#870660000000
0!
0'
0/
#870670000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#870680000000
0!
0'
0/
#870690000000
1!
1'
1/
#870700000000
0!
0'
0/
#870710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#870720000000
0!
0'
0/
#870730000000
1!
1'
1/
#870740000000
0!
0'
0/
#870750000000
#870760000000
1!
1'
1/
#870770000000
0!
0'
0/
#870780000000
1!
1'
1/
#870790000000
0!
1"
0'
1(
0/
10
#870800000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#870810000000
0!
0'
0/
#870820000000
1!
1'
1/
#870830000000
0!
0'
0/
#870840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#870850000000
0!
0'
0/
#870860000000
1!
1'
1/
#870870000000
0!
1"
0'
1(
0/
10
#870880000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#870890000000
0!
1$
0'
1+
0/
#870900000000
1!
1'
1/
#870910000000
0!
0'
0/
#870920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#870930000000
0!
0'
0/
#870940000000
1!
1'
1/
#870950000000
0!
0'
0/
#870960000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#870970000000
0!
0'
0/
#870980000000
1!
1'
1/
#870990000000
0!
0'
0/
#871000000000
1!
1'
1/
#871010000000
0!
0'
0/
#871020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#871030000000
0!
0'
0/
#871040000000
1!
1'
1/
#871050000000
0!
0'
0/
#871060000000
1!
1'
1/
#871070000000
0!
0'
0/
#871080000000
1!
1'
1/
#871090000000
0!
0'
0/
#871100000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#871110000000
0!
0'
0/
#871120000000
1!
1'
1/
#871130000000
0!
0'
0/
#871140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#871150000000
0!
0'
0/
#871160000000
1!
1'
1/
#871170000000
0!
0'
0/
#871180000000
#871190000000
1!
1'
1/
#871200000000
0!
0'
0/
#871210000000
1!
1'
1/
#871220000000
0!
1"
0'
1(
0/
10
#871230000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#871240000000
0!
0'
0/
#871250000000
1!
1'
1/
#871260000000
0!
0'
0/
#871270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#871280000000
0!
0'
0/
#871290000000
1!
1'
1/
#871300000000
0!
1"
0'
1(
0/
10
#871310000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#871320000000
0!
1$
0'
1+
0/
#871330000000
1!
1'
1/
#871340000000
0!
0'
0/
#871350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#871360000000
0!
0'
0/
#871370000000
1!
1'
1/
#871380000000
0!
0'
0/
#871390000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#871400000000
0!
0'
0/
#871410000000
1!
1'
1/
#871420000000
0!
0'
0/
#871430000000
1!
1'
1/
#871440000000
0!
0'
0/
#871450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#871460000000
0!
0'
0/
#871470000000
1!
1'
1/
#871480000000
0!
0'
0/
#871490000000
1!
1'
1/
#871500000000
0!
0'
0/
#871510000000
1!
1'
1/
#871520000000
0!
0'
0/
#871530000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#871540000000
0!
0'
0/
#871550000000
1!
1'
1/
#871560000000
0!
0'
0/
#871570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#871580000000
0!
0'
0/
#871590000000
1!
1'
1/
#871600000000
0!
0'
0/
#871610000000
#871620000000
1!
1'
1/
#871630000000
0!
0'
0/
#871640000000
1!
1'
1/
#871650000000
0!
1"
0'
1(
0/
10
#871660000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#871670000000
0!
0'
0/
#871680000000
1!
1'
1/
#871690000000
0!
0'
0/
#871700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#871710000000
0!
0'
0/
#871720000000
1!
1'
1/
#871730000000
0!
1"
0'
1(
0/
10
#871740000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#871750000000
0!
1$
0'
1+
0/
#871760000000
1!
1'
1/
#871770000000
0!
0'
0/
#871780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#871790000000
0!
0'
0/
#871800000000
1!
1'
1/
#871810000000
0!
0'
0/
#871820000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#871830000000
0!
0'
0/
#871840000000
1!
1'
1/
#871850000000
0!
0'
0/
#871860000000
1!
1'
1/
#871870000000
0!
0'
0/
#871880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#871890000000
0!
0'
0/
#871900000000
1!
1'
1/
#871910000000
0!
0'
0/
#871920000000
1!
1'
1/
#871930000000
0!
0'
0/
#871940000000
1!
1'
1/
#871950000000
0!
0'
0/
#871960000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#871970000000
0!
0'
0/
#871980000000
1!
1'
1/
#871990000000
0!
0'
0/
#872000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#872010000000
0!
0'
0/
#872020000000
1!
1'
1/
#872030000000
0!
0'
0/
#872040000000
#872050000000
1!
1'
1/
#872060000000
0!
0'
0/
#872070000000
1!
1'
1/
#872080000000
0!
1"
0'
1(
0/
10
#872090000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#872100000000
0!
0'
0/
#872110000000
1!
1'
1/
#872120000000
0!
0'
0/
#872130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#872140000000
0!
0'
0/
#872150000000
1!
1'
1/
#872160000000
0!
1"
0'
1(
0/
10
#872170000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#872180000000
0!
1$
0'
1+
0/
#872190000000
1!
1'
1/
#872200000000
0!
0'
0/
#872210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#872220000000
0!
0'
0/
#872230000000
1!
1'
1/
#872240000000
0!
0'
0/
#872250000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#872260000000
0!
0'
0/
#872270000000
1!
1'
1/
#872280000000
0!
0'
0/
#872290000000
1!
1'
1/
#872300000000
0!
0'
0/
#872310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#872320000000
0!
0'
0/
#872330000000
1!
1'
1/
#872340000000
0!
0'
0/
#872350000000
1!
1'
1/
#872360000000
0!
0'
0/
#872370000000
1!
1'
1/
#872380000000
0!
0'
0/
#872390000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#872400000000
0!
0'
0/
#872410000000
1!
1'
1/
#872420000000
0!
0'
0/
#872430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#872440000000
0!
0'
0/
#872450000000
1!
1'
1/
#872460000000
0!
0'
0/
#872470000000
#872480000000
1!
1'
1/
#872490000000
0!
0'
0/
#872500000000
1!
1'
1/
#872510000000
0!
1"
0'
1(
0/
10
#872520000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#872530000000
0!
0'
0/
#872540000000
1!
1'
1/
#872550000000
0!
0'
0/
#872560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#872570000000
0!
0'
0/
#872580000000
1!
1'
1/
#872590000000
0!
1"
0'
1(
0/
10
#872600000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#872610000000
0!
1$
0'
1+
0/
#872620000000
1!
1'
1/
#872630000000
0!
0'
0/
#872640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#872650000000
0!
0'
0/
#872660000000
1!
1'
1/
#872670000000
0!
0'
0/
#872680000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#872690000000
0!
0'
0/
#872700000000
1!
1'
1/
#872710000000
0!
0'
0/
#872720000000
1!
1'
1/
#872730000000
0!
0'
0/
#872740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#872750000000
0!
0'
0/
#872760000000
1!
1'
1/
#872770000000
0!
0'
0/
#872780000000
1!
1'
1/
#872790000000
0!
0'
0/
#872800000000
1!
1'
1/
#872810000000
0!
0'
0/
#872820000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#872830000000
0!
0'
0/
#872840000000
1!
1'
1/
#872850000000
0!
0'
0/
#872860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#872870000000
0!
0'
0/
#872880000000
1!
1'
1/
#872890000000
0!
0'
0/
#872900000000
#872910000000
1!
1'
1/
#872920000000
0!
0'
0/
#872930000000
1!
1'
1/
#872940000000
0!
1"
0'
1(
0/
10
#872950000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#872960000000
0!
0'
0/
#872970000000
1!
1'
1/
#872980000000
0!
0'
0/
#872990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#873000000000
0!
0'
0/
#873010000000
1!
1'
1/
#873020000000
0!
1"
0'
1(
0/
10
#873030000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#873040000000
0!
1$
0'
1+
0/
#873050000000
1!
1'
1/
#873060000000
0!
0'
0/
#873070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#873080000000
0!
0'
0/
#873090000000
1!
1'
1/
#873100000000
0!
0'
0/
#873110000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#873120000000
0!
0'
0/
#873130000000
1!
1'
1/
#873140000000
0!
0'
0/
#873150000000
1!
1'
1/
#873160000000
0!
0'
0/
#873170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#873180000000
0!
0'
0/
#873190000000
1!
1'
1/
#873200000000
0!
0'
0/
#873210000000
1!
1'
1/
#873220000000
0!
0'
0/
#873230000000
1!
1'
1/
#873240000000
0!
0'
0/
#873250000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#873260000000
0!
0'
0/
#873270000000
1!
1'
1/
#873280000000
0!
0'
0/
#873290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#873300000000
0!
0'
0/
#873310000000
1!
1'
1/
#873320000000
0!
0'
0/
#873330000000
#873340000000
1!
1'
1/
#873350000000
0!
0'
0/
#873360000000
1!
1'
1/
#873370000000
0!
1"
0'
1(
0/
10
#873380000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#873390000000
0!
0'
0/
#873400000000
1!
1'
1/
#873410000000
0!
0'
0/
#873420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#873430000000
0!
0'
0/
#873440000000
1!
1'
1/
#873450000000
0!
1"
0'
1(
0/
10
#873460000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#873470000000
0!
1$
0'
1+
0/
#873480000000
1!
1'
1/
#873490000000
0!
0'
0/
#873500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#873510000000
0!
0'
0/
#873520000000
1!
1'
1/
#873530000000
0!
0'
0/
#873540000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#873550000000
0!
0'
0/
#873560000000
1!
1'
1/
#873570000000
0!
0'
0/
#873580000000
1!
1'
1/
#873590000000
0!
0'
0/
#873600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#873610000000
0!
0'
0/
#873620000000
1!
1'
1/
#873630000000
0!
0'
0/
#873640000000
1!
1'
1/
#873650000000
0!
0'
0/
#873660000000
1!
1'
1/
#873670000000
0!
0'
0/
#873680000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#873690000000
0!
0'
0/
#873700000000
1!
1'
1/
#873710000000
0!
0'
0/
#873720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#873730000000
0!
0'
0/
#873740000000
1!
1'
1/
#873750000000
0!
0'
0/
#873760000000
#873770000000
1!
1'
1/
#873780000000
0!
0'
0/
#873790000000
1!
1'
1/
#873800000000
0!
1"
0'
1(
0/
10
#873810000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#873820000000
0!
0'
0/
#873830000000
1!
1'
1/
#873840000000
0!
0'
0/
#873850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#873860000000
0!
0'
0/
#873870000000
1!
1'
1/
#873880000000
0!
1"
0'
1(
0/
10
#873890000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#873900000000
0!
1$
0'
1+
0/
#873910000000
1!
1'
1/
#873920000000
0!
0'
0/
#873930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#873940000000
0!
0'
0/
#873950000000
1!
1'
1/
#873960000000
0!
0'
0/
#873970000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#873980000000
0!
0'
0/
#873990000000
1!
1'
1/
#874000000000
0!
0'
0/
#874010000000
1!
1'
1/
#874020000000
0!
0'
0/
#874030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#874040000000
0!
0'
0/
#874050000000
1!
1'
1/
#874060000000
0!
0'
0/
#874070000000
1!
1'
1/
#874080000000
0!
0'
0/
#874090000000
1!
1'
1/
#874100000000
0!
0'
0/
#874110000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#874120000000
0!
0'
0/
#874130000000
1!
1'
1/
#874140000000
0!
0'
0/
#874150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#874160000000
0!
0'
0/
#874170000000
1!
1'
1/
#874180000000
0!
0'
0/
#874190000000
#874200000000
1!
1'
1/
#874210000000
0!
0'
0/
#874220000000
1!
1'
1/
#874230000000
0!
1"
0'
1(
0/
10
#874240000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#874250000000
0!
0'
0/
#874260000000
1!
1'
1/
#874270000000
0!
0'
0/
#874280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#874290000000
0!
0'
0/
#874300000000
1!
1'
1/
#874310000000
0!
1"
0'
1(
0/
10
#874320000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#874330000000
0!
1$
0'
1+
0/
#874340000000
1!
1'
1/
#874350000000
0!
0'
0/
#874360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#874370000000
0!
0'
0/
#874380000000
1!
1'
1/
#874390000000
0!
0'
0/
#874400000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#874410000000
0!
0'
0/
#874420000000
1!
1'
1/
#874430000000
0!
0'
0/
#874440000000
1!
1'
1/
#874450000000
0!
0'
0/
#874460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#874470000000
0!
0'
0/
#874480000000
1!
1'
1/
#874490000000
0!
0'
0/
#874500000000
1!
1'
1/
#874510000000
0!
0'
0/
#874520000000
1!
1'
1/
#874530000000
0!
0'
0/
#874540000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#874550000000
0!
0'
0/
#874560000000
1!
1'
1/
#874570000000
0!
0'
0/
#874580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#874590000000
0!
0'
0/
#874600000000
1!
1'
1/
#874610000000
0!
0'
0/
#874620000000
#874630000000
1!
1'
1/
#874640000000
0!
0'
0/
#874650000000
1!
1'
1/
#874660000000
0!
1"
0'
1(
0/
10
#874670000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#874680000000
0!
0'
0/
#874690000000
1!
1'
1/
#874700000000
0!
0'
0/
#874710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#874720000000
0!
0'
0/
#874730000000
1!
1'
1/
#874740000000
0!
1"
0'
1(
0/
10
#874750000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#874760000000
0!
1$
0'
1+
0/
#874770000000
1!
1'
1/
#874780000000
0!
0'
0/
#874790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#874800000000
0!
0'
0/
#874810000000
1!
1'
1/
#874820000000
0!
0'
0/
#874830000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#874840000000
0!
0'
0/
#874850000000
1!
1'
1/
#874860000000
0!
0'
0/
#874870000000
1!
1'
1/
#874880000000
0!
0'
0/
#874890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#874900000000
0!
0'
0/
#874910000000
1!
1'
1/
#874920000000
0!
0'
0/
#874930000000
1!
1'
1/
#874940000000
0!
0'
0/
#874950000000
1!
1'
1/
#874960000000
0!
0'
0/
#874970000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#874980000000
0!
0'
0/
#874990000000
1!
1'
1/
#875000000000
0!
0'
0/
#875010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#875020000000
0!
0'
0/
#875030000000
1!
1'
1/
#875040000000
0!
0'
0/
#875050000000
#875060000000
1!
1'
1/
#875070000000
0!
0'
0/
#875080000000
1!
1'
1/
#875090000000
0!
1"
0'
1(
0/
10
#875100000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#875110000000
0!
0'
0/
#875120000000
1!
1'
1/
#875130000000
0!
0'
0/
#875140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#875150000000
0!
0'
0/
#875160000000
1!
1'
1/
#875170000000
0!
1"
0'
1(
0/
10
#875180000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#875190000000
0!
1$
0'
1+
0/
#875200000000
1!
1'
1/
#875210000000
0!
0'
0/
#875220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#875230000000
0!
0'
0/
#875240000000
1!
1'
1/
#875250000000
0!
0'
0/
#875260000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#875270000000
0!
0'
0/
#875280000000
1!
1'
1/
#875290000000
0!
0'
0/
#875300000000
1!
1'
1/
#875310000000
0!
0'
0/
#875320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#875330000000
0!
0'
0/
#875340000000
1!
1'
1/
#875350000000
0!
0'
0/
#875360000000
1!
1'
1/
#875370000000
0!
0'
0/
#875380000000
1!
1'
1/
#875390000000
0!
0'
0/
#875400000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#875410000000
0!
0'
0/
#875420000000
1!
1'
1/
#875430000000
0!
0'
0/
#875440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#875450000000
0!
0'
0/
#875460000000
1!
1'
1/
#875470000000
0!
0'
0/
#875480000000
#875490000000
1!
1'
1/
#875500000000
0!
0'
0/
#875510000000
1!
1'
1/
#875520000000
0!
1"
0'
1(
0/
10
#875530000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#875540000000
0!
0'
0/
#875550000000
1!
1'
1/
#875560000000
0!
0'
0/
#875570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#875580000000
0!
0'
0/
#875590000000
1!
1'
1/
#875600000000
0!
1"
0'
1(
0/
10
#875610000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#875620000000
0!
1$
0'
1+
0/
#875630000000
1!
1'
1/
#875640000000
0!
0'
0/
#875650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#875660000000
0!
0'
0/
#875670000000
1!
1'
1/
#875680000000
0!
0'
0/
#875690000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#875700000000
0!
0'
0/
#875710000000
1!
1'
1/
#875720000000
0!
0'
0/
#875730000000
1!
1'
1/
#875740000000
0!
0'
0/
#875750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#875760000000
0!
0'
0/
#875770000000
1!
1'
1/
#875780000000
0!
0'
0/
#875790000000
1!
1'
1/
#875800000000
0!
0'
0/
#875810000000
1!
1'
1/
#875820000000
0!
0'
0/
#875830000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#875840000000
0!
0'
0/
#875850000000
1!
1'
1/
#875860000000
0!
0'
0/
#875870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#875880000000
0!
0'
0/
#875890000000
1!
1'
1/
#875900000000
0!
0'
0/
#875910000000
#875920000000
1!
1'
1/
#875930000000
0!
0'
0/
#875940000000
1!
1'
1/
#875950000000
0!
1"
0'
1(
0/
10
#875960000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#875970000000
0!
0'
0/
#875980000000
1!
1'
1/
#875990000000
0!
0'
0/
#876000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#876010000000
0!
0'
0/
#876020000000
1!
1'
1/
#876030000000
0!
1"
0'
1(
0/
10
#876040000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#876050000000
0!
1$
0'
1+
0/
#876060000000
1!
1'
1/
#876070000000
0!
0'
0/
#876080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#876090000000
0!
0'
0/
#876100000000
1!
1'
1/
#876110000000
0!
0'
0/
#876120000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#876130000000
0!
0'
0/
#876140000000
1!
1'
1/
#876150000000
0!
0'
0/
#876160000000
1!
1'
1/
#876170000000
0!
0'
0/
#876180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#876190000000
0!
0'
0/
#876200000000
1!
1'
1/
#876210000000
0!
0'
0/
#876220000000
1!
1'
1/
#876230000000
0!
0'
0/
#876240000000
1!
1'
1/
#876250000000
0!
0'
0/
#876260000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#876270000000
0!
0'
0/
#876280000000
1!
1'
1/
#876290000000
0!
0'
0/
#876300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#876310000000
0!
0'
0/
#876320000000
1!
1'
1/
#876330000000
0!
0'
0/
#876340000000
#876350000000
1!
1'
1/
#876360000000
0!
0'
0/
#876370000000
1!
1'
1/
#876380000000
0!
1"
0'
1(
0/
10
#876390000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#876400000000
0!
0'
0/
#876410000000
1!
1'
1/
#876420000000
0!
0'
0/
#876430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#876440000000
0!
0'
0/
#876450000000
1!
1'
1/
#876460000000
0!
1"
0'
1(
0/
10
#876470000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#876480000000
0!
1$
0'
1+
0/
#876490000000
1!
1'
1/
#876500000000
0!
0'
0/
#876510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#876520000000
0!
0'
0/
#876530000000
1!
1'
1/
#876540000000
0!
0'
0/
#876550000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#876560000000
0!
0'
0/
#876570000000
1!
1'
1/
#876580000000
0!
0'
0/
#876590000000
1!
1'
1/
#876600000000
0!
0'
0/
#876610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#876620000000
0!
0'
0/
#876630000000
1!
1'
1/
#876640000000
0!
0'
0/
#876650000000
1!
1'
1/
#876660000000
0!
0'
0/
#876670000000
1!
1'
1/
#876680000000
0!
0'
0/
#876690000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#876700000000
0!
0'
0/
#876710000000
1!
1'
1/
#876720000000
0!
0'
0/
#876730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#876740000000
0!
0'
0/
#876750000000
1!
1'
1/
#876760000000
0!
0'
0/
#876770000000
#876780000000
1!
1'
1/
#876790000000
0!
0'
0/
#876800000000
1!
1'
1/
#876810000000
0!
1"
0'
1(
0/
10
#876820000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#876830000000
0!
0'
0/
#876840000000
1!
1'
1/
#876850000000
0!
0'
0/
#876860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#876870000000
0!
0'
0/
#876880000000
1!
1'
1/
#876890000000
0!
1"
0'
1(
0/
10
#876900000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#876910000000
0!
1$
0'
1+
0/
#876920000000
1!
1'
1/
#876930000000
0!
0'
0/
#876940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#876950000000
0!
0'
0/
#876960000000
1!
1'
1/
#876970000000
0!
0'
0/
#876980000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#876990000000
0!
0'
0/
#877000000000
1!
1'
1/
#877010000000
0!
0'
0/
#877020000000
1!
1'
1/
#877030000000
0!
0'
0/
#877040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#877050000000
0!
0'
0/
#877060000000
1!
1'
1/
#877070000000
0!
0'
0/
#877080000000
1!
1'
1/
#877090000000
0!
0'
0/
#877100000000
1!
1'
1/
#877110000000
0!
0'
0/
#877120000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#877130000000
0!
0'
0/
#877140000000
1!
1'
1/
#877150000000
0!
0'
0/
#877160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#877170000000
0!
0'
0/
#877180000000
1!
1'
1/
#877190000000
0!
0'
0/
#877200000000
#877210000000
1!
1'
1/
#877220000000
0!
0'
0/
#877230000000
1!
1'
1/
#877240000000
0!
1"
0'
1(
0/
10
#877250000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#877260000000
0!
0'
0/
#877270000000
1!
1'
1/
#877280000000
0!
0'
0/
#877290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#877300000000
0!
0'
0/
#877310000000
1!
1'
1/
#877320000000
0!
1"
0'
1(
0/
10
#877330000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#877340000000
0!
1$
0'
1+
0/
#877350000000
1!
1'
1/
#877360000000
0!
0'
0/
#877370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#877380000000
0!
0'
0/
#877390000000
1!
1'
1/
#877400000000
0!
0'
0/
#877410000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#877420000000
0!
0'
0/
#877430000000
1!
1'
1/
#877440000000
0!
0'
0/
#877450000000
1!
1'
1/
#877460000000
0!
0'
0/
#877470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#877480000000
0!
0'
0/
#877490000000
1!
1'
1/
#877500000000
0!
0'
0/
#877510000000
1!
1'
1/
#877520000000
0!
0'
0/
#877530000000
1!
1'
1/
#877540000000
0!
0'
0/
#877550000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#877560000000
0!
0'
0/
#877570000000
1!
1'
1/
#877580000000
0!
0'
0/
#877590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#877600000000
0!
0'
0/
#877610000000
1!
1'
1/
#877620000000
0!
0'
0/
#877630000000
#877640000000
1!
1'
1/
#877650000000
0!
0'
0/
#877660000000
1!
1'
1/
#877670000000
0!
1"
0'
1(
0/
10
#877680000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#877690000000
0!
0'
0/
#877700000000
1!
1'
1/
#877710000000
0!
0'
0/
#877720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#877730000000
0!
0'
0/
#877740000000
1!
1'
1/
#877750000000
0!
1"
0'
1(
0/
10
#877760000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#877770000000
0!
1$
0'
1+
0/
#877780000000
1!
1'
1/
#877790000000
0!
0'
0/
#877800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#877810000000
0!
0'
0/
#877820000000
1!
1'
1/
#877830000000
0!
0'
0/
#877840000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#877850000000
0!
0'
0/
#877860000000
1!
1'
1/
#877870000000
0!
0'
0/
#877880000000
1!
1'
1/
#877890000000
0!
0'
0/
#877900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#877910000000
0!
0'
0/
#877920000000
1!
1'
1/
#877930000000
0!
0'
0/
#877940000000
1!
1'
1/
#877950000000
0!
0'
0/
#877960000000
1!
1'
1/
#877970000000
0!
0'
0/
#877980000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#877990000000
0!
0'
0/
#878000000000
1!
1'
1/
#878010000000
0!
0'
0/
#878020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#878030000000
0!
0'
0/
#878040000000
1!
1'
1/
#878050000000
0!
0'
0/
#878060000000
#878070000000
1!
1'
1/
#878080000000
0!
0'
0/
#878090000000
1!
1'
1/
#878100000000
0!
1"
0'
1(
0/
10
#878110000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#878120000000
0!
0'
0/
#878130000000
1!
1'
1/
#878140000000
0!
0'
0/
#878150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#878160000000
0!
0'
0/
#878170000000
1!
1'
1/
#878180000000
0!
1"
0'
1(
0/
10
#878190000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#878200000000
0!
1$
0'
1+
0/
#878210000000
1!
1'
1/
#878220000000
0!
0'
0/
#878230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#878240000000
0!
0'
0/
#878250000000
1!
1'
1/
#878260000000
0!
0'
0/
#878270000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#878280000000
0!
0'
0/
#878290000000
1!
1'
1/
#878300000000
0!
0'
0/
#878310000000
1!
1'
1/
#878320000000
0!
0'
0/
#878330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#878340000000
0!
0'
0/
#878350000000
1!
1'
1/
#878360000000
0!
0'
0/
#878370000000
1!
1'
1/
#878380000000
0!
0'
0/
#878390000000
1!
1'
1/
#878400000000
0!
0'
0/
#878410000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#878420000000
0!
0'
0/
#878430000000
1!
1'
1/
#878440000000
0!
0'
0/
#878450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#878460000000
0!
0'
0/
#878470000000
1!
1'
1/
#878480000000
0!
0'
0/
#878490000000
#878500000000
1!
1'
1/
#878510000000
0!
0'
0/
#878520000000
1!
1'
1/
#878530000000
0!
1"
0'
1(
0/
10
#878540000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#878550000000
0!
0'
0/
#878560000000
1!
1'
1/
#878570000000
0!
0'
0/
#878580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#878590000000
0!
0'
0/
#878600000000
1!
1'
1/
#878610000000
0!
1"
0'
1(
0/
10
#878620000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#878630000000
0!
1$
0'
1+
0/
#878640000000
1!
1'
1/
#878650000000
0!
0'
0/
#878660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#878670000000
0!
0'
0/
#878680000000
1!
1'
1/
#878690000000
0!
0'
0/
#878700000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#878710000000
0!
0'
0/
#878720000000
1!
1'
1/
#878730000000
0!
0'
0/
#878740000000
1!
1'
1/
#878750000000
0!
0'
0/
#878760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#878770000000
0!
0'
0/
#878780000000
1!
1'
1/
#878790000000
0!
0'
0/
#878800000000
1!
1'
1/
#878810000000
0!
0'
0/
#878820000000
1!
1'
1/
#878830000000
0!
0'
0/
#878840000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#878850000000
0!
0'
0/
#878860000000
1!
1'
1/
#878870000000
0!
0'
0/
#878880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#878890000000
0!
0'
0/
#878900000000
1!
1'
1/
#878910000000
0!
0'
0/
#878920000000
#878930000000
1!
1'
1/
#878940000000
0!
0'
0/
#878950000000
1!
1'
1/
#878960000000
0!
1"
0'
1(
0/
10
#878970000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#878980000000
0!
0'
0/
#878990000000
1!
1'
1/
#879000000000
0!
0'
0/
#879010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#879020000000
0!
0'
0/
#879030000000
1!
1'
1/
#879040000000
0!
1"
0'
1(
0/
10
#879050000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#879060000000
0!
1$
0'
1+
0/
#879070000000
1!
1'
1/
#879080000000
0!
0'
0/
#879090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#879100000000
0!
0'
0/
#879110000000
1!
1'
1/
#879120000000
0!
0'
0/
#879130000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#879140000000
0!
0'
0/
#879150000000
1!
1'
1/
#879160000000
0!
0'
0/
#879170000000
1!
1'
1/
#879180000000
0!
0'
0/
#879190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#879200000000
0!
0'
0/
#879210000000
1!
1'
1/
#879220000000
0!
0'
0/
#879230000000
1!
1'
1/
#879240000000
0!
0'
0/
#879250000000
1!
1'
1/
#879260000000
0!
0'
0/
#879270000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#879280000000
0!
0'
0/
#879290000000
1!
1'
1/
#879300000000
0!
0'
0/
#879310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#879320000000
0!
0'
0/
#879330000000
1!
1'
1/
#879340000000
0!
0'
0/
#879350000000
#879360000000
1!
1'
1/
#879370000000
0!
0'
0/
#879380000000
1!
1'
1/
#879390000000
0!
1"
0'
1(
0/
10
#879400000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#879410000000
0!
0'
0/
#879420000000
1!
1'
1/
#879430000000
0!
0'
0/
#879440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#879450000000
0!
0'
0/
#879460000000
1!
1'
1/
#879470000000
0!
1"
0'
1(
0/
10
#879480000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#879490000000
0!
1$
0'
1+
0/
#879500000000
1!
1'
1/
#879510000000
0!
0'
0/
#879520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#879530000000
0!
0'
0/
#879540000000
1!
1'
1/
#879550000000
0!
0'
0/
#879560000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#879570000000
0!
0'
0/
#879580000000
1!
1'
1/
#879590000000
0!
0'
0/
#879600000000
1!
1'
1/
#879610000000
0!
0'
0/
#879620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#879630000000
0!
0'
0/
#879640000000
1!
1'
1/
#879650000000
0!
0'
0/
#879660000000
1!
1'
1/
#879670000000
0!
0'
0/
#879680000000
1!
1'
1/
#879690000000
0!
0'
0/
#879700000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#879710000000
0!
0'
0/
#879720000000
1!
1'
1/
#879730000000
0!
0'
0/
#879740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#879750000000
0!
0'
0/
#879760000000
1!
1'
1/
#879770000000
0!
0'
0/
#879780000000
#879790000000
1!
1'
1/
#879800000000
0!
0'
0/
#879810000000
1!
1'
1/
#879820000000
0!
1"
0'
1(
0/
10
#879830000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#879840000000
0!
0'
0/
#879850000000
1!
1'
1/
#879860000000
0!
0'
0/
#879870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#879880000000
0!
0'
0/
#879890000000
1!
1'
1/
#879900000000
0!
1"
0'
1(
0/
10
#879910000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#879920000000
0!
1$
0'
1+
0/
#879930000000
1!
1'
1/
#879940000000
0!
0'
0/
#879950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#879960000000
0!
0'
0/
#879970000000
1!
1'
1/
#879980000000
0!
0'
0/
#879990000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#880000000000
0!
0'
0/
#880010000000
1!
1'
1/
#880020000000
0!
0'
0/
#880030000000
1!
1'
1/
#880040000000
0!
0'
0/
#880050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#880060000000
0!
0'
0/
#880070000000
1!
1'
1/
#880080000000
0!
0'
0/
#880090000000
1!
1'
1/
#880100000000
0!
0'
0/
#880110000000
1!
1'
1/
#880120000000
0!
0'
0/
#880130000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#880140000000
0!
0'
0/
#880150000000
1!
1'
1/
#880160000000
0!
0'
0/
#880170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#880180000000
0!
0'
0/
#880190000000
1!
1'
1/
#880200000000
0!
0'
0/
#880210000000
#880220000000
1!
1'
1/
#880230000000
0!
0'
0/
#880240000000
1!
1'
1/
#880250000000
0!
1"
0'
1(
0/
10
#880260000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#880270000000
0!
0'
0/
#880280000000
1!
1'
1/
#880290000000
0!
0'
0/
#880300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#880310000000
0!
0'
0/
#880320000000
1!
1'
1/
#880330000000
0!
1"
0'
1(
0/
10
#880340000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#880350000000
0!
1$
0'
1+
0/
#880360000000
1!
1'
1/
#880370000000
0!
0'
0/
#880380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#880390000000
0!
0'
0/
#880400000000
1!
1'
1/
#880410000000
0!
0'
0/
#880420000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#880430000000
0!
0'
0/
#880440000000
1!
1'
1/
#880450000000
0!
0'
0/
#880460000000
1!
1'
1/
#880470000000
0!
0'
0/
#880480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#880490000000
0!
0'
0/
#880500000000
1!
1'
1/
#880510000000
0!
0'
0/
#880520000000
1!
1'
1/
#880530000000
0!
0'
0/
#880540000000
1!
1'
1/
#880550000000
0!
0'
0/
#880560000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#880570000000
0!
0'
0/
#880580000000
1!
1'
1/
#880590000000
0!
0'
0/
#880600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#880610000000
0!
0'
0/
#880620000000
1!
1'
1/
#880630000000
0!
0'
0/
#880640000000
#880650000000
1!
1'
1/
#880660000000
0!
0'
0/
#880670000000
1!
1'
1/
#880680000000
0!
1"
0'
1(
0/
10
#880690000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#880700000000
0!
0'
0/
#880710000000
1!
1'
1/
#880720000000
0!
0'
0/
#880730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#880740000000
0!
0'
0/
#880750000000
1!
1'
1/
#880760000000
0!
1"
0'
1(
0/
10
#880770000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#880780000000
0!
1$
0'
1+
0/
#880790000000
1!
1'
1/
#880800000000
0!
0'
0/
#880810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#880820000000
0!
0'
0/
#880830000000
1!
1'
1/
#880840000000
0!
0'
0/
#880850000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#880860000000
0!
0'
0/
#880870000000
1!
1'
1/
#880880000000
0!
0'
0/
#880890000000
1!
1'
1/
#880900000000
0!
0'
0/
#880910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#880920000000
0!
0'
0/
#880930000000
1!
1'
1/
#880940000000
0!
0'
0/
#880950000000
1!
1'
1/
#880960000000
0!
0'
0/
#880970000000
1!
1'
1/
#880980000000
0!
0'
0/
#880990000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#881000000000
0!
0'
0/
#881010000000
1!
1'
1/
#881020000000
0!
0'
0/
#881030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#881040000000
0!
0'
0/
#881050000000
1!
1'
1/
#881060000000
0!
0'
0/
#881070000000
#881080000000
1!
1'
1/
#881090000000
0!
0'
0/
#881100000000
1!
1'
1/
#881110000000
0!
1"
0'
1(
0/
10
#881120000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#881130000000
0!
0'
0/
#881140000000
1!
1'
1/
#881150000000
0!
0'
0/
#881160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#881170000000
0!
0'
0/
#881180000000
1!
1'
1/
#881190000000
0!
1"
0'
1(
0/
10
#881200000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#881210000000
0!
1$
0'
1+
0/
#881220000000
1!
1'
1/
#881230000000
0!
0'
0/
#881240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#881250000000
0!
0'
0/
#881260000000
1!
1'
1/
#881270000000
0!
0'
0/
#881280000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#881290000000
0!
0'
0/
#881300000000
1!
1'
1/
#881310000000
0!
0'
0/
#881320000000
1!
1'
1/
#881330000000
0!
0'
0/
#881340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#881350000000
0!
0'
0/
#881360000000
1!
1'
1/
#881370000000
0!
0'
0/
#881380000000
1!
1'
1/
#881390000000
0!
0'
0/
#881400000000
1!
1'
1/
#881410000000
0!
0'
0/
#881420000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#881430000000
0!
0'
0/
#881440000000
1!
1'
1/
#881450000000
0!
0'
0/
#881460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#881470000000
0!
0'
0/
#881480000000
1!
1'
1/
#881490000000
0!
0'
0/
#881500000000
#881510000000
1!
1'
1/
#881520000000
0!
0'
0/
#881530000000
1!
1'
1/
#881540000000
0!
1"
0'
1(
0/
10
#881550000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#881560000000
0!
0'
0/
#881570000000
1!
1'
1/
#881580000000
0!
0'
0/
#881590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#881600000000
0!
0'
0/
#881610000000
1!
1'
1/
#881620000000
0!
1"
0'
1(
0/
10
#881630000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#881640000000
0!
1$
0'
1+
0/
#881650000000
1!
1'
1/
#881660000000
0!
0'
0/
#881670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#881680000000
0!
0'
0/
#881690000000
1!
1'
1/
#881700000000
0!
0'
0/
#881710000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#881720000000
0!
0'
0/
#881730000000
1!
1'
1/
#881740000000
0!
0'
0/
#881750000000
1!
1'
1/
#881760000000
0!
0'
0/
#881770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#881780000000
0!
0'
0/
#881790000000
1!
1'
1/
#881800000000
0!
0'
0/
#881810000000
1!
1'
1/
#881820000000
0!
0'
0/
#881830000000
1!
1'
1/
#881840000000
0!
0'
0/
#881850000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#881860000000
0!
0'
0/
#881870000000
1!
1'
1/
#881880000000
0!
0'
0/
#881890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#881900000000
0!
0'
0/
#881910000000
1!
1'
1/
#881920000000
0!
0'
0/
#881930000000
#881940000000
1!
1'
1/
#881950000000
0!
0'
0/
#881960000000
1!
1'
1/
#881970000000
0!
1"
0'
1(
0/
10
#881980000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#881990000000
0!
0'
0/
#882000000000
1!
1'
1/
#882010000000
0!
0'
0/
#882020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#882030000000
0!
0'
0/
#882040000000
1!
1'
1/
#882050000000
0!
1"
0'
1(
0/
10
#882060000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#882070000000
0!
1$
0'
1+
0/
#882080000000
1!
1'
1/
#882090000000
0!
0'
0/
#882100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#882110000000
0!
0'
0/
#882120000000
1!
1'
1/
#882130000000
0!
0'
0/
#882140000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#882150000000
0!
0'
0/
#882160000000
1!
1'
1/
#882170000000
0!
0'
0/
#882180000000
1!
1'
1/
#882190000000
0!
0'
0/
#882200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#882210000000
0!
0'
0/
#882220000000
1!
1'
1/
#882230000000
0!
0'
0/
#882240000000
1!
1'
1/
#882250000000
0!
0'
0/
#882260000000
1!
1'
1/
#882270000000
0!
0'
0/
#882280000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#882290000000
0!
0'
0/
#882300000000
1!
1'
1/
#882310000000
0!
0'
0/
#882320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#882330000000
0!
0'
0/
#882340000000
1!
1'
1/
#882350000000
0!
0'
0/
#882360000000
#882370000000
1!
1'
1/
#882380000000
0!
0'
0/
#882390000000
1!
1'
1/
#882400000000
0!
1"
0'
1(
0/
10
#882410000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#882420000000
0!
0'
0/
#882430000000
1!
1'
1/
#882440000000
0!
0'
0/
#882450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#882460000000
0!
0'
0/
#882470000000
1!
1'
1/
#882480000000
0!
1"
0'
1(
0/
10
#882490000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#882500000000
0!
1$
0'
1+
0/
#882510000000
1!
1'
1/
#882520000000
0!
0'
0/
#882530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#882540000000
0!
0'
0/
#882550000000
1!
1'
1/
#882560000000
0!
0'
0/
#882570000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#882580000000
0!
0'
0/
#882590000000
1!
1'
1/
#882600000000
0!
0'
0/
#882610000000
1!
1'
1/
#882620000000
0!
0'
0/
#882630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#882640000000
0!
0'
0/
#882650000000
1!
1'
1/
#882660000000
0!
0'
0/
#882670000000
1!
1'
1/
#882680000000
0!
0'
0/
#882690000000
1!
1'
1/
#882700000000
0!
0'
0/
#882710000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#882720000000
0!
0'
0/
#882730000000
1!
1'
1/
#882740000000
0!
0'
0/
#882750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#882760000000
0!
0'
0/
#882770000000
1!
1'
1/
#882780000000
0!
0'
0/
#882790000000
#882800000000
1!
1'
1/
#882810000000
0!
0'
0/
#882820000000
1!
1'
1/
#882830000000
0!
1"
0'
1(
0/
10
#882840000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#882850000000
0!
0'
0/
#882860000000
1!
1'
1/
#882870000000
0!
0'
0/
#882880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#882890000000
0!
0'
0/
#882900000000
1!
1'
1/
#882910000000
0!
1"
0'
1(
0/
10
#882920000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#882930000000
0!
1$
0'
1+
0/
#882940000000
1!
1'
1/
#882950000000
0!
0'
0/
#882960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#882970000000
0!
0'
0/
#882980000000
1!
1'
1/
#882990000000
0!
0'
0/
#883000000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#883010000000
0!
0'
0/
#883020000000
1!
1'
1/
#883030000000
0!
0'
0/
#883040000000
1!
1'
1/
#883050000000
0!
0'
0/
#883060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#883070000000
0!
0'
0/
#883080000000
1!
1'
1/
#883090000000
0!
0'
0/
#883100000000
1!
1'
1/
#883110000000
0!
0'
0/
#883120000000
1!
1'
1/
#883130000000
0!
0'
0/
#883140000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#883150000000
0!
0'
0/
#883160000000
1!
1'
1/
#883170000000
0!
0'
0/
#883180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#883190000000
0!
0'
0/
#883200000000
1!
1'
1/
#883210000000
0!
0'
0/
#883220000000
#883230000000
1!
1'
1/
#883240000000
0!
0'
0/
#883250000000
1!
1'
1/
#883260000000
0!
1"
0'
1(
0/
10
#883270000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#883280000000
0!
0'
0/
#883290000000
1!
1'
1/
#883300000000
0!
0'
0/
#883310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#883320000000
0!
0'
0/
#883330000000
1!
1'
1/
#883340000000
0!
1"
0'
1(
0/
10
#883350000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#883360000000
0!
1$
0'
1+
0/
#883370000000
1!
1'
1/
#883380000000
0!
0'
0/
#883390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#883400000000
0!
0'
0/
#883410000000
1!
1'
1/
#883420000000
0!
0'
0/
#883430000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#883440000000
0!
0'
0/
#883450000000
1!
1'
1/
#883460000000
0!
0'
0/
#883470000000
1!
1'
1/
#883480000000
0!
0'
0/
#883490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#883500000000
0!
0'
0/
#883510000000
1!
1'
1/
#883520000000
0!
0'
0/
#883530000000
1!
1'
1/
#883540000000
0!
0'
0/
#883550000000
1!
1'
1/
#883560000000
0!
0'
0/
#883570000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#883580000000
0!
0'
0/
#883590000000
1!
1'
1/
#883600000000
0!
0'
0/
#883610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#883620000000
0!
0'
0/
#883630000000
1!
1'
1/
#883640000000
0!
0'
0/
#883650000000
#883660000000
1!
1'
1/
#883670000000
0!
0'
0/
#883680000000
1!
1'
1/
#883690000000
0!
1"
0'
1(
0/
10
#883700000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#883710000000
0!
0'
0/
#883720000000
1!
1'
1/
#883730000000
0!
0'
0/
#883740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#883750000000
0!
0'
0/
#883760000000
1!
1'
1/
#883770000000
0!
1"
0'
1(
0/
10
#883780000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#883790000000
0!
1$
0'
1+
0/
#883800000000
1!
1'
1/
#883810000000
0!
0'
0/
#883820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#883830000000
0!
0'
0/
#883840000000
1!
1'
1/
#883850000000
0!
0'
0/
#883860000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#883870000000
0!
0'
0/
#883880000000
1!
1'
1/
#883890000000
0!
0'
0/
#883900000000
1!
1'
1/
#883910000000
0!
0'
0/
#883920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#883930000000
0!
0'
0/
#883940000000
1!
1'
1/
#883950000000
0!
0'
0/
#883960000000
1!
1'
1/
#883970000000
0!
0'
0/
#883980000000
1!
1'
1/
#883990000000
0!
0'
0/
#884000000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#884010000000
0!
0'
0/
#884020000000
1!
1'
1/
#884030000000
0!
0'
0/
#884040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#884050000000
0!
0'
0/
#884060000000
1!
1'
1/
#884070000000
0!
0'
0/
#884080000000
#884090000000
1!
1'
1/
#884100000000
0!
0'
0/
#884110000000
1!
1'
1/
#884120000000
0!
1"
0'
1(
0/
10
#884130000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#884140000000
0!
0'
0/
#884150000000
1!
1'
1/
#884160000000
0!
0'
0/
#884170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#884180000000
0!
0'
0/
#884190000000
1!
1'
1/
#884200000000
0!
1"
0'
1(
0/
10
#884210000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#884220000000
0!
1$
0'
1+
0/
#884230000000
1!
1'
1/
#884240000000
0!
0'
0/
#884250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#884260000000
0!
0'
0/
#884270000000
1!
1'
1/
#884280000000
0!
0'
0/
#884290000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#884300000000
0!
0'
0/
#884310000000
1!
1'
1/
#884320000000
0!
0'
0/
#884330000000
1!
1'
1/
#884340000000
0!
0'
0/
#884350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#884360000000
0!
0'
0/
#884370000000
1!
1'
1/
#884380000000
0!
0'
0/
#884390000000
1!
1'
1/
#884400000000
0!
0'
0/
#884410000000
1!
1'
1/
#884420000000
0!
0'
0/
#884430000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#884440000000
0!
0'
0/
#884450000000
1!
1'
1/
#884460000000
0!
0'
0/
#884470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#884480000000
0!
0'
0/
#884490000000
1!
1'
1/
#884500000000
0!
0'
0/
#884510000000
#884520000000
1!
1'
1/
#884530000000
0!
0'
0/
#884540000000
1!
1'
1/
#884550000000
0!
1"
0'
1(
0/
10
#884560000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#884570000000
0!
0'
0/
#884580000000
1!
1'
1/
#884590000000
0!
0'
0/
#884600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#884610000000
0!
0'
0/
#884620000000
1!
1'
1/
#884630000000
0!
1"
0'
1(
0/
10
#884640000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#884650000000
0!
1$
0'
1+
0/
#884660000000
1!
1'
1/
#884670000000
0!
0'
0/
#884680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#884690000000
0!
0'
0/
#884700000000
1!
1'
1/
#884710000000
0!
0'
0/
#884720000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#884730000000
0!
0'
0/
#884740000000
1!
1'
1/
#884750000000
0!
0'
0/
#884760000000
1!
1'
1/
#884770000000
0!
0'
0/
#884780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#884790000000
0!
0'
0/
#884800000000
1!
1'
1/
#884810000000
0!
0'
0/
#884820000000
1!
1'
1/
#884830000000
0!
0'
0/
#884840000000
1!
1'
1/
#884850000000
0!
0'
0/
#884860000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#884870000000
0!
0'
0/
#884880000000
1!
1'
1/
#884890000000
0!
0'
0/
#884900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#884910000000
0!
0'
0/
#884920000000
1!
1'
1/
#884930000000
0!
0'
0/
#884940000000
#884950000000
1!
1'
1/
#884960000000
0!
0'
0/
#884970000000
1!
1'
1/
#884980000000
0!
1"
0'
1(
0/
10
#884990000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#885000000000
0!
0'
0/
#885010000000
1!
1'
1/
#885020000000
0!
0'
0/
#885030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#885040000000
0!
0'
0/
#885050000000
1!
1'
1/
#885060000000
0!
1"
0'
1(
0/
10
#885070000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#885080000000
0!
1$
0'
1+
0/
#885090000000
1!
1'
1/
#885100000000
0!
0'
0/
#885110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#885120000000
0!
0'
0/
#885130000000
1!
1'
1/
#885140000000
0!
0'
0/
#885150000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#885160000000
0!
0'
0/
#885170000000
1!
1'
1/
#885180000000
0!
0'
0/
#885190000000
1!
1'
1/
#885200000000
0!
0'
0/
#885210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#885220000000
0!
0'
0/
#885230000000
1!
1'
1/
#885240000000
0!
0'
0/
#885250000000
1!
1'
1/
#885260000000
0!
0'
0/
#885270000000
1!
1'
1/
#885280000000
0!
0'
0/
#885290000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#885300000000
0!
0'
0/
#885310000000
1!
1'
1/
#885320000000
0!
0'
0/
#885330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#885340000000
0!
0'
0/
#885350000000
1!
1'
1/
#885360000000
0!
0'
0/
#885370000000
#885380000000
1!
1'
1/
#885390000000
0!
0'
0/
#885400000000
1!
1'
1/
#885410000000
0!
1"
0'
1(
0/
10
#885420000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#885430000000
0!
0'
0/
#885440000000
1!
1'
1/
#885450000000
0!
0'
0/
#885460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#885470000000
0!
0'
0/
#885480000000
1!
1'
1/
#885490000000
0!
1"
0'
1(
0/
10
#885500000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#885510000000
0!
1$
0'
1+
0/
#885520000000
1!
1'
1/
#885530000000
0!
0'
0/
#885540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#885550000000
0!
0'
0/
#885560000000
1!
1'
1/
#885570000000
0!
0'
0/
#885580000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#885590000000
0!
0'
0/
#885600000000
1!
1'
1/
#885610000000
0!
0'
0/
#885620000000
1!
1'
1/
#885630000000
0!
0'
0/
#885640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#885650000000
0!
0'
0/
#885660000000
1!
1'
1/
#885670000000
0!
0'
0/
#885680000000
1!
1'
1/
#885690000000
0!
0'
0/
#885700000000
1!
1'
1/
#885710000000
0!
0'
0/
#885720000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#885730000000
0!
0'
0/
#885740000000
1!
1'
1/
#885750000000
0!
0'
0/
#885760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#885770000000
0!
0'
0/
#885780000000
1!
1'
1/
#885790000000
0!
0'
0/
#885800000000
#885810000000
1!
1'
1/
#885820000000
0!
0'
0/
#885830000000
1!
1'
1/
#885840000000
0!
1"
0'
1(
0/
10
#885850000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#885860000000
0!
0'
0/
#885870000000
1!
1'
1/
#885880000000
0!
0'
0/
#885890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#885900000000
0!
0'
0/
#885910000000
1!
1'
1/
#885920000000
0!
1"
0'
1(
0/
10
#885930000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#885940000000
0!
1$
0'
1+
0/
#885950000000
1!
1'
1/
#885960000000
0!
0'
0/
#885970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#885980000000
0!
0'
0/
#885990000000
1!
1'
1/
#886000000000
0!
0'
0/
#886010000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#886020000000
0!
0'
0/
#886030000000
1!
1'
1/
#886040000000
0!
0'
0/
#886050000000
1!
1'
1/
#886060000000
0!
0'
0/
#886070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#886080000000
0!
0'
0/
#886090000000
1!
1'
1/
#886100000000
0!
0'
0/
#886110000000
1!
1'
1/
#886120000000
0!
0'
0/
#886130000000
1!
1'
1/
#886140000000
0!
0'
0/
#886150000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#886160000000
0!
0'
0/
#886170000000
1!
1'
1/
#886180000000
0!
0'
0/
#886190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#886200000000
0!
0'
0/
#886210000000
1!
1'
1/
#886220000000
0!
0'
0/
#886230000000
#886240000000
1!
1'
1/
#886250000000
0!
0'
0/
#886260000000
1!
1'
1/
#886270000000
0!
1"
0'
1(
0/
10
#886280000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#886290000000
0!
0'
0/
#886300000000
1!
1'
1/
#886310000000
0!
0'
0/
#886320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#886330000000
0!
0'
0/
#886340000000
1!
1'
1/
#886350000000
0!
1"
0'
1(
0/
10
#886360000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#886370000000
0!
1$
0'
1+
0/
#886380000000
1!
1'
1/
#886390000000
0!
0'
0/
#886400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#886410000000
0!
0'
0/
#886420000000
1!
1'
1/
#886430000000
0!
0'
0/
#886440000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#886450000000
0!
0'
0/
#886460000000
1!
1'
1/
#886470000000
0!
0'
0/
#886480000000
1!
1'
1/
#886490000000
0!
0'
0/
#886500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#886510000000
0!
0'
0/
#886520000000
1!
1'
1/
#886530000000
0!
0'
0/
#886540000000
1!
1'
1/
#886550000000
0!
0'
0/
#886560000000
1!
1'
1/
#886570000000
0!
0'
0/
#886580000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#886590000000
0!
0'
0/
#886600000000
1!
1'
1/
#886610000000
0!
0'
0/
#886620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#886630000000
0!
0'
0/
#886640000000
1!
1'
1/
#886650000000
0!
0'
0/
#886660000000
#886670000000
1!
1'
1/
#886680000000
0!
0'
0/
#886690000000
1!
1'
1/
#886700000000
0!
1"
0'
1(
0/
10
#886710000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#886720000000
0!
0'
0/
#886730000000
1!
1'
1/
#886740000000
0!
0'
0/
#886750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#886760000000
0!
0'
0/
#886770000000
1!
1'
1/
#886780000000
0!
1"
0'
1(
0/
10
#886790000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#886800000000
0!
1$
0'
1+
0/
#886810000000
1!
1'
1/
#886820000000
0!
0'
0/
#886830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#886840000000
0!
0'
0/
#886850000000
1!
1'
1/
#886860000000
0!
0'
0/
#886870000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#886880000000
0!
0'
0/
#886890000000
1!
1'
1/
#886900000000
0!
0'
0/
#886910000000
1!
1'
1/
#886920000000
0!
0'
0/
#886930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#886940000000
0!
0'
0/
#886950000000
1!
1'
1/
#886960000000
0!
0'
0/
#886970000000
1!
1'
1/
#886980000000
0!
0'
0/
#886990000000
1!
1'
1/
#887000000000
0!
0'
0/
#887010000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#887020000000
0!
0'
0/
#887030000000
1!
1'
1/
#887040000000
0!
0'
0/
#887050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#887060000000
0!
0'
0/
#887070000000
1!
1'
1/
#887080000000
0!
0'
0/
#887090000000
#887100000000
1!
1'
1/
#887110000000
0!
0'
0/
#887120000000
1!
1'
1/
#887130000000
0!
1"
0'
1(
0/
10
#887140000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#887150000000
0!
0'
0/
#887160000000
1!
1'
1/
#887170000000
0!
0'
0/
#887180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#887190000000
0!
0'
0/
#887200000000
1!
1'
1/
#887210000000
0!
1"
0'
1(
0/
10
#887220000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#887230000000
0!
1$
0'
1+
0/
#887240000000
1!
1'
1/
#887250000000
0!
0'
0/
#887260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#887270000000
0!
0'
0/
#887280000000
1!
1'
1/
#887290000000
0!
0'
0/
#887300000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#887310000000
0!
0'
0/
#887320000000
1!
1'
1/
#887330000000
0!
0'
0/
#887340000000
1!
1'
1/
#887350000000
0!
0'
0/
#887360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#887370000000
0!
0'
0/
#887380000000
1!
1'
1/
#887390000000
0!
0'
0/
#887400000000
1!
1'
1/
#887410000000
0!
0'
0/
#887420000000
1!
1'
1/
#887430000000
0!
0'
0/
#887440000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#887450000000
0!
0'
0/
#887460000000
1!
1'
1/
#887470000000
0!
0'
0/
#887480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#887490000000
0!
0'
0/
#887500000000
1!
1'
1/
#887510000000
0!
0'
0/
#887520000000
#887530000000
1!
1'
1/
#887540000000
0!
0'
0/
#887550000000
1!
1'
1/
#887560000000
0!
1"
0'
1(
0/
10
#887570000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#887580000000
0!
0'
0/
#887590000000
1!
1'
1/
#887600000000
0!
0'
0/
#887610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#887620000000
0!
0'
0/
#887630000000
1!
1'
1/
#887640000000
0!
1"
0'
1(
0/
10
#887650000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#887660000000
0!
1$
0'
1+
0/
#887670000000
1!
1'
1/
#887680000000
0!
0'
0/
#887690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#887700000000
0!
0'
0/
#887710000000
1!
1'
1/
#887720000000
0!
0'
0/
#887730000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#887740000000
0!
0'
0/
#887750000000
1!
1'
1/
#887760000000
0!
0'
0/
#887770000000
1!
1'
1/
#887780000000
0!
0'
0/
#887790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#887800000000
0!
0'
0/
#887810000000
1!
1'
1/
#887820000000
0!
0'
0/
#887830000000
1!
1'
1/
#887840000000
0!
0'
0/
#887850000000
1!
1'
1/
#887860000000
0!
0'
0/
#887870000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#887880000000
0!
0'
0/
#887890000000
1!
1'
1/
#887900000000
0!
0'
0/
#887910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#887920000000
0!
0'
0/
#887930000000
1!
1'
1/
#887940000000
0!
0'
0/
#887950000000
#887960000000
1!
1'
1/
#887970000000
0!
0'
0/
#887980000000
1!
1'
1/
#887990000000
0!
1"
0'
1(
0/
10
#888000000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#888010000000
0!
0'
0/
#888020000000
1!
1'
1/
#888030000000
0!
0'
0/
#888040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#888050000000
0!
0'
0/
#888060000000
1!
1'
1/
#888070000000
0!
1"
0'
1(
0/
10
#888080000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#888090000000
0!
1$
0'
1+
0/
#888100000000
1!
1'
1/
#888110000000
0!
0'
0/
#888120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#888130000000
0!
0'
0/
#888140000000
1!
1'
1/
#888150000000
0!
0'
0/
#888160000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#888170000000
0!
0'
0/
#888180000000
1!
1'
1/
#888190000000
0!
0'
0/
#888200000000
1!
1'
1/
#888210000000
0!
0'
0/
#888220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#888230000000
0!
0'
0/
#888240000000
1!
1'
1/
#888250000000
0!
0'
0/
#888260000000
1!
1'
1/
#888270000000
0!
0'
0/
#888280000000
1!
1'
1/
#888290000000
0!
0'
0/
#888300000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#888310000000
0!
0'
0/
#888320000000
1!
1'
1/
#888330000000
0!
0'
0/
#888340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#888350000000
0!
0'
0/
#888360000000
1!
1'
1/
#888370000000
0!
0'
0/
#888380000000
#888390000000
1!
1'
1/
#888400000000
0!
0'
0/
#888410000000
1!
1'
1/
#888420000000
0!
1"
0'
1(
0/
10
#888430000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#888440000000
0!
0'
0/
#888450000000
1!
1'
1/
#888460000000
0!
0'
0/
#888470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#888480000000
0!
0'
0/
#888490000000
1!
1'
1/
#888500000000
0!
1"
0'
1(
0/
10
#888510000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#888520000000
0!
1$
0'
1+
0/
#888530000000
1!
1'
1/
#888540000000
0!
0'
0/
#888550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#888560000000
0!
0'
0/
#888570000000
1!
1'
1/
#888580000000
0!
0'
0/
#888590000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#888600000000
0!
0'
0/
#888610000000
1!
1'
1/
#888620000000
0!
0'
0/
#888630000000
1!
1'
1/
#888640000000
0!
0'
0/
#888650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#888660000000
0!
0'
0/
#888670000000
1!
1'
1/
#888680000000
0!
0'
0/
#888690000000
1!
1'
1/
#888700000000
0!
0'
0/
#888710000000
1!
1'
1/
#888720000000
0!
0'
0/
#888730000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#888740000000
0!
0'
0/
#888750000000
1!
1'
1/
#888760000000
0!
0'
0/
#888770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#888780000000
0!
0'
0/
#888790000000
1!
1'
1/
#888800000000
0!
0'
0/
#888810000000
#888820000000
1!
1'
1/
#888830000000
0!
0'
0/
#888840000000
1!
1'
1/
#888850000000
0!
1"
0'
1(
0/
10
#888860000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#888870000000
0!
0'
0/
#888880000000
1!
1'
1/
#888890000000
0!
0'
0/
#888900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#888910000000
0!
0'
0/
#888920000000
1!
1'
1/
#888930000000
0!
1"
0'
1(
0/
10
#888940000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#888950000000
0!
1$
0'
1+
0/
#888960000000
1!
1'
1/
#888970000000
0!
0'
0/
#888980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#888990000000
0!
0'
0/
#889000000000
1!
1'
1/
#889010000000
0!
0'
0/
#889020000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#889030000000
0!
0'
0/
#889040000000
1!
1'
1/
#889050000000
0!
0'
0/
#889060000000
1!
1'
1/
#889070000000
0!
0'
0/
#889080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#889090000000
0!
0'
0/
#889100000000
1!
1'
1/
#889110000000
0!
0'
0/
#889120000000
1!
1'
1/
#889130000000
0!
0'
0/
#889140000000
1!
1'
1/
#889150000000
0!
0'
0/
#889160000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#889170000000
0!
0'
0/
#889180000000
1!
1'
1/
#889190000000
0!
0'
0/
#889200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#889210000000
0!
0'
0/
#889220000000
1!
1'
1/
#889230000000
0!
0'
0/
#889240000000
#889250000000
1!
1'
1/
#889260000000
0!
0'
0/
#889270000000
1!
1'
1/
#889280000000
0!
1"
0'
1(
0/
10
#889290000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#889300000000
0!
0'
0/
#889310000000
1!
1'
1/
#889320000000
0!
0'
0/
#889330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#889340000000
0!
0'
0/
#889350000000
1!
1'
1/
#889360000000
0!
1"
0'
1(
0/
10
#889370000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#889380000000
0!
1$
0'
1+
0/
#889390000000
1!
1'
1/
#889400000000
0!
0'
0/
#889410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#889420000000
0!
0'
0/
#889430000000
1!
1'
1/
#889440000000
0!
0'
0/
#889450000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#889460000000
0!
0'
0/
#889470000000
1!
1'
1/
#889480000000
0!
0'
0/
#889490000000
1!
1'
1/
#889500000000
0!
0'
0/
#889510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#889520000000
0!
0'
0/
#889530000000
1!
1'
1/
#889540000000
0!
0'
0/
#889550000000
1!
1'
1/
#889560000000
0!
0'
0/
#889570000000
1!
1'
1/
#889580000000
0!
0'
0/
#889590000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#889600000000
0!
0'
0/
#889610000000
1!
1'
1/
#889620000000
0!
0'
0/
#889630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#889640000000
0!
0'
0/
#889650000000
1!
1'
1/
#889660000000
0!
0'
0/
#889670000000
#889680000000
1!
1'
1/
#889690000000
0!
0'
0/
#889700000000
1!
1'
1/
#889710000000
0!
1"
0'
1(
0/
10
#889720000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#889730000000
0!
0'
0/
#889740000000
1!
1'
1/
#889750000000
0!
0'
0/
#889760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#889770000000
0!
0'
0/
#889780000000
1!
1'
1/
#889790000000
0!
1"
0'
1(
0/
10
#889800000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#889810000000
0!
1$
0'
1+
0/
#889820000000
1!
1'
1/
#889830000000
0!
0'
0/
#889840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#889850000000
0!
0'
0/
#889860000000
1!
1'
1/
#889870000000
0!
0'
0/
#889880000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#889890000000
0!
0'
0/
#889900000000
1!
1'
1/
#889910000000
0!
0'
0/
#889920000000
1!
1'
1/
#889930000000
0!
0'
0/
#889940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#889950000000
0!
0'
0/
#889960000000
1!
1'
1/
#889970000000
0!
0'
0/
#889980000000
1!
1'
1/
#889990000000
0!
0'
0/
#890000000000
1!
1'
1/
#890010000000
0!
0'
0/
#890020000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#890030000000
0!
0'
0/
#890040000000
1!
1'
1/
#890050000000
0!
0'
0/
#890060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#890070000000
0!
0'
0/
#890080000000
1!
1'
1/
#890090000000
0!
0'
0/
#890100000000
#890110000000
1!
1'
1/
#890120000000
0!
0'
0/
#890130000000
1!
1'
1/
#890140000000
0!
1"
0'
1(
0/
10
#890150000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#890160000000
0!
0'
0/
#890170000000
1!
1'
1/
#890180000000
0!
0'
0/
#890190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#890200000000
0!
0'
0/
#890210000000
1!
1'
1/
#890220000000
0!
1"
0'
1(
0/
10
#890230000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#890240000000
0!
1$
0'
1+
0/
#890250000000
1!
1'
1/
#890260000000
0!
0'
0/
#890270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#890280000000
0!
0'
0/
#890290000000
1!
1'
1/
#890300000000
0!
0'
0/
#890310000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#890320000000
0!
0'
0/
#890330000000
1!
1'
1/
#890340000000
0!
0'
0/
#890350000000
1!
1'
1/
#890360000000
0!
0'
0/
#890370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#890380000000
0!
0'
0/
#890390000000
1!
1'
1/
#890400000000
0!
0'
0/
#890410000000
1!
1'
1/
#890420000000
0!
0'
0/
#890430000000
1!
1'
1/
#890440000000
0!
0'
0/
#890450000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#890460000000
0!
0'
0/
#890470000000
1!
1'
1/
#890480000000
0!
0'
0/
#890490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#890500000000
0!
0'
0/
#890510000000
1!
1'
1/
#890520000000
0!
0'
0/
#890530000000
#890540000000
1!
1'
1/
#890550000000
0!
0'
0/
#890560000000
1!
1'
1/
#890570000000
0!
1"
0'
1(
0/
10
#890580000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#890590000000
0!
0'
0/
#890600000000
1!
1'
1/
#890610000000
0!
0'
0/
#890620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#890630000000
0!
0'
0/
#890640000000
1!
1'
1/
#890650000000
0!
1"
0'
1(
0/
10
#890660000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#890670000000
0!
1$
0'
1+
0/
#890680000000
1!
1'
1/
#890690000000
0!
0'
0/
#890700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#890710000000
0!
0'
0/
#890720000000
1!
1'
1/
#890730000000
0!
0'
0/
#890740000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#890750000000
0!
0'
0/
#890760000000
1!
1'
1/
#890770000000
0!
0'
0/
#890780000000
1!
1'
1/
#890790000000
0!
0'
0/
#890800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#890810000000
0!
0'
0/
#890820000000
1!
1'
1/
#890830000000
0!
0'
0/
#890840000000
1!
1'
1/
#890850000000
0!
0'
0/
#890860000000
1!
1'
1/
#890870000000
0!
0'
0/
#890880000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#890890000000
0!
0'
0/
#890900000000
1!
1'
1/
#890910000000
0!
0'
0/
#890920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#890930000000
0!
0'
0/
#890940000000
1!
1'
1/
#890950000000
0!
0'
0/
#890960000000
#890970000000
1!
1'
1/
#890980000000
0!
0'
0/
#890990000000
1!
1'
1/
#891000000000
0!
1"
0'
1(
0/
10
#891010000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#891020000000
0!
0'
0/
#891030000000
1!
1'
1/
#891040000000
0!
0'
0/
#891050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#891060000000
0!
0'
0/
#891070000000
1!
1'
1/
#891080000000
0!
1"
0'
1(
0/
10
#891090000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#891100000000
0!
1$
0'
1+
0/
#891110000000
1!
1'
1/
#891120000000
0!
0'
0/
#891130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#891140000000
0!
0'
0/
#891150000000
1!
1'
1/
#891160000000
0!
0'
0/
#891170000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#891180000000
0!
0'
0/
#891190000000
1!
1'
1/
#891200000000
0!
0'
0/
#891210000000
1!
1'
1/
#891220000000
0!
0'
0/
#891230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#891240000000
0!
0'
0/
#891250000000
1!
1'
1/
#891260000000
0!
0'
0/
#891270000000
1!
1'
1/
#891280000000
0!
0'
0/
#891290000000
1!
1'
1/
#891300000000
0!
0'
0/
#891310000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#891320000000
0!
0'
0/
#891330000000
1!
1'
1/
#891340000000
0!
0'
0/
#891350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#891360000000
0!
0'
0/
#891370000000
1!
1'
1/
#891380000000
0!
0'
0/
#891390000000
#891400000000
1!
1'
1/
#891410000000
0!
0'
0/
#891420000000
1!
1'
1/
#891430000000
0!
1"
0'
1(
0/
10
#891440000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#891450000000
0!
0'
0/
#891460000000
1!
1'
1/
#891470000000
0!
0'
0/
#891480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#891490000000
0!
0'
0/
#891500000000
1!
1'
1/
#891510000000
0!
1"
0'
1(
0/
10
#891520000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#891530000000
0!
1$
0'
1+
0/
#891540000000
1!
1'
1/
#891550000000
0!
0'
0/
#891560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#891570000000
0!
0'
0/
#891580000000
1!
1'
1/
#891590000000
0!
0'
0/
#891600000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#891610000000
0!
0'
0/
#891620000000
1!
1'
1/
#891630000000
0!
0'
0/
#891640000000
1!
1'
1/
#891650000000
0!
0'
0/
#891660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#891670000000
0!
0'
0/
#891680000000
1!
1'
1/
#891690000000
0!
0'
0/
#891700000000
1!
1'
1/
#891710000000
0!
0'
0/
#891720000000
1!
1'
1/
#891730000000
0!
0'
0/
#891740000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#891750000000
0!
0'
0/
#891760000000
1!
1'
1/
#891770000000
0!
0'
0/
#891780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#891790000000
0!
0'
0/
#891800000000
1!
1'
1/
#891810000000
0!
0'
0/
#891820000000
#891830000000
1!
1'
1/
#891840000000
0!
0'
0/
#891850000000
1!
1'
1/
#891860000000
0!
1"
0'
1(
0/
10
#891870000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#891880000000
0!
0'
0/
#891890000000
1!
1'
1/
#891900000000
0!
0'
0/
#891910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#891920000000
0!
0'
0/
#891930000000
1!
1'
1/
#891940000000
0!
1"
0'
1(
0/
10
#891950000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#891960000000
0!
1$
0'
1+
0/
#891970000000
1!
1'
1/
#891980000000
0!
0'
0/
#891990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#892000000000
0!
0'
0/
#892010000000
1!
1'
1/
#892020000000
0!
0'
0/
#892030000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#892040000000
0!
0'
0/
#892050000000
1!
1'
1/
#892060000000
0!
0'
0/
#892070000000
1!
1'
1/
#892080000000
0!
0'
0/
#892090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#892100000000
0!
0'
0/
#892110000000
1!
1'
1/
#892120000000
0!
0'
0/
#892130000000
1!
1'
1/
#892140000000
0!
0'
0/
#892150000000
1!
1'
1/
#892160000000
0!
0'
0/
#892170000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#892180000000
0!
0'
0/
#892190000000
1!
1'
1/
#892200000000
0!
0'
0/
#892210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#892220000000
0!
0'
0/
#892230000000
1!
1'
1/
#892240000000
0!
0'
0/
#892250000000
#892260000000
1!
1'
1/
#892270000000
0!
0'
0/
#892280000000
1!
1'
1/
#892290000000
0!
1"
0'
1(
0/
10
#892300000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#892310000000
0!
0'
0/
#892320000000
1!
1'
1/
#892330000000
0!
0'
0/
#892340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#892350000000
0!
0'
0/
#892360000000
1!
1'
1/
#892370000000
0!
1"
0'
1(
0/
10
#892380000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#892390000000
0!
1$
0'
1+
0/
#892400000000
1!
1'
1/
#892410000000
0!
0'
0/
#892420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#892430000000
0!
0'
0/
#892440000000
1!
1'
1/
#892450000000
0!
0'
0/
#892460000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#892470000000
0!
0'
0/
#892480000000
1!
1'
1/
#892490000000
0!
0'
0/
#892500000000
1!
1'
1/
#892510000000
0!
0'
0/
#892520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#892530000000
0!
0'
0/
#892540000000
1!
1'
1/
#892550000000
0!
0'
0/
#892560000000
1!
1'
1/
#892570000000
0!
0'
0/
#892580000000
1!
1'
1/
#892590000000
0!
0'
0/
#892600000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#892610000000
0!
0'
0/
#892620000000
1!
1'
1/
#892630000000
0!
0'
0/
#892640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#892650000000
0!
0'
0/
#892660000000
1!
1'
1/
#892670000000
0!
0'
0/
#892680000000
#892690000000
1!
1'
1/
#892700000000
0!
0'
0/
#892710000000
1!
1'
1/
#892720000000
0!
1"
0'
1(
0/
10
#892730000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#892740000000
0!
0'
0/
#892750000000
1!
1'
1/
#892760000000
0!
0'
0/
#892770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#892780000000
0!
0'
0/
#892790000000
1!
1'
1/
#892800000000
0!
1"
0'
1(
0/
10
#892810000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#892820000000
0!
1$
0'
1+
0/
#892830000000
1!
1'
1/
#892840000000
0!
0'
0/
#892850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#892860000000
0!
0'
0/
#892870000000
1!
1'
1/
#892880000000
0!
0'
0/
#892890000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#892900000000
0!
0'
0/
#892910000000
1!
1'
1/
#892920000000
0!
0'
0/
#892930000000
1!
1'
1/
#892940000000
0!
0'
0/
#892950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#892960000000
0!
0'
0/
#892970000000
1!
1'
1/
#892980000000
0!
0'
0/
#892990000000
1!
1'
1/
#893000000000
0!
0'
0/
#893010000000
1!
1'
1/
#893020000000
0!
0'
0/
#893030000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#893040000000
0!
0'
0/
#893050000000
1!
1'
1/
#893060000000
0!
0'
0/
#893070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#893080000000
0!
0'
0/
#893090000000
1!
1'
1/
#893100000000
0!
0'
0/
#893110000000
#893120000000
1!
1'
1/
#893130000000
0!
0'
0/
#893140000000
1!
1'
1/
#893150000000
0!
1"
0'
1(
0/
10
#893160000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#893170000000
0!
0'
0/
#893180000000
1!
1'
1/
#893190000000
0!
0'
0/
#893200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#893210000000
0!
0'
0/
#893220000000
1!
1'
1/
#893230000000
0!
1"
0'
1(
0/
10
#893240000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#893250000000
0!
1$
0'
1+
0/
#893260000000
1!
1'
1/
#893270000000
0!
0'
0/
#893280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#893290000000
0!
0'
0/
#893300000000
1!
1'
1/
#893310000000
0!
0'
0/
#893320000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#893330000000
0!
0'
0/
#893340000000
1!
1'
1/
#893350000000
0!
0'
0/
#893360000000
1!
1'
1/
#893370000000
0!
0'
0/
#893380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#893390000000
0!
0'
0/
#893400000000
1!
1'
1/
#893410000000
0!
0'
0/
#893420000000
1!
1'
1/
#893430000000
0!
0'
0/
#893440000000
1!
1'
1/
#893450000000
0!
0'
0/
#893460000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#893470000000
0!
0'
0/
#893480000000
1!
1'
1/
#893490000000
0!
0'
0/
#893500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#893510000000
0!
0'
0/
#893520000000
1!
1'
1/
#893530000000
0!
0'
0/
#893540000000
#893550000000
1!
1'
1/
#893560000000
0!
0'
0/
#893570000000
1!
1'
1/
#893580000000
0!
1"
0'
1(
0/
10
#893590000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#893600000000
0!
0'
0/
#893610000000
1!
1'
1/
#893620000000
0!
0'
0/
#893630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#893640000000
0!
0'
0/
#893650000000
1!
1'
1/
#893660000000
0!
1"
0'
1(
0/
10
#893670000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#893680000000
0!
1$
0'
1+
0/
#893690000000
1!
1'
1/
#893700000000
0!
0'
0/
#893710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#893720000000
0!
0'
0/
#893730000000
1!
1'
1/
#893740000000
0!
0'
0/
#893750000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#893760000000
0!
0'
0/
#893770000000
1!
1'
1/
#893780000000
0!
0'
0/
#893790000000
1!
1'
1/
#893800000000
0!
0'
0/
#893810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#893820000000
0!
0'
0/
#893830000000
1!
1'
1/
#893840000000
0!
0'
0/
#893850000000
1!
1'
1/
#893860000000
0!
0'
0/
#893870000000
1!
1'
1/
#893880000000
0!
0'
0/
#893890000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#893900000000
0!
0'
0/
#893910000000
1!
1'
1/
#893920000000
0!
0'
0/
#893930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#893940000000
0!
0'
0/
#893950000000
1!
1'
1/
#893960000000
0!
0'
0/
#893970000000
#893980000000
1!
1'
1/
#893990000000
0!
0'
0/
#894000000000
1!
1'
1/
#894010000000
0!
1"
0'
1(
0/
10
#894020000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#894030000000
0!
0'
0/
#894040000000
1!
1'
1/
#894050000000
0!
0'
0/
#894060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#894070000000
0!
0'
0/
#894080000000
1!
1'
1/
#894090000000
0!
1"
0'
1(
0/
10
#894100000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#894110000000
0!
1$
0'
1+
0/
#894120000000
1!
1'
1/
#894130000000
0!
0'
0/
#894140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#894150000000
0!
0'
0/
#894160000000
1!
1'
1/
#894170000000
0!
0'
0/
#894180000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#894190000000
0!
0'
0/
#894200000000
1!
1'
1/
#894210000000
0!
0'
0/
#894220000000
1!
1'
1/
#894230000000
0!
0'
0/
#894240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#894250000000
0!
0'
0/
#894260000000
1!
1'
1/
#894270000000
0!
0'
0/
#894280000000
1!
1'
1/
#894290000000
0!
0'
0/
#894300000000
1!
1'
1/
#894310000000
0!
0'
0/
#894320000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#894330000000
0!
0'
0/
#894340000000
1!
1'
1/
#894350000000
0!
0'
0/
#894360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#894370000000
0!
0'
0/
#894380000000
1!
1'
1/
#894390000000
0!
0'
0/
#894400000000
#894410000000
1!
1'
1/
#894420000000
0!
0'
0/
#894430000000
1!
1'
1/
#894440000000
0!
1"
0'
1(
0/
10
#894450000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#894460000000
0!
0'
0/
#894470000000
1!
1'
1/
#894480000000
0!
0'
0/
#894490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#894500000000
0!
0'
0/
#894510000000
1!
1'
1/
#894520000000
0!
1"
0'
1(
0/
10
#894530000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#894540000000
0!
1$
0'
1+
0/
#894550000000
1!
1'
1/
#894560000000
0!
0'
0/
#894570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#894580000000
0!
0'
0/
#894590000000
1!
1'
1/
#894600000000
0!
0'
0/
#894610000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#894620000000
0!
0'
0/
#894630000000
1!
1'
1/
#894640000000
0!
0'
0/
#894650000000
1!
1'
1/
#894660000000
0!
0'
0/
#894670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#894680000000
0!
0'
0/
#894690000000
1!
1'
1/
#894700000000
0!
0'
0/
#894710000000
1!
1'
1/
#894720000000
0!
0'
0/
#894730000000
1!
1'
1/
#894740000000
0!
0'
0/
#894750000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#894760000000
0!
0'
0/
#894770000000
1!
1'
1/
#894780000000
0!
0'
0/
#894790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#894800000000
0!
0'
0/
#894810000000
1!
1'
1/
#894820000000
0!
0'
0/
#894830000000
#894840000000
1!
1'
1/
#894850000000
0!
0'
0/
#894860000000
1!
1'
1/
#894870000000
0!
1"
0'
1(
0/
10
#894880000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#894890000000
0!
0'
0/
#894900000000
1!
1'
1/
#894910000000
0!
0'
0/
#894920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#894930000000
0!
0'
0/
#894940000000
1!
1'
1/
#894950000000
0!
1"
0'
1(
0/
10
#894960000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#894970000000
0!
1$
0'
1+
0/
#894980000000
1!
1'
1/
#894990000000
0!
0'
0/
#895000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#895010000000
0!
0'
0/
#895020000000
1!
1'
1/
#895030000000
0!
0'
0/
#895040000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#895050000000
0!
0'
0/
#895060000000
1!
1'
1/
#895070000000
0!
0'
0/
#895080000000
1!
1'
1/
#895090000000
0!
0'
0/
#895100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#895110000000
0!
0'
0/
#895120000000
1!
1'
1/
#895130000000
0!
0'
0/
#895140000000
1!
1'
1/
#895150000000
0!
0'
0/
#895160000000
1!
1'
1/
#895170000000
0!
0'
0/
#895180000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#895190000000
0!
0'
0/
#895200000000
1!
1'
1/
#895210000000
0!
0'
0/
#895220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#895230000000
0!
0'
0/
#895240000000
1!
1'
1/
#895250000000
0!
0'
0/
#895260000000
#895270000000
1!
1'
1/
#895280000000
0!
0'
0/
#895290000000
1!
1'
1/
#895300000000
0!
1"
0'
1(
0/
10
#895310000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#895320000000
0!
0'
0/
#895330000000
1!
1'
1/
#895340000000
0!
0'
0/
#895350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#895360000000
0!
0'
0/
#895370000000
1!
1'
1/
#895380000000
0!
1"
0'
1(
0/
10
#895390000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#895400000000
0!
1$
0'
1+
0/
#895410000000
1!
1'
1/
#895420000000
0!
0'
0/
#895430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#895440000000
0!
0'
0/
#895450000000
1!
1'
1/
#895460000000
0!
0'
0/
#895470000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#895480000000
0!
0'
0/
#895490000000
1!
1'
1/
#895500000000
0!
0'
0/
#895510000000
1!
1'
1/
#895520000000
0!
0'
0/
#895530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#895540000000
0!
0'
0/
#895550000000
1!
1'
1/
#895560000000
0!
0'
0/
#895570000000
1!
1'
1/
#895580000000
0!
0'
0/
#895590000000
1!
1'
1/
#895600000000
0!
0'
0/
#895610000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#895620000000
0!
0'
0/
#895630000000
1!
1'
1/
#895640000000
0!
0'
0/
#895650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#895660000000
0!
0'
0/
#895670000000
1!
1'
1/
#895680000000
0!
0'
0/
#895690000000
#895700000000
1!
1'
1/
#895710000000
0!
0'
0/
#895720000000
1!
1'
1/
#895730000000
0!
1"
0'
1(
0/
10
#895740000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#895750000000
0!
0'
0/
#895760000000
1!
1'
1/
#895770000000
0!
0'
0/
#895780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#895790000000
0!
0'
0/
#895800000000
1!
1'
1/
#895810000000
0!
1"
0'
1(
0/
10
#895820000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#895830000000
0!
1$
0'
1+
0/
#895840000000
1!
1'
1/
#895850000000
0!
0'
0/
#895860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#895870000000
0!
0'
0/
#895880000000
1!
1'
1/
#895890000000
0!
0'
0/
#895900000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#895910000000
0!
0'
0/
#895920000000
1!
1'
1/
#895930000000
0!
0'
0/
#895940000000
1!
1'
1/
#895950000000
0!
0'
0/
#895960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#895970000000
0!
0'
0/
#895980000000
1!
1'
1/
#895990000000
0!
0'
0/
#896000000000
1!
1'
1/
#896010000000
0!
0'
0/
#896020000000
1!
1'
1/
#896030000000
0!
0'
0/
#896040000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#896050000000
0!
0'
0/
#896060000000
1!
1'
1/
#896070000000
0!
0'
0/
#896080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#896090000000
0!
0'
0/
#896100000000
1!
1'
1/
#896110000000
0!
0'
0/
#896120000000
#896130000000
1!
1'
1/
#896140000000
0!
0'
0/
#896150000000
1!
1'
1/
#896160000000
0!
1"
0'
1(
0/
10
#896170000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#896180000000
0!
0'
0/
#896190000000
1!
1'
1/
#896200000000
0!
0'
0/
#896210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#896220000000
0!
0'
0/
#896230000000
1!
1'
1/
#896240000000
0!
1"
0'
1(
0/
10
#896250000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#896260000000
0!
1$
0'
1+
0/
#896270000000
1!
1'
1/
#896280000000
0!
0'
0/
#896290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#896300000000
0!
0'
0/
#896310000000
1!
1'
1/
#896320000000
0!
0'
0/
#896330000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#896340000000
0!
0'
0/
#896350000000
1!
1'
1/
#896360000000
0!
0'
0/
#896370000000
1!
1'
1/
#896380000000
0!
0'
0/
#896390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#896400000000
0!
0'
0/
#896410000000
1!
1'
1/
#896420000000
0!
0'
0/
#896430000000
1!
1'
1/
#896440000000
0!
0'
0/
#896450000000
1!
1'
1/
#896460000000
0!
0'
0/
#896470000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#896480000000
0!
0'
0/
#896490000000
1!
1'
1/
#896500000000
0!
0'
0/
#896510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#896520000000
0!
0'
0/
#896530000000
1!
1'
1/
#896540000000
0!
0'
0/
#896550000000
#896560000000
1!
1'
1/
#896570000000
0!
0'
0/
#896580000000
1!
1'
1/
#896590000000
0!
1"
0'
1(
0/
10
#896600000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#896610000000
0!
0'
0/
#896620000000
1!
1'
1/
#896630000000
0!
0'
0/
#896640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#896650000000
0!
0'
0/
#896660000000
1!
1'
1/
#896670000000
0!
1"
0'
1(
0/
10
#896680000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#896690000000
0!
1$
0'
1+
0/
#896700000000
1!
1'
1/
#896710000000
0!
0'
0/
#896720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#896730000000
0!
0'
0/
#896740000000
1!
1'
1/
#896750000000
0!
0'
0/
#896760000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#896770000000
0!
0'
0/
#896780000000
1!
1'
1/
#896790000000
0!
0'
0/
#896800000000
1!
1'
1/
#896810000000
0!
0'
0/
#896820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#896830000000
0!
0'
0/
#896840000000
1!
1'
1/
#896850000000
0!
0'
0/
#896860000000
1!
1'
1/
#896870000000
0!
0'
0/
#896880000000
1!
1'
1/
#896890000000
0!
0'
0/
#896900000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#896910000000
0!
0'
0/
#896920000000
1!
1'
1/
#896930000000
0!
0'
0/
#896940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#896950000000
0!
0'
0/
#896960000000
1!
1'
1/
#896970000000
0!
0'
0/
#896980000000
#896990000000
1!
1'
1/
#897000000000
0!
0'
0/
#897010000000
1!
1'
1/
#897020000000
0!
1"
0'
1(
0/
10
#897030000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#897040000000
0!
0'
0/
#897050000000
1!
1'
1/
#897060000000
0!
0'
0/
#897070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#897080000000
0!
0'
0/
#897090000000
1!
1'
1/
#897100000000
0!
1"
0'
1(
0/
10
#897110000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#897120000000
0!
1$
0'
1+
0/
#897130000000
1!
1'
1/
#897140000000
0!
0'
0/
#897150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#897160000000
0!
0'
0/
#897170000000
1!
1'
1/
#897180000000
0!
0'
0/
#897190000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#897200000000
0!
0'
0/
#897210000000
1!
1'
1/
#897220000000
0!
0'
0/
#897230000000
1!
1'
1/
#897240000000
0!
0'
0/
#897250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#897260000000
0!
0'
0/
#897270000000
1!
1'
1/
#897280000000
0!
0'
0/
#897290000000
1!
1'
1/
#897300000000
0!
0'
0/
#897310000000
1!
1'
1/
#897320000000
0!
0'
0/
#897330000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#897340000000
0!
0'
0/
#897350000000
1!
1'
1/
#897360000000
0!
0'
0/
#897370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#897380000000
0!
0'
0/
#897390000000
1!
1'
1/
#897400000000
0!
0'
0/
#897410000000
#897420000000
1!
1'
1/
#897430000000
0!
0'
0/
#897440000000
1!
1'
1/
#897450000000
0!
1"
0'
1(
0/
10
#897460000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#897470000000
0!
0'
0/
#897480000000
1!
1'
1/
#897490000000
0!
0'
0/
#897500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#897510000000
0!
0'
0/
#897520000000
1!
1'
1/
#897530000000
0!
1"
0'
1(
0/
10
#897540000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#897550000000
0!
1$
0'
1+
0/
#897560000000
1!
1'
1/
#897570000000
0!
0'
0/
#897580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#897590000000
0!
0'
0/
#897600000000
1!
1'
1/
#897610000000
0!
0'
0/
#897620000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#897630000000
0!
0'
0/
#897640000000
1!
1'
1/
#897650000000
0!
0'
0/
#897660000000
1!
1'
1/
#897670000000
0!
0'
0/
#897680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#897690000000
0!
0'
0/
#897700000000
1!
1'
1/
#897710000000
0!
0'
0/
#897720000000
1!
1'
1/
#897730000000
0!
0'
0/
#897740000000
1!
1'
1/
#897750000000
0!
0'
0/
#897760000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#897770000000
0!
0'
0/
#897780000000
1!
1'
1/
#897790000000
0!
0'
0/
#897800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#897810000000
0!
0'
0/
#897820000000
1!
1'
1/
#897830000000
0!
0'
0/
#897840000000
#897850000000
1!
1'
1/
#897860000000
0!
0'
0/
#897870000000
1!
1'
1/
#897880000000
0!
1"
0'
1(
0/
10
#897890000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#897900000000
0!
0'
0/
#897910000000
1!
1'
1/
#897920000000
0!
0'
0/
#897930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#897940000000
0!
0'
0/
#897950000000
1!
1'
1/
#897960000000
0!
1"
0'
1(
0/
10
#897970000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#897980000000
0!
1$
0'
1+
0/
#897990000000
1!
1'
1/
#898000000000
0!
0'
0/
#898010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#898020000000
0!
0'
0/
#898030000000
1!
1'
1/
#898040000000
0!
0'
0/
#898050000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#898060000000
0!
0'
0/
#898070000000
1!
1'
1/
#898080000000
0!
0'
0/
#898090000000
1!
1'
1/
#898100000000
0!
0'
0/
#898110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#898120000000
0!
0'
0/
#898130000000
1!
1'
1/
#898140000000
0!
0'
0/
#898150000000
1!
1'
1/
#898160000000
0!
0'
0/
#898170000000
1!
1'
1/
#898180000000
0!
0'
0/
#898190000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#898200000000
0!
0'
0/
#898210000000
1!
1'
1/
#898220000000
0!
0'
0/
#898230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#898240000000
0!
0'
0/
#898250000000
1!
1'
1/
#898260000000
0!
0'
0/
#898270000000
#898280000000
1!
1'
1/
#898290000000
0!
0'
0/
#898300000000
1!
1'
1/
#898310000000
0!
1"
0'
1(
0/
10
#898320000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#898330000000
0!
0'
0/
#898340000000
1!
1'
1/
#898350000000
0!
0'
0/
#898360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#898370000000
0!
0'
0/
#898380000000
1!
1'
1/
#898390000000
0!
1"
0'
1(
0/
10
#898400000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#898410000000
0!
1$
0'
1+
0/
#898420000000
1!
1'
1/
#898430000000
0!
0'
0/
#898440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#898450000000
0!
0'
0/
#898460000000
1!
1'
1/
#898470000000
0!
0'
0/
#898480000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#898490000000
0!
0'
0/
#898500000000
1!
1'
1/
#898510000000
0!
0'
0/
#898520000000
1!
1'
1/
#898530000000
0!
0'
0/
#898540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#898550000000
0!
0'
0/
#898560000000
1!
1'
1/
#898570000000
0!
0'
0/
#898580000000
1!
1'
1/
#898590000000
0!
0'
0/
#898600000000
1!
1'
1/
#898610000000
0!
0'
0/
#898620000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#898630000000
0!
0'
0/
#898640000000
1!
1'
1/
#898650000000
0!
0'
0/
#898660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#898670000000
0!
0'
0/
#898680000000
1!
1'
1/
#898690000000
0!
0'
0/
#898700000000
#898710000000
1!
1'
1/
#898720000000
0!
0'
0/
#898730000000
1!
1'
1/
#898740000000
0!
1"
0'
1(
0/
10
#898750000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#898760000000
0!
0'
0/
#898770000000
1!
1'
1/
#898780000000
0!
0'
0/
#898790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#898800000000
0!
0'
0/
#898810000000
1!
1'
1/
#898820000000
0!
1"
0'
1(
0/
10
#898830000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#898840000000
0!
1$
0'
1+
0/
#898850000000
1!
1'
1/
#898860000000
0!
0'
0/
#898870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#898880000000
0!
0'
0/
#898890000000
1!
1'
1/
#898900000000
0!
0'
0/
#898910000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#898920000000
0!
0'
0/
#898930000000
1!
1'
1/
#898940000000
0!
0'
0/
#898950000000
1!
1'
1/
#898960000000
0!
0'
0/
#898970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#898980000000
0!
0'
0/
#898990000000
1!
1'
1/
#899000000000
0!
0'
0/
#899010000000
1!
1'
1/
#899020000000
0!
0'
0/
#899030000000
1!
1'
1/
#899040000000
0!
0'
0/
#899050000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#899060000000
0!
0'
0/
#899070000000
1!
1'
1/
#899080000000
0!
0'
0/
#899090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#899100000000
0!
0'
0/
#899110000000
1!
1'
1/
#899120000000
0!
0'
0/
#899130000000
#899140000000
1!
1'
1/
#899150000000
0!
0'
0/
#899160000000
1!
1'
1/
#899170000000
0!
1"
0'
1(
0/
10
#899180000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#899190000000
0!
0'
0/
#899200000000
1!
1'
1/
#899210000000
0!
0'
0/
#899220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#899230000000
0!
0'
0/
#899240000000
1!
1'
1/
#899250000000
0!
1"
0'
1(
0/
10
#899260000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#899270000000
0!
1$
0'
1+
0/
#899280000000
1!
1'
1/
#899290000000
0!
0'
0/
#899300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#899310000000
0!
0'
0/
#899320000000
1!
1'
1/
#899330000000
0!
0'
0/
#899340000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#899350000000
0!
0'
0/
#899360000000
1!
1'
1/
#899370000000
0!
0'
0/
#899380000000
1!
1'
1/
#899390000000
0!
0'
0/
#899400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#899410000000
0!
0'
0/
#899420000000
1!
1'
1/
#899430000000
0!
0'
0/
#899440000000
1!
1'
1/
#899450000000
0!
0'
0/
#899460000000
1!
1'
1/
#899470000000
0!
0'
0/
#899480000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#899490000000
0!
0'
0/
#899500000000
1!
1'
1/
#899510000000
0!
0'
0/
#899520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#899530000000
0!
0'
0/
#899540000000
1!
1'
1/
#899550000000
0!
0'
0/
#899560000000
#899570000000
1!
1'
1/
#899580000000
0!
0'
0/
#899590000000
1!
1'
1/
#899600000000
0!
1"
0'
1(
0/
10
#899610000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#899620000000
0!
0'
0/
#899630000000
1!
1'
1/
#899640000000
0!
0'
0/
#899650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#899660000000
0!
0'
0/
#899670000000
1!
1'
1/
#899680000000
0!
1"
0'
1(
0/
10
#899690000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#899700000000
0!
1$
0'
1+
0/
#899710000000
1!
1'
1/
#899720000000
0!
0'
0/
#899730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#899740000000
0!
0'
0/
#899750000000
1!
1'
1/
#899760000000
0!
0'
0/
#899770000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#899780000000
0!
0'
0/
#899790000000
1!
1'
1/
#899800000000
0!
0'
0/
#899810000000
1!
1'
1/
#899820000000
0!
0'
0/
#899830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#899840000000
0!
0'
0/
#899850000000
1!
1'
1/
#899860000000
0!
0'
0/
#899870000000
1!
1'
1/
#899880000000
0!
0'
0/
#899890000000
1!
1'
1/
#899900000000
0!
0'
0/
#899910000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#899920000000
0!
0'
0/
#899930000000
1!
1'
1/
#899940000000
0!
0'
0/
#899950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#899960000000
0!
0'
0/
#899970000000
1!
1'
1/
#899980000000
0!
0'
0/
#899990000000
#900000000000
1!
1'
1/
#900010000000
0!
0'
0/
#900020000000
1!
1'
1/
#900030000000
0!
1"
0'
1(
0/
10
#900040000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#900050000000
0!
0'
0/
#900060000000
1!
1'
1/
#900070000000
0!
0'
0/
#900080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#900090000000
0!
0'
0/
#900100000000
1!
1'
1/
#900110000000
0!
1"
0'
1(
0/
10
#900120000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#900130000000
0!
1$
0'
1+
0/
#900140000000
1!
1'
1/
#900150000000
0!
0'
0/
#900160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#900170000000
0!
0'
0/
#900180000000
1!
1'
1/
#900190000000
0!
0'
0/
#900200000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#900210000000
0!
0'
0/
#900220000000
1!
1'
1/
#900230000000
0!
0'
0/
#900240000000
1!
1'
1/
#900250000000
0!
0'
0/
#900260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#900270000000
0!
0'
0/
#900280000000
1!
1'
1/
#900290000000
0!
0'
0/
#900300000000
1!
1'
1/
#900310000000
0!
0'
0/
#900320000000
1!
1'
1/
#900330000000
0!
0'
0/
#900340000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#900350000000
0!
0'
0/
#900360000000
1!
1'
1/
#900370000000
0!
0'
0/
#900380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#900390000000
0!
0'
0/
#900400000000
1!
1'
1/
#900410000000
0!
0'
0/
#900420000000
#900430000000
1!
1'
1/
#900440000000
0!
0'
0/
#900450000000
1!
1'
1/
#900460000000
0!
1"
0'
1(
0/
10
#900470000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#900480000000
0!
0'
0/
#900490000000
1!
1'
1/
#900500000000
0!
0'
0/
#900510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#900520000000
0!
0'
0/
#900530000000
1!
1'
1/
#900540000000
0!
1"
0'
1(
0/
10
#900550000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#900560000000
0!
1$
0'
1+
0/
#900570000000
1!
1'
1/
#900580000000
0!
0'
0/
#900590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#900600000000
0!
0'
0/
#900610000000
1!
1'
1/
#900620000000
0!
0'
0/
#900630000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#900640000000
0!
0'
0/
#900650000000
1!
1'
1/
#900660000000
0!
0'
0/
#900670000000
1!
1'
1/
#900680000000
0!
0'
0/
#900690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#900700000000
0!
0'
0/
#900710000000
1!
1'
1/
#900720000000
0!
0'
0/
#900730000000
1!
1'
1/
#900740000000
0!
0'
0/
#900750000000
1!
1'
1/
#900760000000
0!
0'
0/
#900770000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#900780000000
0!
0'
0/
#900790000000
1!
1'
1/
#900800000000
0!
0'
0/
#900810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#900820000000
0!
0'
0/
#900830000000
1!
1'
1/
#900840000000
0!
0'
0/
#900850000000
#900860000000
1!
1'
1/
#900870000000
0!
0'
0/
#900880000000
1!
1'
1/
#900890000000
0!
1"
0'
1(
0/
10
#900900000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#900910000000
0!
0'
0/
#900920000000
1!
1'
1/
#900930000000
0!
0'
0/
#900940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#900950000000
0!
0'
0/
#900960000000
1!
1'
1/
#900970000000
0!
1"
0'
1(
0/
10
#900980000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#900990000000
0!
1$
0'
1+
0/
#901000000000
1!
1'
1/
#901010000000
0!
0'
0/
#901020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#901030000000
0!
0'
0/
#901040000000
1!
1'
1/
#901050000000
0!
0'
0/
#901060000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#901070000000
0!
0'
0/
#901080000000
1!
1'
1/
#901090000000
0!
0'
0/
#901100000000
1!
1'
1/
#901110000000
0!
0'
0/
#901120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#901130000000
0!
0'
0/
#901140000000
1!
1'
1/
#901150000000
0!
0'
0/
#901160000000
1!
1'
1/
#901170000000
0!
0'
0/
#901180000000
1!
1'
1/
#901190000000
0!
0'
0/
#901200000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#901210000000
0!
0'
0/
#901220000000
1!
1'
1/
#901230000000
0!
0'
0/
#901240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#901250000000
0!
0'
0/
#901260000000
1!
1'
1/
#901270000000
0!
0'
0/
#901280000000
#901290000000
1!
1'
1/
#901300000000
0!
0'
0/
#901310000000
1!
1'
1/
#901320000000
0!
1"
0'
1(
0/
10
#901330000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#901340000000
0!
0'
0/
#901350000000
1!
1'
1/
#901360000000
0!
0'
0/
#901370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#901380000000
0!
0'
0/
#901390000000
1!
1'
1/
#901400000000
0!
1"
0'
1(
0/
10
#901410000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#901420000000
0!
1$
0'
1+
0/
#901430000000
1!
1'
1/
#901440000000
0!
0'
0/
#901450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#901460000000
0!
0'
0/
#901470000000
1!
1'
1/
#901480000000
0!
0'
0/
#901490000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#901500000000
0!
0'
0/
#901510000000
1!
1'
1/
#901520000000
0!
0'
0/
#901530000000
1!
1'
1/
#901540000000
0!
0'
0/
#901550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#901560000000
0!
0'
0/
#901570000000
1!
1'
1/
#901580000000
0!
0'
0/
#901590000000
1!
1'
1/
#901600000000
0!
0'
0/
#901610000000
1!
1'
1/
#901620000000
0!
0'
0/
#901630000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#901640000000
0!
0'
0/
#901650000000
1!
1'
1/
#901660000000
0!
0'
0/
#901670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#901680000000
0!
0'
0/
#901690000000
1!
1'
1/
#901700000000
0!
0'
0/
#901710000000
#901720000000
1!
1'
1/
#901730000000
0!
0'
0/
#901740000000
1!
1'
1/
#901750000000
0!
1"
0'
1(
0/
10
#901760000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#901770000000
0!
0'
0/
#901780000000
1!
1'
1/
#901790000000
0!
0'
0/
#901800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#901810000000
0!
0'
0/
#901820000000
1!
1'
1/
#901830000000
0!
1"
0'
1(
0/
10
#901840000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#901850000000
0!
1$
0'
1+
0/
#901860000000
1!
1'
1/
#901870000000
0!
0'
0/
#901880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#901890000000
0!
0'
0/
#901900000000
1!
1'
1/
#901910000000
0!
0'
0/
#901920000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#901930000000
0!
0'
0/
#901940000000
1!
1'
1/
#901950000000
0!
0'
0/
#901960000000
1!
1'
1/
#901970000000
0!
0'
0/
#901980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#901990000000
0!
0'
0/
#902000000000
1!
1'
1/
#902010000000
0!
0'
0/
#902020000000
1!
1'
1/
#902030000000
0!
0'
0/
#902040000000
1!
1'
1/
#902050000000
0!
0'
0/
#902060000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#902070000000
0!
0'
0/
#902080000000
1!
1'
1/
#902090000000
0!
0'
0/
#902100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#902110000000
0!
0'
0/
#902120000000
1!
1'
1/
#902130000000
0!
0'
0/
#902140000000
#902150000000
1!
1'
1/
#902160000000
0!
0'
0/
#902170000000
1!
1'
1/
#902180000000
0!
1"
0'
1(
0/
10
#902190000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#902200000000
0!
0'
0/
#902210000000
1!
1'
1/
#902220000000
0!
0'
0/
#902230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#902240000000
0!
0'
0/
#902250000000
1!
1'
1/
#902260000000
0!
1"
0'
1(
0/
10
#902270000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#902280000000
0!
1$
0'
1+
0/
#902290000000
1!
1'
1/
#902300000000
0!
0'
0/
#902310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#902320000000
0!
0'
0/
#902330000000
1!
1'
1/
#902340000000
0!
0'
0/
#902350000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#902360000000
0!
0'
0/
#902370000000
1!
1'
1/
#902380000000
0!
0'
0/
#902390000000
1!
1'
1/
#902400000000
0!
0'
0/
#902410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#902420000000
0!
0'
0/
#902430000000
1!
1'
1/
#902440000000
0!
0'
0/
#902450000000
1!
1'
1/
#902460000000
0!
0'
0/
#902470000000
1!
1'
1/
#902480000000
0!
0'
0/
#902490000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#902500000000
0!
0'
0/
#902510000000
1!
1'
1/
#902520000000
0!
0'
0/
#902530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#902540000000
0!
0'
0/
#902550000000
1!
1'
1/
#902560000000
0!
0'
0/
#902570000000
#902580000000
1!
1'
1/
#902590000000
0!
0'
0/
#902600000000
1!
1'
1/
#902610000000
0!
1"
0'
1(
0/
10
#902620000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#902630000000
0!
0'
0/
#902640000000
1!
1'
1/
#902650000000
0!
0'
0/
#902660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#902670000000
0!
0'
0/
#902680000000
1!
1'
1/
#902690000000
0!
1"
0'
1(
0/
10
#902700000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#902710000000
0!
1$
0'
1+
0/
#902720000000
1!
1'
1/
#902730000000
0!
0'
0/
#902740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#902750000000
0!
0'
0/
#902760000000
1!
1'
1/
#902770000000
0!
0'
0/
#902780000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#902790000000
0!
0'
0/
#902800000000
1!
1'
1/
#902810000000
0!
0'
0/
#902820000000
1!
1'
1/
#902830000000
0!
0'
0/
#902840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#902850000000
0!
0'
0/
#902860000000
1!
1'
1/
#902870000000
0!
0'
0/
#902880000000
1!
1'
1/
#902890000000
0!
0'
0/
#902900000000
1!
1'
1/
#902910000000
0!
0'
0/
#902920000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#902930000000
0!
0'
0/
#902940000000
1!
1'
1/
#902950000000
0!
0'
0/
#902960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#902970000000
0!
0'
0/
#902980000000
1!
1'
1/
#902990000000
0!
0'
0/
#903000000000
#903010000000
1!
1'
1/
#903020000000
0!
0'
0/
#903030000000
1!
1'
1/
#903040000000
0!
1"
0'
1(
0/
10
#903050000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#903060000000
0!
0'
0/
#903070000000
1!
1'
1/
#903080000000
0!
0'
0/
#903090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#903100000000
0!
0'
0/
#903110000000
1!
1'
1/
#903120000000
0!
1"
0'
1(
0/
10
#903130000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#903140000000
0!
1$
0'
1+
0/
#903150000000
1!
1'
1/
#903160000000
0!
0'
0/
#903170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#903180000000
0!
0'
0/
#903190000000
1!
1'
1/
#903200000000
0!
0'
0/
#903210000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#903220000000
0!
0'
0/
#903230000000
1!
1'
1/
#903240000000
0!
0'
0/
#903250000000
1!
1'
1/
#903260000000
0!
0'
0/
#903270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#903280000000
0!
0'
0/
#903290000000
1!
1'
1/
#903300000000
0!
0'
0/
#903310000000
1!
1'
1/
#903320000000
0!
0'
0/
#903330000000
1!
1'
1/
#903340000000
0!
0'
0/
#903350000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#903360000000
0!
0'
0/
#903370000000
1!
1'
1/
#903380000000
0!
0'
0/
#903390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#903400000000
0!
0'
0/
#903410000000
1!
1'
1/
#903420000000
0!
0'
0/
#903430000000
#903440000000
1!
1'
1/
#903450000000
0!
0'
0/
#903460000000
1!
1'
1/
#903470000000
0!
1"
0'
1(
0/
10
#903480000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#903490000000
0!
0'
0/
#903500000000
1!
1'
1/
#903510000000
0!
0'
0/
#903520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#903530000000
0!
0'
0/
#903540000000
1!
1'
1/
#903550000000
0!
1"
0'
1(
0/
10
#903560000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#903570000000
0!
1$
0'
1+
0/
#903580000000
1!
1'
1/
#903590000000
0!
0'
0/
#903600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#903610000000
0!
0'
0/
#903620000000
1!
1'
1/
#903630000000
0!
0'
0/
#903640000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#903650000000
0!
0'
0/
#903660000000
1!
1'
1/
#903670000000
0!
0'
0/
#903680000000
1!
1'
1/
#903690000000
0!
0'
0/
#903700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#903710000000
0!
0'
0/
#903720000000
1!
1'
1/
#903730000000
0!
0'
0/
#903740000000
1!
1'
1/
#903750000000
0!
0'
0/
#903760000000
1!
1'
1/
#903770000000
0!
0'
0/
#903780000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#903790000000
0!
0'
0/
#903800000000
1!
1'
1/
#903810000000
0!
0'
0/
#903820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#903830000000
0!
0'
0/
#903840000000
1!
1'
1/
#903850000000
0!
0'
0/
#903860000000
#903870000000
1!
1'
1/
#903880000000
0!
0'
0/
#903890000000
1!
1'
1/
#903900000000
0!
1"
0'
1(
0/
10
#903910000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#903920000000
0!
0'
0/
#903930000000
1!
1'
1/
#903940000000
0!
0'
0/
#903950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#903960000000
0!
0'
0/
#903970000000
1!
1'
1/
#903980000000
0!
1"
0'
1(
0/
10
#903990000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#904000000000
0!
1$
0'
1+
0/
#904010000000
1!
1'
1/
#904020000000
0!
0'
0/
#904030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#904040000000
0!
0'
0/
#904050000000
1!
1'
1/
#904060000000
0!
0'
0/
#904070000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#904080000000
0!
0'
0/
#904090000000
1!
1'
1/
#904100000000
0!
0'
0/
#904110000000
1!
1'
1/
#904120000000
0!
0'
0/
#904130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#904140000000
0!
0'
0/
#904150000000
1!
1'
1/
#904160000000
0!
0'
0/
#904170000000
1!
1'
1/
#904180000000
0!
0'
0/
#904190000000
1!
1'
1/
#904200000000
0!
0'
0/
#904210000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#904220000000
0!
0'
0/
#904230000000
1!
1'
1/
#904240000000
0!
0'
0/
#904250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#904260000000
0!
0'
0/
#904270000000
1!
1'
1/
#904280000000
0!
0'
0/
#904290000000
#904300000000
1!
1'
1/
#904310000000
0!
0'
0/
#904320000000
1!
1'
1/
#904330000000
0!
1"
0'
1(
0/
10
#904340000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#904350000000
0!
0'
0/
#904360000000
1!
1'
1/
#904370000000
0!
0'
0/
#904380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#904390000000
0!
0'
0/
#904400000000
1!
1'
1/
#904410000000
0!
1"
0'
1(
0/
10
#904420000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#904430000000
0!
1$
0'
1+
0/
#904440000000
1!
1'
1/
#904450000000
0!
0'
0/
#904460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#904470000000
0!
0'
0/
#904480000000
1!
1'
1/
#904490000000
0!
0'
0/
#904500000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#904510000000
0!
0'
0/
#904520000000
1!
1'
1/
#904530000000
0!
0'
0/
#904540000000
1!
1'
1/
#904550000000
0!
0'
0/
#904560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#904570000000
0!
0'
0/
#904580000000
1!
1'
1/
#904590000000
0!
0'
0/
#904600000000
1!
1'
1/
#904610000000
0!
0'
0/
#904620000000
1!
1'
1/
#904630000000
0!
0'
0/
#904640000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#904650000000
0!
0'
0/
#904660000000
1!
1'
1/
#904670000000
0!
0'
0/
#904680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#904690000000
0!
0'
0/
#904700000000
1!
1'
1/
#904710000000
0!
0'
0/
#904720000000
#904730000000
1!
1'
1/
#904740000000
0!
0'
0/
#904750000000
1!
1'
1/
#904760000000
0!
1"
0'
1(
0/
10
#904770000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#904780000000
0!
0'
0/
#904790000000
1!
1'
1/
#904800000000
0!
0'
0/
#904810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#904820000000
0!
0'
0/
#904830000000
1!
1'
1/
#904840000000
0!
1"
0'
1(
0/
10
#904850000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#904860000000
0!
1$
0'
1+
0/
#904870000000
1!
1'
1/
#904880000000
0!
0'
0/
#904890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#904900000000
0!
0'
0/
#904910000000
1!
1'
1/
#904920000000
0!
0'
0/
#904930000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#904940000000
0!
0'
0/
#904950000000
1!
1'
1/
#904960000000
0!
0'
0/
#904970000000
1!
1'
1/
#904980000000
0!
0'
0/
#904990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#905000000000
0!
0'
0/
#905010000000
1!
1'
1/
#905020000000
0!
0'
0/
#905030000000
1!
1'
1/
#905040000000
0!
0'
0/
#905050000000
1!
1'
1/
#905060000000
0!
0'
0/
#905070000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#905080000000
0!
0'
0/
#905090000000
1!
1'
1/
#905100000000
0!
0'
0/
#905110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#905120000000
0!
0'
0/
#905130000000
1!
1'
1/
#905140000000
0!
0'
0/
#905150000000
#905160000000
1!
1'
1/
#905170000000
0!
0'
0/
#905180000000
1!
1'
1/
#905190000000
0!
1"
0'
1(
0/
10
#905200000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#905210000000
0!
0'
0/
#905220000000
1!
1'
1/
#905230000000
0!
0'
0/
#905240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#905250000000
0!
0'
0/
#905260000000
1!
1'
1/
#905270000000
0!
1"
0'
1(
0/
10
#905280000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#905290000000
0!
1$
0'
1+
0/
#905300000000
1!
1'
1/
#905310000000
0!
0'
0/
#905320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#905330000000
0!
0'
0/
#905340000000
1!
1'
1/
#905350000000
0!
0'
0/
#905360000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#905370000000
0!
0'
0/
#905380000000
1!
1'
1/
#905390000000
0!
0'
0/
#905400000000
1!
1'
1/
#905410000000
0!
0'
0/
#905420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#905430000000
0!
0'
0/
#905440000000
1!
1'
1/
#905450000000
0!
0'
0/
#905460000000
1!
1'
1/
#905470000000
0!
0'
0/
#905480000000
1!
1'
1/
#905490000000
0!
0'
0/
#905500000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#905510000000
0!
0'
0/
#905520000000
1!
1'
1/
#905530000000
0!
0'
0/
#905540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#905550000000
0!
0'
0/
#905560000000
1!
1'
1/
#905570000000
0!
0'
0/
#905580000000
#905590000000
1!
1'
1/
#905600000000
0!
0'
0/
#905610000000
1!
1'
1/
#905620000000
0!
1"
0'
1(
0/
10
#905630000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#905640000000
0!
0'
0/
#905650000000
1!
1'
1/
#905660000000
0!
0'
0/
#905670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#905680000000
0!
0'
0/
#905690000000
1!
1'
1/
#905700000000
0!
1"
0'
1(
0/
10
#905710000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#905720000000
0!
1$
0'
1+
0/
#905730000000
1!
1'
1/
#905740000000
0!
0'
0/
#905750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#905760000000
0!
0'
0/
#905770000000
1!
1'
1/
#905780000000
0!
0'
0/
#905790000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#905800000000
0!
0'
0/
#905810000000
1!
1'
1/
#905820000000
0!
0'
0/
#905830000000
1!
1'
1/
#905840000000
0!
0'
0/
#905850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#905860000000
0!
0'
0/
#905870000000
1!
1'
1/
#905880000000
0!
0'
0/
#905890000000
1!
1'
1/
#905900000000
0!
0'
0/
#905910000000
1!
1'
1/
#905920000000
0!
0'
0/
#905930000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#905940000000
0!
0'
0/
#905950000000
1!
1'
1/
#905960000000
0!
0'
0/
#905970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#905980000000
0!
0'
0/
#905990000000
1!
1'
1/
#906000000000
0!
0'
0/
#906010000000
#906020000000
1!
1'
1/
#906030000000
0!
0'
0/
#906040000000
1!
1'
1/
#906050000000
0!
1"
0'
1(
0/
10
#906060000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#906070000000
0!
0'
0/
#906080000000
1!
1'
1/
#906090000000
0!
0'
0/
#906100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#906110000000
0!
0'
0/
#906120000000
1!
1'
1/
#906130000000
0!
1"
0'
1(
0/
10
#906140000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#906150000000
0!
1$
0'
1+
0/
#906160000000
1!
1'
1/
#906170000000
0!
0'
0/
#906180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#906190000000
0!
0'
0/
#906200000000
1!
1'
1/
#906210000000
0!
0'
0/
#906220000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#906230000000
0!
0'
0/
#906240000000
1!
1'
1/
#906250000000
0!
0'
0/
#906260000000
1!
1'
1/
#906270000000
0!
0'
0/
#906280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#906290000000
0!
0'
0/
#906300000000
1!
1'
1/
#906310000000
0!
0'
0/
#906320000000
1!
1'
1/
#906330000000
0!
0'
0/
#906340000000
1!
1'
1/
#906350000000
0!
0'
0/
#906360000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#906370000000
0!
0'
0/
#906380000000
1!
1'
1/
#906390000000
0!
0'
0/
#906400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#906410000000
0!
0'
0/
#906420000000
1!
1'
1/
#906430000000
0!
0'
0/
#906440000000
#906450000000
1!
1'
1/
#906460000000
0!
0'
0/
#906470000000
1!
1'
1/
#906480000000
0!
1"
0'
1(
0/
10
#906490000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#906500000000
0!
0'
0/
#906510000000
1!
1'
1/
#906520000000
0!
0'
0/
#906530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#906540000000
0!
0'
0/
#906550000000
1!
1'
1/
#906560000000
0!
1"
0'
1(
0/
10
#906570000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#906580000000
0!
1$
0'
1+
0/
#906590000000
1!
1'
1/
#906600000000
0!
0'
0/
#906610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#906620000000
0!
0'
0/
#906630000000
1!
1'
1/
#906640000000
0!
0'
0/
#906650000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#906660000000
0!
0'
0/
#906670000000
1!
1'
1/
#906680000000
0!
0'
0/
#906690000000
1!
1'
1/
#906700000000
0!
0'
0/
#906710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#906720000000
0!
0'
0/
#906730000000
1!
1'
1/
#906740000000
0!
0'
0/
#906750000000
1!
1'
1/
#906760000000
0!
0'
0/
#906770000000
1!
1'
1/
#906780000000
0!
0'
0/
#906790000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#906800000000
0!
0'
0/
#906810000000
1!
1'
1/
#906820000000
0!
0'
0/
#906830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#906840000000
0!
0'
0/
#906850000000
1!
1'
1/
#906860000000
0!
0'
0/
#906870000000
#906880000000
1!
1'
1/
#906890000000
0!
0'
0/
#906900000000
1!
1'
1/
#906910000000
0!
1"
0'
1(
0/
10
#906920000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#906930000000
0!
0'
0/
#906940000000
1!
1'
1/
#906950000000
0!
0'
0/
#906960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#906970000000
0!
0'
0/
#906980000000
1!
1'
1/
#906990000000
0!
1"
0'
1(
0/
10
#907000000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#907010000000
0!
1$
0'
1+
0/
#907020000000
1!
1'
1/
#907030000000
0!
0'
0/
#907040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#907050000000
0!
0'
0/
#907060000000
1!
1'
1/
#907070000000
0!
0'
0/
#907080000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#907090000000
0!
0'
0/
#907100000000
1!
1'
1/
#907110000000
0!
0'
0/
#907120000000
1!
1'
1/
#907130000000
0!
0'
0/
#907140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#907150000000
0!
0'
0/
#907160000000
1!
1'
1/
#907170000000
0!
0'
0/
#907180000000
1!
1'
1/
#907190000000
0!
0'
0/
#907200000000
1!
1'
1/
#907210000000
0!
0'
0/
#907220000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#907230000000
0!
0'
0/
#907240000000
1!
1'
1/
#907250000000
0!
0'
0/
#907260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#907270000000
0!
0'
0/
#907280000000
1!
1'
1/
#907290000000
0!
0'
0/
#907300000000
#907310000000
1!
1'
1/
#907320000000
0!
0'
0/
#907330000000
1!
1'
1/
#907340000000
0!
1"
0'
1(
0/
10
#907350000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#907360000000
0!
0'
0/
#907370000000
1!
1'
1/
#907380000000
0!
0'
0/
#907390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#907400000000
0!
0'
0/
#907410000000
1!
1'
1/
#907420000000
0!
1"
0'
1(
0/
10
#907430000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#907440000000
0!
1$
0'
1+
0/
#907450000000
1!
1'
1/
#907460000000
0!
0'
0/
#907470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#907480000000
0!
0'
0/
#907490000000
1!
1'
1/
#907500000000
0!
0'
0/
#907510000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#907520000000
0!
0'
0/
#907530000000
1!
1'
1/
#907540000000
0!
0'
0/
#907550000000
1!
1'
1/
#907560000000
0!
0'
0/
#907570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#907580000000
0!
0'
0/
#907590000000
1!
1'
1/
#907600000000
0!
0'
0/
#907610000000
1!
1'
1/
#907620000000
0!
0'
0/
#907630000000
1!
1'
1/
#907640000000
0!
0'
0/
#907650000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#907660000000
0!
0'
0/
#907670000000
1!
1'
1/
#907680000000
0!
0'
0/
#907690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#907700000000
0!
0'
0/
#907710000000
1!
1'
1/
#907720000000
0!
0'
0/
#907730000000
#907740000000
1!
1'
1/
#907750000000
0!
0'
0/
#907760000000
1!
1'
1/
#907770000000
0!
1"
0'
1(
0/
10
#907780000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#907790000000
0!
0'
0/
#907800000000
1!
1'
1/
#907810000000
0!
0'
0/
#907820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#907830000000
0!
0'
0/
#907840000000
1!
1'
1/
#907850000000
0!
1"
0'
1(
0/
10
#907860000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#907870000000
0!
1$
0'
1+
0/
#907880000000
1!
1'
1/
#907890000000
0!
0'
0/
#907900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#907910000000
0!
0'
0/
#907920000000
1!
1'
1/
#907930000000
0!
0'
0/
#907940000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#907950000000
0!
0'
0/
#907960000000
1!
1'
1/
#907970000000
0!
0'
0/
#907980000000
1!
1'
1/
#907990000000
0!
0'
0/
#908000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#908010000000
0!
0'
0/
#908020000000
1!
1'
1/
#908030000000
0!
0'
0/
#908040000000
1!
1'
1/
#908050000000
0!
0'
0/
#908060000000
1!
1'
1/
#908070000000
0!
0'
0/
#908080000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#908090000000
0!
0'
0/
#908100000000
1!
1'
1/
#908110000000
0!
0'
0/
#908120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#908130000000
0!
0'
0/
#908140000000
1!
1'
1/
#908150000000
0!
0'
0/
#908160000000
#908170000000
1!
1'
1/
#908180000000
0!
0'
0/
#908190000000
1!
1'
1/
#908200000000
0!
1"
0'
1(
0/
10
#908210000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#908220000000
0!
0'
0/
#908230000000
1!
1'
1/
#908240000000
0!
0'
0/
#908250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#908260000000
0!
0'
0/
#908270000000
1!
1'
1/
#908280000000
0!
1"
0'
1(
0/
10
#908290000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#908300000000
0!
1$
0'
1+
0/
#908310000000
1!
1'
1/
#908320000000
0!
0'
0/
#908330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#908340000000
0!
0'
0/
#908350000000
1!
1'
1/
#908360000000
0!
0'
0/
#908370000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#908380000000
0!
0'
0/
#908390000000
1!
1'
1/
#908400000000
0!
0'
0/
#908410000000
1!
1'
1/
#908420000000
0!
0'
0/
#908430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#908440000000
0!
0'
0/
#908450000000
1!
1'
1/
#908460000000
0!
0'
0/
#908470000000
1!
1'
1/
#908480000000
0!
0'
0/
#908490000000
1!
1'
1/
#908500000000
0!
0'
0/
#908510000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#908520000000
0!
0'
0/
#908530000000
1!
1'
1/
#908540000000
0!
0'
0/
#908550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#908560000000
0!
0'
0/
#908570000000
1!
1'
1/
#908580000000
0!
0'
0/
#908590000000
#908600000000
1!
1'
1/
#908610000000
0!
0'
0/
#908620000000
1!
1'
1/
#908630000000
0!
1"
0'
1(
0/
10
#908640000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#908650000000
0!
0'
0/
#908660000000
1!
1'
1/
#908670000000
0!
0'
0/
#908680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#908690000000
0!
0'
0/
#908700000000
1!
1'
1/
#908710000000
0!
1"
0'
1(
0/
10
#908720000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#908730000000
0!
1$
0'
1+
0/
#908740000000
1!
1'
1/
#908750000000
0!
0'
0/
#908760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#908770000000
0!
0'
0/
#908780000000
1!
1'
1/
#908790000000
0!
0'
0/
#908800000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#908810000000
0!
0'
0/
#908820000000
1!
1'
1/
#908830000000
0!
0'
0/
#908840000000
1!
1'
1/
#908850000000
0!
0'
0/
#908860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#908870000000
0!
0'
0/
#908880000000
1!
1'
1/
#908890000000
0!
0'
0/
#908900000000
1!
1'
1/
#908910000000
0!
0'
0/
#908920000000
1!
1'
1/
#908930000000
0!
0'
0/
#908940000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#908950000000
0!
0'
0/
#908960000000
1!
1'
1/
#908970000000
0!
0'
0/
#908980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#908990000000
0!
0'
0/
#909000000000
1!
1'
1/
#909010000000
0!
0'
0/
#909020000000
#909030000000
1!
1'
1/
#909040000000
0!
0'
0/
#909050000000
1!
1'
1/
#909060000000
0!
1"
0'
1(
0/
10
#909070000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#909080000000
0!
0'
0/
#909090000000
1!
1'
1/
#909100000000
0!
0'
0/
#909110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#909120000000
0!
0'
0/
#909130000000
1!
1'
1/
#909140000000
0!
1"
0'
1(
0/
10
#909150000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#909160000000
0!
1$
0'
1+
0/
#909170000000
1!
1'
1/
#909180000000
0!
0'
0/
#909190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#909200000000
0!
0'
0/
#909210000000
1!
1'
1/
#909220000000
0!
0'
0/
#909230000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#909240000000
0!
0'
0/
#909250000000
1!
1'
1/
#909260000000
0!
0'
0/
#909270000000
1!
1'
1/
#909280000000
0!
0'
0/
#909290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#909300000000
0!
0'
0/
#909310000000
1!
1'
1/
#909320000000
0!
0'
0/
#909330000000
1!
1'
1/
#909340000000
0!
0'
0/
#909350000000
1!
1'
1/
#909360000000
0!
0'
0/
#909370000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#909380000000
0!
0'
0/
#909390000000
1!
1'
1/
#909400000000
0!
0'
0/
#909410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#909420000000
0!
0'
0/
#909430000000
1!
1'
1/
#909440000000
0!
0'
0/
#909450000000
#909460000000
1!
1'
1/
#909470000000
0!
0'
0/
#909480000000
1!
1'
1/
#909490000000
0!
1"
0'
1(
0/
10
#909500000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#909510000000
0!
0'
0/
#909520000000
1!
1'
1/
#909530000000
0!
0'
0/
#909540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#909550000000
0!
0'
0/
#909560000000
1!
1'
1/
#909570000000
0!
1"
0'
1(
0/
10
#909580000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#909590000000
0!
1$
0'
1+
0/
#909600000000
1!
1'
1/
#909610000000
0!
0'
0/
#909620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#909630000000
0!
0'
0/
#909640000000
1!
1'
1/
#909650000000
0!
0'
0/
#909660000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#909670000000
0!
0'
0/
#909680000000
1!
1'
1/
#909690000000
0!
0'
0/
#909700000000
1!
1'
1/
#909710000000
0!
0'
0/
#909720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#909730000000
0!
0'
0/
#909740000000
1!
1'
1/
#909750000000
0!
0'
0/
#909760000000
1!
1'
1/
#909770000000
0!
0'
0/
#909780000000
1!
1'
1/
#909790000000
0!
0'
0/
#909800000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#909810000000
0!
0'
0/
#909820000000
1!
1'
1/
#909830000000
0!
0'
0/
#909840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#909850000000
0!
0'
0/
#909860000000
1!
1'
1/
#909870000000
0!
0'
0/
#909880000000
#909890000000
1!
1'
1/
#909900000000
0!
0'
0/
#909910000000
1!
1'
1/
#909920000000
0!
1"
0'
1(
0/
10
#909930000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#909940000000
0!
0'
0/
#909950000000
1!
1'
1/
#909960000000
0!
0'
0/
#909970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#909980000000
0!
0'
0/
#909990000000
1!
1'
1/
#910000000000
0!
1"
0'
1(
0/
10
#910010000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#910020000000
0!
1$
0'
1+
0/
#910030000000
1!
1'
1/
#910040000000
0!
0'
0/
#910050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#910060000000
0!
0'
0/
#910070000000
1!
1'
1/
#910080000000
0!
0'
0/
#910090000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#910100000000
0!
0'
0/
#910110000000
1!
1'
1/
#910120000000
0!
0'
0/
#910130000000
1!
1'
1/
#910140000000
0!
0'
0/
#910150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#910160000000
0!
0'
0/
#910170000000
1!
1'
1/
#910180000000
0!
0'
0/
#910190000000
1!
1'
1/
#910200000000
0!
0'
0/
#910210000000
1!
1'
1/
#910220000000
0!
0'
0/
#910230000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#910240000000
0!
0'
0/
#910250000000
1!
1'
1/
#910260000000
0!
0'
0/
#910270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#910280000000
0!
0'
0/
#910290000000
1!
1'
1/
#910300000000
0!
0'
0/
#910310000000
#910320000000
1!
1'
1/
#910330000000
0!
0'
0/
#910340000000
1!
1'
1/
#910350000000
0!
1"
0'
1(
0/
10
#910360000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#910370000000
0!
0'
0/
#910380000000
1!
1'
1/
#910390000000
0!
0'
0/
#910400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#910410000000
0!
0'
0/
#910420000000
1!
1'
1/
#910430000000
0!
1"
0'
1(
0/
10
#910440000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#910450000000
0!
1$
0'
1+
0/
#910460000000
1!
1'
1/
#910470000000
0!
0'
0/
#910480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#910490000000
0!
0'
0/
#910500000000
1!
1'
1/
#910510000000
0!
0'
0/
#910520000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#910530000000
0!
0'
0/
#910540000000
1!
1'
1/
#910550000000
0!
0'
0/
#910560000000
1!
1'
1/
#910570000000
0!
0'
0/
#910580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#910590000000
0!
0'
0/
#910600000000
1!
1'
1/
#910610000000
0!
0'
0/
#910620000000
1!
1'
1/
#910630000000
0!
0'
0/
#910640000000
1!
1'
1/
#910650000000
0!
0'
0/
#910660000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#910670000000
0!
0'
0/
#910680000000
1!
1'
1/
#910690000000
0!
0'
0/
#910700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#910710000000
0!
0'
0/
#910720000000
1!
1'
1/
#910730000000
0!
0'
0/
#910740000000
#910750000000
1!
1'
1/
#910760000000
0!
0'
0/
#910770000000
1!
1'
1/
#910780000000
0!
1"
0'
1(
0/
10
#910790000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#910800000000
0!
0'
0/
#910810000000
1!
1'
1/
#910820000000
0!
0'
0/
#910830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#910840000000
0!
0'
0/
#910850000000
1!
1'
1/
#910860000000
0!
1"
0'
1(
0/
10
#910870000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#910880000000
0!
1$
0'
1+
0/
#910890000000
1!
1'
1/
#910900000000
0!
0'
0/
#910910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#910920000000
0!
0'
0/
#910930000000
1!
1'
1/
#910940000000
0!
0'
0/
#910950000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#910960000000
0!
0'
0/
#910970000000
1!
1'
1/
#910980000000
0!
0'
0/
#910990000000
1!
1'
1/
#911000000000
0!
0'
0/
#911010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#911020000000
0!
0'
0/
#911030000000
1!
1'
1/
#911040000000
0!
0'
0/
#911050000000
1!
1'
1/
#911060000000
0!
0'
0/
#911070000000
1!
1'
1/
#911080000000
0!
0'
0/
#911090000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#911100000000
0!
0'
0/
#911110000000
1!
1'
1/
#911120000000
0!
0'
0/
#911130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#911140000000
0!
0'
0/
#911150000000
1!
1'
1/
#911160000000
0!
0'
0/
#911170000000
#911180000000
1!
1'
1/
#911190000000
0!
0'
0/
#911200000000
1!
1'
1/
#911210000000
0!
1"
0'
1(
0/
10
#911220000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#911230000000
0!
0'
0/
#911240000000
1!
1'
1/
#911250000000
0!
0'
0/
#911260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#911270000000
0!
0'
0/
#911280000000
1!
1'
1/
#911290000000
0!
1"
0'
1(
0/
10
#911300000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#911310000000
0!
1$
0'
1+
0/
#911320000000
1!
1'
1/
#911330000000
0!
0'
0/
#911340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#911350000000
0!
0'
0/
#911360000000
1!
1'
1/
#911370000000
0!
0'
0/
#911380000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#911390000000
0!
0'
0/
#911400000000
1!
1'
1/
#911410000000
0!
0'
0/
#911420000000
1!
1'
1/
#911430000000
0!
0'
0/
#911440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#911450000000
0!
0'
0/
#911460000000
1!
1'
1/
#911470000000
0!
0'
0/
#911480000000
1!
1'
1/
#911490000000
0!
0'
0/
#911500000000
1!
1'
1/
#911510000000
0!
0'
0/
#911520000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#911530000000
0!
0'
0/
#911540000000
1!
1'
1/
#911550000000
0!
0'
0/
#911560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#911570000000
0!
0'
0/
#911580000000
1!
1'
1/
#911590000000
0!
0'
0/
#911600000000
#911610000000
1!
1'
1/
#911620000000
0!
0'
0/
#911630000000
1!
1'
1/
#911640000000
0!
1"
0'
1(
0/
10
#911650000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#911660000000
0!
0'
0/
#911670000000
1!
1'
1/
#911680000000
0!
0'
0/
#911690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#911700000000
0!
0'
0/
#911710000000
1!
1'
1/
#911720000000
0!
1"
0'
1(
0/
10
#911730000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#911740000000
0!
1$
0'
1+
0/
#911750000000
1!
1'
1/
#911760000000
0!
0'
0/
#911770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#911780000000
0!
0'
0/
#911790000000
1!
1'
1/
#911800000000
0!
0'
0/
#911810000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#911820000000
0!
0'
0/
#911830000000
1!
1'
1/
#911840000000
0!
0'
0/
#911850000000
1!
1'
1/
#911860000000
0!
0'
0/
#911870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#911880000000
0!
0'
0/
#911890000000
1!
1'
1/
#911900000000
0!
0'
0/
#911910000000
1!
1'
1/
#911920000000
0!
0'
0/
#911930000000
1!
1'
1/
#911940000000
0!
0'
0/
#911950000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#911960000000
0!
0'
0/
#911970000000
1!
1'
1/
#911980000000
0!
0'
0/
#911990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#912000000000
0!
0'
0/
#912010000000
1!
1'
1/
#912020000000
0!
0'
0/
#912030000000
#912040000000
1!
1'
1/
#912050000000
0!
0'
0/
#912060000000
1!
1'
1/
#912070000000
0!
1"
0'
1(
0/
10
#912080000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#912090000000
0!
0'
0/
#912100000000
1!
1'
1/
#912110000000
0!
0'
0/
#912120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#912130000000
0!
0'
0/
#912140000000
1!
1'
1/
#912150000000
0!
1"
0'
1(
0/
10
#912160000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#912170000000
0!
1$
0'
1+
0/
#912180000000
1!
1'
1/
#912190000000
0!
0'
0/
#912200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#912210000000
0!
0'
0/
#912220000000
1!
1'
1/
#912230000000
0!
0'
0/
#912240000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#912250000000
0!
0'
0/
#912260000000
1!
1'
1/
#912270000000
0!
0'
0/
#912280000000
1!
1'
1/
#912290000000
0!
0'
0/
#912300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#912310000000
0!
0'
0/
#912320000000
1!
1'
1/
#912330000000
0!
0'
0/
#912340000000
1!
1'
1/
#912350000000
0!
0'
0/
#912360000000
1!
1'
1/
#912370000000
0!
0'
0/
#912380000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#912390000000
0!
0'
0/
#912400000000
1!
1'
1/
#912410000000
0!
0'
0/
#912420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#912430000000
0!
0'
0/
#912440000000
1!
1'
1/
#912450000000
0!
0'
0/
#912460000000
#912470000000
1!
1'
1/
#912480000000
0!
0'
0/
#912490000000
1!
1'
1/
#912500000000
0!
1"
0'
1(
0/
10
#912510000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#912520000000
0!
0'
0/
#912530000000
1!
1'
1/
#912540000000
0!
0'
0/
#912550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#912560000000
0!
0'
0/
#912570000000
1!
1'
1/
#912580000000
0!
1"
0'
1(
0/
10
#912590000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#912600000000
0!
1$
0'
1+
0/
#912610000000
1!
1'
1/
#912620000000
0!
0'
0/
#912630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#912640000000
0!
0'
0/
#912650000000
1!
1'
1/
#912660000000
0!
0'
0/
#912670000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#912680000000
0!
0'
0/
#912690000000
1!
1'
1/
#912700000000
0!
0'
0/
#912710000000
1!
1'
1/
#912720000000
0!
0'
0/
#912730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#912740000000
0!
0'
0/
#912750000000
1!
1'
1/
#912760000000
0!
0'
0/
#912770000000
1!
1'
1/
#912780000000
0!
0'
0/
#912790000000
1!
1'
1/
#912800000000
0!
0'
0/
#912810000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#912820000000
0!
0'
0/
#912830000000
1!
1'
1/
#912840000000
0!
0'
0/
#912850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#912860000000
0!
0'
0/
#912870000000
1!
1'
1/
#912880000000
0!
0'
0/
#912890000000
#912900000000
1!
1'
1/
#912910000000
0!
0'
0/
#912920000000
1!
1'
1/
#912930000000
0!
1"
0'
1(
0/
10
#912940000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#912950000000
0!
0'
0/
#912960000000
1!
1'
1/
#912970000000
0!
0'
0/
#912980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#912990000000
0!
0'
0/
#913000000000
1!
1'
1/
#913010000000
0!
1"
0'
1(
0/
10
#913020000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#913030000000
0!
1$
0'
1+
0/
#913040000000
1!
1'
1/
#913050000000
0!
0'
0/
#913060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#913070000000
0!
0'
0/
#913080000000
1!
1'
1/
#913090000000
0!
0'
0/
#913100000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#913110000000
0!
0'
0/
#913120000000
1!
1'
1/
#913130000000
0!
0'
0/
#913140000000
1!
1'
1/
#913150000000
0!
0'
0/
#913160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#913170000000
0!
0'
0/
#913180000000
1!
1'
1/
#913190000000
0!
0'
0/
#913200000000
1!
1'
1/
#913210000000
0!
0'
0/
#913220000000
1!
1'
1/
#913230000000
0!
0'
0/
#913240000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#913250000000
0!
0'
0/
#913260000000
1!
1'
1/
#913270000000
0!
0'
0/
#913280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#913290000000
0!
0'
0/
#913300000000
1!
1'
1/
#913310000000
0!
0'
0/
#913320000000
#913330000000
1!
1'
1/
#913340000000
0!
0'
0/
#913350000000
1!
1'
1/
#913360000000
0!
1"
0'
1(
0/
10
#913370000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#913380000000
0!
0'
0/
#913390000000
1!
1'
1/
#913400000000
0!
0'
0/
#913410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#913420000000
0!
0'
0/
#913430000000
1!
1'
1/
#913440000000
0!
1"
0'
1(
0/
10
#913450000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#913460000000
0!
1$
0'
1+
0/
#913470000000
1!
1'
1/
#913480000000
0!
0'
0/
#913490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#913500000000
0!
0'
0/
#913510000000
1!
1'
1/
#913520000000
0!
0'
0/
#913530000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#913540000000
0!
0'
0/
#913550000000
1!
1'
1/
#913560000000
0!
0'
0/
#913570000000
1!
1'
1/
#913580000000
0!
0'
0/
#913590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#913600000000
0!
0'
0/
#913610000000
1!
1'
1/
#913620000000
0!
0'
0/
#913630000000
1!
1'
1/
#913640000000
0!
0'
0/
#913650000000
1!
1'
1/
#913660000000
0!
0'
0/
#913670000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#913680000000
0!
0'
0/
#913690000000
1!
1'
1/
#913700000000
0!
0'
0/
#913710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#913720000000
0!
0'
0/
#913730000000
1!
1'
1/
#913740000000
0!
0'
0/
#913750000000
#913760000000
1!
1'
1/
#913770000000
0!
0'
0/
#913780000000
1!
1'
1/
#913790000000
0!
1"
0'
1(
0/
10
#913800000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#913810000000
0!
0'
0/
#913820000000
1!
1'
1/
#913830000000
0!
0'
0/
#913840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#913850000000
0!
0'
0/
#913860000000
1!
1'
1/
#913870000000
0!
1"
0'
1(
0/
10
#913880000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#913890000000
0!
1$
0'
1+
0/
#913900000000
1!
1'
1/
#913910000000
0!
0'
0/
#913920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#913930000000
0!
0'
0/
#913940000000
1!
1'
1/
#913950000000
0!
0'
0/
#913960000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#913970000000
0!
0'
0/
#913980000000
1!
1'
1/
#913990000000
0!
0'
0/
#914000000000
1!
1'
1/
#914010000000
0!
0'
0/
#914020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#914030000000
0!
0'
0/
#914040000000
1!
1'
1/
#914050000000
0!
0'
0/
#914060000000
1!
1'
1/
#914070000000
0!
0'
0/
#914080000000
1!
1'
1/
#914090000000
0!
0'
0/
#914100000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#914110000000
0!
0'
0/
#914120000000
1!
1'
1/
#914130000000
0!
0'
0/
#914140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#914150000000
0!
0'
0/
#914160000000
1!
1'
1/
#914170000000
0!
0'
0/
#914180000000
#914190000000
1!
1'
1/
#914200000000
0!
0'
0/
#914210000000
1!
1'
1/
#914220000000
0!
1"
0'
1(
0/
10
#914230000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#914240000000
0!
0'
0/
#914250000000
1!
1'
1/
#914260000000
0!
0'
0/
#914270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#914280000000
0!
0'
0/
#914290000000
1!
1'
1/
#914300000000
0!
1"
0'
1(
0/
10
#914310000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#914320000000
0!
1$
0'
1+
0/
#914330000000
1!
1'
1/
#914340000000
0!
0'
0/
#914350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#914360000000
0!
0'
0/
#914370000000
1!
1'
1/
#914380000000
0!
0'
0/
#914390000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#914400000000
0!
0'
0/
#914410000000
1!
1'
1/
#914420000000
0!
0'
0/
#914430000000
1!
1'
1/
#914440000000
0!
0'
0/
#914450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#914460000000
0!
0'
0/
#914470000000
1!
1'
1/
#914480000000
0!
0'
0/
#914490000000
1!
1'
1/
#914500000000
0!
0'
0/
#914510000000
1!
1'
1/
#914520000000
0!
0'
0/
#914530000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#914540000000
0!
0'
0/
#914550000000
1!
1'
1/
#914560000000
0!
0'
0/
#914570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#914580000000
0!
0'
0/
#914590000000
1!
1'
1/
#914600000000
0!
0'
0/
#914610000000
#914620000000
1!
1'
1/
#914630000000
0!
0'
0/
#914640000000
1!
1'
1/
#914650000000
0!
1"
0'
1(
0/
10
#914660000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#914670000000
0!
0'
0/
#914680000000
1!
1'
1/
#914690000000
0!
0'
0/
#914700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#914710000000
0!
0'
0/
#914720000000
1!
1'
1/
#914730000000
0!
1"
0'
1(
0/
10
#914740000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#914750000000
0!
1$
0'
1+
0/
#914760000000
1!
1'
1/
#914770000000
0!
0'
0/
#914780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#914790000000
0!
0'
0/
#914800000000
1!
1'
1/
#914810000000
0!
0'
0/
#914820000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#914830000000
0!
0'
0/
#914840000000
1!
1'
1/
#914850000000
0!
0'
0/
#914860000000
1!
1'
1/
#914870000000
0!
0'
0/
#914880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#914890000000
0!
0'
0/
#914900000000
1!
1'
1/
#914910000000
0!
0'
0/
#914920000000
1!
1'
1/
#914930000000
0!
0'
0/
#914940000000
1!
1'
1/
#914950000000
0!
0'
0/
#914960000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#914970000000
0!
0'
0/
#914980000000
1!
1'
1/
#914990000000
0!
0'
0/
#915000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#915010000000
0!
0'
0/
#915020000000
1!
1'
1/
#915030000000
0!
0'
0/
#915040000000
#915050000000
1!
1'
1/
#915060000000
0!
0'
0/
#915070000000
1!
1'
1/
#915080000000
0!
1"
0'
1(
0/
10
#915090000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#915100000000
0!
0'
0/
#915110000000
1!
1'
1/
#915120000000
0!
0'
0/
#915130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#915140000000
0!
0'
0/
#915150000000
1!
1'
1/
#915160000000
0!
1"
0'
1(
0/
10
#915170000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#915180000000
0!
1$
0'
1+
0/
#915190000000
1!
1'
1/
#915200000000
0!
0'
0/
#915210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#915220000000
0!
0'
0/
#915230000000
1!
1'
1/
#915240000000
0!
0'
0/
#915250000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#915260000000
0!
0'
0/
#915270000000
1!
1'
1/
#915280000000
0!
0'
0/
#915290000000
1!
1'
1/
#915300000000
0!
0'
0/
#915310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#915320000000
0!
0'
0/
#915330000000
1!
1'
1/
#915340000000
0!
0'
0/
#915350000000
1!
1'
1/
#915360000000
0!
0'
0/
#915370000000
1!
1'
1/
#915380000000
0!
0'
0/
#915390000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#915400000000
0!
0'
0/
#915410000000
1!
1'
1/
#915420000000
0!
0'
0/
#915430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#915440000000
0!
0'
0/
#915450000000
1!
1'
1/
#915460000000
0!
0'
0/
#915470000000
#915480000000
1!
1'
1/
#915490000000
0!
0'
0/
#915500000000
1!
1'
1/
#915510000000
0!
1"
0'
1(
0/
10
#915520000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#915530000000
0!
0'
0/
#915540000000
1!
1'
1/
#915550000000
0!
0'
0/
#915560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#915570000000
0!
0'
0/
#915580000000
1!
1'
1/
#915590000000
0!
1"
0'
1(
0/
10
#915600000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#915610000000
0!
1$
0'
1+
0/
#915620000000
1!
1'
1/
#915630000000
0!
0'
0/
#915640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#915650000000
0!
0'
0/
#915660000000
1!
1'
1/
#915670000000
0!
0'
0/
#915680000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#915690000000
0!
0'
0/
#915700000000
1!
1'
1/
#915710000000
0!
0'
0/
#915720000000
1!
1'
1/
#915730000000
0!
0'
0/
#915740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#915750000000
0!
0'
0/
#915760000000
1!
1'
1/
#915770000000
0!
0'
0/
#915780000000
1!
1'
1/
#915790000000
0!
0'
0/
#915800000000
1!
1'
1/
#915810000000
0!
0'
0/
#915820000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#915830000000
0!
0'
0/
#915840000000
1!
1'
1/
#915850000000
0!
0'
0/
#915860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#915870000000
0!
0'
0/
#915880000000
1!
1'
1/
#915890000000
0!
0'
0/
#915900000000
#915910000000
1!
1'
1/
#915920000000
0!
0'
0/
#915930000000
1!
1'
1/
#915940000000
0!
1"
0'
1(
0/
10
#915950000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#915960000000
0!
0'
0/
#915970000000
1!
1'
1/
#915980000000
0!
0'
0/
#915990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#916000000000
0!
0'
0/
#916010000000
1!
1'
1/
#916020000000
0!
1"
0'
1(
0/
10
#916030000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#916040000000
0!
1$
0'
1+
0/
#916050000000
1!
1'
1/
#916060000000
0!
0'
0/
#916070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#916080000000
0!
0'
0/
#916090000000
1!
1'
1/
#916100000000
0!
0'
0/
#916110000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#916120000000
0!
0'
0/
#916130000000
1!
1'
1/
#916140000000
0!
0'
0/
#916150000000
1!
1'
1/
#916160000000
0!
0'
0/
#916170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#916180000000
0!
0'
0/
#916190000000
1!
1'
1/
#916200000000
0!
0'
0/
#916210000000
1!
1'
1/
#916220000000
0!
0'
0/
#916230000000
1!
1'
1/
#916240000000
0!
0'
0/
#916250000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#916260000000
0!
0'
0/
#916270000000
1!
1'
1/
#916280000000
0!
0'
0/
#916290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#916300000000
0!
0'
0/
#916310000000
1!
1'
1/
#916320000000
0!
0'
0/
#916330000000
#916340000000
1!
1'
1/
#916350000000
0!
0'
0/
#916360000000
1!
1'
1/
#916370000000
0!
1"
0'
1(
0/
10
#916380000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#916390000000
0!
0'
0/
#916400000000
1!
1'
1/
#916410000000
0!
0'
0/
#916420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#916430000000
0!
0'
0/
#916440000000
1!
1'
1/
#916450000000
0!
1"
0'
1(
0/
10
#916460000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#916470000000
0!
1$
0'
1+
0/
#916480000000
1!
1'
1/
#916490000000
0!
0'
0/
#916500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#916510000000
0!
0'
0/
#916520000000
1!
1'
1/
#916530000000
0!
0'
0/
#916540000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#916550000000
0!
0'
0/
#916560000000
1!
1'
1/
#916570000000
0!
0'
0/
#916580000000
1!
1'
1/
#916590000000
0!
0'
0/
#916600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#916610000000
0!
0'
0/
#916620000000
1!
1'
1/
#916630000000
0!
0'
0/
#916640000000
1!
1'
1/
#916650000000
0!
0'
0/
#916660000000
1!
1'
1/
#916670000000
0!
0'
0/
#916680000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#916690000000
0!
0'
0/
#916700000000
1!
1'
1/
#916710000000
0!
0'
0/
#916720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#916730000000
0!
0'
0/
#916740000000
1!
1'
1/
#916750000000
0!
0'
0/
#916760000000
#916770000000
1!
1'
1/
#916780000000
0!
0'
0/
#916790000000
1!
1'
1/
#916800000000
0!
1"
0'
1(
0/
10
#916810000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#916820000000
0!
0'
0/
#916830000000
1!
1'
1/
#916840000000
0!
0'
0/
#916850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#916860000000
0!
0'
0/
#916870000000
1!
1'
1/
#916880000000
0!
1"
0'
1(
0/
10
#916890000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#916900000000
0!
1$
0'
1+
0/
#916910000000
1!
1'
1/
#916920000000
0!
0'
0/
#916930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#916940000000
0!
0'
0/
#916950000000
1!
1'
1/
#916960000000
0!
0'
0/
#916970000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#916980000000
0!
0'
0/
#916990000000
1!
1'
1/
#917000000000
0!
0'
0/
#917010000000
1!
1'
1/
#917020000000
0!
0'
0/
#917030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#917040000000
0!
0'
0/
#917050000000
1!
1'
1/
#917060000000
0!
0'
0/
#917070000000
1!
1'
1/
#917080000000
0!
0'
0/
#917090000000
1!
1'
1/
#917100000000
0!
0'
0/
#917110000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#917120000000
0!
0'
0/
#917130000000
1!
1'
1/
#917140000000
0!
0'
0/
#917150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#917160000000
0!
0'
0/
#917170000000
1!
1'
1/
#917180000000
0!
0'
0/
#917190000000
#917200000000
1!
1'
1/
#917210000000
0!
0'
0/
#917220000000
1!
1'
1/
#917230000000
0!
1"
0'
1(
0/
10
#917240000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#917250000000
0!
0'
0/
#917260000000
1!
1'
1/
#917270000000
0!
0'
0/
#917280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#917290000000
0!
0'
0/
#917300000000
1!
1'
1/
#917310000000
0!
1"
0'
1(
0/
10
#917320000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#917330000000
0!
1$
0'
1+
0/
#917340000000
1!
1'
1/
#917350000000
0!
0'
0/
#917360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#917370000000
0!
0'
0/
#917380000000
1!
1'
1/
#917390000000
0!
0'
0/
#917400000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#917410000000
0!
0'
0/
#917420000000
1!
1'
1/
#917430000000
0!
0'
0/
#917440000000
1!
1'
1/
#917450000000
0!
0'
0/
#917460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#917470000000
0!
0'
0/
#917480000000
1!
1'
1/
#917490000000
0!
0'
0/
#917500000000
1!
1'
1/
#917510000000
0!
0'
0/
#917520000000
1!
1'
1/
#917530000000
0!
0'
0/
#917540000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#917550000000
0!
0'
0/
#917560000000
1!
1'
1/
#917570000000
0!
0'
0/
#917580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#917590000000
0!
0'
0/
#917600000000
1!
1'
1/
#917610000000
0!
0'
0/
#917620000000
#917630000000
1!
1'
1/
#917640000000
0!
0'
0/
#917650000000
1!
1'
1/
#917660000000
0!
1"
0'
1(
0/
10
#917670000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#917680000000
0!
0'
0/
#917690000000
1!
1'
1/
#917700000000
0!
0'
0/
#917710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#917720000000
0!
0'
0/
#917730000000
1!
1'
1/
#917740000000
0!
1"
0'
1(
0/
10
#917750000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#917760000000
0!
1$
0'
1+
0/
#917770000000
1!
1'
1/
#917780000000
0!
0'
0/
#917790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#917800000000
0!
0'
0/
#917810000000
1!
1'
1/
#917820000000
0!
0'
0/
#917830000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#917840000000
0!
0'
0/
#917850000000
1!
1'
1/
#917860000000
0!
0'
0/
#917870000000
1!
1'
1/
#917880000000
0!
0'
0/
#917890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#917900000000
0!
0'
0/
#917910000000
1!
1'
1/
#917920000000
0!
0'
0/
#917930000000
1!
1'
1/
#917940000000
0!
0'
0/
#917950000000
1!
1'
1/
#917960000000
0!
0'
0/
#917970000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#917980000000
0!
0'
0/
#917990000000
1!
1'
1/
#918000000000
0!
0'
0/
#918010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#918020000000
0!
0'
0/
#918030000000
1!
1'
1/
#918040000000
0!
0'
0/
#918050000000
#918060000000
1!
1'
1/
#918070000000
0!
0'
0/
#918080000000
1!
1'
1/
#918090000000
0!
1"
0'
1(
0/
10
#918100000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#918110000000
0!
0'
0/
#918120000000
1!
1'
1/
#918130000000
0!
0'
0/
#918140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#918150000000
0!
0'
0/
#918160000000
1!
1'
1/
#918170000000
0!
1"
0'
1(
0/
10
#918180000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#918190000000
0!
1$
0'
1+
0/
#918200000000
1!
1'
1/
#918210000000
0!
0'
0/
#918220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#918230000000
0!
0'
0/
#918240000000
1!
1'
1/
#918250000000
0!
0'
0/
#918260000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#918270000000
0!
0'
0/
#918280000000
1!
1'
1/
#918290000000
0!
0'
0/
#918300000000
1!
1'
1/
#918310000000
0!
0'
0/
#918320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#918330000000
0!
0'
0/
#918340000000
1!
1'
1/
#918350000000
0!
0'
0/
#918360000000
1!
1'
1/
#918370000000
0!
0'
0/
#918380000000
1!
1'
1/
#918390000000
0!
0'
0/
#918400000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#918410000000
0!
0'
0/
#918420000000
1!
1'
1/
#918430000000
0!
0'
0/
#918440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#918450000000
0!
0'
0/
#918460000000
1!
1'
1/
#918470000000
0!
0'
0/
#918480000000
#918490000000
1!
1'
1/
#918500000000
0!
0'
0/
#918510000000
1!
1'
1/
#918520000000
0!
1"
0'
1(
0/
10
#918530000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#918540000000
0!
0'
0/
#918550000000
1!
1'
1/
#918560000000
0!
0'
0/
#918570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#918580000000
0!
0'
0/
#918590000000
1!
1'
1/
#918600000000
0!
1"
0'
1(
0/
10
#918610000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#918620000000
0!
1$
0'
1+
0/
#918630000000
1!
1'
1/
#918640000000
0!
0'
0/
#918650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#918660000000
0!
0'
0/
#918670000000
1!
1'
1/
#918680000000
0!
0'
0/
#918690000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#918700000000
0!
0'
0/
#918710000000
1!
1'
1/
#918720000000
0!
0'
0/
#918730000000
1!
1'
1/
#918740000000
0!
0'
0/
#918750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#918760000000
0!
0'
0/
#918770000000
1!
1'
1/
#918780000000
0!
0'
0/
#918790000000
1!
1'
1/
#918800000000
0!
0'
0/
#918810000000
1!
1'
1/
#918820000000
0!
0'
0/
#918830000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#918840000000
0!
0'
0/
#918850000000
1!
1'
1/
#918860000000
0!
0'
0/
#918870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#918880000000
0!
0'
0/
#918890000000
1!
1'
1/
#918900000000
0!
0'
0/
#918910000000
#918920000000
1!
1'
1/
#918930000000
0!
0'
0/
#918940000000
1!
1'
1/
#918950000000
0!
1"
0'
1(
0/
10
#918960000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#918970000000
0!
0'
0/
#918980000000
1!
1'
1/
#918990000000
0!
0'
0/
#919000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#919010000000
0!
0'
0/
#919020000000
1!
1'
1/
#919030000000
0!
1"
0'
1(
0/
10
#919040000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#919050000000
0!
1$
0'
1+
0/
#919060000000
1!
1'
1/
#919070000000
0!
0'
0/
#919080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#919090000000
0!
0'
0/
#919100000000
1!
1'
1/
#919110000000
0!
0'
0/
#919120000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#919130000000
0!
0'
0/
#919140000000
1!
1'
1/
#919150000000
0!
0'
0/
#919160000000
1!
1'
1/
#919170000000
0!
0'
0/
#919180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#919190000000
0!
0'
0/
#919200000000
1!
1'
1/
#919210000000
0!
0'
0/
#919220000000
1!
1'
1/
#919230000000
0!
0'
0/
#919240000000
1!
1'
1/
#919250000000
0!
0'
0/
#919260000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#919270000000
0!
0'
0/
#919280000000
1!
1'
1/
#919290000000
0!
0'
0/
#919300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#919310000000
0!
0'
0/
#919320000000
1!
1'
1/
#919330000000
0!
0'
0/
#919340000000
#919350000000
1!
1'
1/
#919360000000
0!
0'
0/
#919370000000
1!
1'
1/
#919380000000
0!
1"
0'
1(
0/
10
#919390000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#919400000000
0!
0'
0/
#919410000000
1!
1'
1/
#919420000000
0!
0'
0/
#919430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#919440000000
0!
0'
0/
#919450000000
1!
1'
1/
#919460000000
0!
1"
0'
1(
0/
10
#919470000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#919480000000
0!
1$
0'
1+
0/
#919490000000
1!
1'
1/
#919500000000
0!
0'
0/
#919510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#919520000000
0!
0'
0/
#919530000000
1!
1'
1/
#919540000000
0!
0'
0/
#919550000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#919560000000
0!
0'
0/
#919570000000
1!
1'
1/
#919580000000
0!
0'
0/
#919590000000
1!
1'
1/
#919600000000
0!
0'
0/
#919610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#919620000000
0!
0'
0/
#919630000000
1!
1'
1/
#919640000000
0!
0'
0/
#919650000000
1!
1'
1/
#919660000000
0!
0'
0/
#919670000000
1!
1'
1/
#919680000000
0!
0'
0/
#919690000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#919700000000
0!
0'
0/
#919710000000
1!
1'
1/
#919720000000
0!
0'
0/
#919730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#919740000000
0!
0'
0/
#919750000000
1!
1'
1/
#919760000000
0!
0'
0/
#919770000000
#919780000000
1!
1'
1/
#919790000000
0!
0'
0/
#919800000000
1!
1'
1/
#919810000000
0!
1"
0'
1(
0/
10
#919820000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#919830000000
0!
0'
0/
#919840000000
1!
1'
1/
#919850000000
0!
0'
0/
#919860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#919870000000
0!
0'
0/
#919880000000
1!
1'
1/
#919890000000
0!
1"
0'
1(
0/
10
#919900000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#919910000000
0!
1$
0'
1+
0/
#919920000000
1!
1'
1/
#919930000000
0!
0'
0/
#919940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#919950000000
0!
0'
0/
#919960000000
1!
1'
1/
#919970000000
0!
0'
0/
#919980000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#919990000000
0!
0'
0/
#920000000000
1!
1'
1/
#920010000000
0!
0'
0/
#920020000000
1!
1'
1/
#920030000000
0!
0'
0/
#920040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#920050000000
0!
0'
0/
#920060000000
1!
1'
1/
#920070000000
0!
0'
0/
#920080000000
1!
1'
1/
#920090000000
0!
0'
0/
#920100000000
1!
1'
1/
#920110000000
0!
0'
0/
#920120000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#920130000000
0!
0'
0/
#920140000000
1!
1'
1/
#920150000000
0!
0'
0/
#920160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#920170000000
0!
0'
0/
#920180000000
1!
1'
1/
#920190000000
0!
0'
0/
#920200000000
#920210000000
1!
1'
1/
#920220000000
0!
0'
0/
#920230000000
1!
1'
1/
#920240000000
0!
1"
0'
1(
0/
10
#920250000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#920260000000
0!
0'
0/
#920270000000
1!
1'
1/
#920280000000
0!
0'
0/
#920290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#920300000000
0!
0'
0/
#920310000000
1!
1'
1/
#920320000000
0!
1"
0'
1(
0/
10
#920330000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#920340000000
0!
1$
0'
1+
0/
#920350000000
1!
1'
1/
#920360000000
0!
0'
0/
#920370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#920380000000
0!
0'
0/
#920390000000
1!
1'
1/
#920400000000
0!
0'
0/
#920410000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#920420000000
0!
0'
0/
#920430000000
1!
1'
1/
#920440000000
0!
0'
0/
#920450000000
1!
1'
1/
#920460000000
0!
0'
0/
#920470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#920480000000
0!
0'
0/
#920490000000
1!
1'
1/
#920500000000
0!
0'
0/
#920510000000
1!
1'
1/
#920520000000
0!
0'
0/
#920530000000
1!
1'
1/
#920540000000
0!
0'
0/
#920550000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#920560000000
0!
0'
0/
#920570000000
1!
1'
1/
#920580000000
0!
0'
0/
#920590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#920600000000
0!
0'
0/
#920610000000
1!
1'
1/
#920620000000
0!
0'
0/
#920630000000
#920640000000
1!
1'
1/
#920650000000
0!
0'
0/
#920660000000
1!
1'
1/
#920670000000
0!
1"
0'
1(
0/
10
#920680000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#920690000000
0!
0'
0/
#920700000000
1!
1'
1/
#920710000000
0!
0'
0/
#920720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#920730000000
0!
0'
0/
#920740000000
1!
1'
1/
#920750000000
0!
1"
0'
1(
0/
10
#920760000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#920770000000
0!
1$
0'
1+
0/
#920780000000
1!
1'
1/
#920790000000
0!
0'
0/
#920800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#920810000000
0!
0'
0/
#920820000000
1!
1'
1/
#920830000000
0!
0'
0/
#920840000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#920850000000
0!
0'
0/
#920860000000
1!
1'
1/
#920870000000
0!
0'
0/
#920880000000
1!
1'
1/
#920890000000
0!
0'
0/
#920900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#920910000000
0!
0'
0/
#920920000000
1!
1'
1/
#920930000000
0!
0'
0/
#920940000000
1!
1'
1/
#920950000000
0!
0'
0/
#920960000000
1!
1'
1/
#920970000000
0!
0'
0/
#920980000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#920990000000
0!
0'
0/
#921000000000
1!
1'
1/
#921010000000
0!
0'
0/
#921020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#921030000000
0!
0'
0/
#921040000000
1!
1'
1/
#921050000000
0!
0'
0/
#921060000000
#921070000000
1!
1'
1/
#921080000000
0!
0'
0/
#921090000000
1!
1'
1/
#921100000000
0!
1"
0'
1(
0/
10
#921110000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#921120000000
0!
0'
0/
#921130000000
1!
1'
1/
#921140000000
0!
0'
0/
#921150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#921160000000
0!
0'
0/
#921170000000
1!
1'
1/
#921180000000
0!
1"
0'
1(
0/
10
#921190000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#921200000000
0!
1$
0'
1+
0/
#921210000000
1!
1'
1/
#921220000000
0!
0'
0/
#921230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#921240000000
0!
0'
0/
#921250000000
1!
1'
1/
#921260000000
0!
0'
0/
#921270000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#921280000000
0!
0'
0/
#921290000000
1!
1'
1/
#921300000000
0!
0'
0/
#921310000000
1!
1'
1/
#921320000000
0!
0'
0/
#921330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#921340000000
0!
0'
0/
#921350000000
1!
1'
1/
#921360000000
0!
0'
0/
#921370000000
1!
1'
1/
#921380000000
0!
0'
0/
#921390000000
1!
1'
1/
#921400000000
0!
0'
0/
#921410000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#921420000000
0!
0'
0/
#921430000000
1!
1'
1/
#921440000000
0!
0'
0/
#921450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#921460000000
0!
0'
0/
#921470000000
1!
1'
1/
#921480000000
0!
0'
0/
#921490000000
#921500000000
1!
1'
1/
#921510000000
0!
0'
0/
#921520000000
1!
1'
1/
#921530000000
0!
1"
0'
1(
0/
10
#921540000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#921550000000
0!
0'
0/
#921560000000
1!
1'
1/
#921570000000
0!
0'
0/
#921580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#921590000000
0!
0'
0/
#921600000000
1!
1'
1/
#921610000000
0!
1"
0'
1(
0/
10
#921620000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#921630000000
0!
1$
0'
1+
0/
#921640000000
1!
1'
1/
#921650000000
0!
0'
0/
#921660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#921670000000
0!
0'
0/
#921680000000
1!
1'
1/
#921690000000
0!
0'
0/
#921700000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#921710000000
0!
0'
0/
#921720000000
1!
1'
1/
#921730000000
0!
0'
0/
#921740000000
1!
1'
1/
#921750000000
0!
0'
0/
#921760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#921770000000
0!
0'
0/
#921780000000
1!
1'
1/
#921790000000
0!
0'
0/
#921800000000
1!
1'
1/
#921810000000
0!
0'
0/
#921820000000
1!
1'
1/
#921830000000
0!
0'
0/
#921840000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#921850000000
0!
0'
0/
#921860000000
1!
1'
1/
#921870000000
0!
0'
0/
#921880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#921890000000
0!
0'
0/
#921900000000
1!
1'
1/
#921910000000
0!
0'
0/
#921920000000
#921930000000
1!
1'
1/
#921940000000
0!
0'
0/
#921950000000
1!
1'
1/
#921960000000
0!
1"
0'
1(
0/
10
#921970000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#921980000000
0!
0'
0/
#921990000000
1!
1'
1/
#922000000000
0!
0'
0/
#922010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#922020000000
0!
0'
0/
#922030000000
1!
1'
1/
#922040000000
0!
1"
0'
1(
0/
10
#922050000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#922060000000
0!
1$
0'
1+
0/
#922070000000
1!
1'
1/
#922080000000
0!
0'
0/
#922090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#922100000000
0!
0'
0/
#922110000000
1!
1'
1/
#922120000000
0!
0'
0/
#922130000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#922140000000
0!
0'
0/
#922150000000
1!
1'
1/
#922160000000
0!
0'
0/
#922170000000
1!
1'
1/
#922180000000
0!
0'
0/
#922190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#922200000000
0!
0'
0/
#922210000000
1!
1'
1/
#922220000000
0!
0'
0/
#922230000000
1!
1'
1/
#922240000000
0!
0'
0/
#922250000000
1!
1'
1/
#922260000000
0!
0'
0/
#922270000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#922280000000
0!
0'
0/
#922290000000
1!
1'
1/
#922300000000
0!
0'
0/
#922310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#922320000000
0!
0'
0/
#922330000000
1!
1'
1/
#922340000000
0!
0'
0/
#922350000000
#922360000000
1!
1'
1/
#922370000000
0!
0'
0/
#922380000000
1!
1'
1/
#922390000000
0!
1"
0'
1(
0/
10
#922400000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#922410000000
0!
0'
0/
#922420000000
1!
1'
1/
#922430000000
0!
0'
0/
#922440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#922450000000
0!
0'
0/
#922460000000
1!
1'
1/
#922470000000
0!
1"
0'
1(
0/
10
#922480000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#922490000000
0!
1$
0'
1+
0/
#922500000000
1!
1'
1/
#922510000000
0!
0'
0/
#922520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#922530000000
0!
0'
0/
#922540000000
1!
1'
1/
#922550000000
0!
0'
0/
#922560000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#922570000000
0!
0'
0/
#922580000000
1!
1'
1/
#922590000000
0!
0'
0/
#922600000000
1!
1'
1/
#922610000000
0!
0'
0/
#922620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#922630000000
0!
0'
0/
#922640000000
1!
1'
1/
#922650000000
0!
0'
0/
#922660000000
1!
1'
1/
#922670000000
0!
0'
0/
#922680000000
1!
1'
1/
#922690000000
0!
0'
0/
#922700000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#922710000000
0!
0'
0/
#922720000000
1!
1'
1/
#922730000000
0!
0'
0/
#922740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#922750000000
0!
0'
0/
#922760000000
1!
1'
1/
#922770000000
0!
0'
0/
#922780000000
#922790000000
1!
1'
1/
#922800000000
0!
0'
0/
#922810000000
1!
1'
1/
#922820000000
0!
1"
0'
1(
0/
10
#922830000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#922840000000
0!
0'
0/
#922850000000
1!
1'
1/
#922860000000
0!
0'
0/
#922870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#922880000000
0!
0'
0/
#922890000000
1!
1'
1/
#922900000000
0!
1"
0'
1(
0/
10
#922910000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#922920000000
0!
1$
0'
1+
0/
#922930000000
1!
1'
1/
#922940000000
0!
0'
0/
#922950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#922960000000
0!
0'
0/
#922970000000
1!
1'
1/
#922980000000
0!
0'
0/
#922990000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#923000000000
0!
0'
0/
#923010000000
1!
1'
1/
#923020000000
0!
0'
0/
#923030000000
1!
1'
1/
#923040000000
0!
0'
0/
#923050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#923060000000
0!
0'
0/
#923070000000
1!
1'
1/
#923080000000
0!
0'
0/
#923090000000
1!
1'
1/
#923100000000
0!
0'
0/
#923110000000
1!
1'
1/
#923120000000
0!
0'
0/
#923130000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#923140000000
0!
0'
0/
#923150000000
1!
1'
1/
#923160000000
0!
0'
0/
#923170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#923180000000
0!
0'
0/
#923190000000
1!
1'
1/
#923200000000
0!
0'
0/
#923210000000
#923220000000
1!
1'
1/
#923230000000
0!
0'
0/
#923240000000
1!
1'
1/
#923250000000
0!
1"
0'
1(
0/
10
#923260000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#923270000000
0!
0'
0/
#923280000000
1!
1'
1/
#923290000000
0!
0'
0/
#923300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#923310000000
0!
0'
0/
#923320000000
1!
1'
1/
#923330000000
0!
1"
0'
1(
0/
10
#923340000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#923350000000
0!
1$
0'
1+
0/
#923360000000
1!
1'
1/
#923370000000
0!
0'
0/
#923380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#923390000000
0!
0'
0/
#923400000000
1!
1'
1/
#923410000000
0!
0'
0/
#923420000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#923430000000
0!
0'
0/
#923440000000
1!
1'
1/
#923450000000
0!
0'
0/
#923460000000
1!
1'
1/
#923470000000
0!
0'
0/
#923480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#923490000000
0!
0'
0/
#923500000000
1!
1'
1/
#923510000000
0!
0'
0/
#923520000000
1!
1'
1/
#923530000000
0!
0'
0/
#923540000000
1!
1'
1/
#923550000000
0!
0'
0/
#923560000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#923570000000
0!
0'
0/
#923580000000
1!
1'
1/
#923590000000
0!
0'
0/
#923600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#923610000000
0!
0'
0/
#923620000000
1!
1'
1/
#923630000000
0!
0'
0/
#923640000000
#923650000000
1!
1'
1/
#923660000000
0!
0'
0/
#923670000000
1!
1'
1/
#923680000000
0!
1"
0'
1(
0/
10
#923690000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#923700000000
0!
0'
0/
#923710000000
1!
1'
1/
#923720000000
0!
0'
0/
#923730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#923740000000
0!
0'
0/
#923750000000
1!
1'
1/
#923760000000
0!
1"
0'
1(
0/
10
#923770000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#923780000000
0!
1$
0'
1+
0/
#923790000000
1!
1'
1/
#923800000000
0!
0'
0/
#923810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#923820000000
0!
0'
0/
#923830000000
1!
1'
1/
#923840000000
0!
0'
0/
#923850000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#923860000000
0!
0'
0/
#923870000000
1!
1'
1/
#923880000000
0!
0'
0/
#923890000000
1!
1'
1/
#923900000000
0!
0'
0/
#923910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#923920000000
0!
0'
0/
#923930000000
1!
1'
1/
#923940000000
0!
0'
0/
#923950000000
1!
1'
1/
#923960000000
0!
0'
0/
#923970000000
1!
1'
1/
#923980000000
0!
0'
0/
#923990000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#924000000000
0!
0'
0/
#924010000000
1!
1'
1/
#924020000000
0!
0'
0/
#924030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#924040000000
0!
0'
0/
#924050000000
1!
1'
1/
#924060000000
0!
0'
0/
#924070000000
#924080000000
1!
1'
1/
#924090000000
0!
0'
0/
#924100000000
1!
1'
1/
#924110000000
0!
1"
0'
1(
0/
10
#924120000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#924130000000
0!
0'
0/
#924140000000
1!
1'
1/
#924150000000
0!
0'
0/
#924160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#924170000000
0!
0'
0/
#924180000000
1!
1'
1/
#924190000000
0!
1"
0'
1(
0/
10
#924200000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#924210000000
0!
1$
0'
1+
0/
#924220000000
1!
1'
1/
#924230000000
0!
0'
0/
#924240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#924250000000
0!
0'
0/
#924260000000
1!
1'
1/
#924270000000
0!
0'
0/
#924280000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#924290000000
0!
0'
0/
#924300000000
1!
1'
1/
#924310000000
0!
0'
0/
#924320000000
1!
1'
1/
#924330000000
0!
0'
0/
#924340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#924350000000
0!
0'
0/
#924360000000
1!
1'
1/
#924370000000
0!
0'
0/
#924380000000
1!
1'
1/
#924390000000
0!
0'
0/
#924400000000
1!
1'
1/
#924410000000
0!
0'
0/
#924420000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#924430000000
0!
0'
0/
#924440000000
1!
1'
1/
#924450000000
0!
0'
0/
#924460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#924470000000
0!
0'
0/
#924480000000
1!
1'
1/
#924490000000
0!
0'
0/
#924500000000
#924510000000
1!
1'
1/
#924520000000
0!
0'
0/
#924530000000
1!
1'
1/
#924540000000
0!
1"
0'
1(
0/
10
#924550000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#924560000000
0!
0'
0/
#924570000000
1!
1'
1/
#924580000000
0!
0'
0/
#924590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#924600000000
0!
0'
0/
#924610000000
1!
1'
1/
#924620000000
0!
1"
0'
1(
0/
10
#924630000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#924640000000
0!
1$
0'
1+
0/
#924650000000
1!
1'
1/
#924660000000
0!
0'
0/
#924670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#924680000000
0!
0'
0/
#924690000000
1!
1'
1/
#924700000000
0!
0'
0/
#924710000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#924720000000
0!
0'
0/
#924730000000
1!
1'
1/
#924740000000
0!
0'
0/
#924750000000
1!
1'
1/
#924760000000
0!
0'
0/
#924770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#924780000000
0!
0'
0/
#924790000000
1!
1'
1/
#924800000000
0!
0'
0/
#924810000000
1!
1'
1/
#924820000000
0!
0'
0/
#924830000000
1!
1'
1/
#924840000000
0!
0'
0/
#924850000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#924860000000
0!
0'
0/
#924870000000
1!
1'
1/
#924880000000
0!
0'
0/
#924890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#924900000000
0!
0'
0/
#924910000000
1!
1'
1/
#924920000000
0!
0'
0/
#924930000000
#924940000000
1!
1'
1/
#924950000000
0!
0'
0/
#924960000000
1!
1'
1/
#924970000000
0!
1"
0'
1(
0/
10
#924980000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#924990000000
0!
0'
0/
#925000000000
1!
1'
1/
#925010000000
0!
0'
0/
#925020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#925030000000
0!
0'
0/
#925040000000
1!
1'
1/
#925050000000
0!
1"
0'
1(
0/
10
#925060000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#925070000000
0!
1$
0'
1+
0/
#925080000000
1!
1'
1/
#925090000000
0!
0'
0/
#925100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#925110000000
0!
0'
0/
#925120000000
1!
1'
1/
#925130000000
0!
0'
0/
#925140000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#925150000000
0!
0'
0/
#925160000000
1!
1'
1/
#925170000000
0!
0'
0/
#925180000000
1!
1'
1/
#925190000000
0!
0'
0/
#925200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#925210000000
0!
0'
0/
#925220000000
1!
1'
1/
#925230000000
0!
0'
0/
#925240000000
1!
1'
1/
#925250000000
0!
0'
0/
#925260000000
1!
1'
1/
#925270000000
0!
0'
0/
#925280000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#925290000000
0!
0'
0/
#925300000000
1!
1'
1/
#925310000000
0!
0'
0/
#925320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#925330000000
0!
0'
0/
#925340000000
1!
1'
1/
#925350000000
0!
0'
0/
#925360000000
#925370000000
1!
1'
1/
#925380000000
0!
0'
0/
#925390000000
1!
1'
1/
#925400000000
0!
1"
0'
1(
0/
10
#925410000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#925420000000
0!
0'
0/
#925430000000
1!
1'
1/
#925440000000
0!
0'
0/
#925450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#925460000000
0!
0'
0/
#925470000000
1!
1'
1/
#925480000000
0!
1"
0'
1(
0/
10
#925490000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#925500000000
0!
1$
0'
1+
0/
#925510000000
1!
1'
1/
#925520000000
0!
0'
0/
#925530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#925540000000
0!
0'
0/
#925550000000
1!
1'
1/
#925560000000
0!
0'
0/
#925570000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#925580000000
0!
0'
0/
#925590000000
1!
1'
1/
#925600000000
0!
0'
0/
#925610000000
1!
1'
1/
#925620000000
0!
0'
0/
#925630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#925640000000
0!
0'
0/
#925650000000
1!
1'
1/
#925660000000
0!
0'
0/
#925670000000
1!
1'
1/
#925680000000
0!
0'
0/
#925690000000
1!
1'
1/
#925700000000
0!
0'
0/
#925710000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#925720000000
0!
0'
0/
#925730000000
1!
1'
1/
#925740000000
0!
0'
0/
#925750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#925760000000
0!
0'
0/
#925770000000
1!
1'
1/
#925780000000
0!
0'
0/
#925790000000
#925800000000
1!
1'
1/
#925810000000
0!
0'
0/
#925820000000
1!
1'
1/
#925830000000
0!
1"
0'
1(
0/
10
#925840000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#925850000000
0!
0'
0/
#925860000000
1!
1'
1/
#925870000000
0!
0'
0/
#925880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#925890000000
0!
0'
0/
#925900000000
1!
1'
1/
#925910000000
0!
1"
0'
1(
0/
10
#925920000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#925930000000
0!
1$
0'
1+
0/
#925940000000
1!
1'
1/
#925950000000
0!
0'
0/
#925960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#925970000000
0!
0'
0/
#925980000000
1!
1'
1/
#925990000000
0!
0'
0/
#926000000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#926010000000
0!
0'
0/
#926020000000
1!
1'
1/
#926030000000
0!
0'
0/
#926040000000
1!
1'
1/
#926050000000
0!
0'
0/
#926060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#926070000000
0!
0'
0/
#926080000000
1!
1'
1/
#926090000000
0!
0'
0/
#926100000000
1!
1'
1/
#926110000000
0!
0'
0/
#926120000000
1!
1'
1/
#926130000000
0!
0'
0/
#926140000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#926150000000
0!
0'
0/
#926160000000
1!
1'
1/
#926170000000
0!
0'
0/
#926180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#926190000000
0!
0'
0/
#926200000000
1!
1'
1/
#926210000000
0!
0'
0/
#926220000000
#926230000000
1!
1'
1/
#926240000000
0!
0'
0/
#926250000000
1!
1'
1/
#926260000000
0!
1"
0'
1(
0/
10
#926270000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#926280000000
0!
0'
0/
#926290000000
1!
1'
1/
#926300000000
0!
0'
0/
#926310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#926320000000
0!
0'
0/
#926330000000
1!
1'
1/
#926340000000
0!
1"
0'
1(
0/
10
#926350000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#926360000000
0!
1$
0'
1+
0/
#926370000000
1!
1'
1/
#926380000000
0!
0'
0/
#926390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#926400000000
0!
0'
0/
#926410000000
1!
1'
1/
#926420000000
0!
0'
0/
#926430000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#926440000000
0!
0'
0/
#926450000000
1!
1'
1/
#926460000000
0!
0'
0/
#926470000000
1!
1'
1/
#926480000000
0!
0'
0/
#926490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#926500000000
0!
0'
0/
#926510000000
1!
1'
1/
#926520000000
0!
0'
0/
#926530000000
1!
1'
1/
#926540000000
0!
0'
0/
#926550000000
1!
1'
1/
#926560000000
0!
0'
0/
#926570000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#926580000000
0!
0'
0/
#926590000000
1!
1'
1/
#926600000000
0!
0'
0/
#926610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#926620000000
0!
0'
0/
#926630000000
1!
1'
1/
#926640000000
0!
0'
0/
#926650000000
#926660000000
1!
1'
1/
#926670000000
0!
0'
0/
#926680000000
1!
1'
1/
#926690000000
0!
1"
0'
1(
0/
10
#926700000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#926710000000
0!
0'
0/
#926720000000
1!
1'
1/
#926730000000
0!
0'
0/
#926740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#926750000000
0!
0'
0/
#926760000000
1!
1'
1/
#926770000000
0!
1"
0'
1(
0/
10
#926780000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#926790000000
0!
1$
0'
1+
0/
#926800000000
1!
1'
1/
#926810000000
0!
0'
0/
#926820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#926830000000
0!
0'
0/
#926840000000
1!
1'
1/
#926850000000
0!
0'
0/
#926860000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#926870000000
0!
0'
0/
#926880000000
1!
1'
1/
#926890000000
0!
0'
0/
#926900000000
1!
1'
1/
#926910000000
0!
0'
0/
#926920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#926930000000
0!
0'
0/
#926940000000
1!
1'
1/
#926950000000
0!
0'
0/
#926960000000
1!
1'
1/
#926970000000
0!
0'
0/
#926980000000
1!
1'
1/
#926990000000
0!
0'
0/
#927000000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#927010000000
0!
0'
0/
#927020000000
1!
1'
1/
#927030000000
0!
0'
0/
#927040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#927050000000
0!
0'
0/
#927060000000
1!
1'
1/
#927070000000
0!
0'
0/
#927080000000
#927090000000
1!
1'
1/
#927100000000
0!
0'
0/
#927110000000
1!
1'
1/
#927120000000
0!
1"
0'
1(
0/
10
#927130000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#927140000000
0!
0'
0/
#927150000000
1!
1'
1/
#927160000000
0!
0'
0/
#927170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#927180000000
0!
0'
0/
#927190000000
1!
1'
1/
#927200000000
0!
1"
0'
1(
0/
10
#927210000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#927220000000
0!
1$
0'
1+
0/
#927230000000
1!
1'
1/
#927240000000
0!
0'
0/
#927250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#927260000000
0!
0'
0/
#927270000000
1!
1'
1/
#927280000000
0!
0'
0/
#927290000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#927300000000
0!
0'
0/
#927310000000
1!
1'
1/
#927320000000
0!
0'
0/
#927330000000
1!
1'
1/
#927340000000
0!
0'
0/
#927350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#927360000000
0!
0'
0/
#927370000000
1!
1'
1/
#927380000000
0!
0'
0/
#927390000000
1!
1'
1/
#927400000000
0!
0'
0/
#927410000000
1!
1'
1/
#927420000000
0!
0'
0/
#927430000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#927440000000
0!
0'
0/
#927450000000
1!
1'
1/
#927460000000
0!
0'
0/
#927470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#927480000000
0!
0'
0/
#927490000000
1!
1'
1/
#927500000000
0!
0'
0/
#927510000000
#927520000000
1!
1'
1/
#927530000000
0!
0'
0/
#927540000000
1!
1'
1/
#927550000000
0!
1"
0'
1(
0/
10
#927560000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#927570000000
0!
0'
0/
#927580000000
1!
1'
1/
#927590000000
0!
0'
0/
#927600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#927610000000
0!
0'
0/
#927620000000
1!
1'
1/
#927630000000
0!
1"
0'
1(
0/
10
#927640000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#927650000000
0!
1$
0'
1+
0/
#927660000000
1!
1'
1/
#927670000000
0!
0'
0/
#927680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#927690000000
0!
0'
0/
#927700000000
1!
1'
1/
#927710000000
0!
0'
0/
#927720000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#927730000000
0!
0'
0/
#927740000000
1!
1'
1/
#927750000000
0!
0'
0/
#927760000000
1!
1'
1/
#927770000000
0!
0'
0/
#927780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#927790000000
0!
0'
0/
#927800000000
1!
1'
1/
#927810000000
0!
0'
0/
#927820000000
1!
1'
1/
#927830000000
0!
0'
0/
#927840000000
1!
1'
1/
#927850000000
0!
0'
0/
#927860000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#927870000000
0!
0'
0/
#927880000000
1!
1'
1/
#927890000000
0!
0'
0/
#927900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#927910000000
0!
0'
0/
#927920000000
1!
1'
1/
#927930000000
0!
0'
0/
#927940000000
#927950000000
1!
1'
1/
#927960000000
0!
0'
0/
#927970000000
1!
1'
1/
#927980000000
0!
1"
0'
1(
0/
10
#927990000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#928000000000
0!
0'
0/
#928010000000
1!
1'
1/
#928020000000
0!
0'
0/
#928030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#928040000000
0!
0'
0/
#928050000000
1!
1'
1/
#928060000000
0!
1"
0'
1(
0/
10
#928070000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#928080000000
0!
1$
0'
1+
0/
#928090000000
1!
1'
1/
#928100000000
0!
0'
0/
#928110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#928120000000
0!
0'
0/
#928130000000
1!
1'
1/
#928140000000
0!
0'
0/
#928150000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#928160000000
0!
0'
0/
#928170000000
1!
1'
1/
#928180000000
0!
0'
0/
#928190000000
1!
1'
1/
#928200000000
0!
0'
0/
#928210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#928220000000
0!
0'
0/
#928230000000
1!
1'
1/
#928240000000
0!
0'
0/
#928250000000
1!
1'
1/
#928260000000
0!
0'
0/
#928270000000
1!
1'
1/
#928280000000
0!
0'
0/
#928290000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#928300000000
0!
0'
0/
#928310000000
1!
1'
1/
#928320000000
0!
0'
0/
#928330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#928340000000
0!
0'
0/
#928350000000
1!
1'
1/
#928360000000
0!
0'
0/
#928370000000
#928380000000
1!
1'
1/
#928390000000
0!
0'
0/
#928400000000
1!
1'
1/
#928410000000
0!
1"
0'
1(
0/
10
#928420000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#928430000000
0!
0'
0/
#928440000000
1!
1'
1/
#928450000000
0!
0'
0/
#928460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#928470000000
0!
0'
0/
#928480000000
1!
1'
1/
#928490000000
0!
1"
0'
1(
0/
10
#928500000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#928510000000
0!
1$
0'
1+
0/
#928520000000
1!
1'
1/
#928530000000
0!
0'
0/
#928540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#928550000000
0!
0'
0/
#928560000000
1!
1'
1/
#928570000000
0!
0'
0/
#928580000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#928590000000
0!
0'
0/
#928600000000
1!
1'
1/
#928610000000
0!
0'
0/
#928620000000
1!
1'
1/
#928630000000
0!
0'
0/
#928640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#928650000000
0!
0'
0/
#928660000000
1!
1'
1/
#928670000000
0!
0'
0/
#928680000000
1!
1'
1/
#928690000000
0!
0'
0/
#928700000000
1!
1'
1/
#928710000000
0!
0'
0/
#928720000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#928730000000
0!
0'
0/
#928740000000
1!
1'
1/
#928750000000
0!
0'
0/
#928760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#928770000000
0!
0'
0/
#928780000000
1!
1'
1/
#928790000000
0!
0'
0/
#928800000000
#928810000000
1!
1'
1/
#928820000000
0!
0'
0/
#928830000000
1!
1'
1/
#928840000000
0!
1"
0'
1(
0/
10
#928850000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#928860000000
0!
0'
0/
#928870000000
1!
1'
1/
#928880000000
0!
0'
0/
#928890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#928900000000
0!
0'
0/
#928910000000
1!
1'
1/
#928920000000
0!
1"
0'
1(
0/
10
#928930000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#928940000000
0!
1$
0'
1+
0/
#928950000000
1!
1'
1/
#928960000000
0!
0'
0/
#928970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#928980000000
0!
0'
0/
#928990000000
1!
1'
1/
#929000000000
0!
0'
0/
#929010000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#929020000000
0!
0'
0/
#929030000000
1!
1'
1/
#929040000000
0!
0'
0/
#929050000000
1!
1'
1/
#929060000000
0!
0'
0/
#929070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#929080000000
0!
0'
0/
#929090000000
1!
1'
1/
#929100000000
0!
0'
0/
#929110000000
1!
1'
1/
#929120000000
0!
0'
0/
#929130000000
1!
1'
1/
#929140000000
0!
0'
0/
#929150000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#929160000000
0!
0'
0/
#929170000000
1!
1'
1/
#929180000000
0!
0'
0/
#929190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#929200000000
0!
0'
0/
#929210000000
1!
1'
1/
#929220000000
0!
0'
0/
#929230000000
#929240000000
1!
1'
1/
#929250000000
0!
0'
0/
#929260000000
1!
1'
1/
#929270000000
0!
1"
0'
1(
0/
10
#929280000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#929290000000
0!
0'
0/
#929300000000
1!
1'
1/
#929310000000
0!
0'
0/
#929320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#929330000000
0!
0'
0/
#929340000000
1!
1'
1/
#929350000000
0!
1"
0'
1(
0/
10
#929360000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#929370000000
0!
1$
0'
1+
0/
#929380000000
1!
1'
1/
#929390000000
0!
0'
0/
#929400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#929410000000
0!
0'
0/
#929420000000
1!
1'
1/
#929430000000
0!
0'
0/
#929440000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#929450000000
0!
0'
0/
#929460000000
1!
1'
1/
#929470000000
0!
0'
0/
#929480000000
1!
1'
1/
#929490000000
0!
0'
0/
#929500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#929510000000
0!
0'
0/
#929520000000
1!
1'
1/
#929530000000
0!
0'
0/
#929540000000
1!
1'
1/
#929550000000
0!
0'
0/
#929560000000
1!
1'
1/
#929570000000
0!
0'
0/
#929580000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#929590000000
0!
0'
0/
#929600000000
1!
1'
1/
#929610000000
0!
0'
0/
#929620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#929630000000
0!
0'
0/
#929640000000
1!
1'
1/
#929650000000
0!
0'
0/
#929660000000
#929670000000
1!
1'
1/
#929680000000
0!
0'
0/
#929690000000
1!
1'
1/
#929700000000
0!
1"
0'
1(
0/
10
#929710000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#929720000000
0!
0'
0/
#929730000000
1!
1'
1/
#929740000000
0!
0'
0/
#929750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#929760000000
0!
0'
0/
#929770000000
1!
1'
1/
#929780000000
0!
1"
0'
1(
0/
10
#929790000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#929800000000
0!
1$
0'
1+
0/
#929810000000
1!
1'
1/
#929820000000
0!
0'
0/
#929830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#929840000000
0!
0'
0/
#929850000000
1!
1'
1/
#929860000000
0!
0'
0/
#929870000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#929880000000
0!
0'
0/
#929890000000
1!
1'
1/
#929900000000
0!
0'
0/
#929910000000
1!
1'
1/
#929920000000
0!
0'
0/
#929930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#929940000000
0!
0'
0/
#929950000000
1!
1'
1/
#929960000000
0!
0'
0/
#929970000000
1!
1'
1/
#929980000000
0!
0'
0/
#929990000000
1!
1'
1/
#930000000000
0!
0'
0/
#930010000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#930020000000
0!
0'
0/
#930030000000
1!
1'
1/
#930040000000
0!
0'
0/
#930050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#930060000000
0!
0'
0/
#930070000000
1!
1'
1/
#930080000000
0!
0'
0/
#930090000000
#930100000000
1!
1'
1/
#930110000000
0!
0'
0/
#930120000000
1!
1'
1/
#930130000000
0!
1"
0'
1(
0/
10
#930140000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#930150000000
0!
0'
0/
#930160000000
1!
1'
1/
#930170000000
0!
0'
0/
#930180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#930190000000
0!
0'
0/
#930200000000
1!
1'
1/
#930210000000
0!
1"
0'
1(
0/
10
#930220000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#930230000000
0!
1$
0'
1+
0/
#930240000000
1!
1'
1/
#930250000000
0!
0'
0/
#930260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#930270000000
0!
0'
0/
#930280000000
1!
1'
1/
#930290000000
0!
0'
0/
#930300000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#930310000000
0!
0'
0/
#930320000000
1!
1'
1/
#930330000000
0!
0'
0/
#930340000000
1!
1'
1/
#930350000000
0!
0'
0/
#930360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#930370000000
0!
0'
0/
#930380000000
1!
1'
1/
#930390000000
0!
0'
0/
#930400000000
1!
1'
1/
#930410000000
0!
0'
0/
#930420000000
1!
1'
1/
#930430000000
0!
0'
0/
#930440000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#930450000000
0!
0'
0/
#930460000000
1!
1'
1/
#930470000000
0!
0'
0/
#930480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#930490000000
0!
0'
0/
#930500000000
1!
1'
1/
#930510000000
0!
0'
0/
#930520000000
#930530000000
1!
1'
1/
#930540000000
0!
0'
0/
#930550000000
1!
1'
1/
#930560000000
0!
1"
0'
1(
0/
10
#930570000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#930580000000
0!
0'
0/
#930590000000
1!
1'
1/
#930600000000
0!
0'
0/
#930610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#930620000000
0!
0'
0/
#930630000000
1!
1'
1/
#930640000000
0!
1"
0'
1(
0/
10
#930650000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#930660000000
0!
1$
0'
1+
0/
#930670000000
1!
1'
1/
#930680000000
0!
0'
0/
#930690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#930700000000
0!
0'
0/
#930710000000
1!
1'
1/
#930720000000
0!
0'
0/
#930730000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#930740000000
0!
0'
0/
#930750000000
1!
1'
1/
#930760000000
0!
0'
0/
#930770000000
1!
1'
1/
#930780000000
0!
0'
0/
#930790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#930800000000
0!
0'
0/
#930810000000
1!
1'
1/
#930820000000
0!
0'
0/
#930830000000
1!
1'
1/
#930840000000
0!
0'
0/
#930850000000
1!
1'
1/
#930860000000
0!
0'
0/
#930870000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#930880000000
0!
0'
0/
#930890000000
1!
1'
1/
#930900000000
0!
0'
0/
#930910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#930920000000
0!
0'
0/
#930930000000
1!
1'
1/
#930940000000
0!
0'
0/
#930950000000
#930960000000
1!
1'
1/
#930970000000
0!
0'
0/
#930980000000
1!
1'
1/
#930990000000
0!
1"
0'
1(
0/
10
#931000000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#931010000000
0!
0'
0/
#931020000000
1!
1'
1/
#931030000000
0!
0'
0/
#931040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#931050000000
0!
0'
0/
#931060000000
1!
1'
1/
#931070000000
0!
1"
0'
1(
0/
10
#931080000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#931090000000
0!
1$
0'
1+
0/
#931100000000
1!
1'
1/
#931110000000
0!
0'
0/
#931120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#931130000000
0!
0'
0/
#931140000000
1!
1'
1/
#931150000000
0!
0'
0/
#931160000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#931170000000
0!
0'
0/
#931180000000
1!
1'
1/
#931190000000
0!
0'
0/
#931200000000
1!
1'
1/
#931210000000
0!
0'
0/
#931220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#931230000000
0!
0'
0/
#931240000000
1!
1'
1/
#931250000000
0!
0'
0/
#931260000000
1!
1'
1/
#931270000000
0!
0'
0/
#931280000000
1!
1'
1/
#931290000000
0!
0'
0/
#931300000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#931310000000
0!
0'
0/
#931320000000
1!
1'
1/
#931330000000
0!
0'
0/
#931340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#931350000000
0!
0'
0/
#931360000000
1!
1'
1/
#931370000000
0!
0'
0/
#931380000000
#931390000000
1!
1'
1/
#931400000000
0!
0'
0/
#931410000000
1!
1'
1/
#931420000000
0!
1"
0'
1(
0/
10
#931430000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#931440000000
0!
0'
0/
#931450000000
1!
1'
1/
#931460000000
0!
0'
0/
#931470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#931480000000
0!
0'
0/
#931490000000
1!
1'
1/
#931500000000
0!
1"
0'
1(
0/
10
#931510000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#931520000000
0!
1$
0'
1+
0/
#931530000000
1!
1'
1/
#931540000000
0!
0'
0/
#931550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#931560000000
0!
0'
0/
#931570000000
1!
1'
1/
#931580000000
0!
0'
0/
#931590000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#931600000000
0!
0'
0/
#931610000000
1!
1'
1/
#931620000000
0!
0'
0/
#931630000000
1!
1'
1/
#931640000000
0!
0'
0/
#931650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#931660000000
0!
0'
0/
#931670000000
1!
1'
1/
#931680000000
0!
0'
0/
#931690000000
1!
1'
1/
#931700000000
0!
0'
0/
#931710000000
1!
1'
1/
#931720000000
0!
0'
0/
#931730000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#931740000000
0!
0'
0/
#931750000000
1!
1'
1/
#931760000000
0!
0'
0/
#931770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#931780000000
0!
0'
0/
#931790000000
1!
1'
1/
#931800000000
0!
0'
0/
#931810000000
#931820000000
1!
1'
1/
#931830000000
0!
0'
0/
#931840000000
1!
1'
1/
#931850000000
0!
1"
0'
1(
0/
10
#931860000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#931870000000
0!
0'
0/
#931880000000
1!
1'
1/
#931890000000
0!
0'
0/
#931900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#931910000000
0!
0'
0/
#931920000000
1!
1'
1/
#931930000000
0!
1"
0'
1(
0/
10
#931940000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#931950000000
0!
1$
0'
1+
0/
#931960000000
1!
1'
1/
#931970000000
0!
0'
0/
#931980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#931990000000
0!
0'
0/
#932000000000
1!
1'
1/
#932010000000
0!
0'
0/
#932020000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#932030000000
0!
0'
0/
#932040000000
1!
1'
1/
#932050000000
0!
0'
0/
#932060000000
1!
1'
1/
#932070000000
0!
0'
0/
#932080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#932090000000
0!
0'
0/
#932100000000
1!
1'
1/
#932110000000
0!
0'
0/
#932120000000
1!
1'
1/
#932130000000
0!
0'
0/
#932140000000
1!
1'
1/
#932150000000
0!
0'
0/
#932160000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#932170000000
0!
0'
0/
#932180000000
1!
1'
1/
#932190000000
0!
0'
0/
#932200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#932210000000
0!
0'
0/
#932220000000
1!
1'
1/
#932230000000
0!
0'
0/
#932240000000
#932250000000
1!
1'
1/
#932260000000
0!
0'
0/
#932270000000
1!
1'
1/
#932280000000
0!
1"
0'
1(
0/
10
#932290000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#932300000000
0!
0'
0/
#932310000000
1!
1'
1/
#932320000000
0!
0'
0/
#932330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#932340000000
0!
0'
0/
#932350000000
1!
1'
1/
#932360000000
0!
1"
0'
1(
0/
10
#932370000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#932380000000
0!
1$
0'
1+
0/
#932390000000
1!
1'
1/
#932400000000
0!
0'
0/
#932410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#932420000000
0!
0'
0/
#932430000000
1!
1'
1/
#932440000000
0!
0'
0/
#932450000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#932460000000
0!
0'
0/
#932470000000
1!
1'
1/
#932480000000
0!
0'
0/
#932490000000
1!
1'
1/
#932500000000
0!
0'
0/
#932510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#932520000000
0!
0'
0/
#932530000000
1!
1'
1/
#932540000000
0!
0'
0/
#932550000000
1!
1'
1/
#932560000000
0!
0'
0/
#932570000000
1!
1'
1/
#932580000000
0!
0'
0/
#932590000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#932600000000
0!
0'
0/
#932610000000
1!
1'
1/
#932620000000
0!
0'
0/
#932630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#932640000000
0!
0'
0/
#932650000000
1!
1'
1/
#932660000000
0!
0'
0/
#932670000000
#932680000000
1!
1'
1/
#932690000000
0!
0'
0/
#932700000000
1!
1'
1/
#932710000000
0!
1"
0'
1(
0/
10
#932720000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#932730000000
0!
0'
0/
#932740000000
1!
1'
1/
#932750000000
0!
0'
0/
#932760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#932770000000
0!
0'
0/
#932780000000
1!
1'
1/
#932790000000
0!
1"
0'
1(
0/
10
#932800000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#932810000000
0!
1$
0'
1+
0/
#932820000000
1!
1'
1/
#932830000000
0!
0'
0/
#932840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#932850000000
0!
0'
0/
#932860000000
1!
1'
1/
#932870000000
0!
0'
0/
#932880000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#932890000000
0!
0'
0/
#932900000000
1!
1'
1/
#932910000000
0!
0'
0/
#932920000000
1!
1'
1/
#932930000000
0!
0'
0/
#932940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#932950000000
0!
0'
0/
#932960000000
1!
1'
1/
#932970000000
0!
0'
0/
#932980000000
1!
1'
1/
#932990000000
0!
0'
0/
#933000000000
1!
1'
1/
#933010000000
0!
0'
0/
#933020000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#933030000000
0!
0'
0/
#933040000000
1!
1'
1/
#933050000000
0!
0'
0/
#933060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#933070000000
0!
0'
0/
#933080000000
1!
1'
1/
#933090000000
0!
0'
0/
#933100000000
#933110000000
1!
1'
1/
#933120000000
0!
0'
0/
#933130000000
1!
1'
1/
#933140000000
0!
1"
0'
1(
0/
10
#933150000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#933160000000
0!
0'
0/
#933170000000
1!
1'
1/
#933180000000
0!
0'
0/
#933190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#933200000000
0!
0'
0/
#933210000000
1!
1'
1/
#933220000000
0!
1"
0'
1(
0/
10
#933230000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#933240000000
0!
1$
0'
1+
0/
#933250000000
1!
1'
1/
#933260000000
0!
0'
0/
#933270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#933280000000
0!
0'
0/
#933290000000
1!
1'
1/
#933300000000
0!
0'
0/
#933310000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#933320000000
0!
0'
0/
#933330000000
1!
1'
1/
#933340000000
0!
0'
0/
#933350000000
1!
1'
1/
#933360000000
0!
0'
0/
#933370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#933380000000
0!
0'
0/
#933390000000
1!
1'
1/
#933400000000
0!
0'
0/
#933410000000
1!
1'
1/
#933420000000
0!
0'
0/
#933430000000
1!
1'
1/
#933440000000
0!
0'
0/
#933450000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#933460000000
0!
0'
0/
#933470000000
1!
1'
1/
#933480000000
0!
0'
0/
#933490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#933500000000
0!
0'
0/
#933510000000
1!
1'
1/
#933520000000
0!
0'
0/
#933530000000
#933540000000
1!
1'
1/
#933550000000
0!
0'
0/
#933560000000
1!
1'
1/
#933570000000
0!
1"
0'
1(
0/
10
#933580000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#933590000000
0!
0'
0/
#933600000000
1!
1'
1/
#933610000000
0!
0'
0/
#933620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#933630000000
0!
0'
0/
#933640000000
1!
1'
1/
#933650000000
0!
1"
0'
1(
0/
10
#933660000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#933670000000
0!
1$
0'
1+
0/
#933680000000
1!
1'
1/
#933690000000
0!
0'
0/
#933700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#933710000000
0!
0'
0/
#933720000000
1!
1'
1/
#933730000000
0!
0'
0/
#933740000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#933750000000
0!
0'
0/
#933760000000
1!
1'
1/
#933770000000
0!
0'
0/
#933780000000
1!
1'
1/
#933790000000
0!
0'
0/
#933800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#933810000000
0!
0'
0/
#933820000000
1!
1'
1/
#933830000000
0!
0'
0/
#933840000000
1!
1'
1/
#933850000000
0!
0'
0/
#933860000000
1!
1'
1/
#933870000000
0!
0'
0/
#933880000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#933890000000
0!
0'
0/
#933900000000
1!
1'
1/
#933910000000
0!
0'
0/
#933920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#933930000000
0!
0'
0/
#933940000000
1!
1'
1/
#933950000000
0!
0'
0/
#933960000000
#933970000000
1!
1'
1/
#933980000000
0!
0'
0/
#933990000000
1!
1'
1/
#934000000000
0!
1"
0'
1(
0/
10
#934010000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#934020000000
0!
0'
0/
#934030000000
1!
1'
1/
#934040000000
0!
0'
0/
#934050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#934060000000
0!
0'
0/
#934070000000
1!
1'
1/
#934080000000
0!
1"
0'
1(
0/
10
#934090000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#934100000000
0!
1$
0'
1+
0/
#934110000000
1!
1'
1/
#934120000000
0!
0'
0/
#934130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#934140000000
0!
0'
0/
#934150000000
1!
1'
1/
#934160000000
0!
0'
0/
#934170000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#934180000000
0!
0'
0/
#934190000000
1!
1'
1/
#934200000000
0!
0'
0/
#934210000000
1!
1'
1/
#934220000000
0!
0'
0/
#934230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#934240000000
0!
0'
0/
#934250000000
1!
1'
1/
#934260000000
0!
0'
0/
#934270000000
1!
1'
1/
#934280000000
0!
0'
0/
#934290000000
1!
1'
1/
#934300000000
0!
0'
0/
#934310000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#934320000000
0!
0'
0/
#934330000000
1!
1'
1/
#934340000000
0!
0'
0/
#934350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#934360000000
0!
0'
0/
#934370000000
1!
1'
1/
#934380000000
0!
0'
0/
#934390000000
#934400000000
1!
1'
1/
#934410000000
0!
0'
0/
#934420000000
1!
1'
1/
#934430000000
0!
1"
0'
1(
0/
10
#934440000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#934450000000
0!
0'
0/
#934460000000
1!
1'
1/
#934470000000
0!
0'
0/
#934480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#934490000000
0!
0'
0/
#934500000000
1!
1'
1/
#934510000000
0!
1"
0'
1(
0/
10
#934520000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#934530000000
0!
1$
0'
1+
0/
#934540000000
1!
1'
1/
#934550000000
0!
0'
0/
#934560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#934570000000
0!
0'
0/
#934580000000
1!
1'
1/
#934590000000
0!
0'
0/
#934600000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#934610000000
0!
0'
0/
#934620000000
1!
1'
1/
#934630000000
0!
0'
0/
#934640000000
1!
1'
1/
#934650000000
0!
0'
0/
#934660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#934670000000
0!
0'
0/
#934680000000
1!
1'
1/
#934690000000
0!
0'
0/
#934700000000
1!
1'
1/
#934710000000
0!
0'
0/
#934720000000
1!
1'
1/
#934730000000
0!
0'
0/
#934740000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#934750000000
0!
0'
0/
#934760000000
1!
1'
1/
#934770000000
0!
0'
0/
#934780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#934790000000
0!
0'
0/
#934800000000
1!
1'
1/
#934810000000
0!
0'
0/
#934820000000
#934830000000
1!
1'
1/
#934840000000
0!
0'
0/
#934850000000
1!
1'
1/
#934860000000
0!
1"
0'
1(
0/
10
#934870000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#934880000000
0!
0'
0/
#934890000000
1!
1'
1/
#934900000000
0!
0'
0/
#934910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#934920000000
0!
0'
0/
#934930000000
1!
1'
1/
#934940000000
0!
1"
0'
1(
0/
10
#934950000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#934960000000
0!
1$
0'
1+
0/
#934970000000
1!
1'
1/
#934980000000
0!
0'
0/
#934990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#935000000000
0!
0'
0/
#935010000000
1!
1'
1/
#935020000000
0!
0'
0/
#935030000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#935040000000
0!
0'
0/
#935050000000
1!
1'
1/
#935060000000
0!
0'
0/
#935070000000
1!
1'
1/
#935080000000
0!
0'
0/
#935090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#935100000000
0!
0'
0/
#935110000000
1!
1'
1/
#935120000000
0!
0'
0/
#935130000000
1!
1'
1/
#935140000000
0!
0'
0/
#935150000000
1!
1'
1/
#935160000000
0!
0'
0/
#935170000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#935180000000
0!
0'
0/
#935190000000
1!
1'
1/
#935200000000
0!
0'
0/
#935210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#935220000000
0!
0'
0/
#935230000000
1!
1'
1/
#935240000000
0!
0'
0/
#935250000000
#935260000000
1!
1'
1/
#935270000000
0!
0'
0/
#935280000000
1!
1'
1/
#935290000000
0!
1"
0'
1(
0/
10
#935300000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#935310000000
0!
0'
0/
#935320000000
1!
1'
1/
#935330000000
0!
0'
0/
#935340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#935350000000
0!
0'
0/
#935360000000
1!
1'
1/
#935370000000
0!
1"
0'
1(
0/
10
#935380000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#935390000000
0!
1$
0'
1+
0/
#935400000000
1!
1'
1/
#935410000000
0!
0'
0/
#935420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#935430000000
0!
0'
0/
#935440000000
1!
1'
1/
#935450000000
0!
0'
0/
#935460000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#935470000000
0!
0'
0/
#935480000000
1!
1'
1/
#935490000000
0!
0'
0/
#935500000000
1!
1'
1/
#935510000000
0!
0'
0/
#935520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#935530000000
0!
0'
0/
#935540000000
1!
1'
1/
#935550000000
0!
0'
0/
#935560000000
1!
1'
1/
#935570000000
0!
0'
0/
#935580000000
1!
1'
1/
#935590000000
0!
0'
0/
#935600000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#935610000000
0!
0'
0/
#935620000000
1!
1'
1/
#935630000000
0!
0'
0/
#935640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#935650000000
0!
0'
0/
#935660000000
1!
1'
1/
#935670000000
0!
0'
0/
#935680000000
#935690000000
1!
1'
1/
#935700000000
0!
0'
0/
#935710000000
1!
1'
1/
#935720000000
0!
1"
0'
1(
0/
10
#935730000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#935740000000
0!
0'
0/
#935750000000
1!
1'
1/
#935760000000
0!
0'
0/
#935770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#935780000000
0!
0'
0/
#935790000000
1!
1'
1/
#935800000000
0!
1"
0'
1(
0/
10
#935810000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#935820000000
0!
1$
0'
1+
0/
#935830000000
1!
1'
1/
#935840000000
0!
0'
0/
#935850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#935860000000
0!
0'
0/
#935870000000
1!
1'
1/
#935880000000
0!
0'
0/
#935890000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#935900000000
0!
0'
0/
#935910000000
1!
1'
1/
#935920000000
0!
0'
0/
#935930000000
1!
1'
1/
#935940000000
0!
0'
0/
#935950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#935960000000
0!
0'
0/
#935970000000
1!
1'
1/
#935980000000
0!
0'
0/
#935990000000
1!
1'
1/
#936000000000
0!
0'
0/
#936010000000
1!
1'
1/
#936020000000
0!
0'
0/
#936030000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#936040000000
0!
0'
0/
#936050000000
1!
1'
1/
#936060000000
0!
0'
0/
#936070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#936080000000
0!
0'
0/
#936090000000
1!
1'
1/
#936100000000
0!
0'
0/
#936110000000
#936120000000
1!
1'
1/
#936130000000
0!
0'
0/
#936140000000
1!
1'
1/
#936150000000
0!
1"
0'
1(
0/
10
#936160000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#936170000000
0!
0'
0/
#936180000000
1!
1'
1/
#936190000000
0!
0'
0/
#936200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#936210000000
0!
0'
0/
#936220000000
1!
1'
1/
#936230000000
0!
1"
0'
1(
0/
10
#936240000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#936250000000
0!
1$
0'
1+
0/
#936260000000
1!
1'
1/
#936270000000
0!
0'
0/
#936280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#936290000000
0!
0'
0/
#936300000000
1!
1'
1/
#936310000000
0!
0'
0/
#936320000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#936330000000
0!
0'
0/
#936340000000
1!
1'
1/
#936350000000
0!
0'
0/
#936360000000
1!
1'
1/
#936370000000
0!
0'
0/
#936380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#936390000000
0!
0'
0/
#936400000000
1!
1'
1/
#936410000000
0!
0'
0/
#936420000000
1!
1'
1/
#936430000000
0!
0'
0/
#936440000000
1!
1'
1/
#936450000000
0!
0'
0/
#936460000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#936470000000
0!
0'
0/
#936480000000
1!
1'
1/
#936490000000
0!
0'
0/
#936500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#936510000000
0!
0'
0/
#936520000000
1!
1'
1/
#936530000000
0!
0'
0/
#936540000000
#936550000000
1!
1'
1/
#936560000000
0!
0'
0/
#936570000000
1!
1'
1/
#936580000000
0!
1"
0'
1(
0/
10
#936590000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#936600000000
0!
0'
0/
#936610000000
1!
1'
1/
#936620000000
0!
0'
0/
#936630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#936640000000
0!
0'
0/
#936650000000
1!
1'
1/
#936660000000
0!
1"
0'
1(
0/
10
#936670000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#936680000000
0!
1$
0'
1+
0/
#936690000000
1!
1'
1/
#936700000000
0!
0'
0/
#936710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#936720000000
0!
0'
0/
#936730000000
1!
1'
1/
#936740000000
0!
0'
0/
#936750000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#936760000000
0!
0'
0/
#936770000000
1!
1'
1/
#936780000000
0!
0'
0/
#936790000000
1!
1'
1/
#936800000000
0!
0'
0/
#936810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#936820000000
0!
0'
0/
#936830000000
1!
1'
1/
#936840000000
0!
0'
0/
#936850000000
1!
1'
1/
#936860000000
0!
0'
0/
#936870000000
1!
1'
1/
#936880000000
0!
0'
0/
#936890000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#936900000000
0!
0'
0/
#936910000000
1!
1'
1/
#936920000000
0!
0'
0/
#936930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#936940000000
0!
0'
0/
#936950000000
1!
1'
1/
#936960000000
0!
0'
0/
#936970000000
#936980000000
1!
1'
1/
#936990000000
0!
0'
0/
#937000000000
1!
1'
1/
#937010000000
0!
1"
0'
1(
0/
10
#937020000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#937030000000
0!
0'
0/
#937040000000
1!
1'
1/
#937050000000
0!
0'
0/
#937060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#937070000000
0!
0'
0/
#937080000000
1!
1'
1/
#937090000000
0!
1"
0'
1(
0/
10
#937100000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#937110000000
0!
1$
0'
1+
0/
#937120000000
1!
1'
1/
#937130000000
0!
0'
0/
#937140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#937150000000
0!
0'
0/
#937160000000
1!
1'
1/
#937170000000
0!
0'
0/
#937180000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#937190000000
0!
0'
0/
#937200000000
1!
1'
1/
#937210000000
0!
0'
0/
#937220000000
1!
1'
1/
#937230000000
0!
0'
0/
#937240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#937250000000
0!
0'
0/
#937260000000
1!
1'
1/
#937270000000
0!
0'
0/
#937280000000
1!
1'
1/
#937290000000
0!
0'
0/
#937300000000
1!
1'
1/
#937310000000
0!
0'
0/
#937320000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#937330000000
0!
0'
0/
#937340000000
1!
1'
1/
#937350000000
0!
0'
0/
#937360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#937370000000
0!
0'
0/
#937380000000
1!
1'
1/
#937390000000
0!
0'
0/
#937400000000
#937410000000
1!
1'
1/
#937420000000
0!
0'
0/
#937430000000
1!
1'
1/
#937440000000
0!
1"
0'
1(
0/
10
#937450000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#937460000000
0!
0'
0/
#937470000000
1!
1'
1/
#937480000000
0!
0'
0/
#937490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#937500000000
0!
0'
0/
#937510000000
1!
1'
1/
#937520000000
0!
1"
0'
1(
0/
10
#937530000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#937540000000
0!
1$
0'
1+
0/
#937550000000
1!
1'
1/
#937560000000
0!
0'
0/
#937570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#937580000000
0!
0'
0/
#937590000000
1!
1'
1/
#937600000000
0!
0'
0/
#937610000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#937620000000
0!
0'
0/
#937630000000
1!
1'
1/
#937640000000
0!
0'
0/
#937650000000
1!
1'
1/
#937660000000
0!
0'
0/
#937670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#937680000000
0!
0'
0/
#937690000000
1!
1'
1/
#937700000000
0!
0'
0/
#937710000000
1!
1'
1/
#937720000000
0!
0'
0/
#937730000000
1!
1'
1/
#937740000000
0!
0'
0/
#937750000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#937760000000
0!
0'
0/
#937770000000
1!
1'
1/
#937780000000
0!
0'
0/
#937790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#937800000000
0!
0'
0/
#937810000000
1!
1'
1/
#937820000000
0!
0'
0/
#937830000000
#937840000000
1!
1'
1/
#937850000000
0!
0'
0/
#937860000000
1!
1'
1/
#937870000000
0!
1"
0'
1(
0/
10
#937880000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#937890000000
0!
0'
0/
#937900000000
1!
1'
1/
#937910000000
0!
0'
0/
#937920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#937930000000
0!
0'
0/
#937940000000
1!
1'
1/
#937950000000
0!
1"
0'
1(
0/
10
#937960000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#937970000000
0!
1$
0'
1+
0/
#937980000000
1!
1'
1/
#937990000000
0!
0'
0/
#938000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#938010000000
0!
0'
0/
#938020000000
1!
1'
1/
#938030000000
0!
0'
0/
#938040000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#938050000000
0!
0'
0/
#938060000000
1!
1'
1/
#938070000000
0!
0'
0/
#938080000000
1!
1'
1/
#938090000000
0!
0'
0/
#938100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#938110000000
0!
0'
0/
#938120000000
1!
1'
1/
#938130000000
0!
0'
0/
#938140000000
1!
1'
1/
#938150000000
0!
0'
0/
#938160000000
1!
1'
1/
#938170000000
0!
0'
0/
#938180000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#938190000000
0!
0'
0/
#938200000000
1!
1'
1/
#938210000000
0!
0'
0/
#938220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#938230000000
0!
0'
0/
#938240000000
1!
1'
1/
#938250000000
0!
0'
0/
#938260000000
#938270000000
1!
1'
1/
#938280000000
0!
0'
0/
#938290000000
1!
1'
1/
#938300000000
0!
1"
0'
1(
0/
10
#938310000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#938320000000
0!
0'
0/
#938330000000
1!
1'
1/
#938340000000
0!
0'
0/
#938350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#938360000000
0!
0'
0/
#938370000000
1!
1'
1/
#938380000000
0!
1"
0'
1(
0/
10
#938390000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#938400000000
0!
1$
0'
1+
0/
#938410000000
1!
1'
1/
#938420000000
0!
0'
0/
#938430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#938440000000
0!
0'
0/
#938450000000
1!
1'
1/
#938460000000
0!
0'
0/
#938470000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#938480000000
0!
0'
0/
#938490000000
1!
1'
1/
#938500000000
0!
0'
0/
#938510000000
1!
1'
1/
#938520000000
0!
0'
0/
#938530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#938540000000
0!
0'
0/
#938550000000
1!
1'
1/
#938560000000
0!
0'
0/
#938570000000
1!
1'
1/
#938580000000
0!
0'
0/
#938590000000
1!
1'
1/
#938600000000
0!
0'
0/
#938610000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#938620000000
0!
0'
0/
#938630000000
1!
1'
1/
#938640000000
0!
0'
0/
#938650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#938660000000
0!
0'
0/
#938670000000
1!
1'
1/
#938680000000
0!
0'
0/
#938690000000
#938700000000
1!
1'
1/
#938710000000
0!
0'
0/
#938720000000
1!
1'
1/
#938730000000
0!
1"
0'
1(
0/
10
#938740000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#938750000000
0!
0'
0/
#938760000000
1!
1'
1/
#938770000000
0!
0'
0/
#938780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#938790000000
0!
0'
0/
#938800000000
1!
1'
1/
#938810000000
0!
1"
0'
1(
0/
10
#938820000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#938830000000
0!
1$
0'
1+
0/
#938840000000
1!
1'
1/
#938850000000
0!
0'
0/
#938860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#938870000000
0!
0'
0/
#938880000000
1!
1'
1/
#938890000000
0!
0'
0/
#938900000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#938910000000
0!
0'
0/
#938920000000
1!
1'
1/
#938930000000
0!
0'
0/
#938940000000
1!
1'
1/
#938950000000
0!
0'
0/
#938960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#938970000000
0!
0'
0/
#938980000000
1!
1'
1/
#938990000000
0!
0'
0/
#939000000000
1!
1'
1/
#939010000000
0!
0'
0/
#939020000000
1!
1'
1/
#939030000000
0!
0'
0/
#939040000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#939050000000
0!
0'
0/
#939060000000
1!
1'
1/
#939070000000
0!
0'
0/
#939080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#939090000000
0!
0'
0/
#939100000000
1!
1'
1/
#939110000000
0!
0'
0/
#939120000000
#939130000000
1!
1'
1/
#939140000000
0!
0'
0/
#939150000000
1!
1'
1/
#939160000000
0!
1"
0'
1(
0/
10
#939170000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#939180000000
0!
0'
0/
#939190000000
1!
1'
1/
#939200000000
0!
0'
0/
#939210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#939220000000
0!
0'
0/
#939230000000
1!
1'
1/
#939240000000
0!
1"
0'
1(
0/
10
#939250000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#939260000000
0!
1$
0'
1+
0/
#939270000000
1!
1'
1/
#939280000000
0!
0'
0/
#939290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#939300000000
0!
0'
0/
#939310000000
1!
1'
1/
#939320000000
0!
0'
0/
#939330000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#939340000000
0!
0'
0/
#939350000000
1!
1'
1/
#939360000000
0!
0'
0/
#939370000000
1!
1'
1/
#939380000000
0!
0'
0/
#939390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#939400000000
0!
0'
0/
#939410000000
1!
1'
1/
#939420000000
0!
0'
0/
#939430000000
1!
1'
1/
#939440000000
0!
0'
0/
#939450000000
1!
1'
1/
#939460000000
0!
0'
0/
#939470000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#939480000000
0!
0'
0/
#939490000000
1!
1'
1/
#939500000000
0!
0'
0/
#939510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#939520000000
0!
0'
0/
#939530000000
1!
1'
1/
#939540000000
0!
0'
0/
#939550000000
#939560000000
1!
1'
1/
#939570000000
0!
0'
0/
#939580000000
1!
1'
1/
#939590000000
0!
1"
0'
1(
0/
10
#939600000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#939610000000
0!
0'
0/
#939620000000
1!
1'
1/
#939630000000
0!
0'
0/
#939640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#939650000000
0!
0'
0/
#939660000000
1!
1'
1/
#939670000000
0!
1"
0'
1(
0/
10
#939680000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#939690000000
0!
1$
0'
1+
0/
#939700000000
1!
1'
1/
#939710000000
0!
0'
0/
#939720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#939730000000
0!
0'
0/
#939740000000
1!
1'
1/
#939750000000
0!
0'
0/
#939760000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#939770000000
0!
0'
0/
#939780000000
1!
1'
1/
#939790000000
0!
0'
0/
#939800000000
1!
1'
1/
#939810000000
0!
0'
0/
#939820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#939830000000
0!
0'
0/
#939840000000
1!
1'
1/
#939850000000
0!
0'
0/
#939860000000
1!
1'
1/
#939870000000
0!
0'
0/
#939880000000
1!
1'
1/
#939890000000
0!
0'
0/
#939900000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#939910000000
0!
0'
0/
#939920000000
1!
1'
1/
#939930000000
0!
0'
0/
#939940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#939950000000
0!
0'
0/
#939960000000
1!
1'
1/
#939970000000
0!
0'
0/
#939980000000
#939990000000
1!
1'
1/
#940000000000
0!
0'
0/
#940010000000
1!
1'
1/
#940020000000
0!
1"
0'
1(
0/
10
#940030000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#940040000000
0!
0'
0/
#940050000000
1!
1'
1/
#940060000000
0!
0'
0/
#940070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#940080000000
0!
0'
0/
#940090000000
1!
1'
1/
#940100000000
0!
1"
0'
1(
0/
10
#940110000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#940120000000
0!
1$
0'
1+
0/
#940130000000
1!
1'
1/
#940140000000
0!
0'
0/
#940150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#940160000000
0!
0'
0/
#940170000000
1!
1'
1/
#940180000000
0!
0'
0/
#940190000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#940200000000
0!
0'
0/
#940210000000
1!
1'
1/
#940220000000
0!
0'
0/
#940230000000
1!
1'
1/
#940240000000
0!
0'
0/
#940250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#940260000000
0!
0'
0/
#940270000000
1!
1'
1/
#940280000000
0!
0'
0/
#940290000000
1!
1'
1/
#940300000000
0!
0'
0/
#940310000000
1!
1'
1/
#940320000000
0!
0'
0/
#940330000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#940340000000
0!
0'
0/
#940350000000
1!
1'
1/
#940360000000
0!
0'
0/
#940370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#940380000000
0!
0'
0/
#940390000000
1!
1'
1/
#940400000000
0!
0'
0/
#940410000000
#940420000000
1!
1'
1/
#940430000000
0!
0'
0/
#940440000000
1!
1'
1/
#940450000000
0!
1"
0'
1(
0/
10
#940460000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#940470000000
0!
0'
0/
#940480000000
1!
1'
1/
#940490000000
0!
0'
0/
#940500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#940510000000
0!
0'
0/
#940520000000
1!
1'
1/
#940530000000
0!
1"
0'
1(
0/
10
#940540000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#940550000000
0!
1$
0'
1+
0/
#940560000000
1!
1'
1/
#940570000000
0!
0'
0/
#940580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#940590000000
0!
0'
0/
#940600000000
1!
1'
1/
#940610000000
0!
0'
0/
#940620000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#940630000000
0!
0'
0/
#940640000000
1!
1'
1/
#940650000000
0!
0'
0/
#940660000000
1!
1'
1/
#940670000000
0!
0'
0/
#940680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#940690000000
0!
0'
0/
#940700000000
1!
1'
1/
#940710000000
0!
0'
0/
#940720000000
1!
1'
1/
#940730000000
0!
0'
0/
#940740000000
1!
1'
1/
#940750000000
0!
0'
0/
#940760000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#940770000000
0!
0'
0/
#940780000000
1!
1'
1/
#940790000000
0!
0'
0/
#940800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#940810000000
0!
0'
0/
#940820000000
1!
1'
1/
#940830000000
0!
0'
0/
#940840000000
#940850000000
1!
1'
1/
#940860000000
0!
0'
0/
#940870000000
1!
1'
1/
#940880000000
0!
1"
0'
1(
0/
10
#940890000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#940900000000
0!
0'
0/
#940910000000
1!
1'
1/
#940920000000
0!
0'
0/
#940930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#940940000000
0!
0'
0/
#940950000000
1!
1'
1/
#940960000000
0!
1"
0'
1(
0/
10
#940970000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#940980000000
0!
1$
0'
1+
0/
#940990000000
1!
1'
1/
#941000000000
0!
0'
0/
#941010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#941020000000
0!
0'
0/
#941030000000
1!
1'
1/
#941040000000
0!
0'
0/
#941050000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#941060000000
0!
0'
0/
#941070000000
1!
1'
1/
#941080000000
0!
0'
0/
#941090000000
1!
1'
1/
#941100000000
0!
0'
0/
#941110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#941120000000
0!
0'
0/
#941130000000
1!
1'
1/
#941140000000
0!
0'
0/
#941150000000
1!
1'
1/
#941160000000
0!
0'
0/
#941170000000
1!
1'
1/
#941180000000
0!
0'
0/
#941190000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#941200000000
0!
0'
0/
#941210000000
1!
1'
1/
#941220000000
0!
0'
0/
#941230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#941240000000
0!
0'
0/
#941250000000
1!
1'
1/
#941260000000
0!
0'
0/
#941270000000
#941280000000
1!
1'
1/
#941290000000
0!
0'
0/
#941300000000
1!
1'
1/
#941310000000
0!
1"
0'
1(
0/
10
#941320000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#941330000000
0!
0'
0/
#941340000000
1!
1'
1/
#941350000000
0!
0'
0/
#941360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#941370000000
0!
0'
0/
#941380000000
1!
1'
1/
#941390000000
0!
1"
0'
1(
0/
10
#941400000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#941410000000
0!
1$
0'
1+
0/
#941420000000
1!
1'
1/
#941430000000
0!
0'
0/
#941440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#941450000000
0!
0'
0/
#941460000000
1!
1'
1/
#941470000000
0!
0'
0/
#941480000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#941490000000
0!
0'
0/
#941500000000
1!
1'
1/
#941510000000
0!
0'
0/
#941520000000
1!
1'
1/
#941530000000
0!
0'
0/
#941540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#941550000000
0!
0'
0/
#941560000000
1!
1'
1/
#941570000000
0!
0'
0/
#941580000000
1!
1'
1/
#941590000000
0!
0'
0/
#941600000000
1!
1'
1/
#941610000000
0!
0'
0/
#941620000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#941630000000
0!
0'
0/
#941640000000
1!
1'
1/
#941650000000
0!
0'
0/
#941660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#941670000000
0!
0'
0/
#941680000000
1!
1'
1/
#941690000000
0!
0'
0/
#941700000000
#941710000000
1!
1'
1/
#941720000000
0!
0'
0/
#941730000000
1!
1'
1/
#941740000000
0!
1"
0'
1(
0/
10
#941750000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#941760000000
0!
0'
0/
#941770000000
1!
1'
1/
#941780000000
0!
0'
0/
#941790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#941800000000
0!
0'
0/
#941810000000
1!
1'
1/
#941820000000
0!
1"
0'
1(
0/
10
#941830000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#941840000000
0!
1$
0'
1+
0/
#941850000000
1!
1'
1/
#941860000000
0!
0'
0/
#941870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#941880000000
0!
0'
0/
#941890000000
1!
1'
1/
#941900000000
0!
0'
0/
#941910000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#941920000000
0!
0'
0/
#941930000000
1!
1'
1/
#941940000000
0!
0'
0/
#941950000000
1!
1'
1/
#941960000000
0!
0'
0/
#941970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#941980000000
0!
0'
0/
#941990000000
1!
1'
1/
#942000000000
0!
0'
0/
#942010000000
1!
1'
1/
#942020000000
0!
0'
0/
#942030000000
1!
1'
1/
#942040000000
0!
0'
0/
#942050000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#942060000000
0!
0'
0/
#942070000000
1!
1'
1/
#942080000000
0!
0'
0/
#942090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#942100000000
0!
0'
0/
#942110000000
1!
1'
1/
#942120000000
0!
0'
0/
#942130000000
#942140000000
1!
1'
1/
#942150000000
0!
0'
0/
#942160000000
1!
1'
1/
#942170000000
0!
1"
0'
1(
0/
10
#942180000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#942190000000
0!
0'
0/
#942200000000
1!
1'
1/
#942210000000
0!
0'
0/
#942220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#942230000000
0!
0'
0/
#942240000000
1!
1'
1/
#942250000000
0!
1"
0'
1(
0/
10
#942260000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#942270000000
0!
1$
0'
1+
0/
#942280000000
1!
1'
1/
#942290000000
0!
0'
0/
#942300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#942310000000
0!
0'
0/
#942320000000
1!
1'
1/
#942330000000
0!
0'
0/
#942340000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#942350000000
0!
0'
0/
#942360000000
1!
1'
1/
#942370000000
0!
0'
0/
#942380000000
1!
1'
1/
#942390000000
0!
0'
0/
#942400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#942410000000
0!
0'
0/
#942420000000
1!
1'
1/
#942430000000
0!
0'
0/
#942440000000
1!
1'
1/
#942450000000
0!
0'
0/
#942460000000
1!
1'
1/
#942470000000
0!
0'
0/
#942480000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#942490000000
0!
0'
0/
#942500000000
1!
1'
1/
#942510000000
0!
0'
0/
#942520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#942530000000
0!
0'
0/
#942540000000
1!
1'
1/
#942550000000
0!
0'
0/
#942560000000
#942570000000
1!
1'
1/
#942580000000
0!
0'
0/
#942590000000
1!
1'
1/
#942600000000
0!
1"
0'
1(
0/
10
#942610000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#942620000000
0!
0'
0/
#942630000000
1!
1'
1/
#942640000000
0!
0'
0/
#942650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#942660000000
0!
0'
0/
#942670000000
1!
1'
1/
#942680000000
0!
1"
0'
1(
0/
10
#942690000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#942700000000
0!
1$
0'
1+
0/
#942710000000
1!
1'
1/
#942720000000
0!
0'
0/
#942730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#942740000000
0!
0'
0/
#942750000000
1!
1'
1/
#942760000000
0!
0'
0/
#942770000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#942780000000
0!
0'
0/
#942790000000
1!
1'
1/
#942800000000
0!
0'
0/
#942810000000
1!
1'
1/
#942820000000
0!
0'
0/
#942830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#942840000000
0!
0'
0/
#942850000000
1!
1'
1/
#942860000000
0!
0'
0/
#942870000000
1!
1'
1/
#942880000000
0!
0'
0/
#942890000000
1!
1'
1/
#942900000000
0!
0'
0/
#942910000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#942920000000
0!
0'
0/
#942930000000
1!
1'
1/
#942940000000
0!
0'
0/
#942950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#942960000000
0!
0'
0/
#942970000000
1!
1'
1/
#942980000000
0!
0'
0/
#942990000000
#943000000000
1!
1'
1/
#943010000000
0!
0'
0/
#943020000000
1!
1'
1/
#943030000000
0!
1"
0'
1(
0/
10
#943040000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#943050000000
0!
0'
0/
#943060000000
1!
1'
1/
#943070000000
0!
0'
0/
#943080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#943090000000
0!
0'
0/
#943100000000
1!
1'
1/
#943110000000
0!
1"
0'
1(
0/
10
#943120000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#943130000000
0!
1$
0'
1+
0/
#943140000000
1!
1'
1/
#943150000000
0!
0'
0/
#943160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#943170000000
0!
0'
0/
#943180000000
1!
1'
1/
#943190000000
0!
0'
0/
#943200000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#943210000000
0!
0'
0/
#943220000000
1!
1'
1/
#943230000000
0!
0'
0/
#943240000000
1!
1'
1/
#943250000000
0!
0'
0/
#943260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#943270000000
0!
0'
0/
#943280000000
1!
1'
1/
#943290000000
0!
0'
0/
#943300000000
1!
1'
1/
#943310000000
0!
0'
0/
#943320000000
1!
1'
1/
#943330000000
0!
0'
0/
#943340000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#943350000000
0!
0'
0/
#943360000000
1!
1'
1/
#943370000000
0!
0'
0/
#943380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#943390000000
0!
0'
0/
#943400000000
1!
1'
1/
#943410000000
0!
0'
0/
#943420000000
#943430000000
1!
1'
1/
#943440000000
0!
0'
0/
#943450000000
1!
1'
1/
#943460000000
0!
1"
0'
1(
0/
10
#943470000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#943480000000
0!
0'
0/
#943490000000
1!
1'
1/
#943500000000
0!
0'
0/
#943510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#943520000000
0!
0'
0/
#943530000000
1!
1'
1/
#943540000000
0!
1"
0'
1(
0/
10
#943550000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#943560000000
0!
1$
0'
1+
0/
#943570000000
1!
1'
1/
#943580000000
0!
0'
0/
#943590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#943600000000
0!
0'
0/
#943610000000
1!
1'
1/
#943620000000
0!
0'
0/
#943630000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#943640000000
0!
0'
0/
#943650000000
1!
1'
1/
#943660000000
0!
0'
0/
#943670000000
1!
1'
1/
#943680000000
0!
0'
0/
#943690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#943700000000
0!
0'
0/
#943710000000
1!
1'
1/
#943720000000
0!
0'
0/
#943730000000
1!
1'
1/
#943740000000
0!
0'
0/
#943750000000
1!
1'
1/
#943760000000
0!
0'
0/
#943770000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#943780000000
0!
0'
0/
#943790000000
1!
1'
1/
#943800000000
0!
0'
0/
#943810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#943820000000
0!
0'
0/
#943830000000
1!
1'
1/
#943840000000
0!
0'
0/
#943850000000
#943860000000
1!
1'
1/
#943870000000
0!
0'
0/
#943880000000
1!
1'
1/
#943890000000
0!
1"
0'
1(
0/
10
#943900000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#943910000000
0!
0'
0/
#943920000000
1!
1'
1/
#943930000000
0!
0'
0/
#943940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#943950000000
0!
0'
0/
#943960000000
1!
1'
1/
#943970000000
0!
1"
0'
1(
0/
10
#943980000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#943990000000
0!
1$
0'
1+
0/
#944000000000
1!
1'
1/
#944010000000
0!
0'
0/
#944020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#944030000000
0!
0'
0/
#944040000000
1!
1'
1/
#944050000000
0!
0'
0/
#944060000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#944070000000
0!
0'
0/
#944080000000
1!
1'
1/
#944090000000
0!
0'
0/
#944100000000
1!
1'
1/
#944110000000
0!
0'
0/
#944120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#944130000000
0!
0'
0/
#944140000000
1!
1'
1/
#944150000000
0!
0'
0/
#944160000000
1!
1'
1/
#944170000000
0!
0'
0/
#944180000000
1!
1'
1/
#944190000000
0!
0'
0/
#944200000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#944210000000
0!
0'
0/
#944220000000
1!
1'
1/
#944230000000
0!
0'
0/
#944240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#944250000000
0!
0'
0/
#944260000000
1!
1'
1/
#944270000000
0!
0'
0/
#944280000000
#944290000000
1!
1'
1/
#944300000000
0!
0'
0/
#944310000000
1!
1'
1/
#944320000000
0!
1"
0'
1(
0/
10
#944330000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#944340000000
0!
0'
0/
#944350000000
1!
1'
1/
#944360000000
0!
0'
0/
#944370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#944380000000
0!
0'
0/
#944390000000
1!
1'
1/
#944400000000
0!
1"
0'
1(
0/
10
#944410000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#944420000000
0!
1$
0'
1+
0/
#944430000000
1!
1'
1/
#944440000000
0!
0'
0/
#944450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#944460000000
0!
0'
0/
#944470000000
1!
1'
1/
#944480000000
0!
0'
0/
#944490000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#944500000000
0!
0'
0/
#944510000000
1!
1'
1/
#944520000000
0!
0'
0/
#944530000000
1!
1'
1/
#944540000000
0!
0'
0/
#944550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#944560000000
0!
0'
0/
#944570000000
1!
1'
1/
#944580000000
0!
0'
0/
#944590000000
1!
1'
1/
#944600000000
0!
0'
0/
#944610000000
1!
1'
1/
#944620000000
0!
0'
0/
#944630000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#944640000000
0!
0'
0/
#944650000000
1!
1'
1/
#944660000000
0!
0'
0/
#944670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#944680000000
0!
0'
0/
#944690000000
1!
1'
1/
#944700000000
0!
0'
0/
#944710000000
#944720000000
1!
1'
1/
#944730000000
0!
0'
0/
#944740000000
1!
1'
1/
#944750000000
0!
1"
0'
1(
0/
10
#944760000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#944770000000
0!
0'
0/
#944780000000
1!
1'
1/
#944790000000
0!
0'
0/
#944800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#944810000000
0!
0'
0/
#944820000000
1!
1'
1/
#944830000000
0!
1"
0'
1(
0/
10
#944840000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#944850000000
0!
1$
0'
1+
0/
#944860000000
1!
1'
1/
#944870000000
0!
0'
0/
#944880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#944890000000
0!
0'
0/
#944900000000
1!
1'
1/
#944910000000
0!
0'
0/
#944920000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#944930000000
0!
0'
0/
#944940000000
1!
1'
1/
#944950000000
0!
0'
0/
#944960000000
1!
1'
1/
#944970000000
0!
0'
0/
#944980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#944990000000
0!
0'
0/
#945000000000
1!
1'
1/
#945010000000
0!
0'
0/
#945020000000
1!
1'
1/
#945030000000
0!
0'
0/
#945040000000
1!
1'
1/
#945050000000
0!
0'
0/
#945060000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#945070000000
0!
0'
0/
#945080000000
1!
1'
1/
#945090000000
0!
0'
0/
#945100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#945110000000
0!
0'
0/
#945120000000
1!
1'
1/
#945130000000
0!
0'
0/
#945140000000
#945150000000
1!
1'
1/
#945160000000
0!
0'
0/
#945170000000
1!
1'
1/
#945180000000
0!
1"
0'
1(
0/
10
#945190000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#945200000000
0!
0'
0/
#945210000000
1!
1'
1/
#945220000000
0!
0'
0/
#945230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#945240000000
0!
0'
0/
#945250000000
1!
1'
1/
#945260000000
0!
1"
0'
1(
0/
10
#945270000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#945280000000
0!
1$
0'
1+
0/
#945290000000
1!
1'
1/
#945300000000
0!
0'
0/
#945310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#945320000000
0!
0'
0/
#945330000000
1!
1'
1/
#945340000000
0!
0'
0/
#945350000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#945360000000
0!
0'
0/
#945370000000
1!
1'
1/
#945380000000
0!
0'
0/
#945390000000
1!
1'
1/
#945400000000
0!
0'
0/
#945410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#945420000000
0!
0'
0/
#945430000000
1!
1'
1/
#945440000000
0!
0'
0/
#945450000000
1!
1'
1/
#945460000000
0!
0'
0/
#945470000000
1!
1'
1/
#945480000000
0!
0'
0/
#945490000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#945500000000
0!
0'
0/
#945510000000
1!
1'
1/
#945520000000
0!
0'
0/
#945530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#945540000000
0!
0'
0/
#945550000000
1!
1'
1/
#945560000000
0!
0'
0/
#945570000000
#945580000000
1!
1'
1/
#945590000000
0!
0'
0/
#945600000000
1!
1'
1/
#945610000000
0!
1"
0'
1(
0/
10
#945620000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#945630000000
0!
0'
0/
#945640000000
1!
1'
1/
#945650000000
0!
0'
0/
#945660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#945670000000
0!
0'
0/
#945680000000
1!
1'
1/
#945690000000
0!
1"
0'
1(
0/
10
#945700000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#945710000000
0!
1$
0'
1+
0/
#945720000000
1!
1'
1/
#945730000000
0!
0'
0/
#945740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#945750000000
0!
0'
0/
#945760000000
1!
1'
1/
#945770000000
0!
0'
0/
#945780000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#945790000000
0!
0'
0/
#945800000000
1!
1'
1/
#945810000000
0!
0'
0/
#945820000000
1!
1'
1/
#945830000000
0!
0'
0/
#945840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#945850000000
0!
0'
0/
#945860000000
1!
1'
1/
#945870000000
0!
0'
0/
#945880000000
1!
1'
1/
#945890000000
0!
0'
0/
#945900000000
1!
1'
1/
#945910000000
0!
0'
0/
#945920000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#945930000000
0!
0'
0/
#945940000000
1!
1'
1/
#945950000000
0!
0'
0/
#945960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#945970000000
0!
0'
0/
#945980000000
1!
1'
1/
#945990000000
0!
0'
0/
#946000000000
#946010000000
1!
1'
1/
#946020000000
0!
0'
0/
#946030000000
1!
1'
1/
#946040000000
0!
1"
0'
1(
0/
10
#946050000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#946060000000
0!
0'
0/
#946070000000
1!
1'
1/
#946080000000
0!
0'
0/
#946090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#946100000000
0!
0'
0/
#946110000000
1!
1'
1/
#946120000000
0!
1"
0'
1(
0/
10
#946130000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#946140000000
0!
1$
0'
1+
0/
#946150000000
1!
1'
1/
#946160000000
0!
0'
0/
#946170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#946180000000
0!
0'
0/
#946190000000
1!
1'
1/
#946200000000
0!
0'
0/
#946210000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#946220000000
0!
0'
0/
#946230000000
1!
1'
1/
#946240000000
0!
0'
0/
#946250000000
1!
1'
1/
#946260000000
0!
0'
0/
#946270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#946280000000
0!
0'
0/
#946290000000
1!
1'
1/
#946300000000
0!
0'
0/
#946310000000
1!
1'
1/
#946320000000
0!
0'
0/
#946330000000
1!
1'
1/
#946340000000
0!
0'
0/
#946350000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#946360000000
0!
0'
0/
#946370000000
1!
1'
1/
#946380000000
0!
0'
0/
#946390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#946400000000
0!
0'
0/
#946410000000
1!
1'
1/
#946420000000
0!
0'
0/
#946430000000
#946440000000
1!
1'
1/
#946450000000
0!
0'
0/
#946460000000
1!
1'
1/
#946470000000
0!
1"
0'
1(
0/
10
#946480000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#946490000000
0!
0'
0/
#946500000000
1!
1'
1/
#946510000000
0!
0'
0/
#946520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#946530000000
0!
0'
0/
#946540000000
1!
1'
1/
#946550000000
0!
1"
0'
1(
0/
10
#946560000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#946570000000
0!
1$
0'
1+
0/
#946580000000
1!
1'
1/
#946590000000
0!
0'
0/
#946600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#946610000000
0!
0'
0/
#946620000000
1!
1'
1/
#946630000000
0!
0'
0/
#946640000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#946650000000
0!
0'
0/
#946660000000
1!
1'
1/
#946670000000
0!
0'
0/
#946680000000
1!
1'
1/
#946690000000
0!
0'
0/
#946700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#946710000000
0!
0'
0/
#946720000000
1!
1'
1/
#946730000000
0!
0'
0/
#946740000000
1!
1'
1/
#946750000000
0!
0'
0/
#946760000000
1!
1'
1/
#946770000000
0!
0'
0/
#946780000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#946790000000
0!
0'
0/
#946800000000
1!
1'
1/
#946810000000
0!
0'
0/
#946820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#946830000000
0!
0'
0/
#946840000000
1!
1'
1/
#946850000000
0!
0'
0/
#946860000000
#946870000000
1!
1'
1/
#946880000000
0!
0'
0/
#946890000000
1!
1'
1/
#946900000000
0!
1"
0'
1(
0/
10
#946910000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#946920000000
0!
0'
0/
#946930000000
1!
1'
1/
#946940000000
0!
0'
0/
#946950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#946960000000
0!
0'
0/
#946970000000
1!
1'
1/
#946980000000
0!
1"
0'
1(
0/
10
#946990000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#947000000000
0!
1$
0'
1+
0/
#947010000000
1!
1'
1/
#947020000000
0!
0'
0/
#947030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#947040000000
0!
0'
0/
#947050000000
1!
1'
1/
#947060000000
0!
0'
0/
#947070000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#947080000000
0!
0'
0/
#947090000000
1!
1'
1/
#947100000000
0!
0'
0/
#947110000000
1!
1'
1/
#947120000000
0!
0'
0/
#947130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#947140000000
0!
0'
0/
#947150000000
1!
1'
1/
#947160000000
0!
0'
0/
#947170000000
1!
1'
1/
#947180000000
0!
0'
0/
#947190000000
1!
1'
1/
#947200000000
0!
0'
0/
#947210000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#947220000000
0!
0'
0/
#947230000000
1!
1'
1/
#947240000000
0!
0'
0/
#947250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#947260000000
0!
0'
0/
#947270000000
1!
1'
1/
#947280000000
0!
0'
0/
#947290000000
#947300000000
1!
1'
1/
#947310000000
0!
0'
0/
#947320000000
1!
1'
1/
#947330000000
0!
1"
0'
1(
0/
10
#947340000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#947350000000
0!
0'
0/
#947360000000
1!
1'
1/
#947370000000
0!
0'
0/
#947380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#947390000000
0!
0'
0/
#947400000000
1!
1'
1/
#947410000000
0!
1"
0'
1(
0/
10
#947420000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#947430000000
0!
1$
0'
1+
0/
#947440000000
1!
1'
1/
#947450000000
0!
0'
0/
#947460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#947470000000
0!
0'
0/
#947480000000
1!
1'
1/
#947490000000
0!
0'
0/
#947500000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#947510000000
0!
0'
0/
#947520000000
1!
1'
1/
#947530000000
0!
0'
0/
#947540000000
1!
1'
1/
#947550000000
0!
0'
0/
#947560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#947570000000
0!
0'
0/
#947580000000
1!
1'
1/
#947590000000
0!
0'
0/
#947600000000
1!
1'
1/
#947610000000
0!
0'
0/
#947620000000
1!
1'
1/
#947630000000
0!
0'
0/
#947640000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#947650000000
0!
0'
0/
#947660000000
1!
1'
1/
#947670000000
0!
0'
0/
#947680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#947690000000
0!
0'
0/
#947700000000
1!
1'
1/
#947710000000
0!
0'
0/
#947720000000
#947730000000
1!
1'
1/
#947740000000
0!
0'
0/
#947750000000
1!
1'
1/
#947760000000
0!
1"
0'
1(
0/
10
#947770000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#947780000000
0!
0'
0/
#947790000000
1!
1'
1/
#947800000000
0!
0'
0/
#947810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#947820000000
0!
0'
0/
#947830000000
1!
1'
1/
#947840000000
0!
1"
0'
1(
0/
10
#947850000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#947860000000
0!
1$
0'
1+
0/
#947870000000
1!
1'
1/
#947880000000
0!
0'
0/
#947890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#947900000000
0!
0'
0/
#947910000000
1!
1'
1/
#947920000000
0!
0'
0/
#947930000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#947940000000
0!
0'
0/
#947950000000
1!
1'
1/
#947960000000
0!
0'
0/
#947970000000
1!
1'
1/
#947980000000
0!
0'
0/
#947990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#948000000000
0!
0'
0/
#948010000000
1!
1'
1/
#948020000000
0!
0'
0/
#948030000000
1!
1'
1/
#948040000000
0!
0'
0/
#948050000000
1!
1'
1/
#948060000000
0!
0'
0/
#948070000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#948080000000
0!
0'
0/
#948090000000
1!
1'
1/
#948100000000
0!
0'
0/
#948110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#948120000000
0!
0'
0/
#948130000000
1!
1'
1/
#948140000000
0!
0'
0/
#948150000000
#948160000000
1!
1'
1/
#948170000000
0!
0'
0/
#948180000000
1!
1'
1/
#948190000000
0!
1"
0'
1(
0/
10
#948200000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#948210000000
0!
0'
0/
#948220000000
1!
1'
1/
#948230000000
0!
0'
0/
#948240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#948250000000
0!
0'
0/
#948260000000
1!
1'
1/
#948270000000
0!
1"
0'
1(
0/
10
#948280000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#948290000000
0!
1$
0'
1+
0/
#948300000000
1!
1'
1/
#948310000000
0!
0'
0/
#948320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#948330000000
0!
0'
0/
#948340000000
1!
1'
1/
#948350000000
0!
0'
0/
#948360000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#948370000000
0!
0'
0/
#948380000000
1!
1'
1/
#948390000000
0!
0'
0/
#948400000000
1!
1'
1/
#948410000000
0!
0'
0/
#948420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#948430000000
0!
0'
0/
#948440000000
1!
1'
1/
#948450000000
0!
0'
0/
#948460000000
1!
1'
1/
#948470000000
0!
0'
0/
#948480000000
1!
1'
1/
#948490000000
0!
0'
0/
#948500000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#948510000000
0!
0'
0/
#948520000000
1!
1'
1/
#948530000000
0!
0'
0/
#948540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#948550000000
0!
0'
0/
#948560000000
1!
1'
1/
#948570000000
0!
0'
0/
#948580000000
#948590000000
1!
1'
1/
#948600000000
0!
0'
0/
#948610000000
1!
1'
1/
#948620000000
0!
1"
0'
1(
0/
10
#948630000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#948640000000
0!
0'
0/
#948650000000
1!
1'
1/
#948660000000
0!
0'
0/
#948670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#948680000000
0!
0'
0/
#948690000000
1!
1'
1/
#948700000000
0!
1"
0'
1(
0/
10
#948710000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#948720000000
0!
1$
0'
1+
0/
#948730000000
1!
1'
1/
#948740000000
0!
0'
0/
#948750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#948760000000
0!
0'
0/
#948770000000
1!
1'
1/
#948780000000
0!
0'
0/
#948790000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#948800000000
0!
0'
0/
#948810000000
1!
1'
1/
#948820000000
0!
0'
0/
#948830000000
1!
1'
1/
#948840000000
0!
0'
0/
#948850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#948860000000
0!
0'
0/
#948870000000
1!
1'
1/
#948880000000
0!
0'
0/
#948890000000
1!
1'
1/
#948900000000
0!
0'
0/
#948910000000
1!
1'
1/
#948920000000
0!
0'
0/
#948930000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#948940000000
0!
0'
0/
#948950000000
1!
1'
1/
#948960000000
0!
0'
0/
#948970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#948980000000
0!
0'
0/
#948990000000
1!
1'
1/
#949000000000
0!
0'
0/
#949010000000
#949020000000
1!
1'
1/
#949030000000
0!
0'
0/
#949040000000
1!
1'
1/
#949050000000
0!
1"
0'
1(
0/
10
#949060000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#949070000000
0!
0'
0/
#949080000000
1!
1'
1/
#949090000000
0!
0'
0/
#949100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#949110000000
0!
0'
0/
#949120000000
1!
1'
1/
#949130000000
0!
1"
0'
1(
0/
10
#949140000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#949150000000
0!
1$
0'
1+
0/
#949160000000
1!
1'
1/
#949170000000
0!
0'
0/
#949180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#949190000000
0!
0'
0/
#949200000000
1!
1'
1/
#949210000000
0!
0'
0/
#949220000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#949230000000
0!
0'
0/
#949240000000
1!
1'
1/
#949250000000
0!
0'
0/
#949260000000
1!
1'
1/
#949270000000
0!
0'
0/
#949280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#949290000000
0!
0'
0/
#949300000000
1!
1'
1/
#949310000000
0!
0'
0/
#949320000000
1!
1'
1/
#949330000000
0!
0'
0/
#949340000000
1!
1'
1/
#949350000000
0!
0'
0/
#949360000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#949370000000
0!
0'
0/
#949380000000
1!
1'
1/
#949390000000
0!
0'
0/
#949400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#949410000000
0!
0'
0/
#949420000000
1!
1'
1/
#949430000000
0!
0'
0/
#949440000000
#949450000000
1!
1'
1/
#949460000000
0!
0'
0/
#949470000000
1!
1'
1/
#949480000000
0!
1"
0'
1(
0/
10
#949490000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#949500000000
0!
0'
0/
#949510000000
1!
1'
1/
#949520000000
0!
0'
0/
#949530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#949540000000
0!
0'
0/
#949550000000
1!
1'
1/
#949560000000
0!
1"
0'
1(
0/
10
#949570000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#949580000000
0!
1$
0'
1+
0/
#949590000000
1!
1'
1/
#949600000000
0!
0'
0/
#949610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#949620000000
0!
0'
0/
#949630000000
1!
1'
1/
#949640000000
0!
0'
0/
#949650000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#949660000000
0!
0'
0/
#949670000000
1!
1'
1/
#949680000000
0!
0'
0/
#949690000000
1!
1'
1/
#949700000000
0!
0'
0/
#949710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#949720000000
0!
0'
0/
#949730000000
1!
1'
1/
#949740000000
0!
0'
0/
#949750000000
1!
1'
1/
#949760000000
0!
0'
0/
#949770000000
1!
1'
1/
#949780000000
0!
0'
0/
#949790000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#949800000000
0!
0'
0/
#949810000000
1!
1'
1/
#949820000000
0!
0'
0/
#949830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#949840000000
0!
0'
0/
#949850000000
1!
1'
1/
#949860000000
0!
0'
0/
#949870000000
#949880000000
1!
1'
1/
#949890000000
0!
0'
0/
#949900000000
1!
1'
1/
#949910000000
0!
1"
0'
1(
0/
10
#949920000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#949930000000
0!
0'
0/
#949940000000
1!
1'
1/
#949950000000
0!
0'
0/
#949960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#949970000000
0!
0'
0/
#949980000000
1!
1'
1/
#949990000000
0!
1"
0'
1(
0/
10
#950000000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#950010000000
0!
1$
0'
1+
0/
#950020000000
1!
1'
1/
#950030000000
0!
0'
0/
#950040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#950050000000
0!
0'
0/
#950060000000
1!
1'
1/
#950070000000
0!
0'
0/
#950080000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#950090000000
0!
0'
0/
#950100000000
1!
1'
1/
#950110000000
0!
0'
0/
#950120000000
1!
1'
1/
#950130000000
0!
0'
0/
#950140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#950150000000
0!
0'
0/
#950160000000
1!
1'
1/
#950170000000
0!
0'
0/
#950180000000
1!
1'
1/
#950190000000
0!
0'
0/
#950200000000
1!
1'
1/
#950210000000
0!
0'
0/
#950220000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#950230000000
0!
0'
0/
#950240000000
1!
1'
1/
#950250000000
0!
0'
0/
#950260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#950270000000
0!
0'
0/
#950280000000
1!
1'
1/
#950290000000
0!
0'
0/
#950300000000
#950310000000
1!
1'
1/
#950320000000
0!
0'
0/
#950330000000
1!
1'
1/
#950340000000
0!
1"
0'
1(
0/
10
#950350000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#950360000000
0!
0'
0/
#950370000000
1!
1'
1/
#950380000000
0!
0'
0/
#950390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#950400000000
0!
0'
0/
#950410000000
1!
1'
1/
#950420000000
0!
1"
0'
1(
0/
10
#950430000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#950440000000
0!
1$
0'
1+
0/
#950450000000
1!
1'
1/
#950460000000
0!
0'
0/
#950470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#950480000000
0!
0'
0/
#950490000000
1!
1'
1/
#950500000000
0!
0'
0/
#950510000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#950520000000
0!
0'
0/
#950530000000
1!
1'
1/
#950540000000
0!
0'
0/
#950550000000
1!
1'
1/
#950560000000
0!
0'
0/
#950570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#950580000000
0!
0'
0/
#950590000000
1!
1'
1/
#950600000000
0!
0'
0/
#950610000000
1!
1'
1/
#950620000000
0!
0'
0/
#950630000000
1!
1'
1/
#950640000000
0!
0'
0/
#950650000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#950660000000
0!
0'
0/
#950670000000
1!
1'
1/
#950680000000
0!
0'
0/
#950690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#950700000000
0!
0'
0/
#950710000000
1!
1'
1/
#950720000000
0!
0'
0/
#950730000000
#950740000000
1!
1'
1/
#950750000000
0!
0'
0/
#950760000000
1!
1'
1/
#950770000000
0!
1"
0'
1(
0/
10
#950780000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#950790000000
0!
0'
0/
#950800000000
1!
1'
1/
#950810000000
0!
0'
0/
#950820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#950830000000
0!
0'
0/
#950840000000
1!
1'
1/
#950850000000
0!
1"
0'
1(
0/
10
#950860000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#950870000000
0!
1$
0'
1+
0/
#950880000000
1!
1'
1/
#950890000000
0!
0'
0/
#950900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#950910000000
0!
0'
0/
#950920000000
1!
1'
1/
#950930000000
0!
0'
0/
#950940000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#950950000000
0!
0'
0/
#950960000000
1!
1'
1/
#950970000000
0!
0'
0/
#950980000000
1!
1'
1/
#950990000000
0!
0'
0/
#951000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#951010000000
0!
0'
0/
#951020000000
1!
1'
1/
#951030000000
0!
0'
0/
#951040000000
1!
1'
1/
#951050000000
0!
0'
0/
#951060000000
1!
1'
1/
#951070000000
0!
0'
0/
#951080000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#951090000000
0!
0'
0/
#951100000000
1!
1'
1/
#951110000000
0!
0'
0/
#951120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#951130000000
0!
0'
0/
#951140000000
1!
1'
1/
#951150000000
0!
0'
0/
#951160000000
#951170000000
1!
1'
1/
#951180000000
0!
0'
0/
#951190000000
1!
1'
1/
#951200000000
0!
1"
0'
1(
0/
10
#951210000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#951220000000
0!
0'
0/
#951230000000
1!
1'
1/
#951240000000
0!
0'
0/
#951250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#951260000000
0!
0'
0/
#951270000000
1!
1'
1/
#951280000000
0!
1"
0'
1(
0/
10
#951290000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#951300000000
0!
1$
0'
1+
0/
#951310000000
1!
1'
1/
#951320000000
0!
0'
0/
#951330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#951340000000
0!
0'
0/
#951350000000
1!
1'
1/
#951360000000
0!
0'
0/
#951370000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#951380000000
0!
0'
0/
#951390000000
1!
1'
1/
#951400000000
0!
0'
0/
#951410000000
1!
1'
1/
#951420000000
0!
0'
0/
#951430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#951440000000
0!
0'
0/
#951450000000
1!
1'
1/
#951460000000
0!
0'
0/
#951470000000
1!
1'
1/
#951480000000
0!
0'
0/
#951490000000
1!
1'
1/
#951500000000
0!
0'
0/
#951510000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#951520000000
0!
0'
0/
#951530000000
1!
1'
1/
#951540000000
0!
0'
0/
#951550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#951560000000
0!
0'
0/
#951570000000
1!
1'
1/
#951580000000
0!
0'
0/
#951590000000
#951600000000
1!
1'
1/
#951610000000
0!
0'
0/
#951620000000
1!
1'
1/
#951630000000
0!
1"
0'
1(
0/
10
#951640000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#951650000000
0!
0'
0/
#951660000000
1!
1'
1/
#951670000000
0!
0'
0/
#951680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#951690000000
0!
0'
0/
#951700000000
1!
1'
1/
#951710000000
0!
1"
0'
1(
0/
10
#951720000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#951730000000
0!
1$
0'
1+
0/
#951740000000
1!
1'
1/
#951750000000
0!
0'
0/
#951760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#951770000000
0!
0'
0/
#951780000000
1!
1'
1/
#951790000000
0!
0'
0/
#951800000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#951810000000
0!
0'
0/
#951820000000
1!
1'
1/
#951830000000
0!
0'
0/
#951840000000
1!
1'
1/
#951850000000
0!
0'
0/
#951860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#951870000000
0!
0'
0/
#951880000000
1!
1'
1/
#951890000000
0!
0'
0/
#951900000000
1!
1'
1/
#951910000000
0!
0'
0/
#951920000000
1!
1'
1/
#951930000000
0!
0'
0/
#951940000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#951950000000
0!
0'
0/
#951960000000
1!
1'
1/
#951970000000
0!
0'
0/
#951980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#951990000000
0!
0'
0/
#952000000000
1!
1'
1/
#952010000000
0!
0'
0/
#952020000000
#952030000000
1!
1'
1/
#952040000000
0!
0'
0/
#952050000000
1!
1'
1/
#952060000000
0!
1"
0'
1(
0/
10
#952070000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#952080000000
0!
0'
0/
#952090000000
1!
1'
1/
#952100000000
0!
0'
0/
#952110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#952120000000
0!
0'
0/
#952130000000
1!
1'
1/
#952140000000
0!
1"
0'
1(
0/
10
#952150000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#952160000000
0!
1$
0'
1+
0/
#952170000000
1!
1'
1/
#952180000000
0!
0'
0/
#952190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#952200000000
0!
0'
0/
#952210000000
1!
1'
1/
#952220000000
0!
0'
0/
#952230000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#952240000000
0!
0'
0/
#952250000000
1!
1'
1/
#952260000000
0!
0'
0/
#952270000000
1!
1'
1/
#952280000000
0!
0'
0/
#952290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#952300000000
0!
0'
0/
#952310000000
1!
1'
1/
#952320000000
0!
0'
0/
#952330000000
1!
1'
1/
#952340000000
0!
0'
0/
#952350000000
1!
1'
1/
#952360000000
0!
0'
0/
#952370000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#952380000000
0!
0'
0/
#952390000000
1!
1'
1/
#952400000000
0!
0'
0/
#952410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#952420000000
0!
0'
0/
#952430000000
1!
1'
1/
#952440000000
0!
0'
0/
#952450000000
#952460000000
1!
1'
1/
#952470000000
0!
0'
0/
#952480000000
1!
1'
1/
#952490000000
0!
1"
0'
1(
0/
10
#952500000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#952510000000
0!
0'
0/
#952520000000
1!
1'
1/
#952530000000
0!
0'
0/
#952540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#952550000000
0!
0'
0/
#952560000000
1!
1'
1/
#952570000000
0!
1"
0'
1(
0/
10
#952580000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#952590000000
0!
1$
0'
1+
0/
#952600000000
1!
1'
1/
#952610000000
0!
0'
0/
#952620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#952630000000
0!
0'
0/
#952640000000
1!
1'
1/
#952650000000
0!
0'
0/
#952660000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#952670000000
0!
0'
0/
#952680000000
1!
1'
1/
#952690000000
0!
0'
0/
#952700000000
1!
1'
1/
#952710000000
0!
0'
0/
#952720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#952730000000
0!
0'
0/
#952740000000
1!
1'
1/
#952750000000
0!
0'
0/
#952760000000
1!
1'
1/
#952770000000
0!
0'
0/
#952780000000
1!
1'
1/
#952790000000
0!
0'
0/
#952800000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#952810000000
0!
0'
0/
#952820000000
1!
1'
1/
#952830000000
0!
0'
0/
#952840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#952850000000
0!
0'
0/
#952860000000
1!
1'
1/
#952870000000
0!
0'
0/
#952880000000
#952890000000
1!
1'
1/
#952900000000
0!
0'
0/
#952910000000
1!
1'
1/
#952920000000
0!
1"
0'
1(
0/
10
#952930000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#952940000000
0!
0'
0/
#952950000000
1!
1'
1/
#952960000000
0!
0'
0/
#952970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#952980000000
0!
0'
0/
#952990000000
1!
1'
1/
#953000000000
0!
1"
0'
1(
0/
10
#953010000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#953020000000
0!
1$
0'
1+
0/
#953030000000
1!
1'
1/
#953040000000
0!
0'
0/
#953050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#953060000000
0!
0'
0/
#953070000000
1!
1'
1/
#953080000000
0!
0'
0/
#953090000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#953100000000
0!
0'
0/
#953110000000
1!
1'
1/
#953120000000
0!
0'
0/
#953130000000
1!
1'
1/
#953140000000
0!
0'
0/
#953150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#953160000000
0!
0'
0/
#953170000000
1!
1'
1/
#953180000000
0!
0'
0/
#953190000000
1!
1'
1/
#953200000000
0!
0'
0/
#953210000000
1!
1'
1/
#953220000000
0!
0'
0/
#953230000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#953240000000
0!
0'
0/
#953250000000
1!
1'
1/
#953260000000
0!
0'
0/
#953270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#953280000000
0!
0'
0/
#953290000000
1!
1'
1/
#953300000000
0!
0'
0/
#953310000000
#953320000000
1!
1'
1/
#953330000000
0!
0'
0/
#953340000000
1!
1'
1/
#953350000000
0!
1"
0'
1(
0/
10
#953360000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#953370000000
0!
0'
0/
#953380000000
1!
1'
1/
#953390000000
0!
0'
0/
#953400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#953410000000
0!
0'
0/
#953420000000
1!
1'
1/
#953430000000
0!
1"
0'
1(
0/
10
#953440000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#953450000000
0!
1$
0'
1+
0/
#953460000000
1!
1'
1/
#953470000000
0!
0'
0/
#953480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#953490000000
0!
0'
0/
#953500000000
1!
1'
1/
#953510000000
0!
0'
0/
#953520000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#953530000000
0!
0'
0/
#953540000000
1!
1'
1/
#953550000000
0!
0'
0/
#953560000000
1!
1'
1/
#953570000000
0!
0'
0/
#953580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#953590000000
0!
0'
0/
#953600000000
1!
1'
1/
#953610000000
0!
0'
0/
#953620000000
1!
1'
1/
#953630000000
0!
0'
0/
#953640000000
1!
1'
1/
#953650000000
0!
0'
0/
#953660000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#953670000000
0!
0'
0/
#953680000000
1!
1'
1/
#953690000000
0!
0'
0/
#953700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#953710000000
0!
0'
0/
#953720000000
1!
1'
1/
#953730000000
0!
0'
0/
#953740000000
#953750000000
1!
1'
1/
#953760000000
0!
0'
0/
#953770000000
1!
1'
1/
#953780000000
0!
1"
0'
1(
0/
10
#953790000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#953800000000
0!
0'
0/
#953810000000
1!
1'
1/
#953820000000
0!
0'
0/
#953830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#953840000000
0!
0'
0/
#953850000000
1!
1'
1/
#953860000000
0!
1"
0'
1(
0/
10
#953870000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#953880000000
0!
1$
0'
1+
0/
#953890000000
1!
1'
1/
#953900000000
0!
0'
0/
#953910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#953920000000
0!
0'
0/
#953930000000
1!
1'
1/
#953940000000
0!
0'
0/
#953950000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#953960000000
0!
0'
0/
#953970000000
1!
1'
1/
#953980000000
0!
0'
0/
#953990000000
1!
1'
1/
#954000000000
0!
0'
0/
#954010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#954020000000
0!
0'
0/
#954030000000
1!
1'
1/
#954040000000
0!
0'
0/
#954050000000
1!
1'
1/
#954060000000
0!
0'
0/
#954070000000
1!
1'
1/
#954080000000
0!
0'
0/
#954090000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#954100000000
0!
0'
0/
#954110000000
1!
1'
1/
#954120000000
0!
0'
0/
#954130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#954140000000
0!
0'
0/
#954150000000
1!
1'
1/
#954160000000
0!
0'
0/
#954170000000
#954180000000
1!
1'
1/
#954190000000
0!
0'
0/
#954200000000
1!
1'
1/
#954210000000
0!
1"
0'
1(
0/
10
#954220000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#954230000000
0!
0'
0/
#954240000000
1!
1'
1/
#954250000000
0!
0'
0/
#954260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#954270000000
0!
0'
0/
#954280000000
1!
1'
1/
#954290000000
0!
1"
0'
1(
0/
10
#954300000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#954310000000
0!
1$
0'
1+
0/
#954320000000
1!
1'
1/
#954330000000
0!
0'
0/
#954340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#954350000000
0!
0'
0/
#954360000000
1!
1'
1/
#954370000000
0!
0'
0/
#954380000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#954390000000
0!
0'
0/
#954400000000
1!
1'
1/
#954410000000
0!
0'
0/
#954420000000
1!
1'
1/
#954430000000
0!
0'
0/
#954440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#954450000000
0!
0'
0/
#954460000000
1!
1'
1/
#954470000000
0!
0'
0/
#954480000000
1!
1'
1/
#954490000000
0!
0'
0/
#954500000000
1!
1'
1/
#954510000000
0!
0'
0/
#954520000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#954530000000
0!
0'
0/
#954540000000
1!
1'
1/
#954550000000
0!
0'
0/
#954560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#954570000000
0!
0'
0/
#954580000000
1!
1'
1/
#954590000000
0!
0'
0/
#954600000000
#954610000000
1!
1'
1/
#954620000000
0!
0'
0/
#954630000000
1!
1'
1/
#954640000000
0!
1"
0'
1(
0/
10
#954650000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#954660000000
0!
0'
0/
#954670000000
1!
1'
1/
#954680000000
0!
0'
0/
#954690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#954700000000
0!
0'
0/
#954710000000
1!
1'
1/
#954720000000
0!
1"
0'
1(
0/
10
#954730000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#954740000000
0!
1$
0'
1+
0/
#954750000000
1!
1'
1/
#954760000000
0!
0'
0/
#954770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#954780000000
0!
0'
0/
#954790000000
1!
1'
1/
#954800000000
0!
0'
0/
#954810000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#954820000000
0!
0'
0/
#954830000000
1!
1'
1/
#954840000000
0!
0'
0/
#954850000000
1!
1'
1/
#954860000000
0!
0'
0/
#954870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#954880000000
0!
0'
0/
#954890000000
1!
1'
1/
#954900000000
0!
0'
0/
#954910000000
1!
1'
1/
#954920000000
0!
0'
0/
#954930000000
1!
1'
1/
#954940000000
0!
0'
0/
#954950000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#954960000000
0!
0'
0/
#954970000000
1!
1'
1/
#954980000000
0!
0'
0/
#954990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#955000000000
0!
0'
0/
#955010000000
1!
1'
1/
#955020000000
0!
0'
0/
#955030000000
#955040000000
1!
1'
1/
#955050000000
0!
0'
0/
#955060000000
1!
1'
1/
#955070000000
0!
1"
0'
1(
0/
10
#955080000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#955090000000
0!
0'
0/
#955100000000
1!
1'
1/
#955110000000
0!
0'
0/
#955120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#955130000000
0!
0'
0/
#955140000000
1!
1'
1/
#955150000000
0!
1"
0'
1(
0/
10
#955160000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#955170000000
0!
1$
0'
1+
0/
#955180000000
1!
1'
1/
#955190000000
0!
0'
0/
#955200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#955210000000
0!
0'
0/
#955220000000
1!
1'
1/
#955230000000
0!
0'
0/
#955240000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#955250000000
0!
0'
0/
#955260000000
1!
1'
1/
#955270000000
0!
0'
0/
#955280000000
1!
1'
1/
#955290000000
0!
0'
0/
#955300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#955310000000
0!
0'
0/
#955320000000
1!
1'
1/
#955330000000
0!
0'
0/
#955340000000
1!
1'
1/
#955350000000
0!
0'
0/
#955360000000
1!
1'
1/
#955370000000
0!
0'
0/
#955380000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#955390000000
0!
0'
0/
#955400000000
1!
1'
1/
#955410000000
0!
0'
0/
#955420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#955430000000
0!
0'
0/
#955440000000
1!
1'
1/
#955450000000
0!
0'
0/
#955460000000
#955470000000
1!
1'
1/
#955480000000
0!
0'
0/
#955490000000
1!
1'
1/
#955500000000
0!
1"
0'
1(
0/
10
#955510000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#955520000000
0!
0'
0/
#955530000000
1!
1'
1/
#955540000000
0!
0'
0/
#955550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#955560000000
0!
0'
0/
#955570000000
1!
1'
1/
#955580000000
0!
1"
0'
1(
0/
10
#955590000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#955600000000
0!
1$
0'
1+
0/
#955610000000
1!
1'
1/
#955620000000
0!
0'
0/
#955630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#955640000000
0!
0'
0/
#955650000000
1!
1'
1/
#955660000000
0!
0'
0/
#955670000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#955680000000
0!
0'
0/
#955690000000
1!
1'
1/
#955700000000
0!
0'
0/
#955710000000
1!
1'
1/
#955720000000
0!
0'
0/
#955730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#955740000000
0!
0'
0/
#955750000000
1!
1'
1/
#955760000000
0!
0'
0/
#955770000000
1!
1'
1/
#955780000000
0!
0'
0/
#955790000000
1!
1'
1/
#955800000000
0!
0'
0/
#955810000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#955820000000
0!
0'
0/
#955830000000
1!
1'
1/
#955840000000
0!
0'
0/
#955850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#955860000000
0!
0'
0/
#955870000000
1!
1'
1/
#955880000000
0!
0'
0/
#955890000000
#955900000000
1!
1'
1/
#955910000000
0!
0'
0/
#955920000000
1!
1'
1/
#955930000000
0!
1"
0'
1(
0/
10
#955940000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#955950000000
0!
0'
0/
#955960000000
1!
1'
1/
#955970000000
0!
0'
0/
#955980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#955990000000
0!
0'
0/
#956000000000
1!
1'
1/
#956010000000
0!
1"
0'
1(
0/
10
#956020000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#956030000000
0!
1$
0'
1+
0/
#956040000000
1!
1'
1/
#956050000000
0!
0'
0/
#956060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#956070000000
0!
0'
0/
#956080000000
1!
1'
1/
#956090000000
0!
0'
0/
#956100000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#956110000000
0!
0'
0/
#956120000000
1!
1'
1/
#956130000000
0!
0'
0/
#956140000000
1!
1'
1/
#956150000000
0!
0'
0/
#956160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#956170000000
0!
0'
0/
#956180000000
1!
1'
1/
#956190000000
0!
0'
0/
#956200000000
1!
1'
1/
#956210000000
0!
0'
0/
#956220000000
1!
1'
1/
#956230000000
0!
0'
0/
#956240000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#956250000000
0!
0'
0/
#956260000000
1!
1'
1/
#956270000000
0!
0'
0/
#956280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#956290000000
0!
0'
0/
#956300000000
1!
1'
1/
#956310000000
0!
0'
0/
#956320000000
#956330000000
1!
1'
1/
#956340000000
0!
0'
0/
#956350000000
1!
1'
1/
#956360000000
0!
1"
0'
1(
0/
10
#956370000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#956380000000
0!
0'
0/
#956390000000
1!
1'
1/
#956400000000
0!
0'
0/
#956410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#956420000000
0!
0'
0/
#956430000000
1!
1'
1/
#956440000000
0!
1"
0'
1(
0/
10
#956450000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#956460000000
0!
1$
0'
1+
0/
#956470000000
1!
1'
1/
#956480000000
0!
0'
0/
#956490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#956500000000
0!
0'
0/
#956510000000
1!
1'
1/
#956520000000
0!
0'
0/
#956530000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#956540000000
0!
0'
0/
#956550000000
1!
1'
1/
#956560000000
0!
0'
0/
#956570000000
1!
1'
1/
#956580000000
0!
0'
0/
#956590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#956600000000
0!
0'
0/
#956610000000
1!
1'
1/
#956620000000
0!
0'
0/
#956630000000
1!
1'
1/
#956640000000
0!
0'
0/
#956650000000
1!
1'
1/
#956660000000
0!
0'
0/
#956670000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#956680000000
0!
0'
0/
#956690000000
1!
1'
1/
#956700000000
0!
0'
0/
#956710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#956720000000
0!
0'
0/
#956730000000
1!
1'
1/
#956740000000
0!
0'
0/
#956750000000
#956760000000
1!
1'
1/
#956770000000
0!
0'
0/
#956780000000
1!
1'
1/
#956790000000
0!
1"
0'
1(
0/
10
#956800000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#956810000000
0!
0'
0/
#956820000000
1!
1'
1/
#956830000000
0!
0'
0/
#956840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#956850000000
0!
0'
0/
#956860000000
1!
1'
1/
#956870000000
0!
1"
0'
1(
0/
10
#956880000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#956890000000
0!
1$
0'
1+
0/
#956900000000
1!
1'
1/
#956910000000
0!
0'
0/
#956920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#956930000000
0!
0'
0/
#956940000000
1!
1'
1/
#956950000000
0!
0'
0/
#956960000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#956970000000
0!
0'
0/
#956980000000
1!
1'
1/
#956990000000
0!
0'
0/
#957000000000
1!
1'
1/
#957010000000
0!
0'
0/
#957020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#957030000000
0!
0'
0/
#957040000000
1!
1'
1/
#957050000000
0!
0'
0/
#957060000000
1!
1'
1/
#957070000000
0!
0'
0/
#957080000000
1!
1'
1/
#957090000000
0!
0'
0/
#957100000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#957110000000
0!
0'
0/
#957120000000
1!
1'
1/
#957130000000
0!
0'
0/
#957140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#957150000000
0!
0'
0/
#957160000000
1!
1'
1/
#957170000000
0!
0'
0/
#957180000000
#957190000000
1!
1'
1/
#957200000000
0!
0'
0/
#957210000000
1!
1'
1/
#957220000000
0!
1"
0'
1(
0/
10
#957230000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#957240000000
0!
0'
0/
#957250000000
1!
1'
1/
#957260000000
0!
0'
0/
#957270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#957280000000
0!
0'
0/
#957290000000
1!
1'
1/
#957300000000
0!
1"
0'
1(
0/
10
#957310000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#957320000000
0!
1$
0'
1+
0/
#957330000000
1!
1'
1/
#957340000000
0!
0'
0/
#957350000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#957360000000
0!
0'
0/
#957370000000
1!
1'
1/
#957380000000
0!
0'
0/
#957390000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#957400000000
0!
0'
0/
#957410000000
1!
1'
1/
#957420000000
0!
0'
0/
#957430000000
1!
1'
1/
#957440000000
0!
0'
0/
#957450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#957460000000
0!
0'
0/
#957470000000
1!
1'
1/
#957480000000
0!
0'
0/
#957490000000
1!
1'
1/
#957500000000
0!
0'
0/
#957510000000
1!
1'
1/
#957520000000
0!
0'
0/
#957530000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#957540000000
0!
0'
0/
#957550000000
1!
1'
1/
#957560000000
0!
0'
0/
#957570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#957580000000
0!
0'
0/
#957590000000
1!
1'
1/
#957600000000
0!
0'
0/
#957610000000
#957620000000
1!
1'
1/
#957630000000
0!
0'
0/
#957640000000
1!
1'
1/
#957650000000
0!
1"
0'
1(
0/
10
#957660000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#957670000000
0!
0'
0/
#957680000000
1!
1'
1/
#957690000000
0!
0'
0/
#957700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#957710000000
0!
0'
0/
#957720000000
1!
1'
1/
#957730000000
0!
1"
0'
1(
0/
10
#957740000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#957750000000
0!
1$
0'
1+
0/
#957760000000
1!
1'
1/
#957770000000
0!
0'
0/
#957780000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#957790000000
0!
0'
0/
#957800000000
1!
1'
1/
#957810000000
0!
0'
0/
#957820000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#957830000000
0!
0'
0/
#957840000000
1!
1'
1/
#957850000000
0!
0'
0/
#957860000000
1!
1'
1/
#957870000000
0!
0'
0/
#957880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#957890000000
0!
0'
0/
#957900000000
1!
1'
1/
#957910000000
0!
0'
0/
#957920000000
1!
1'
1/
#957930000000
0!
0'
0/
#957940000000
1!
1'
1/
#957950000000
0!
0'
0/
#957960000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#957970000000
0!
0'
0/
#957980000000
1!
1'
1/
#957990000000
0!
0'
0/
#958000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#958010000000
0!
0'
0/
#958020000000
1!
1'
1/
#958030000000
0!
0'
0/
#958040000000
#958050000000
1!
1'
1/
#958060000000
0!
0'
0/
#958070000000
1!
1'
1/
#958080000000
0!
1"
0'
1(
0/
10
#958090000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#958100000000
0!
0'
0/
#958110000000
1!
1'
1/
#958120000000
0!
0'
0/
#958130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#958140000000
0!
0'
0/
#958150000000
1!
1'
1/
#958160000000
0!
1"
0'
1(
0/
10
#958170000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#958180000000
0!
1$
0'
1+
0/
#958190000000
1!
1'
1/
#958200000000
0!
0'
0/
#958210000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#958220000000
0!
0'
0/
#958230000000
1!
1'
1/
#958240000000
0!
0'
0/
#958250000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#958260000000
0!
0'
0/
#958270000000
1!
1'
1/
#958280000000
0!
0'
0/
#958290000000
1!
1'
1/
#958300000000
0!
0'
0/
#958310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#958320000000
0!
0'
0/
#958330000000
1!
1'
1/
#958340000000
0!
0'
0/
#958350000000
1!
1'
1/
#958360000000
0!
0'
0/
#958370000000
1!
1'
1/
#958380000000
0!
0'
0/
#958390000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#958400000000
0!
0'
0/
#958410000000
1!
1'
1/
#958420000000
0!
0'
0/
#958430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#958440000000
0!
0'
0/
#958450000000
1!
1'
1/
#958460000000
0!
0'
0/
#958470000000
#958480000000
1!
1'
1/
#958490000000
0!
0'
0/
#958500000000
1!
1'
1/
#958510000000
0!
1"
0'
1(
0/
10
#958520000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#958530000000
0!
0'
0/
#958540000000
1!
1'
1/
#958550000000
0!
0'
0/
#958560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#958570000000
0!
0'
0/
#958580000000
1!
1'
1/
#958590000000
0!
1"
0'
1(
0/
10
#958600000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#958610000000
0!
1$
0'
1+
0/
#958620000000
1!
1'
1/
#958630000000
0!
0'
0/
#958640000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#958650000000
0!
0'
0/
#958660000000
1!
1'
1/
#958670000000
0!
0'
0/
#958680000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#958690000000
0!
0'
0/
#958700000000
1!
1'
1/
#958710000000
0!
0'
0/
#958720000000
1!
1'
1/
#958730000000
0!
0'
0/
#958740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#958750000000
0!
0'
0/
#958760000000
1!
1'
1/
#958770000000
0!
0'
0/
#958780000000
1!
1'
1/
#958790000000
0!
0'
0/
#958800000000
1!
1'
1/
#958810000000
0!
0'
0/
#958820000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#958830000000
0!
0'
0/
#958840000000
1!
1'
1/
#958850000000
0!
0'
0/
#958860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#958870000000
0!
0'
0/
#958880000000
1!
1'
1/
#958890000000
0!
0'
0/
#958900000000
#958910000000
1!
1'
1/
#958920000000
0!
0'
0/
#958930000000
1!
1'
1/
#958940000000
0!
1"
0'
1(
0/
10
#958950000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#958960000000
0!
0'
0/
#958970000000
1!
1'
1/
#958980000000
0!
0'
0/
#958990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#959000000000
0!
0'
0/
#959010000000
1!
1'
1/
#959020000000
0!
1"
0'
1(
0/
10
#959030000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#959040000000
0!
1$
0'
1+
0/
#959050000000
1!
1'
1/
#959060000000
0!
0'
0/
#959070000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#959080000000
0!
0'
0/
#959090000000
1!
1'
1/
#959100000000
0!
0'
0/
#959110000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#959120000000
0!
0'
0/
#959130000000
1!
1'
1/
#959140000000
0!
0'
0/
#959150000000
1!
1'
1/
#959160000000
0!
0'
0/
#959170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#959180000000
0!
0'
0/
#959190000000
1!
1'
1/
#959200000000
0!
0'
0/
#959210000000
1!
1'
1/
#959220000000
0!
0'
0/
#959230000000
1!
1'
1/
#959240000000
0!
0'
0/
#959250000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#959260000000
0!
0'
0/
#959270000000
1!
1'
1/
#959280000000
0!
0'
0/
#959290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#959300000000
0!
0'
0/
#959310000000
1!
1'
1/
#959320000000
0!
0'
0/
#959330000000
#959340000000
1!
1'
1/
#959350000000
0!
0'
0/
#959360000000
1!
1'
1/
#959370000000
0!
1"
0'
1(
0/
10
#959380000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#959390000000
0!
0'
0/
#959400000000
1!
1'
1/
#959410000000
0!
0'
0/
#959420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#959430000000
0!
0'
0/
#959440000000
1!
1'
1/
#959450000000
0!
1"
0'
1(
0/
10
#959460000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#959470000000
0!
1$
0'
1+
0/
#959480000000
1!
1'
1/
#959490000000
0!
0'
0/
#959500000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#959510000000
0!
0'
0/
#959520000000
1!
1'
1/
#959530000000
0!
0'
0/
#959540000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#959550000000
0!
0'
0/
#959560000000
1!
1'
1/
#959570000000
0!
0'
0/
#959580000000
1!
1'
1/
#959590000000
0!
0'
0/
#959600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#959610000000
0!
0'
0/
#959620000000
1!
1'
1/
#959630000000
0!
0'
0/
#959640000000
1!
1'
1/
#959650000000
0!
0'
0/
#959660000000
1!
1'
1/
#959670000000
0!
0'
0/
#959680000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#959690000000
0!
0'
0/
#959700000000
1!
1'
1/
#959710000000
0!
0'
0/
#959720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#959730000000
0!
0'
0/
#959740000000
1!
1'
1/
#959750000000
0!
0'
0/
#959760000000
#959770000000
1!
1'
1/
#959780000000
0!
0'
0/
#959790000000
1!
1'
1/
#959800000000
0!
1"
0'
1(
0/
10
#959810000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#959820000000
0!
0'
0/
#959830000000
1!
1'
1/
#959840000000
0!
0'
0/
#959850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#959860000000
0!
0'
0/
#959870000000
1!
1'
1/
#959880000000
0!
1"
0'
1(
0/
10
#959890000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#959900000000
0!
1$
0'
1+
0/
#959910000000
1!
1'
1/
#959920000000
0!
0'
0/
#959930000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#959940000000
0!
0'
0/
#959950000000
1!
1'
1/
#959960000000
0!
0'
0/
#959970000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#959980000000
0!
0'
0/
#959990000000
1!
1'
1/
#960000000000
0!
0'
0/
#960010000000
1!
1'
1/
#960020000000
0!
0'
0/
#960030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#960040000000
0!
0'
0/
#960050000000
1!
1'
1/
#960060000000
0!
0'
0/
#960070000000
1!
1'
1/
#960080000000
0!
0'
0/
#960090000000
1!
1'
1/
#960100000000
0!
0'
0/
#960110000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#960120000000
0!
0'
0/
#960130000000
1!
1'
1/
#960140000000
0!
0'
0/
#960150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#960160000000
0!
0'
0/
#960170000000
1!
1'
1/
#960180000000
0!
0'
0/
#960190000000
#960200000000
1!
1'
1/
#960210000000
0!
0'
0/
#960220000000
1!
1'
1/
#960230000000
0!
1"
0'
1(
0/
10
#960240000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#960250000000
0!
0'
0/
#960260000000
1!
1'
1/
#960270000000
0!
0'
0/
#960280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#960290000000
0!
0'
0/
#960300000000
1!
1'
1/
#960310000000
0!
1"
0'
1(
0/
10
#960320000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#960330000000
0!
1$
0'
1+
0/
#960340000000
1!
1'
1/
#960350000000
0!
0'
0/
#960360000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#960370000000
0!
0'
0/
#960380000000
1!
1'
1/
#960390000000
0!
0'
0/
#960400000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#960410000000
0!
0'
0/
#960420000000
1!
1'
1/
#960430000000
0!
0'
0/
#960440000000
1!
1'
1/
#960450000000
0!
0'
0/
#960460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#960470000000
0!
0'
0/
#960480000000
1!
1'
1/
#960490000000
0!
0'
0/
#960500000000
1!
1'
1/
#960510000000
0!
0'
0/
#960520000000
1!
1'
1/
#960530000000
0!
0'
0/
#960540000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#960550000000
0!
0'
0/
#960560000000
1!
1'
1/
#960570000000
0!
0'
0/
#960580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#960590000000
0!
0'
0/
#960600000000
1!
1'
1/
#960610000000
0!
0'
0/
#960620000000
#960630000000
1!
1'
1/
#960640000000
0!
0'
0/
#960650000000
1!
1'
1/
#960660000000
0!
1"
0'
1(
0/
10
#960670000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#960680000000
0!
0'
0/
#960690000000
1!
1'
1/
#960700000000
0!
0'
0/
#960710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#960720000000
0!
0'
0/
#960730000000
1!
1'
1/
#960740000000
0!
1"
0'
1(
0/
10
#960750000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#960760000000
0!
1$
0'
1+
0/
#960770000000
1!
1'
1/
#960780000000
0!
0'
0/
#960790000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#960800000000
0!
0'
0/
#960810000000
1!
1'
1/
#960820000000
0!
0'
0/
#960830000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#960840000000
0!
0'
0/
#960850000000
1!
1'
1/
#960860000000
0!
0'
0/
#960870000000
1!
1'
1/
#960880000000
0!
0'
0/
#960890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#960900000000
0!
0'
0/
#960910000000
1!
1'
1/
#960920000000
0!
0'
0/
#960930000000
1!
1'
1/
#960940000000
0!
0'
0/
#960950000000
1!
1'
1/
#960960000000
0!
0'
0/
#960970000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#960980000000
0!
0'
0/
#960990000000
1!
1'
1/
#961000000000
0!
0'
0/
#961010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#961020000000
0!
0'
0/
#961030000000
1!
1'
1/
#961040000000
0!
0'
0/
#961050000000
#961060000000
1!
1'
1/
#961070000000
0!
0'
0/
#961080000000
1!
1'
1/
#961090000000
0!
1"
0'
1(
0/
10
#961100000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#961110000000
0!
0'
0/
#961120000000
1!
1'
1/
#961130000000
0!
0'
0/
#961140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#961150000000
0!
0'
0/
#961160000000
1!
1'
1/
#961170000000
0!
1"
0'
1(
0/
10
#961180000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#961190000000
0!
1$
0'
1+
0/
#961200000000
1!
1'
1/
#961210000000
0!
0'
0/
#961220000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#961230000000
0!
0'
0/
#961240000000
1!
1'
1/
#961250000000
0!
0'
0/
#961260000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#961270000000
0!
0'
0/
#961280000000
1!
1'
1/
#961290000000
0!
0'
0/
#961300000000
1!
1'
1/
#961310000000
0!
0'
0/
#961320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#961330000000
0!
0'
0/
#961340000000
1!
1'
1/
#961350000000
0!
0'
0/
#961360000000
1!
1'
1/
#961370000000
0!
0'
0/
#961380000000
1!
1'
1/
#961390000000
0!
0'
0/
#961400000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#961410000000
0!
0'
0/
#961420000000
1!
1'
1/
#961430000000
0!
0'
0/
#961440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#961450000000
0!
0'
0/
#961460000000
1!
1'
1/
#961470000000
0!
0'
0/
#961480000000
#961490000000
1!
1'
1/
#961500000000
0!
0'
0/
#961510000000
1!
1'
1/
#961520000000
0!
1"
0'
1(
0/
10
#961530000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#961540000000
0!
0'
0/
#961550000000
1!
1'
1/
#961560000000
0!
0'
0/
#961570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#961580000000
0!
0'
0/
#961590000000
1!
1'
1/
#961600000000
0!
1"
0'
1(
0/
10
#961610000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#961620000000
0!
1$
0'
1+
0/
#961630000000
1!
1'
1/
#961640000000
0!
0'
0/
#961650000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#961660000000
0!
0'
0/
#961670000000
1!
1'
1/
#961680000000
0!
0'
0/
#961690000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#961700000000
0!
0'
0/
#961710000000
1!
1'
1/
#961720000000
0!
0'
0/
#961730000000
1!
1'
1/
#961740000000
0!
0'
0/
#961750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#961760000000
0!
0'
0/
#961770000000
1!
1'
1/
#961780000000
0!
0'
0/
#961790000000
1!
1'
1/
#961800000000
0!
0'
0/
#961810000000
1!
1'
1/
#961820000000
0!
0'
0/
#961830000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#961840000000
0!
0'
0/
#961850000000
1!
1'
1/
#961860000000
0!
0'
0/
#961870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#961880000000
0!
0'
0/
#961890000000
1!
1'
1/
#961900000000
0!
0'
0/
#961910000000
#961920000000
1!
1'
1/
#961930000000
0!
0'
0/
#961940000000
1!
1'
1/
#961950000000
0!
1"
0'
1(
0/
10
#961960000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#961970000000
0!
0'
0/
#961980000000
1!
1'
1/
#961990000000
0!
0'
0/
#962000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#962010000000
0!
0'
0/
#962020000000
1!
1'
1/
#962030000000
0!
1"
0'
1(
0/
10
#962040000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#962050000000
0!
1$
0'
1+
0/
#962060000000
1!
1'
1/
#962070000000
0!
0'
0/
#962080000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#962090000000
0!
0'
0/
#962100000000
1!
1'
1/
#962110000000
0!
0'
0/
#962120000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#962130000000
0!
0'
0/
#962140000000
1!
1'
1/
#962150000000
0!
0'
0/
#962160000000
1!
1'
1/
#962170000000
0!
0'
0/
#962180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#962190000000
0!
0'
0/
#962200000000
1!
1'
1/
#962210000000
0!
0'
0/
#962220000000
1!
1'
1/
#962230000000
0!
0'
0/
#962240000000
1!
1'
1/
#962250000000
0!
0'
0/
#962260000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#962270000000
0!
0'
0/
#962280000000
1!
1'
1/
#962290000000
0!
0'
0/
#962300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#962310000000
0!
0'
0/
#962320000000
1!
1'
1/
#962330000000
0!
0'
0/
#962340000000
#962350000000
1!
1'
1/
#962360000000
0!
0'
0/
#962370000000
1!
1'
1/
#962380000000
0!
1"
0'
1(
0/
10
#962390000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#962400000000
0!
0'
0/
#962410000000
1!
1'
1/
#962420000000
0!
0'
0/
#962430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#962440000000
0!
0'
0/
#962450000000
1!
1'
1/
#962460000000
0!
1"
0'
1(
0/
10
#962470000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#962480000000
0!
1$
0'
1+
0/
#962490000000
1!
1'
1/
#962500000000
0!
0'
0/
#962510000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#962520000000
0!
0'
0/
#962530000000
1!
1'
1/
#962540000000
0!
0'
0/
#962550000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#962560000000
0!
0'
0/
#962570000000
1!
1'
1/
#962580000000
0!
0'
0/
#962590000000
1!
1'
1/
#962600000000
0!
0'
0/
#962610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#962620000000
0!
0'
0/
#962630000000
1!
1'
1/
#962640000000
0!
0'
0/
#962650000000
1!
1'
1/
#962660000000
0!
0'
0/
#962670000000
1!
1'
1/
#962680000000
0!
0'
0/
#962690000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#962700000000
0!
0'
0/
#962710000000
1!
1'
1/
#962720000000
0!
0'
0/
#962730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#962740000000
0!
0'
0/
#962750000000
1!
1'
1/
#962760000000
0!
0'
0/
#962770000000
#962780000000
1!
1'
1/
#962790000000
0!
0'
0/
#962800000000
1!
1'
1/
#962810000000
0!
1"
0'
1(
0/
10
#962820000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#962830000000
0!
0'
0/
#962840000000
1!
1'
1/
#962850000000
0!
0'
0/
#962860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#962870000000
0!
0'
0/
#962880000000
1!
1'
1/
#962890000000
0!
1"
0'
1(
0/
10
#962900000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#962910000000
0!
1$
0'
1+
0/
#962920000000
1!
1'
1/
#962930000000
0!
0'
0/
#962940000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#962950000000
0!
0'
0/
#962960000000
1!
1'
1/
#962970000000
0!
0'
0/
#962980000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#962990000000
0!
0'
0/
#963000000000
1!
1'
1/
#963010000000
0!
0'
0/
#963020000000
1!
1'
1/
#963030000000
0!
0'
0/
#963040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#963050000000
0!
0'
0/
#963060000000
1!
1'
1/
#963070000000
0!
0'
0/
#963080000000
1!
1'
1/
#963090000000
0!
0'
0/
#963100000000
1!
1'
1/
#963110000000
0!
0'
0/
#963120000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#963130000000
0!
0'
0/
#963140000000
1!
1'
1/
#963150000000
0!
0'
0/
#963160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#963170000000
0!
0'
0/
#963180000000
1!
1'
1/
#963190000000
0!
0'
0/
#963200000000
#963210000000
1!
1'
1/
#963220000000
0!
0'
0/
#963230000000
1!
1'
1/
#963240000000
0!
1"
0'
1(
0/
10
#963250000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#963260000000
0!
0'
0/
#963270000000
1!
1'
1/
#963280000000
0!
0'
0/
#963290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#963300000000
0!
0'
0/
#963310000000
1!
1'
1/
#963320000000
0!
1"
0'
1(
0/
10
#963330000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#963340000000
0!
1$
0'
1+
0/
#963350000000
1!
1'
1/
#963360000000
0!
0'
0/
#963370000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#963380000000
0!
0'
0/
#963390000000
1!
1'
1/
#963400000000
0!
0'
0/
#963410000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#963420000000
0!
0'
0/
#963430000000
1!
1'
1/
#963440000000
0!
0'
0/
#963450000000
1!
1'
1/
#963460000000
0!
0'
0/
#963470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#963480000000
0!
0'
0/
#963490000000
1!
1'
1/
#963500000000
0!
0'
0/
#963510000000
1!
1'
1/
#963520000000
0!
0'
0/
#963530000000
1!
1'
1/
#963540000000
0!
0'
0/
#963550000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#963560000000
0!
0'
0/
#963570000000
1!
1'
1/
#963580000000
0!
0'
0/
#963590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#963600000000
0!
0'
0/
#963610000000
1!
1'
1/
#963620000000
0!
0'
0/
#963630000000
#963640000000
1!
1'
1/
#963650000000
0!
0'
0/
#963660000000
1!
1'
1/
#963670000000
0!
1"
0'
1(
0/
10
#963680000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#963690000000
0!
0'
0/
#963700000000
1!
1'
1/
#963710000000
0!
0'
0/
#963720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#963730000000
0!
0'
0/
#963740000000
1!
1'
1/
#963750000000
0!
1"
0'
1(
0/
10
#963760000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#963770000000
0!
1$
0'
1+
0/
#963780000000
1!
1'
1/
#963790000000
0!
0'
0/
#963800000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#963810000000
0!
0'
0/
#963820000000
1!
1'
1/
#963830000000
0!
0'
0/
#963840000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#963850000000
0!
0'
0/
#963860000000
1!
1'
1/
#963870000000
0!
0'
0/
#963880000000
1!
1'
1/
#963890000000
0!
0'
0/
#963900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#963910000000
0!
0'
0/
#963920000000
1!
1'
1/
#963930000000
0!
0'
0/
#963940000000
1!
1'
1/
#963950000000
0!
0'
0/
#963960000000
1!
1'
1/
#963970000000
0!
0'
0/
#963980000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#963990000000
0!
0'
0/
#964000000000
1!
1'
1/
#964010000000
0!
0'
0/
#964020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#964030000000
0!
0'
0/
#964040000000
1!
1'
1/
#964050000000
0!
0'
0/
#964060000000
#964070000000
1!
1'
1/
#964080000000
0!
0'
0/
#964090000000
1!
1'
1/
#964100000000
0!
1"
0'
1(
0/
10
#964110000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#964120000000
0!
0'
0/
#964130000000
1!
1'
1/
#964140000000
0!
0'
0/
#964150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#964160000000
0!
0'
0/
#964170000000
1!
1'
1/
#964180000000
0!
1"
0'
1(
0/
10
#964190000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#964200000000
0!
1$
0'
1+
0/
#964210000000
1!
1'
1/
#964220000000
0!
0'
0/
#964230000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#964240000000
0!
0'
0/
#964250000000
1!
1'
1/
#964260000000
0!
0'
0/
#964270000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#964280000000
0!
0'
0/
#964290000000
1!
1'
1/
#964300000000
0!
0'
0/
#964310000000
1!
1'
1/
#964320000000
0!
0'
0/
#964330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#964340000000
0!
0'
0/
#964350000000
1!
1'
1/
#964360000000
0!
0'
0/
#964370000000
1!
1'
1/
#964380000000
0!
0'
0/
#964390000000
1!
1'
1/
#964400000000
0!
0'
0/
#964410000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#964420000000
0!
0'
0/
#964430000000
1!
1'
1/
#964440000000
0!
0'
0/
#964450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#964460000000
0!
0'
0/
#964470000000
1!
1'
1/
#964480000000
0!
0'
0/
#964490000000
#964500000000
1!
1'
1/
#964510000000
0!
0'
0/
#964520000000
1!
1'
1/
#964530000000
0!
1"
0'
1(
0/
10
#964540000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#964550000000
0!
0'
0/
#964560000000
1!
1'
1/
#964570000000
0!
0'
0/
#964580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#964590000000
0!
0'
0/
#964600000000
1!
1'
1/
#964610000000
0!
1"
0'
1(
0/
10
#964620000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#964630000000
0!
1$
0'
1+
0/
#964640000000
1!
1'
1/
#964650000000
0!
0'
0/
#964660000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#964670000000
0!
0'
0/
#964680000000
1!
1'
1/
#964690000000
0!
0'
0/
#964700000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#964710000000
0!
0'
0/
#964720000000
1!
1'
1/
#964730000000
0!
0'
0/
#964740000000
1!
1'
1/
#964750000000
0!
0'
0/
#964760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#964770000000
0!
0'
0/
#964780000000
1!
1'
1/
#964790000000
0!
0'
0/
#964800000000
1!
1'
1/
#964810000000
0!
0'
0/
#964820000000
1!
1'
1/
#964830000000
0!
0'
0/
#964840000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#964850000000
0!
0'
0/
#964860000000
1!
1'
1/
#964870000000
0!
0'
0/
#964880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#964890000000
0!
0'
0/
#964900000000
1!
1'
1/
#964910000000
0!
0'
0/
#964920000000
#964930000000
1!
1'
1/
#964940000000
0!
0'
0/
#964950000000
1!
1'
1/
#964960000000
0!
1"
0'
1(
0/
10
#964970000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#964980000000
0!
0'
0/
#964990000000
1!
1'
1/
#965000000000
0!
0'
0/
#965010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#965020000000
0!
0'
0/
#965030000000
1!
1'
1/
#965040000000
0!
1"
0'
1(
0/
10
#965050000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#965060000000
0!
1$
0'
1+
0/
#965070000000
1!
1'
1/
#965080000000
0!
0'
0/
#965090000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#965100000000
0!
0'
0/
#965110000000
1!
1'
1/
#965120000000
0!
0'
0/
#965130000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#965140000000
0!
0'
0/
#965150000000
1!
1'
1/
#965160000000
0!
0'
0/
#965170000000
1!
1'
1/
#965180000000
0!
0'
0/
#965190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#965200000000
0!
0'
0/
#965210000000
1!
1'
1/
#965220000000
0!
0'
0/
#965230000000
1!
1'
1/
#965240000000
0!
0'
0/
#965250000000
1!
1'
1/
#965260000000
0!
0'
0/
#965270000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#965280000000
0!
0'
0/
#965290000000
1!
1'
1/
#965300000000
0!
0'
0/
#965310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#965320000000
0!
0'
0/
#965330000000
1!
1'
1/
#965340000000
0!
0'
0/
#965350000000
#965360000000
1!
1'
1/
#965370000000
0!
0'
0/
#965380000000
1!
1'
1/
#965390000000
0!
1"
0'
1(
0/
10
#965400000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#965410000000
0!
0'
0/
#965420000000
1!
1'
1/
#965430000000
0!
0'
0/
#965440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#965450000000
0!
0'
0/
#965460000000
1!
1'
1/
#965470000000
0!
1"
0'
1(
0/
10
#965480000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#965490000000
0!
1$
0'
1+
0/
#965500000000
1!
1'
1/
#965510000000
0!
0'
0/
#965520000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#965530000000
0!
0'
0/
#965540000000
1!
1'
1/
#965550000000
0!
0'
0/
#965560000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#965570000000
0!
0'
0/
#965580000000
1!
1'
1/
#965590000000
0!
0'
0/
#965600000000
1!
1'
1/
#965610000000
0!
0'
0/
#965620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#965630000000
0!
0'
0/
#965640000000
1!
1'
1/
#965650000000
0!
0'
0/
#965660000000
1!
1'
1/
#965670000000
0!
0'
0/
#965680000000
1!
1'
1/
#965690000000
0!
0'
0/
#965700000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#965710000000
0!
0'
0/
#965720000000
1!
1'
1/
#965730000000
0!
0'
0/
#965740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#965750000000
0!
0'
0/
#965760000000
1!
1'
1/
#965770000000
0!
0'
0/
#965780000000
#965790000000
1!
1'
1/
#965800000000
0!
0'
0/
#965810000000
1!
1'
1/
#965820000000
0!
1"
0'
1(
0/
10
#965830000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#965840000000
0!
0'
0/
#965850000000
1!
1'
1/
#965860000000
0!
0'
0/
#965870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#965880000000
0!
0'
0/
#965890000000
1!
1'
1/
#965900000000
0!
1"
0'
1(
0/
10
#965910000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#965920000000
0!
1$
0'
1+
0/
#965930000000
1!
1'
1/
#965940000000
0!
0'
0/
#965950000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#965960000000
0!
0'
0/
#965970000000
1!
1'
1/
#965980000000
0!
0'
0/
#965990000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#966000000000
0!
0'
0/
#966010000000
1!
1'
1/
#966020000000
0!
0'
0/
#966030000000
1!
1'
1/
#966040000000
0!
0'
0/
#966050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#966060000000
0!
0'
0/
#966070000000
1!
1'
1/
#966080000000
0!
0'
0/
#966090000000
1!
1'
1/
#966100000000
0!
0'
0/
#966110000000
1!
1'
1/
#966120000000
0!
0'
0/
#966130000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#966140000000
0!
0'
0/
#966150000000
1!
1'
1/
#966160000000
0!
0'
0/
#966170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#966180000000
0!
0'
0/
#966190000000
1!
1'
1/
#966200000000
0!
0'
0/
#966210000000
#966220000000
1!
1'
1/
#966230000000
0!
0'
0/
#966240000000
1!
1'
1/
#966250000000
0!
1"
0'
1(
0/
10
#966260000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#966270000000
0!
0'
0/
#966280000000
1!
1'
1/
#966290000000
0!
0'
0/
#966300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#966310000000
0!
0'
0/
#966320000000
1!
1'
1/
#966330000000
0!
1"
0'
1(
0/
10
#966340000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#966350000000
0!
1$
0'
1+
0/
#966360000000
1!
1'
1/
#966370000000
0!
0'
0/
#966380000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#966390000000
0!
0'
0/
#966400000000
1!
1'
1/
#966410000000
0!
0'
0/
#966420000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#966430000000
0!
0'
0/
#966440000000
1!
1'
1/
#966450000000
0!
0'
0/
#966460000000
1!
1'
1/
#966470000000
0!
0'
0/
#966480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#966490000000
0!
0'
0/
#966500000000
1!
1'
1/
#966510000000
0!
0'
0/
#966520000000
1!
1'
1/
#966530000000
0!
0'
0/
#966540000000
1!
1'
1/
#966550000000
0!
0'
0/
#966560000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#966570000000
0!
0'
0/
#966580000000
1!
1'
1/
#966590000000
0!
0'
0/
#966600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#966610000000
0!
0'
0/
#966620000000
1!
1'
1/
#966630000000
0!
0'
0/
#966640000000
#966650000000
1!
1'
1/
#966660000000
0!
0'
0/
#966670000000
1!
1'
1/
#966680000000
0!
1"
0'
1(
0/
10
#966690000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#966700000000
0!
0'
0/
#966710000000
1!
1'
1/
#966720000000
0!
0'
0/
#966730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#966740000000
0!
0'
0/
#966750000000
1!
1'
1/
#966760000000
0!
1"
0'
1(
0/
10
#966770000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#966780000000
0!
1$
0'
1+
0/
#966790000000
1!
1'
1/
#966800000000
0!
0'
0/
#966810000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#966820000000
0!
0'
0/
#966830000000
1!
1'
1/
#966840000000
0!
0'
0/
#966850000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#966860000000
0!
0'
0/
#966870000000
1!
1'
1/
#966880000000
0!
0'
0/
#966890000000
1!
1'
1/
#966900000000
0!
0'
0/
#966910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#966920000000
0!
0'
0/
#966930000000
1!
1'
1/
#966940000000
0!
0'
0/
#966950000000
1!
1'
1/
#966960000000
0!
0'
0/
#966970000000
1!
1'
1/
#966980000000
0!
0'
0/
#966990000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#967000000000
0!
0'
0/
#967010000000
1!
1'
1/
#967020000000
0!
0'
0/
#967030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#967040000000
0!
0'
0/
#967050000000
1!
1'
1/
#967060000000
0!
0'
0/
#967070000000
#967080000000
1!
1'
1/
#967090000000
0!
0'
0/
#967100000000
1!
1'
1/
#967110000000
0!
1"
0'
1(
0/
10
#967120000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#967130000000
0!
0'
0/
#967140000000
1!
1'
1/
#967150000000
0!
0'
0/
#967160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#967170000000
0!
0'
0/
#967180000000
1!
1'
1/
#967190000000
0!
1"
0'
1(
0/
10
#967200000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#967210000000
0!
1$
0'
1+
0/
#967220000000
1!
1'
1/
#967230000000
0!
0'
0/
#967240000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#967250000000
0!
0'
0/
#967260000000
1!
1'
1/
#967270000000
0!
0'
0/
#967280000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#967290000000
0!
0'
0/
#967300000000
1!
1'
1/
#967310000000
0!
0'
0/
#967320000000
1!
1'
1/
#967330000000
0!
0'
0/
#967340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#967350000000
0!
0'
0/
#967360000000
1!
1'
1/
#967370000000
0!
0'
0/
#967380000000
1!
1'
1/
#967390000000
0!
0'
0/
#967400000000
1!
1'
1/
#967410000000
0!
0'
0/
#967420000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#967430000000
0!
0'
0/
#967440000000
1!
1'
1/
#967450000000
0!
0'
0/
#967460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#967470000000
0!
0'
0/
#967480000000
1!
1'
1/
#967490000000
0!
0'
0/
#967500000000
#967510000000
1!
1'
1/
#967520000000
0!
0'
0/
#967530000000
1!
1'
1/
#967540000000
0!
1"
0'
1(
0/
10
#967550000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#967560000000
0!
0'
0/
#967570000000
1!
1'
1/
#967580000000
0!
0'
0/
#967590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#967600000000
0!
0'
0/
#967610000000
1!
1'
1/
#967620000000
0!
1"
0'
1(
0/
10
#967630000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#967640000000
0!
1$
0'
1+
0/
#967650000000
1!
1'
1/
#967660000000
0!
0'
0/
#967670000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#967680000000
0!
0'
0/
#967690000000
1!
1'
1/
#967700000000
0!
0'
0/
#967710000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#967720000000
0!
0'
0/
#967730000000
1!
1'
1/
#967740000000
0!
0'
0/
#967750000000
1!
1'
1/
#967760000000
0!
0'
0/
#967770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#967780000000
0!
0'
0/
#967790000000
1!
1'
1/
#967800000000
0!
0'
0/
#967810000000
1!
1'
1/
#967820000000
0!
0'
0/
#967830000000
1!
1'
1/
#967840000000
0!
0'
0/
#967850000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#967860000000
0!
0'
0/
#967870000000
1!
1'
1/
#967880000000
0!
0'
0/
#967890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#967900000000
0!
0'
0/
#967910000000
1!
1'
1/
#967920000000
0!
0'
0/
#967930000000
#967940000000
1!
1'
1/
#967950000000
0!
0'
0/
#967960000000
1!
1'
1/
#967970000000
0!
1"
0'
1(
0/
10
#967980000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#967990000000
0!
0'
0/
#968000000000
1!
1'
1/
#968010000000
0!
0'
0/
#968020000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#968030000000
0!
0'
0/
#968040000000
1!
1'
1/
#968050000000
0!
1"
0'
1(
0/
10
#968060000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#968070000000
0!
1$
0'
1+
0/
#968080000000
1!
1'
1/
#968090000000
0!
0'
0/
#968100000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#968110000000
0!
0'
0/
#968120000000
1!
1'
1/
#968130000000
0!
0'
0/
#968140000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#968150000000
0!
0'
0/
#968160000000
1!
1'
1/
#968170000000
0!
0'
0/
#968180000000
1!
1'
1/
#968190000000
0!
0'
0/
#968200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#968210000000
0!
0'
0/
#968220000000
1!
1'
1/
#968230000000
0!
0'
0/
#968240000000
1!
1'
1/
#968250000000
0!
0'
0/
#968260000000
1!
1'
1/
#968270000000
0!
0'
0/
#968280000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#968290000000
0!
0'
0/
#968300000000
1!
1'
1/
#968310000000
0!
0'
0/
#968320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#968330000000
0!
0'
0/
#968340000000
1!
1'
1/
#968350000000
0!
0'
0/
#968360000000
#968370000000
1!
1'
1/
#968380000000
0!
0'
0/
#968390000000
1!
1'
1/
#968400000000
0!
1"
0'
1(
0/
10
#968410000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#968420000000
0!
0'
0/
#968430000000
1!
1'
1/
#968440000000
0!
0'
0/
#968450000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#968460000000
0!
0'
0/
#968470000000
1!
1'
1/
#968480000000
0!
1"
0'
1(
0/
10
#968490000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#968500000000
0!
1$
0'
1+
0/
#968510000000
1!
1'
1/
#968520000000
0!
0'
0/
#968530000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#968540000000
0!
0'
0/
#968550000000
1!
1'
1/
#968560000000
0!
0'
0/
#968570000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#968580000000
0!
0'
0/
#968590000000
1!
1'
1/
#968600000000
0!
0'
0/
#968610000000
1!
1'
1/
#968620000000
0!
0'
0/
#968630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#968640000000
0!
0'
0/
#968650000000
1!
1'
1/
#968660000000
0!
0'
0/
#968670000000
1!
1'
1/
#968680000000
0!
0'
0/
#968690000000
1!
1'
1/
#968700000000
0!
0'
0/
#968710000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#968720000000
0!
0'
0/
#968730000000
1!
1'
1/
#968740000000
0!
0'
0/
#968750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#968760000000
0!
0'
0/
#968770000000
1!
1'
1/
#968780000000
0!
0'
0/
#968790000000
#968800000000
1!
1'
1/
#968810000000
0!
0'
0/
#968820000000
1!
1'
1/
#968830000000
0!
1"
0'
1(
0/
10
#968840000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#968850000000
0!
0'
0/
#968860000000
1!
1'
1/
#968870000000
0!
0'
0/
#968880000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#968890000000
0!
0'
0/
#968900000000
1!
1'
1/
#968910000000
0!
1"
0'
1(
0/
10
#968920000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#968930000000
0!
1$
0'
1+
0/
#968940000000
1!
1'
1/
#968950000000
0!
0'
0/
#968960000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#968970000000
0!
0'
0/
#968980000000
1!
1'
1/
#968990000000
0!
0'
0/
#969000000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#969010000000
0!
0'
0/
#969020000000
1!
1'
1/
#969030000000
0!
0'
0/
#969040000000
1!
1'
1/
#969050000000
0!
0'
0/
#969060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#969070000000
0!
0'
0/
#969080000000
1!
1'
1/
#969090000000
0!
0'
0/
#969100000000
1!
1'
1/
#969110000000
0!
0'
0/
#969120000000
1!
1'
1/
#969130000000
0!
0'
0/
#969140000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#969150000000
0!
0'
0/
#969160000000
1!
1'
1/
#969170000000
0!
0'
0/
#969180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#969190000000
0!
0'
0/
#969200000000
1!
1'
1/
#969210000000
0!
0'
0/
#969220000000
#969230000000
1!
1'
1/
#969240000000
0!
0'
0/
#969250000000
1!
1'
1/
#969260000000
0!
1"
0'
1(
0/
10
#969270000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#969280000000
0!
0'
0/
#969290000000
1!
1'
1/
#969300000000
0!
0'
0/
#969310000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#969320000000
0!
0'
0/
#969330000000
1!
1'
1/
#969340000000
0!
1"
0'
1(
0/
10
#969350000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#969360000000
0!
1$
0'
1+
0/
#969370000000
1!
1'
1/
#969380000000
0!
0'
0/
#969390000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#969400000000
0!
0'
0/
#969410000000
1!
1'
1/
#969420000000
0!
0'
0/
#969430000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#969440000000
0!
0'
0/
#969450000000
1!
1'
1/
#969460000000
0!
0'
0/
#969470000000
1!
1'
1/
#969480000000
0!
0'
0/
#969490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#969500000000
0!
0'
0/
#969510000000
1!
1'
1/
#969520000000
0!
0'
0/
#969530000000
1!
1'
1/
#969540000000
0!
0'
0/
#969550000000
1!
1'
1/
#969560000000
0!
0'
0/
#969570000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#969580000000
0!
0'
0/
#969590000000
1!
1'
1/
#969600000000
0!
0'
0/
#969610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#969620000000
0!
0'
0/
#969630000000
1!
1'
1/
#969640000000
0!
0'
0/
#969650000000
#969660000000
1!
1'
1/
#969670000000
0!
0'
0/
#969680000000
1!
1'
1/
#969690000000
0!
1"
0'
1(
0/
10
#969700000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#969710000000
0!
0'
0/
#969720000000
1!
1'
1/
#969730000000
0!
0'
0/
#969740000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#969750000000
0!
0'
0/
#969760000000
1!
1'
1/
#969770000000
0!
1"
0'
1(
0/
10
#969780000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#969790000000
0!
1$
0'
1+
0/
#969800000000
1!
1'
1/
#969810000000
0!
0'
0/
#969820000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#969830000000
0!
0'
0/
#969840000000
1!
1'
1/
#969850000000
0!
0'
0/
#969860000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#969870000000
0!
0'
0/
#969880000000
1!
1'
1/
#969890000000
0!
0'
0/
#969900000000
1!
1'
1/
#969910000000
0!
0'
0/
#969920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#969930000000
0!
0'
0/
#969940000000
1!
1'
1/
#969950000000
0!
0'
0/
#969960000000
1!
1'
1/
#969970000000
0!
0'
0/
#969980000000
1!
1'
1/
#969990000000
0!
0'
0/
#970000000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#970010000000
0!
0'
0/
#970020000000
1!
1'
1/
#970030000000
0!
0'
0/
#970040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#970050000000
0!
0'
0/
#970060000000
1!
1'
1/
#970070000000
0!
0'
0/
#970080000000
#970090000000
1!
1'
1/
#970100000000
0!
0'
0/
#970110000000
1!
1'
1/
#970120000000
0!
1"
0'
1(
0/
10
#970130000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#970140000000
0!
0'
0/
#970150000000
1!
1'
1/
#970160000000
0!
0'
0/
#970170000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#970180000000
0!
0'
0/
#970190000000
1!
1'
1/
#970200000000
0!
1"
0'
1(
0/
10
#970210000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#970220000000
0!
1$
0'
1+
0/
#970230000000
1!
1'
1/
#970240000000
0!
0'
0/
#970250000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#970260000000
0!
0'
0/
#970270000000
1!
1'
1/
#970280000000
0!
0'
0/
#970290000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#970300000000
0!
0'
0/
#970310000000
1!
1'
1/
#970320000000
0!
0'
0/
#970330000000
1!
1'
1/
#970340000000
0!
0'
0/
#970350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#970360000000
0!
0'
0/
#970370000000
1!
1'
1/
#970380000000
0!
0'
0/
#970390000000
1!
1'
1/
#970400000000
0!
0'
0/
#970410000000
1!
1'
1/
#970420000000
0!
0'
0/
#970430000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#970440000000
0!
0'
0/
#970450000000
1!
1'
1/
#970460000000
0!
0'
0/
#970470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#970480000000
0!
0'
0/
#970490000000
1!
1'
1/
#970500000000
0!
0'
0/
#970510000000
#970520000000
1!
1'
1/
#970530000000
0!
0'
0/
#970540000000
1!
1'
1/
#970550000000
0!
1"
0'
1(
0/
10
#970560000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#970570000000
0!
0'
0/
#970580000000
1!
1'
1/
#970590000000
0!
0'
0/
#970600000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#970610000000
0!
0'
0/
#970620000000
1!
1'
1/
#970630000000
0!
1"
0'
1(
0/
10
#970640000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#970650000000
0!
1$
0'
1+
0/
#970660000000
1!
1'
1/
#970670000000
0!
0'
0/
#970680000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#970690000000
0!
0'
0/
#970700000000
1!
1'
1/
#970710000000
0!
0'
0/
#970720000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#970730000000
0!
0'
0/
#970740000000
1!
1'
1/
#970750000000
0!
0'
0/
#970760000000
1!
1'
1/
#970770000000
0!
0'
0/
#970780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#970790000000
0!
0'
0/
#970800000000
1!
1'
1/
#970810000000
0!
0'
0/
#970820000000
1!
1'
1/
#970830000000
0!
0'
0/
#970840000000
1!
1'
1/
#970850000000
0!
0'
0/
#970860000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#970870000000
0!
0'
0/
#970880000000
1!
1'
1/
#970890000000
0!
0'
0/
#970900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#970910000000
0!
0'
0/
#970920000000
1!
1'
1/
#970930000000
0!
0'
0/
#970940000000
#970950000000
1!
1'
1/
#970960000000
0!
0'
0/
#970970000000
1!
1'
1/
#970980000000
0!
1"
0'
1(
0/
10
#970990000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#971000000000
0!
0'
0/
#971010000000
1!
1'
1/
#971020000000
0!
0'
0/
#971030000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#971040000000
0!
0'
0/
#971050000000
1!
1'
1/
#971060000000
0!
1"
0'
1(
0/
10
#971070000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#971080000000
0!
1$
0'
1+
0/
#971090000000
1!
1'
1/
#971100000000
0!
0'
0/
#971110000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#971120000000
0!
0'
0/
#971130000000
1!
1'
1/
#971140000000
0!
0'
0/
#971150000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#971160000000
0!
0'
0/
#971170000000
1!
1'
1/
#971180000000
0!
0'
0/
#971190000000
1!
1'
1/
#971200000000
0!
0'
0/
#971210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#971220000000
0!
0'
0/
#971230000000
1!
1'
1/
#971240000000
0!
0'
0/
#971250000000
1!
1'
1/
#971260000000
0!
0'
0/
#971270000000
1!
1'
1/
#971280000000
0!
0'
0/
#971290000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#971300000000
0!
0'
0/
#971310000000
1!
1'
1/
#971320000000
0!
0'
0/
#971330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#971340000000
0!
0'
0/
#971350000000
1!
1'
1/
#971360000000
0!
0'
0/
#971370000000
#971380000000
1!
1'
1/
#971390000000
0!
0'
0/
#971400000000
1!
1'
1/
#971410000000
0!
1"
0'
1(
0/
10
#971420000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#971430000000
0!
0'
0/
#971440000000
1!
1'
1/
#971450000000
0!
0'
0/
#971460000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#971470000000
0!
0'
0/
#971480000000
1!
1'
1/
#971490000000
0!
1"
0'
1(
0/
10
#971500000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#971510000000
0!
1$
0'
1+
0/
#971520000000
1!
1'
1/
#971530000000
0!
0'
0/
#971540000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#971550000000
0!
0'
0/
#971560000000
1!
1'
1/
#971570000000
0!
0'
0/
#971580000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#971590000000
0!
0'
0/
#971600000000
1!
1'
1/
#971610000000
0!
0'
0/
#971620000000
1!
1'
1/
#971630000000
0!
0'
0/
#971640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#971650000000
0!
0'
0/
#971660000000
1!
1'
1/
#971670000000
0!
0'
0/
#971680000000
1!
1'
1/
#971690000000
0!
0'
0/
#971700000000
1!
1'
1/
#971710000000
0!
0'
0/
#971720000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#971730000000
0!
0'
0/
#971740000000
1!
1'
1/
#971750000000
0!
0'
0/
#971760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#971770000000
0!
0'
0/
#971780000000
1!
1'
1/
#971790000000
0!
0'
0/
#971800000000
#971810000000
1!
1'
1/
#971820000000
0!
0'
0/
#971830000000
1!
1'
1/
#971840000000
0!
1"
0'
1(
0/
10
#971850000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#971860000000
0!
0'
0/
#971870000000
1!
1'
1/
#971880000000
0!
0'
0/
#971890000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#971900000000
0!
0'
0/
#971910000000
1!
1'
1/
#971920000000
0!
1"
0'
1(
0/
10
#971930000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#971940000000
0!
1$
0'
1+
0/
#971950000000
1!
1'
1/
#971960000000
0!
0'
0/
#971970000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#971980000000
0!
0'
0/
#971990000000
1!
1'
1/
#972000000000
0!
0'
0/
#972010000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#972020000000
0!
0'
0/
#972030000000
1!
1'
1/
#972040000000
0!
0'
0/
#972050000000
1!
1'
1/
#972060000000
0!
0'
0/
#972070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#972080000000
0!
0'
0/
#972090000000
1!
1'
1/
#972100000000
0!
0'
0/
#972110000000
1!
1'
1/
#972120000000
0!
0'
0/
#972130000000
1!
1'
1/
#972140000000
0!
0'
0/
#972150000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#972160000000
0!
0'
0/
#972170000000
1!
1'
1/
#972180000000
0!
0'
0/
#972190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#972200000000
0!
0'
0/
#972210000000
1!
1'
1/
#972220000000
0!
0'
0/
#972230000000
#972240000000
1!
1'
1/
#972250000000
0!
0'
0/
#972260000000
1!
1'
1/
#972270000000
0!
1"
0'
1(
0/
10
#972280000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#972290000000
0!
0'
0/
#972300000000
1!
1'
1/
#972310000000
0!
0'
0/
#972320000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#972330000000
0!
0'
0/
#972340000000
1!
1'
1/
#972350000000
0!
1"
0'
1(
0/
10
#972360000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#972370000000
0!
1$
0'
1+
0/
#972380000000
1!
1'
1/
#972390000000
0!
0'
0/
#972400000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#972410000000
0!
0'
0/
#972420000000
1!
1'
1/
#972430000000
0!
0'
0/
#972440000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#972450000000
0!
0'
0/
#972460000000
1!
1'
1/
#972470000000
0!
0'
0/
#972480000000
1!
1'
1/
#972490000000
0!
0'
0/
#972500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#972510000000
0!
0'
0/
#972520000000
1!
1'
1/
#972530000000
0!
0'
0/
#972540000000
1!
1'
1/
#972550000000
0!
0'
0/
#972560000000
1!
1'
1/
#972570000000
0!
0'
0/
#972580000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#972590000000
0!
0'
0/
#972600000000
1!
1'
1/
#972610000000
0!
0'
0/
#972620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#972630000000
0!
0'
0/
#972640000000
1!
1'
1/
#972650000000
0!
0'
0/
#972660000000
#972670000000
1!
1'
1/
#972680000000
0!
0'
0/
#972690000000
1!
1'
1/
#972700000000
0!
1"
0'
1(
0/
10
#972710000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#972720000000
0!
0'
0/
#972730000000
1!
1'
1/
#972740000000
0!
0'
0/
#972750000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#972760000000
0!
0'
0/
#972770000000
1!
1'
1/
#972780000000
0!
1"
0'
1(
0/
10
#972790000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#972800000000
0!
1$
0'
1+
0/
#972810000000
1!
1'
1/
#972820000000
0!
0'
0/
#972830000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#972840000000
0!
0'
0/
#972850000000
1!
1'
1/
#972860000000
0!
0'
0/
#972870000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#972880000000
0!
0'
0/
#972890000000
1!
1'
1/
#972900000000
0!
0'
0/
#972910000000
1!
1'
1/
#972920000000
0!
0'
0/
#972930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#972940000000
0!
0'
0/
#972950000000
1!
1'
1/
#972960000000
0!
0'
0/
#972970000000
1!
1'
1/
#972980000000
0!
0'
0/
#972990000000
1!
1'
1/
#973000000000
0!
0'
0/
#973010000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#973020000000
0!
0'
0/
#973030000000
1!
1'
1/
#973040000000
0!
0'
0/
#973050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#973060000000
0!
0'
0/
#973070000000
1!
1'
1/
#973080000000
0!
0'
0/
#973090000000
#973100000000
1!
1'
1/
#973110000000
0!
0'
0/
#973120000000
1!
1'
1/
#973130000000
0!
1"
0'
1(
0/
10
#973140000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#973150000000
0!
0'
0/
#973160000000
1!
1'
1/
#973170000000
0!
0'
0/
#973180000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#973190000000
0!
0'
0/
#973200000000
1!
1'
1/
#973210000000
0!
1"
0'
1(
0/
10
#973220000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#973230000000
0!
1$
0'
1+
0/
#973240000000
1!
1'
1/
#973250000000
0!
0'
0/
#973260000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#973270000000
0!
0'
0/
#973280000000
1!
1'
1/
#973290000000
0!
0'
0/
#973300000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#973310000000
0!
0'
0/
#973320000000
1!
1'
1/
#973330000000
0!
0'
0/
#973340000000
1!
1'
1/
#973350000000
0!
0'
0/
#973360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#973370000000
0!
0'
0/
#973380000000
1!
1'
1/
#973390000000
0!
0'
0/
#973400000000
1!
1'
1/
#973410000000
0!
0'
0/
#973420000000
1!
1'
1/
#973430000000
0!
0'
0/
#973440000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#973450000000
0!
0'
0/
#973460000000
1!
1'
1/
#973470000000
0!
0'
0/
#973480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#973490000000
0!
0'
0/
#973500000000
1!
1'
1/
#973510000000
0!
0'
0/
#973520000000
#973530000000
1!
1'
1/
#973540000000
0!
0'
0/
#973550000000
1!
1'
1/
#973560000000
0!
1"
0'
1(
0/
10
#973570000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#973580000000
0!
0'
0/
#973590000000
1!
1'
1/
#973600000000
0!
0'
0/
#973610000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#973620000000
0!
0'
0/
#973630000000
1!
1'
1/
#973640000000
0!
1"
0'
1(
0/
10
#973650000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#973660000000
0!
1$
0'
1+
0/
#973670000000
1!
1'
1/
#973680000000
0!
0'
0/
#973690000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#973700000000
0!
0'
0/
#973710000000
1!
1'
1/
#973720000000
0!
0'
0/
#973730000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#973740000000
0!
0'
0/
#973750000000
1!
1'
1/
#973760000000
0!
0'
0/
#973770000000
1!
1'
1/
#973780000000
0!
0'
0/
#973790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#973800000000
0!
0'
0/
#973810000000
1!
1'
1/
#973820000000
0!
0'
0/
#973830000000
1!
1'
1/
#973840000000
0!
0'
0/
#973850000000
1!
1'
1/
#973860000000
0!
0'
0/
#973870000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#973880000000
0!
0'
0/
#973890000000
1!
1'
1/
#973900000000
0!
0'
0/
#973910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#973920000000
0!
0'
0/
#973930000000
1!
1'
1/
#973940000000
0!
0'
0/
#973950000000
#973960000000
1!
1'
1/
#973970000000
0!
0'
0/
#973980000000
1!
1'
1/
#973990000000
0!
1"
0'
1(
0/
10
#974000000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#974010000000
0!
0'
0/
#974020000000
1!
1'
1/
#974030000000
0!
0'
0/
#974040000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#974050000000
0!
0'
0/
#974060000000
1!
1'
1/
#974070000000
0!
1"
0'
1(
0/
10
#974080000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#974090000000
0!
1$
0'
1+
0/
#974100000000
1!
1'
1/
#974110000000
0!
0'
0/
#974120000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#974130000000
0!
0'
0/
#974140000000
1!
1'
1/
#974150000000
0!
0'
0/
#974160000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#974170000000
0!
0'
0/
#974180000000
1!
1'
1/
#974190000000
0!
0'
0/
#974200000000
1!
1'
1/
#974210000000
0!
0'
0/
#974220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#974230000000
0!
0'
0/
#974240000000
1!
1'
1/
#974250000000
0!
0'
0/
#974260000000
1!
1'
1/
#974270000000
0!
0'
0/
#974280000000
1!
1'
1/
#974290000000
0!
0'
0/
#974300000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#974310000000
0!
0'
0/
#974320000000
1!
1'
1/
#974330000000
0!
0'
0/
#974340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#974350000000
0!
0'
0/
#974360000000
1!
1'
1/
#974370000000
0!
0'
0/
#974380000000
#974390000000
1!
1'
1/
#974400000000
0!
0'
0/
#974410000000
1!
1'
1/
#974420000000
0!
1"
0'
1(
0/
10
#974430000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#974440000000
0!
0'
0/
#974450000000
1!
1'
1/
#974460000000
0!
0'
0/
#974470000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#974480000000
0!
0'
0/
#974490000000
1!
1'
1/
#974500000000
0!
1"
0'
1(
0/
10
#974510000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#974520000000
0!
1$
0'
1+
0/
#974530000000
1!
1'
1/
#974540000000
0!
0'
0/
#974550000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#974560000000
0!
0'
0/
#974570000000
1!
1'
1/
#974580000000
0!
0'
0/
#974590000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#974600000000
0!
0'
0/
#974610000000
1!
1'
1/
#974620000000
0!
0'
0/
#974630000000
1!
1'
1/
#974640000000
0!
0'
0/
#974650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#974660000000
0!
0'
0/
#974670000000
1!
1'
1/
#974680000000
0!
0'
0/
#974690000000
1!
1'
1/
#974700000000
0!
0'
0/
#974710000000
1!
1'
1/
#974720000000
0!
0'
0/
#974730000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#974740000000
0!
0'
0/
#974750000000
1!
1'
1/
#974760000000
0!
0'
0/
#974770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#974780000000
0!
0'
0/
#974790000000
1!
1'
1/
#974800000000
0!
0'
0/
#974810000000
#974820000000
1!
1'
1/
#974830000000
0!
0'
0/
#974840000000
1!
1'
1/
#974850000000
0!
1"
0'
1(
0/
10
#974860000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#974870000000
0!
0'
0/
#974880000000
1!
1'
1/
#974890000000
0!
0'
0/
#974900000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#974910000000
0!
0'
0/
#974920000000
1!
1'
1/
#974930000000
0!
1"
0'
1(
0/
10
#974940000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#974950000000
0!
1$
0'
1+
0/
#974960000000
1!
1'
1/
#974970000000
0!
0'
0/
#974980000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#974990000000
0!
0'
0/
#975000000000
1!
1'
1/
#975010000000
0!
0'
0/
#975020000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#975030000000
0!
0'
0/
#975040000000
1!
1'
1/
#975050000000
0!
0'
0/
#975060000000
1!
1'
1/
#975070000000
0!
0'
0/
#975080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#975090000000
0!
0'
0/
#975100000000
1!
1'
1/
#975110000000
0!
0'
0/
#975120000000
1!
1'
1/
#975130000000
0!
0'
0/
#975140000000
1!
1'
1/
#975150000000
0!
0'
0/
#975160000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#975170000000
0!
0'
0/
#975180000000
1!
1'
1/
#975190000000
0!
0'
0/
#975200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#975210000000
0!
0'
0/
#975220000000
1!
1'
1/
#975230000000
0!
0'
0/
#975240000000
#975250000000
1!
1'
1/
#975260000000
0!
0'
0/
#975270000000
1!
1'
1/
#975280000000
0!
1"
0'
1(
0/
10
#975290000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#975300000000
0!
0'
0/
#975310000000
1!
1'
1/
#975320000000
0!
0'
0/
#975330000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#975340000000
0!
0'
0/
#975350000000
1!
1'
1/
#975360000000
0!
1"
0'
1(
0/
10
#975370000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#975380000000
0!
1$
0'
1+
0/
#975390000000
1!
1'
1/
#975400000000
0!
0'
0/
#975410000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#975420000000
0!
0'
0/
#975430000000
1!
1'
1/
#975440000000
0!
0'
0/
#975450000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#975460000000
0!
0'
0/
#975470000000
1!
1'
1/
#975480000000
0!
0'
0/
#975490000000
1!
1'
1/
#975500000000
0!
0'
0/
#975510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#975520000000
0!
0'
0/
#975530000000
1!
1'
1/
#975540000000
0!
0'
0/
#975550000000
1!
1'
1/
#975560000000
0!
0'
0/
#975570000000
1!
1'
1/
#975580000000
0!
0'
0/
#975590000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#975600000000
0!
0'
0/
#975610000000
1!
1'
1/
#975620000000
0!
0'
0/
#975630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#975640000000
0!
0'
0/
#975650000000
1!
1'
1/
#975660000000
0!
0'
0/
#975670000000
#975680000000
1!
1'
1/
#975690000000
0!
0'
0/
#975700000000
1!
1'
1/
#975710000000
0!
1"
0'
1(
0/
10
#975720000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#975730000000
0!
0'
0/
#975740000000
1!
1'
1/
#975750000000
0!
0'
0/
#975760000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#975770000000
0!
0'
0/
#975780000000
1!
1'
1/
#975790000000
0!
1"
0'
1(
0/
10
#975800000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#975810000000
0!
1$
0'
1+
0/
#975820000000
1!
1'
1/
#975830000000
0!
0'
0/
#975840000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#975850000000
0!
0'
0/
#975860000000
1!
1'
1/
#975870000000
0!
0'
0/
#975880000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#975890000000
0!
0'
0/
#975900000000
1!
1'
1/
#975910000000
0!
0'
0/
#975920000000
1!
1'
1/
#975930000000
0!
0'
0/
#975940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#975950000000
0!
0'
0/
#975960000000
1!
1'
1/
#975970000000
0!
0'
0/
#975980000000
1!
1'
1/
#975990000000
0!
0'
0/
#976000000000
1!
1'
1/
#976010000000
0!
0'
0/
#976020000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#976030000000
0!
0'
0/
#976040000000
1!
1'
1/
#976050000000
0!
0'
0/
#976060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#976070000000
0!
0'
0/
#976080000000
1!
1'
1/
#976090000000
0!
0'
0/
#976100000000
#976110000000
1!
1'
1/
#976120000000
0!
0'
0/
#976130000000
1!
1'
1/
#976140000000
0!
1"
0'
1(
0/
10
#976150000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#976160000000
0!
0'
0/
#976170000000
1!
1'
1/
#976180000000
0!
0'
0/
#976190000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#976200000000
0!
0'
0/
#976210000000
1!
1'
1/
#976220000000
0!
1"
0'
1(
0/
10
#976230000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#976240000000
0!
1$
0'
1+
0/
#976250000000
1!
1'
1/
#976260000000
0!
0'
0/
#976270000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#976280000000
0!
0'
0/
#976290000000
1!
1'
1/
#976300000000
0!
0'
0/
#976310000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#976320000000
0!
0'
0/
#976330000000
1!
1'
1/
#976340000000
0!
0'
0/
#976350000000
1!
1'
1/
#976360000000
0!
0'
0/
#976370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#976380000000
0!
0'
0/
#976390000000
1!
1'
1/
#976400000000
0!
0'
0/
#976410000000
1!
1'
1/
#976420000000
0!
0'
0/
#976430000000
1!
1'
1/
#976440000000
0!
0'
0/
#976450000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#976460000000
0!
0'
0/
#976470000000
1!
1'
1/
#976480000000
0!
0'
0/
#976490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#976500000000
0!
0'
0/
#976510000000
1!
1'
1/
#976520000000
0!
0'
0/
#976530000000
#976540000000
1!
1'
1/
#976550000000
0!
0'
0/
#976560000000
1!
1'
1/
#976570000000
0!
1"
0'
1(
0/
10
#976580000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#976590000000
0!
0'
0/
#976600000000
1!
1'
1/
#976610000000
0!
0'
0/
#976620000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#976630000000
0!
0'
0/
#976640000000
1!
1'
1/
#976650000000
0!
1"
0'
1(
0/
10
#976660000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#976670000000
0!
1$
0'
1+
0/
#976680000000
1!
1'
1/
#976690000000
0!
0'
0/
#976700000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#976710000000
0!
0'
0/
#976720000000
1!
1'
1/
#976730000000
0!
0'
0/
#976740000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#976750000000
0!
0'
0/
#976760000000
1!
1'
1/
#976770000000
0!
0'
0/
#976780000000
1!
1'
1/
#976790000000
0!
0'
0/
#976800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#976810000000
0!
0'
0/
#976820000000
1!
1'
1/
#976830000000
0!
0'
0/
#976840000000
1!
1'
1/
#976850000000
0!
0'
0/
#976860000000
1!
1'
1/
#976870000000
0!
0'
0/
#976880000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#976890000000
0!
0'
0/
#976900000000
1!
1'
1/
#976910000000
0!
0'
0/
#976920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#976930000000
0!
0'
0/
#976940000000
1!
1'
1/
#976950000000
0!
0'
0/
#976960000000
#976970000000
1!
1'
1/
#976980000000
0!
0'
0/
#976990000000
1!
1'
1/
#977000000000
0!
1"
0'
1(
0/
10
#977010000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#977020000000
0!
0'
0/
#977030000000
1!
1'
1/
#977040000000
0!
0'
0/
#977050000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#977060000000
0!
0'
0/
#977070000000
1!
1'
1/
#977080000000
0!
1"
0'
1(
0/
10
#977090000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#977100000000
0!
1$
0'
1+
0/
#977110000000
1!
1'
1/
#977120000000
0!
0'
0/
#977130000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#977140000000
0!
0'
0/
#977150000000
1!
1'
1/
#977160000000
0!
0'
0/
#977170000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#977180000000
0!
0'
0/
#977190000000
1!
1'
1/
#977200000000
0!
0'
0/
#977210000000
1!
1'
1/
#977220000000
0!
0'
0/
#977230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#977240000000
0!
0'
0/
#977250000000
1!
1'
1/
#977260000000
0!
0'
0/
#977270000000
1!
1'
1/
#977280000000
0!
0'
0/
#977290000000
1!
1'
1/
#977300000000
0!
0'
0/
#977310000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#977320000000
0!
0'
0/
#977330000000
1!
1'
1/
#977340000000
0!
0'
0/
#977350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#977360000000
0!
0'
0/
#977370000000
1!
1'
1/
#977380000000
0!
0'
0/
#977390000000
#977400000000
1!
1'
1/
#977410000000
0!
0'
0/
#977420000000
1!
1'
1/
#977430000000
0!
1"
0'
1(
0/
10
#977440000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#977450000000
0!
0'
0/
#977460000000
1!
1'
1/
#977470000000
0!
0'
0/
#977480000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#977490000000
0!
0'
0/
#977500000000
1!
1'
1/
#977510000000
0!
1"
0'
1(
0/
10
#977520000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#977530000000
0!
1$
0'
1+
0/
#977540000000
1!
1'
1/
#977550000000
0!
0'
0/
#977560000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#977570000000
0!
0'
0/
#977580000000
1!
1'
1/
#977590000000
0!
0'
0/
#977600000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#977610000000
0!
0'
0/
#977620000000
1!
1'
1/
#977630000000
0!
0'
0/
#977640000000
1!
1'
1/
#977650000000
0!
0'
0/
#977660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#977670000000
0!
0'
0/
#977680000000
1!
1'
1/
#977690000000
0!
0'
0/
#977700000000
1!
1'
1/
#977710000000
0!
0'
0/
#977720000000
1!
1'
1/
#977730000000
0!
0'
0/
#977740000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#977750000000
0!
0'
0/
#977760000000
1!
1'
1/
#977770000000
0!
0'
0/
#977780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#977790000000
0!
0'
0/
#977800000000
1!
1'
1/
#977810000000
0!
0'
0/
#977820000000
#977830000000
1!
1'
1/
#977840000000
0!
0'
0/
#977850000000
1!
1'
1/
#977860000000
0!
1"
0'
1(
0/
10
#977870000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#977880000000
0!
0'
0/
#977890000000
1!
1'
1/
#977900000000
0!
0'
0/
#977910000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#977920000000
0!
0'
0/
#977930000000
1!
1'
1/
#977940000000
0!
1"
0'
1(
0/
10
#977950000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#977960000000
0!
1$
0'
1+
0/
#977970000000
1!
1'
1/
#977980000000
0!
0'
0/
#977990000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#978000000000
0!
0'
0/
#978010000000
1!
1'
1/
#978020000000
0!
0'
0/
#978030000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#978040000000
0!
0'
0/
#978050000000
1!
1'
1/
#978060000000
0!
0'
0/
#978070000000
1!
1'
1/
#978080000000
0!
0'
0/
#978090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#978100000000
0!
0'
0/
#978110000000
1!
1'
1/
#978120000000
0!
0'
0/
#978130000000
1!
1'
1/
#978140000000
0!
0'
0/
#978150000000
1!
1'
1/
#978160000000
0!
0'
0/
#978170000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#978180000000
0!
0'
0/
#978190000000
1!
1'
1/
#978200000000
0!
0'
0/
#978210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#978220000000
0!
0'
0/
#978230000000
1!
1'
1/
#978240000000
0!
0'
0/
#978250000000
#978260000000
1!
1'
1/
#978270000000
0!
0'
0/
#978280000000
1!
1'
1/
#978290000000
0!
1"
0'
1(
0/
10
#978300000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#978310000000
0!
0'
0/
#978320000000
1!
1'
1/
#978330000000
0!
0'
0/
#978340000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#978350000000
0!
0'
0/
#978360000000
1!
1'
1/
#978370000000
0!
1"
0'
1(
0/
10
#978380000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#978390000000
0!
1$
0'
1+
0/
#978400000000
1!
1'
1/
#978410000000
0!
0'
0/
#978420000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#978430000000
0!
0'
0/
#978440000000
1!
1'
1/
#978450000000
0!
0'
0/
#978460000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#978470000000
0!
0'
0/
#978480000000
1!
1'
1/
#978490000000
0!
0'
0/
#978500000000
1!
1'
1/
#978510000000
0!
0'
0/
#978520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#978530000000
0!
0'
0/
#978540000000
1!
1'
1/
#978550000000
0!
0'
0/
#978560000000
1!
1'
1/
#978570000000
0!
0'
0/
#978580000000
1!
1'
1/
#978590000000
0!
0'
0/
#978600000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#978610000000
0!
0'
0/
#978620000000
1!
1'
1/
#978630000000
0!
0'
0/
#978640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#978650000000
0!
0'
0/
#978660000000
1!
1'
1/
#978670000000
0!
0'
0/
#978680000000
#978690000000
1!
1'
1/
#978700000000
0!
0'
0/
#978710000000
1!
1'
1/
#978720000000
0!
1"
0'
1(
0/
10
#978730000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#978740000000
0!
0'
0/
#978750000000
1!
1'
1/
#978760000000
0!
0'
0/
#978770000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#978780000000
0!
0'
0/
#978790000000
1!
1'
1/
#978800000000
0!
1"
0'
1(
0/
10
#978810000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#978820000000
0!
1$
0'
1+
0/
#978830000000
1!
1'
1/
#978840000000
0!
0'
0/
#978850000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#978860000000
0!
0'
0/
#978870000000
1!
1'
1/
#978880000000
0!
0'
0/
#978890000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#978900000000
0!
0'
0/
#978910000000
1!
1'
1/
#978920000000
0!
0'
0/
#978930000000
1!
1'
1/
#978940000000
0!
0'
0/
#978950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#978960000000
0!
0'
0/
#978970000000
1!
1'
1/
#978980000000
0!
0'
0/
#978990000000
1!
1'
1/
#979000000000
0!
0'
0/
#979010000000
1!
1'
1/
#979020000000
0!
0'
0/
#979030000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#979040000000
0!
0'
0/
#979050000000
1!
1'
1/
#979060000000
0!
0'
0/
#979070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#979080000000
0!
0'
0/
#979090000000
1!
1'
1/
#979100000000
0!
0'
0/
#979110000000
#979120000000
1!
1'
1/
#979130000000
0!
0'
0/
#979140000000
1!
1'
1/
#979150000000
0!
1"
0'
1(
0/
10
#979160000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#979170000000
0!
0'
0/
#979180000000
1!
1'
1/
#979190000000
0!
0'
0/
#979200000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#979210000000
0!
0'
0/
#979220000000
1!
1'
1/
#979230000000
0!
1"
0'
1(
0/
10
#979240000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#979250000000
0!
1$
0'
1+
0/
#979260000000
1!
1'
1/
#979270000000
0!
0'
0/
#979280000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#979290000000
0!
0'
0/
#979300000000
1!
1'
1/
#979310000000
0!
0'
0/
#979320000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#979330000000
0!
0'
0/
#979340000000
1!
1'
1/
#979350000000
0!
0'
0/
#979360000000
1!
1'
1/
#979370000000
0!
0'
0/
#979380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#979390000000
0!
0'
0/
#979400000000
1!
1'
1/
#979410000000
0!
0'
0/
#979420000000
1!
1'
1/
#979430000000
0!
0'
0/
#979440000000
1!
1'
1/
#979450000000
0!
0'
0/
#979460000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#979470000000
0!
0'
0/
#979480000000
1!
1'
1/
#979490000000
0!
0'
0/
#979500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#979510000000
0!
0'
0/
#979520000000
1!
1'
1/
#979530000000
0!
0'
0/
#979540000000
#979550000000
1!
1'
1/
#979560000000
0!
0'
0/
#979570000000
1!
1'
1/
#979580000000
0!
1"
0'
1(
0/
10
#979590000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#979600000000
0!
0'
0/
#979610000000
1!
1'
1/
#979620000000
0!
0'
0/
#979630000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#979640000000
0!
0'
0/
#979650000000
1!
1'
1/
#979660000000
0!
1"
0'
1(
0/
10
#979670000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#979680000000
0!
1$
0'
1+
0/
#979690000000
1!
1'
1/
#979700000000
0!
0'
0/
#979710000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#979720000000
0!
0'
0/
#979730000000
1!
1'
1/
#979740000000
0!
0'
0/
#979750000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#979760000000
0!
0'
0/
#979770000000
1!
1'
1/
#979780000000
0!
0'
0/
#979790000000
1!
1'
1/
#979800000000
0!
0'
0/
#979810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#979820000000
0!
0'
0/
#979830000000
1!
1'
1/
#979840000000
0!
0'
0/
#979850000000
1!
1'
1/
#979860000000
0!
0'
0/
#979870000000
1!
1'
1/
#979880000000
0!
0'
0/
#979890000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#979900000000
0!
0'
0/
#979910000000
1!
1'
1/
#979920000000
0!
0'
0/
#979930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#979940000000
0!
0'
0/
#979950000000
1!
1'
1/
#979960000000
0!
0'
0/
#979970000000
#979980000000
1!
1'
1/
#979990000000
0!
0'
0/
#980000000000
1!
1'
1/
#980010000000
0!
1"
0'
1(
0/
10
#980020000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#980030000000
0!
0'
0/
#980040000000
1!
1'
1/
#980050000000
0!
0'
0/
#980060000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#980070000000
0!
0'
0/
#980080000000
1!
1'
1/
#980090000000
0!
1"
0'
1(
0/
10
#980100000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#980110000000
0!
1$
0'
1+
0/
#980120000000
1!
1'
1/
#980130000000
0!
0'
0/
#980140000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#980150000000
0!
0'
0/
#980160000000
1!
1'
1/
#980170000000
0!
0'
0/
#980180000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#980190000000
0!
0'
0/
#980200000000
1!
1'
1/
#980210000000
0!
0'
0/
#980220000000
1!
1'
1/
#980230000000
0!
0'
0/
#980240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#980250000000
0!
0'
0/
#980260000000
1!
1'
1/
#980270000000
0!
0'
0/
#980280000000
1!
1'
1/
#980290000000
0!
0'
0/
#980300000000
1!
1'
1/
#980310000000
0!
0'
0/
#980320000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#980330000000
0!
0'
0/
#980340000000
1!
1'
1/
#980350000000
0!
0'
0/
#980360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#980370000000
0!
0'
0/
#980380000000
1!
1'
1/
#980390000000
0!
0'
0/
#980400000000
#980410000000
1!
1'
1/
#980420000000
0!
0'
0/
#980430000000
1!
1'
1/
#980440000000
0!
1"
0'
1(
0/
10
#980450000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#980460000000
0!
0'
0/
#980470000000
1!
1'
1/
#980480000000
0!
0'
0/
#980490000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#980500000000
0!
0'
0/
#980510000000
1!
1'
1/
#980520000000
0!
1"
0'
1(
0/
10
#980530000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#980540000000
0!
1$
0'
1+
0/
#980550000000
1!
1'
1/
#980560000000
0!
0'
0/
#980570000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#980580000000
0!
0'
0/
#980590000000
1!
1'
1/
#980600000000
0!
0'
0/
#980610000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#980620000000
0!
0'
0/
#980630000000
1!
1'
1/
#980640000000
0!
0'
0/
#980650000000
1!
1'
1/
#980660000000
0!
0'
0/
#980670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#980680000000
0!
0'
0/
#980690000000
1!
1'
1/
#980700000000
0!
0'
0/
#980710000000
1!
1'
1/
#980720000000
0!
0'
0/
#980730000000
1!
1'
1/
#980740000000
0!
0'
0/
#980750000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#980760000000
0!
0'
0/
#980770000000
1!
1'
1/
#980780000000
0!
0'
0/
#980790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#980800000000
0!
0'
0/
#980810000000
1!
1'
1/
#980820000000
0!
0'
0/
#980830000000
#980840000000
1!
1'
1/
#980850000000
0!
0'
0/
#980860000000
1!
1'
1/
#980870000000
0!
1"
0'
1(
0/
10
#980880000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#980890000000
0!
0'
0/
#980900000000
1!
1'
1/
#980910000000
0!
0'
0/
#980920000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#980930000000
0!
0'
0/
#980940000000
1!
1'
1/
#980950000000
0!
1"
0'
1(
0/
10
#980960000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#980970000000
0!
1$
0'
1+
0/
#980980000000
1!
1'
1/
#980990000000
0!
0'
0/
#981000000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#981010000000
0!
0'
0/
#981020000000
1!
1'
1/
#981030000000
0!
0'
0/
#981040000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#981050000000
0!
0'
0/
#981060000000
1!
1'
1/
#981070000000
0!
0'
0/
#981080000000
1!
1'
1/
#981090000000
0!
0'
0/
#981100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#981110000000
0!
0'
0/
#981120000000
1!
1'
1/
#981130000000
0!
0'
0/
#981140000000
1!
1'
1/
#981150000000
0!
0'
0/
#981160000000
1!
1'
1/
#981170000000
0!
0'
0/
#981180000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#981190000000
0!
0'
0/
#981200000000
1!
1'
1/
#981210000000
0!
0'
0/
#981220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#981230000000
0!
0'
0/
#981240000000
1!
1'
1/
#981250000000
0!
0'
0/
#981260000000
#981270000000
1!
1'
1/
#981280000000
0!
0'
0/
#981290000000
1!
1'
1/
#981300000000
0!
1"
0'
1(
0/
10
#981310000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#981320000000
0!
0'
0/
#981330000000
1!
1'
1/
#981340000000
0!
0'
0/
#981350000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#981360000000
0!
0'
0/
#981370000000
1!
1'
1/
#981380000000
0!
1"
0'
1(
0/
10
#981390000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#981400000000
0!
1$
0'
1+
0/
#981410000000
1!
1'
1/
#981420000000
0!
0'
0/
#981430000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#981440000000
0!
0'
0/
#981450000000
1!
1'
1/
#981460000000
0!
0'
0/
#981470000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#981480000000
0!
0'
0/
#981490000000
1!
1'
1/
#981500000000
0!
0'
0/
#981510000000
1!
1'
1/
#981520000000
0!
0'
0/
#981530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#981540000000
0!
0'
0/
#981550000000
1!
1'
1/
#981560000000
0!
0'
0/
#981570000000
1!
1'
1/
#981580000000
0!
0'
0/
#981590000000
1!
1'
1/
#981600000000
0!
0'
0/
#981610000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#981620000000
0!
0'
0/
#981630000000
1!
1'
1/
#981640000000
0!
0'
0/
#981650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#981660000000
0!
0'
0/
#981670000000
1!
1'
1/
#981680000000
0!
0'
0/
#981690000000
#981700000000
1!
1'
1/
#981710000000
0!
0'
0/
#981720000000
1!
1'
1/
#981730000000
0!
1"
0'
1(
0/
10
#981740000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#981750000000
0!
0'
0/
#981760000000
1!
1'
1/
#981770000000
0!
0'
0/
#981780000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#981790000000
0!
0'
0/
#981800000000
1!
1'
1/
#981810000000
0!
1"
0'
1(
0/
10
#981820000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#981830000000
0!
1$
0'
1+
0/
#981840000000
1!
1'
1/
#981850000000
0!
0'
0/
#981860000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#981870000000
0!
0'
0/
#981880000000
1!
1'
1/
#981890000000
0!
0'
0/
#981900000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#981910000000
0!
0'
0/
#981920000000
1!
1'
1/
#981930000000
0!
0'
0/
#981940000000
1!
1'
1/
#981950000000
0!
0'
0/
#981960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#981970000000
0!
0'
0/
#981980000000
1!
1'
1/
#981990000000
0!
0'
0/
#982000000000
1!
1'
1/
#982010000000
0!
0'
0/
#982020000000
1!
1'
1/
#982030000000
0!
0'
0/
#982040000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#982050000000
0!
0'
0/
#982060000000
1!
1'
1/
#982070000000
0!
0'
0/
#982080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#982090000000
0!
0'
0/
#982100000000
1!
1'
1/
#982110000000
0!
0'
0/
#982120000000
#982130000000
1!
1'
1/
#982140000000
0!
0'
0/
#982150000000
1!
1'
1/
#982160000000
0!
1"
0'
1(
0/
10
#982170000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#982180000000
0!
0'
0/
#982190000000
1!
1'
1/
#982200000000
0!
0'
0/
#982210000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#982220000000
0!
0'
0/
#982230000000
1!
1'
1/
#982240000000
0!
1"
0'
1(
0/
10
#982250000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#982260000000
0!
1$
0'
1+
0/
#982270000000
1!
1'
1/
#982280000000
0!
0'
0/
#982290000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#982300000000
0!
0'
0/
#982310000000
1!
1'
1/
#982320000000
0!
0'
0/
#982330000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#982340000000
0!
0'
0/
#982350000000
1!
1'
1/
#982360000000
0!
0'
0/
#982370000000
1!
1'
1/
#982380000000
0!
0'
0/
#982390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#982400000000
0!
0'
0/
#982410000000
1!
1'
1/
#982420000000
0!
0'
0/
#982430000000
1!
1'
1/
#982440000000
0!
0'
0/
#982450000000
1!
1'
1/
#982460000000
0!
0'
0/
#982470000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#982480000000
0!
0'
0/
#982490000000
1!
1'
1/
#982500000000
0!
0'
0/
#982510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#982520000000
0!
0'
0/
#982530000000
1!
1'
1/
#982540000000
0!
0'
0/
#982550000000
#982560000000
1!
1'
1/
#982570000000
0!
0'
0/
#982580000000
1!
1'
1/
#982590000000
0!
1"
0'
1(
0/
10
#982600000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#982610000000
0!
0'
0/
#982620000000
1!
1'
1/
#982630000000
0!
0'
0/
#982640000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#982650000000
0!
0'
0/
#982660000000
1!
1'
1/
#982670000000
0!
1"
0'
1(
0/
10
#982680000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#982690000000
0!
1$
0'
1+
0/
#982700000000
1!
1'
1/
#982710000000
0!
0'
0/
#982720000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#982730000000
0!
0'
0/
#982740000000
1!
1'
1/
#982750000000
0!
0'
0/
#982760000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#982770000000
0!
0'
0/
#982780000000
1!
1'
1/
#982790000000
0!
0'
0/
#982800000000
1!
1'
1/
#982810000000
0!
0'
0/
#982820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#982830000000
0!
0'
0/
#982840000000
1!
1'
1/
#982850000000
0!
0'
0/
#982860000000
1!
1'
1/
#982870000000
0!
0'
0/
#982880000000
1!
1'
1/
#982890000000
0!
0'
0/
#982900000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#982910000000
0!
0'
0/
#982920000000
1!
1'
1/
#982930000000
0!
0'
0/
#982940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#982950000000
0!
0'
0/
#982960000000
1!
1'
1/
#982970000000
0!
0'
0/
#982980000000
#982990000000
1!
1'
1/
#983000000000
0!
0'
0/
#983010000000
1!
1'
1/
#983020000000
0!
1"
0'
1(
0/
10
#983030000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#983040000000
0!
0'
0/
#983050000000
1!
1'
1/
#983060000000
0!
0'
0/
#983070000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#983080000000
0!
0'
0/
#983090000000
1!
1'
1/
#983100000000
0!
1"
0'
1(
0/
10
#983110000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#983120000000
0!
1$
0'
1+
0/
#983130000000
1!
1'
1/
#983140000000
0!
0'
0/
#983150000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#983160000000
0!
0'
0/
#983170000000
1!
1'
1/
#983180000000
0!
0'
0/
#983190000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#983200000000
0!
0'
0/
#983210000000
1!
1'
1/
#983220000000
0!
0'
0/
#983230000000
1!
1'
1/
#983240000000
0!
0'
0/
#983250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#983260000000
0!
0'
0/
#983270000000
1!
1'
1/
#983280000000
0!
0'
0/
#983290000000
1!
1'
1/
#983300000000
0!
0'
0/
#983310000000
1!
1'
1/
#983320000000
0!
0'
0/
#983330000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#983340000000
0!
0'
0/
#983350000000
1!
1'
1/
#983360000000
0!
0'
0/
#983370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#983380000000
0!
0'
0/
#983390000000
1!
1'
1/
#983400000000
0!
0'
0/
#983410000000
#983420000000
1!
1'
1/
#983430000000
0!
0'
0/
#983440000000
1!
1'
1/
#983450000000
0!
1"
0'
1(
0/
10
#983460000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#983470000000
0!
0'
0/
#983480000000
1!
1'
1/
#983490000000
0!
0'
0/
#983500000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#983510000000
0!
0'
0/
#983520000000
1!
1'
1/
#983530000000
0!
1"
0'
1(
0/
10
#983540000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#983550000000
0!
1$
0'
1+
0/
#983560000000
1!
1'
1/
#983570000000
0!
0'
0/
#983580000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#983590000000
0!
0'
0/
#983600000000
1!
1'
1/
#983610000000
0!
0'
0/
#983620000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#983630000000
0!
0'
0/
#983640000000
1!
1'
1/
#983650000000
0!
0'
0/
#983660000000
1!
1'
1/
#983670000000
0!
0'
0/
#983680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#983690000000
0!
0'
0/
#983700000000
1!
1'
1/
#983710000000
0!
0'
0/
#983720000000
1!
1'
1/
#983730000000
0!
0'
0/
#983740000000
1!
1'
1/
#983750000000
0!
0'
0/
#983760000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#983770000000
0!
0'
0/
#983780000000
1!
1'
1/
#983790000000
0!
0'
0/
#983800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#983810000000
0!
0'
0/
#983820000000
1!
1'
1/
#983830000000
0!
0'
0/
#983840000000
#983850000000
1!
1'
1/
#983860000000
0!
0'
0/
#983870000000
1!
1'
1/
#983880000000
0!
1"
0'
1(
0/
10
#983890000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#983900000000
0!
0'
0/
#983910000000
1!
1'
1/
#983920000000
0!
0'
0/
#983930000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#983940000000
0!
0'
0/
#983950000000
1!
1'
1/
#983960000000
0!
1"
0'
1(
0/
10
#983970000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#983980000000
0!
1$
0'
1+
0/
#983990000000
1!
1'
1/
#984000000000
0!
0'
0/
#984010000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#984020000000
0!
0'
0/
#984030000000
1!
1'
1/
#984040000000
0!
0'
0/
#984050000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#984060000000
0!
0'
0/
#984070000000
1!
1'
1/
#984080000000
0!
0'
0/
#984090000000
1!
1'
1/
#984100000000
0!
0'
0/
#984110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#984120000000
0!
0'
0/
#984130000000
1!
1'
1/
#984140000000
0!
0'
0/
#984150000000
1!
1'
1/
#984160000000
0!
0'
0/
#984170000000
1!
1'
1/
#984180000000
0!
0'
0/
#984190000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#984200000000
0!
0'
0/
#984210000000
1!
1'
1/
#984220000000
0!
0'
0/
#984230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#984240000000
0!
0'
0/
#984250000000
1!
1'
1/
#984260000000
0!
0'
0/
#984270000000
#984280000000
1!
1'
1/
#984290000000
0!
0'
0/
#984300000000
1!
1'
1/
#984310000000
0!
1"
0'
1(
0/
10
#984320000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#984330000000
0!
0'
0/
#984340000000
1!
1'
1/
#984350000000
0!
0'
0/
#984360000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#984370000000
0!
0'
0/
#984380000000
1!
1'
1/
#984390000000
0!
1"
0'
1(
0/
10
#984400000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#984410000000
0!
1$
0'
1+
0/
#984420000000
1!
1'
1/
#984430000000
0!
0'
0/
#984440000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#984450000000
0!
0'
0/
#984460000000
1!
1'
1/
#984470000000
0!
0'
0/
#984480000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#984490000000
0!
0'
0/
#984500000000
1!
1'
1/
#984510000000
0!
0'
0/
#984520000000
1!
1'
1/
#984530000000
0!
0'
0/
#984540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#984550000000
0!
0'
0/
#984560000000
1!
1'
1/
#984570000000
0!
0'
0/
#984580000000
1!
1'
1/
#984590000000
0!
0'
0/
#984600000000
1!
1'
1/
#984610000000
0!
0'
0/
#984620000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#984630000000
0!
0'
0/
#984640000000
1!
1'
1/
#984650000000
0!
0'
0/
#984660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#984670000000
0!
0'
0/
#984680000000
1!
1'
1/
#984690000000
0!
0'
0/
#984700000000
#984710000000
1!
1'
1/
#984720000000
0!
0'
0/
#984730000000
1!
1'
1/
#984740000000
0!
1"
0'
1(
0/
10
#984750000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#984760000000
0!
0'
0/
#984770000000
1!
1'
1/
#984780000000
0!
0'
0/
#984790000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#984800000000
0!
0'
0/
#984810000000
1!
1'
1/
#984820000000
0!
1"
0'
1(
0/
10
#984830000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#984840000000
0!
1$
0'
1+
0/
#984850000000
1!
1'
1/
#984860000000
0!
0'
0/
#984870000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#984880000000
0!
0'
0/
#984890000000
1!
1'
1/
#984900000000
0!
0'
0/
#984910000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#984920000000
0!
0'
0/
#984930000000
1!
1'
1/
#984940000000
0!
0'
0/
#984950000000
1!
1'
1/
#984960000000
0!
0'
0/
#984970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#984980000000
0!
0'
0/
#984990000000
1!
1'
1/
#985000000000
0!
0'
0/
#985010000000
1!
1'
1/
#985020000000
0!
0'
0/
#985030000000
1!
1'
1/
#985040000000
0!
0'
0/
#985050000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#985060000000
0!
0'
0/
#985070000000
1!
1'
1/
#985080000000
0!
0'
0/
#985090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#985100000000
0!
0'
0/
#985110000000
1!
1'
1/
#985120000000
0!
0'
0/
#985130000000
#985140000000
1!
1'
1/
#985150000000
0!
0'
0/
#985160000000
1!
1'
1/
#985170000000
0!
1"
0'
1(
0/
10
#985180000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#985190000000
0!
0'
0/
#985200000000
1!
1'
1/
#985210000000
0!
0'
0/
#985220000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#985230000000
0!
0'
0/
#985240000000
1!
1'
1/
#985250000000
0!
1"
0'
1(
0/
10
#985260000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#985270000000
0!
1$
0'
1+
0/
#985280000000
1!
1'
1/
#985290000000
0!
0'
0/
#985300000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#985310000000
0!
0'
0/
#985320000000
1!
1'
1/
#985330000000
0!
0'
0/
#985340000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#985350000000
0!
0'
0/
#985360000000
1!
1'
1/
#985370000000
0!
0'
0/
#985380000000
1!
1'
1/
#985390000000
0!
0'
0/
#985400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#985410000000
0!
0'
0/
#985420000000
1!
1'
1/
#985430000000
0!
0'
0/
#985440000000
1!
1'
1/
#985450000000
0!
0'
0/
#985460000000
1!
1'
1/
#985470000000
0!
0'
0/
#985480000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#985490000000
0!
0'
0/
#985500000000
1!
1'
1/
#985510000000
0!
0'
0/
#985520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#985530000000
0!
0'
0/
#985540000000
1!
1'
1/
#985550000000
0!
0'
0/
#985560000000
#985570000000
1!
1'
1/
#985580000000
0!
0'
0/
#985590000000
1!
1'
1/
#985600000000
0!
1"
0'
1(
0/
10
#985610000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#985620000000
0!
0'
0/
#985630000000
1!
1'
1/
#985640000000
0!
0'
0/
#985650000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#985660000000
0!
0'
0/
#985670000000
1!
1'
1/
#985680000000
0!
1"
0'
1(
0/
10
#985690000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#985700000000
0!
1$
0'
1+
0/
#985710000000
1!
1'
1/
#985720000000
0!
0'
0/
#985730000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#985740000000
0!
0'
0/
#985750000000
1!
1'
1/
#985760000000
0!
0'
0/
#985770000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#985780000000
0!
0'
0/
#985790000000
1!
1'
1/
#985800000000
0!
0'
0/
#985810000000
1!
1'
1/
#985820000000
0!
0'
0/
#985830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#985840000000
0!
0'
0/
#985850000000
1!
1'
1/
#985860000000
0!
0'
0/
#985870000000
1!
1'
1/
#985880000000
0!
0'
0/
#985890000000
1!
1'
1/
#985900000000
0!
0'
0/
#985910000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#985920000000
0!
0'
0/
#985930000000
1!
1'
1/
#985940000000
0!
0'
0/
#985950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#985960000000
0!
0'
0/
#985970000000
1!
1'
1/
#985980000000
0!
0'
0/
#985990000000
#986000000000
1!
1'
1/
#986010000000
0!
0'
0/
#986020000000
1!
1'
1/
#986030000000
0!
1"
0'
1(
0/
10
#986040000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#986050000000
0!
0'
0/
#986060000000
1!
1'
1/
#986070000000
0!
0'
0/
#986080000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#986090000000
0!
0'
0/
#986100000000
1!
1'
1/
#986110000000
0!
1"
0'
1(
0/
10
#986120000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#986130000000
0!
1$
0'
1+
0/
#986140000000
1!
1'
1/
#986150000000
0!
0'
0/
#986160000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#986170000000
0!
0'
0/
#986180000000
1!
1'
1/
#986190000000
0!
0'
0/
#986200000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#986210000000
0!
0'
0/
#986220000000
1!
1'
1/
#986230000000
0!
0'
0/
#986240000000
1!
1'
1/
#986250000000
0!
0'
0/
#986260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#986270000000
0!
0'
0/
#986280000000
1!
1'
1/
#986290000000
0!
0'
0/
#986300000000
1!
1'
1/
#986310000000
0!
0'
0/
#986320000000
1!
1'
1/
#986330000000
0!
0'
0/
#986340000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#986350000000
0!
0'
0/
#986360000000
1!
1'
1/
#986370000000
0!
0'
0/
#986380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#986390000000
0!
0'
0/
#986400000000
1!
1'
1/
#986410000000
0!
0'
0/
#986420000000
#986430000000
1!
1'
1/
#986440000000
0!
0'
0/
#986450000000
1!
1'
1/
#986460000000
0!
1"
0'
1(
0/
10
#986470000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#986480000000
0!
0'
0/
#986490000000
1!
1'
1/
#986500000000
0!
0'
0/
#986510000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#986520000000
0!
0'
0/
#986530000000
1!
1'
1/
#986540000000
0!
1"
0'
1(
0/
10
#986550000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#986560000000
0!
1$
0'
1+
0/
#986570000000
1!
1'
1/
#986580000000
0!
0'
0/
#986590000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#986600000000
0!
0'
0/
#986610000000
1!
1'
1/
#986620000000
0!
0'
0/
#986630000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#986640000000
0!
0'
0/
#986650000000
1!
1'
1/
#986660000000
0!
0'
0/
#986670000000
1!
1'
1/
#986680000000
0!
0'
0/
#986690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#986700000000
0!
0'
0/
#986710000000
1!
1'
1/
#986720000000
0!
0'
0/
#986730000000
1!
1'
1/
#986740000000
0!
0'
0/
#986750000000
1!
1'
1/
#986760000000
0!
0'
0/
#986770000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#986780000000
0!
0'
0/
#986790000000
1!
1'
1/
#986800000000
0!
0'
0/
#986810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#986820000000
0!
0'
0/
#986830000000
1!
1'
1/
#986840000000
0!
0'
0/
#986850000000
#986860000000
1!
1'
1/
#986870000000
0!
0'
0/
#986880000000
1!
1'
1/
#986890000000
0!
1"
0'
1(
0/
10
#986900000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#986910000000
0!
0'
0/
#986920000000
1!
1'
1/
#986930000000
0!
0'
0/
#986940000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#986950000000
0!
0'
0/
#986960000000
1!
1'
1/
#986970000000
0!
1"
0'
1(
0/
10
#986980000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#986990000000
0!
1$
0'
1+
0/
#987000000000
1!
1'
1/
#987010000000
0!
0'
0/
#987020000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#987030000000
0!
0'
0/
#987040000000
1!
1'
1/
#987050000000
0!
0'
0/
#987060000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#987070000000
0!
0'
0/
#987080000000
1!
1'
1/
#987090000000
0!
0'
0/
#987100000000
1!
1'
1/
#987110000000
0!
0'
0/
#987120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#987130000000
0!
0'
0/
#987140000000
1!
1'
1/
#987150000000
0!
0'
0/
#987160000000
1!
1'
1/
#987170000000
0!
0'
0/
#987180000000
1!
1'
1/
#987190000000
0!
0'
0/
#987200000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#987210000000
0!
0'
0/
#987220000000
1!
1'
1/
#987230000000
0!
0'
0/
#987240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#987250000000
0!
0'
0/
#987260000000
1!
1'
1/
#987270000000
0!
0'
0/
#987280000000
#987290000000
1!
1'
1/
#987300000000
0!
0'
0/
#987310000000
1!
1'
1/
#987320000000
0!
1"
0'
1(
0/
10
#987330000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#987340000000
0!
0'
0/
#987350000000
1!
1'
1/
#987360000000
0!
0'
0/
#987370000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#987380000000
0!
0'
0/
#987390000000
1!
1'
1/
#987400000000
0!
1"
0'
1(
0/
10
#987410000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#987420000000
0!
1$
0'
1+
0/
#987430000000
1!
1'
1/
#987440000000
0!
0'
0/
#987450000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#987460000000
0!
0'
0/
#987470000000
1!
1'
1/
#987480000000
0!
0'
0/
#987490000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#987500000000
0!
0'
0/
#987510000000
1!
1'
1/
#987520000000
0!
0'
0/
#987530000000
1!
1'
1/
#987540000000
0!
0'
0/
#987550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#987560000000
0!
0'
0/
#987570000000
1!
1'
1/
#987580000000
0!
0'
0/
#987590000000
1!
1'
1/
#987600000000
0!
0'
0/
#987610000000
1!
1'
1/
#987620000000
0!
0'
0/
#987630000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#987640000000
0!
0'
0/
#987650000000
1!
1'
1/
#987660000000
0!
0'
0/
#987670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#987680000000
0!
0'
0/
#987690000000
1!
1'
1/
#987700000000
0!
0'
0/
#987710000000
#987720000000
1!
1'
1/
#987730000000
0!
0'
0/
#987740000000
1!
1'
1/
#987750000000
0!
1"
0'
1(
0/
10
#987760000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#987770000000
0!
0'
0/
#987780000000
1!
1'
1/
#987790000000
0!
0'
0/
#987800000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#987810000000
0!
0'
0/
#987820000000
1!
1'
1/
#987830000000
0!
1"
0'
1(
0/
10
#987840000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#987850000000
0!
1$
0'
1+
0/
#987860000000
1!
1'
1/
#987870000000
0!
0'
0/
#987880000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#987890000000
0!
0'
0/
#987900000000
1!
1'
1/
#987910000000
0!
0'
0/
#987920000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#987930000000
0!
0'
0/
#987940000000
1!
1'
1/
#987950000000
0!
0'
0/
#987960000000
1!
1'
1/
#987970000000
0!
0'
0/
#987980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#987990000000
0!
0'
0/
#988000000000
1!
1'
1/
#988010000000
0!
0'
0/
#988020000000
1!
1'
1/
#988030000000
0!
0'
0/
#988040000000
1!
1'
1/
#988050000000
0!
0'
0/
#988060000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#988070000000
0!
0'
0/
#988080000000
1!
1'
1/
#988090000000
0!
0'
0/
#988100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#988110000000
0!
0'
0/
#988120000000
1!
1'
1/
#988130000000
0!
0'
0/
#988140000000
#988150000000
1!
1'
1/
#988160000000
0!
0'
0/
#988170000000
1!
1'
1/
#988180000000
0!
1"
0'
1(
0/
10
#988190000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#988200000000
0!
0'
0/
#988210000000
1!
1'
1/
#988220000000
0!
0'
0/
#988230000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#988240000000
0!
0'
0/
#988250000000
1!
1'
1/
#988260000000
0!
1"
0'
1(
0/
10
#988270000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#988280000000
0!
1$
0'
1+
0/
#988290000000
1!
1'
1/
#988300000000
0!
0'
0/
#988310000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#988320000000
0!
0'
0/
#988330000000
1!
1'
1/
#988340000000
0!
0'
0/
#988350000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#988360000000
0!
0'
0/
#988370000000
1!
1'
1/
#988380000000
0!
0'
0/
#988390000000
1!
1'
1/
#988400000000
0!
0'
0/
#988410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#988420000000
0!
0'
0/
#988430000000
1!
1'
1/
#988440000000
0!
0'
0/
#988450000000
1!
1'
1/
#988460000000
0!
0'
0/
#988470000000
1!
1'
1/
#988480000000
0!
0'
0/
#988490000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#988500000000
0!
0'
0/
#988510000000
1!
1'
1/
#988520000000
0!
0'
0/
#988530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#988540000000
0!
0'
0/
#988550000000
1!
1'
1/
#988560000000
0!
0'
0/
#988570000000
#988580000000
1!
1'
1/
#988590000000
0!
0'
0/
#988600000000
1!
1'
1/
#988610000000
0!
1"
0'
1(
0/
10
#988620000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#988630000000
0!
0'
0/
#988640000000
1!
1'
1/
#988650000000
0!
0'
0/
#988660000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#988670000000
0!
0'
0/
#988680000000
1!
1'
1/
#988690000000
0!
1"
0'
1(
0/
10
#988700000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#988710000000
0!
1$
0'
1+
0/
#988720000000
1!
1'
1/
#988730000000
0!
0'
0/
#988740000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#988750000000
0!
0'
0/
#988760000000
1!
1'
1/
#988770000000
0!
0'
0/
#988780000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#988790000000
0!
0'
0/
#988800000000
1!
1'
1/
#988810000000
0!
0'
0/
#988820000000
1!
1'
1/
#988830000000
0!
0'
0/
#988840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#988850000000
0!
0'
0/
#988860000000
1!
1'
1/
#988870000000
0!
0'
0/
#988880000000
1!
1'
1/
#988890000000
0!
0'
0/
#988900000000
1!
1'
1/
#988910000000
0!
0'
0/
#988920000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#988930000000
0!
0'
0/
#988940000000
1!
1'
1/
#988950000000
0!
0'
0/
#988960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#988970000000
0!
0'
0/
#988980000000
1!
1'
1/
#988990000000
0!
0'
0/
#989000000000
#989010000000
1!
1'
1/
#989020000000
0!
0'
0/
#989030000000
1!
1'
1/
#989040000000
0!
1"
0'
1(
0/
10
#989050000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#989060000000
0!
0'
0/
#989070000000
1!
1'
1/
#989080000000
0!
0'
0/
#989090000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#989100000000
0!
0'
0/
#989110000000
1!
1'
1/
#989120000000
0!
1"
0'
1(
0/
10
#989130000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#989140000000
0!
1$
0'
1+
0/
#989150000000
1!
1'
1/
#989160000000
0!
0'
0/
#989170000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#989180000000
0!
0'
0/
#989190000000
1!
1'
1/
#989200000000
0!
0'
0/
#989210000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#989220000000
0!
0'
0/
#989230000000
1!
1'
1/
#989240000000
0!
0'
0/
#989250000000
1!
1'
1/
#989260000000
0!
0'
0/
#989270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#989280000000
0!
0'
0/
#989290000000
1!
1'
1/
#989300000000
0!
0'
0/
#989310000000
1!
1'
1/
#989320000000
0!
0'
0/
#989330000000
1!
1'
1/
#989340000000
0!
0'
0/
#989350000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#989360000000
0!
0'
0/
#989370000000
1!
1'
1/
#989380000000
0!
0'
0/
#989390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#989400000000
0!
0'
0/
#989410000000
1!
1'
1/
#989420000000
0!
0'
0/
#989430000000
#989440000000
1!
1'
1/
#989450000000
0!
0'
0/
#989460000000
1!
1'
1/
#989470000000
0!
1"
0'
1(
0/
10
#989480000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#989490000000
0!
0'
0/
#989500000000
1!
1'
1/
#989510000000
0!
0'
0/
#989520000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#989530000000
0!
0'
0/
#989540000000
1!
1'
1/
#989550000000
0!
1"
0'
1(
0/
10
#989560000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#989570000000
0!
1$
0'
1+
0/
#989580000000
1!
1'
1/
#989590000000
0!
0'
0/
#989600000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#989610000000
0!
0'
0/
#989620000000
1!
1'
1/
#989630000000
0!
0'
0/
#989640000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#989650000000
0!
0'
0/
#989660000000
1!
1'
1/
#989670000000
0!
0'
0/
#989680000000
1!
1'
1/
#989690000000
0!
0'
0/
#989700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#989710000000
0!
0'
0/
#989720000000
1!
1'
1/
#989730000000
0!
0'
0/
#989740000000
1!
1'
1/
#989750000000
0!
0'
0/
#989760000000
1!
1'
1/
#989770000000
0!
0'
0/
#989780000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#989790000000
0!
0'
0/
#989800000000
1!
1'
1/
#989810000000
0!
0'
0/
#989820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#989830000000
0!
0'
0/
#989840000000
1!
1'
1/
#989850000000
0!
0'
0/
#989860000000
#989870000000
1!
1'
1/
#989880000000
0!
0'
0/
#989890000000
1!
1'
1/
#989900000000
0!
1"
0'
1(
0/
10
#989910000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#989920000000
0!
0'
0/
#989930000000
1!
1'
1/
#989940000000
0!
0'
0/
#989950000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#989960000000
0!
0'
0/
#989970000000
1!
1'
1/
#989980000000
0!
1"
0'
1(
0/
10
#989990000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#990000000000
0!
1$
0'
1+
0/
#990010000000
1!
1'
1/
#990020000000
0!
0'
0/
#990030000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#990040000000
0!
0'
0/
#990050000000
1!
1'
1/
#990060000000
0!
0'
0/
#990070000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#990080000000
0!
0'
0/
#990090000000
1!
1'
1/
#990100000000
0!
0'
0/
#990110000000
1!
1'
1/
#990120000000
0!
0'
0/
#990130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#990140000000
0!
0'
0/
#990150000000
1!
1'
1/
#990160000000
0!
0'
0/
#990170000000
1!
1'
1/
#990180000000
0!
0'
0/
#990190000000
1!
1'
1/
#990200000000
0!
0'
0/
#990210000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#990220000000
0!
0'
0/
#990230000000
1!
1'
1/
#990240000000
0!
0'
0/
#990250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#990260000000
0!
0'
0/
#990270000000
1!
1'
1/
#990280000000
0!
0'
0/
#990290000000
#990300000000
1!
1'
1/
#990310000000
0!
0'
0/
#990320000000
1!
1'
1/
#990330000000
0!
1"
0'
1(
0/
10
#990340000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#990350000000
0!
0'
0/
#990360000000
1!
1'
1/
#990370000000
0!
0'
0/
#990380000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#990390000000
0!
0'
0/
#990400000000
1!
1'
1/
#990410000000
0!
1"
0'
1(
0/
10
#990420000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#990430000000
0!
1$
0'
1+
0/
#990440000000
1!
1'
1/
#990450000000
0!
0'
0/
#990460000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#990470000000
0!
0'
0/
#990480000000
1!
1'
1/
#990490000000
0!
0'
0/
#990500000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#990510000000
0!
0'
0/
#990520000000
1!
1'
1/
#990530000000
0!
0'
0/
#990540000000
1!
1'
1/
#990550000000
0!
0'
0/
#990560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#990570000000
0!
0'
0/
#990580000000
1!
1'
1/
#990590000000
0!
0'
0/
#990600000000
1!
1'
1/
#990610000000
0!
0'
0/
#990620000000
1!
1'
1/
#990630000000
0!
0'
0/
#990640000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#990650000000
0!
0'
0/
#990660000000
1!
1'
1/
#990670000000
0!
0'
0/
#990680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#990690000000
0!
0'
0/
#990700000000
1!
1'
1/
#990710000000
0!
0'
0/
#990720000000
#990730000000
1!
1'
1/
#990740000000
0!
0'
0/
#990750000000
1!
1'
1/
#990760000000
0!
1"
0'
1(
0/
10
#990770000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#990780000000
0!
0'
0/
#990790000000
1!
1'
1/
#990800000000
0!
0'
0/
#990810000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#990820000000
0!
0'
0/
#990830000000
1!
1'
1/
#990840000000
0!
1"
0'
1(
0/
10
#990850000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#990860000000
0!
1$
0'
1+
0/
#990870000000
1!
1'
1/
#990880000000
0!
0'
0/
#990890000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#990900000000
0!
0'
0/
#990910000000
1!
1'
1/
#990920000000
0!
0'
0/
#990930000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#990940000000
0!
0'
0/
#990950000000
1!
1'
1/
#990960000000
0!
0'
0/
#990970000000
1!
1'
1/
#990980000000
0!
0'
0/
#990990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#991000000000
0!
0'
0/
#991010000000
1!
1'
1/
#991020000000
0!
0'
0/
#991030000000
1!
1'
1/
#991040000000
0!
0'
0/
#991050000000
1!
1'
1/
#991060000000
0!
0'
0/
#991070000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#991080000000
0!
0'
0/
#991090000000
1!
1'
1/
#991100000000
0!
0'
0/
#991110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#991120000000
0!
0'
0/
#991130000000
1!
1'
1/
#991140000000
0!
0'
0/
#991150000000
#991160000000
1!
1'
1/
#991170000000
0!
0'
0/
#991180000000
1!
1'
1/
#991190000000
0!
1"
0'
1(
0/
10
#991200000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#991210000000
0!
0'
0/
#991220000000
1!
1'
1/
#991230000000
0!
0'
0/
#991240000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#991250000000
0!
0'
0/
#991260000000
1!
1'
1/
#991270000000
0!
1"
0'
1(
0/
10
#991280000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#991290000000
0!
1$
0'
1+
0/
#991300000000
1!
1'
1/
#991310000000
0!
0'
0/
#991320000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#991330000000
0!
0'
0/
#991340000000
1!
1'
1/
#991350000000
0!
0'
0/
#991360000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#991370000000
0!
0'
0/
#991380000000
1!
1'
1/
#991390000000
0!
0'
0/
#991400000000
1!
1'
1/
#991410000000
0!
0'
0/
#991420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#991430000000
0!
0'
0/
#991440000000
1!
1'
1/
#991450000000
0!
0'
0/
#991460000000
1!
1'
1/
#991470000000
0!
0'
0/
#991480000000
1!
1'
1/
#991490000000
0!
0'
0/
#991500000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#991510000000
0!
0'
0/
#991520000000
1!
1'
1/
#991530000000
0!
0'
0/
#991540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#991550000000
0!
0'
0/
#991560000000
1!
1'
1/
#991570000000
0!
0'
0/
#991580000000
#991590000000
1!
1'
1/
#991600000000
0!
0'
0/
#991610000000
1!
1'
1/
#991620000000
0!
1"
0'
1(
0/
10
#991630000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#991640000000
0!
0'
0/
#991650000000
1!
1'
1/
#991660000000
0!
0'
0/
#991670000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#991680000000
0!
0'
0/
#991690000000
1!
1'
1/
#991700000000
0!
1"
0'
1(
0/
10
#991710000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#991720000000
0!
1$
0'
1+
0/
#991730000000
1!
1'
1/
#991740000000
0!
0'
0/
#991750000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#991760000000
0!
0'
0/
#991770000000
1!
1'
1/
#991780000000
0!
0'
0/
#991790000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#991800000000
0!
0'
0/
#991810000000
1!
1'
1/
#991820000000
0!
0'
0/
#991830000000
1!
1'
1/
#991840000000
0!
0'
0/
#991850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#991860000000
0!
0'
0/
#991870000000
1!
1'
1/
#991880000000
0!
0'
0/
#991890000000
1!
1'
1/
#991900000000
0!
0'
0/
#991910000000
1!
1'
1/
#991920000000
0!
0'
0/
#991930000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#991940000000
0!
0'
0/
#991950000000
1!
1'
1/
#991960000000
0!
0'
0/
#991970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#991980000000
0!
0'
0/
#991990000000
1!
1'
1/
#992000000000
0!
0'
0/
#992010000000
#992020000000
1!
1'
1/
#992030000000
0!
0'
0/
#992040000000
1!
1'
1/
#992050000000
0!
1"
0'
1(
0/
10
#992060000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#992070000000
0!
0'
0/
#992080000000
1!
1'
1/
#992090000000
0!
0'
0/
#992100000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#992110000000
0!
0'
0/
#992120000000
1!
1'
1/
#992130000000
0!
1"
0'
1(
0/
10
#992140000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#992150000000
0!
1$
0'
1+
0/
#992160000000
1!
1'
1/
#992170000000
0!
0'
0/
#992180000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#992190000000
0!
0'
0/
#992200000000
1!
1'
1/
#992210000000
0!
0'
0/
#992220000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#992230000000
0!
0'
0/
#992240000000
1!
1'
1/
#992250000000
0!
0'
0/
#992260000000
1!
1'
1/
#992270000000
0!
0'
0/
#992280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#992290000000
0!
0'
0/
#992300000000
1!
1'
1/
#992310000000
0!
0'
0/
#992320000000
1!
1'
1/
#992330000000
0!
0'
0/
#992340000000
1!
1'
1/
#992350000000
0!
0'
0/
#992360000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#992370000000
0!
0'
0/
#992380000000
1!
1'
1/
#992390000000
0!
0'
0/
#992400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#992410000000
0!
0'
0/
#992420000000
1!
1'
1/
#992430000000
0!
0'
0/
#992440000000
#992450000000
1!
1'
1/
#992460000000
0!
0'
0/
#992470000000
1!
1'
1/
#992480000000
0!
1"
0'
1(
0/
10
#992490000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#992500000000
0!
0'
0/
#992510000000
1!
1'
1/
#992520000000
0!
0'
0/
#992530000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#992540000000
0!
0'
0/
#992550000000
1!
1'
1/
#992560000000
0!
1"
0'
1(
0/
10
#992570000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#992580000000
0!
1$
0'
1+
0/
#992590000000
1!
1'
1/
#992600000000
0!
0'
0/
#992610000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#992620000000
0!
0'
0/
#992630000000
1!
1'
1/
#992640000000
0!
0'
0/
#992650000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#992660000000
0!
0'
0/
#992670000000
1!
1'
1/
#992680000000
0!
0'
0/
#992690000000
1!
1'
1/
#992700000000
0!
0'
0/
#992710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#992720000000
0!
0'
0/
#992730000000
1!
1'
1/
#992740000000
0!
0'
0/
#992750000000
1!
1'
1/
#992760000000
0!
0'
0/
#992770000000
1!
1'
1/
#992780000000
0!
0'
0/
#992790000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#992800000000
0!
0'
0/
#992810000000
1!
1'
1/
#992820000000
0!
0'
0/
#992830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#992840000000
0!
0'
0/
#992850000000
1!
1'
1/
#992860000000
0!
0'
0/
#992870000000
#992880000000
1!
1'
1/
#992890000000
0!
0'
0/
#992900000000
1!
1'
1/
#992910000000
0!
1"
0'
1(
0/
10
#992920000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#992930000000
0!
0'
0/
#992940000000
1!
1'
1/
#992950000000
0!
0'
0/
#992960000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#992970000000
0!
0'
0/
#992980000000
1!
1'
1/
#992990000000
0!
1"
0'
1(
0/
10
#993000000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#993010000000
0!
1$
0'
1+
0/
#993020000000
1!
1'
1/
#993030000000
0!
0'
0/
#993040000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#993050000000
0!
0'
0/
#993060000000
1!
1'
1/
#993070000000
0!
0'
0/
#993080000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#993090000000
0!
0'
0/
#993100000000
1!
1'
1/
#993110000000
0!
0'
0/
#993120000000
1!
1'
1/
#993130000000
0!
0'
0/
#993140000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#993150000000
0!
0'
0/
#993160000000
1!
1'
1/
#993170000000
0!
0'
0/
#993180000000
1!
1'
1/
#993190000000
0!
0'
0/
#993200000000
1!
1'
1/
#993210000000
0!
0'
0/
#993220000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#993230000000
0!
0'
0/
#993240000000
1!
1'
1/
#993250000000
0!
0'
0/
#993260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#993270000000
0!
0'
0/
#993280000000
1!
1'
1/
#993290000000
0!
0'
0/
#993300000000
#993310000000
1!
1'
1/
#993320000000
0!
0'
0/
#993330000000
1!
1'
1/
#993340000000
0!
1"
0'
1(
0/
10
#993350000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#993360000000
0!
0'
0/
#993370000000
1!
1'
1/
#993380000000
0!
0'
0/
#993390000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#993400000000
0!
0'
0/
#993410000000
1!
1'
1/
#993420000000
0!
1"
0'
1(
0/
10
#993430000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#993440000000
0!
1$
0'
1+
0/
#993450000000
1!
1'
1/
#993460000000
0!
0'
0/
#993470000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#993480000000
0!
0'
0/
#993490000000
1!
1'
1/
#993500000000
0!
0'
0/
#993510000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#993520000000
0!
0'
0/
#993530000000
1!
1'
1/
#993540000000
0!
0'
0/
#993550000000
1!
1'
1/
#993560000000
0!
0'
0/
#993570000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#993580000000
0!
0'
0/
#993590000000
1!
1'
1/
#993600000000
0!
0'
0/
#993610000000
1!
1'
1/
#993620000000
0!
0'
0/
#993630000000
1!
1'
1/
#993640000000
0!
0'
0/
#993650000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#993660000000
0!
0'
0/
#993670000000
1!
1'
1/
#993680000000
0!
0'
0/
#993690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#993700000000
0!
0'
0/
#993710000000
1!
1'
1/
#993720000000
0!
0'
0/
#993730000000
#993740000000
1!
1'
1/
#993750000000
0!
0'
0/
#993760000000
1!
1'
1/
#993770000000
0!
1"
0'
1(
0/
10
#993780000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#993790000000
0!
0'
0/
#993800000000
1!
1'
1/
#993810000000
0!
0'
0/
#993820000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#993830000000
0!
0'
0/
#993840000000
1!
1'
1/
#993850000000
0!
1"
0'
1(
0/
10
#993860000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#993870000000
0!
1$
0'
1+
0/
#993880000000
1!
1'
1/
#993890000000
0!
0'
0/
#993900000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#993910000000
0!
0'
0/
#993920000000
1!
1'
1/
#993930000000
0!
0'
0/
#993940000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#993950000000
0!
0'
0/
#993960000000
1!
1'
1/
#993970000000
0!
0'
0/
#993980000000
1!
1'
1/
#993990000000
0!
0'
0/
#994000000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#994010000000
0!
0'
0/
#994020000000
1!
1'
1/
#994030000000
0!
0'
0/
#994040000000
1!
1'
1/
#994050000000
0!
0'
0/
#994060000000
1!
1'
1/
#994070000000
0!
0'
0/
#994080000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#994090000000
0!
0'
0/
#994100000000
1!
1'
1/
#994110000000
0!
0'
0/
#994120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#994130000000
0!
0'
0/
#994140000000
1!
1'
1/
#994150000000
0!
0'
0/
#994160000000
#994170000000
1!
1'
1/
#994180000000
0!
0'
0/
#994190000000
1!
1'
1/
#994200000000
0!
1"
0'
1(
0/
10
#994210000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#994220000000
0!
0'
0/
#994230000000
1!
1'
1/
#994240000000
0!
0'
0/
#994250000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#994260000000
0!
0'
0/
#994270000000
1!
1'
1/
#994280000000
0!
1"
0'
1(
0/
10
#994290000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#994300000000
0!
1$
0'
1+
0/
#994310000000
1!
1'
1/
#994320000000
0!
0'
0/
#994330000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#994340000000
0!
0'
0/
#994350000000
1!
1'
1/
#994360000000
0!
0'
0/
#994370000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#994380000000
0!
0'
0/
#994390000000
1!
1'
1/
#994400000000
0!
0'
0/
#994410000000
1!
1'
1/
#994420000000
0!
0'
0/
#994430000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#994440000000
0!
0'
0/
#994450000000
1!
1'
1/
#994460000000
0!
0'
0/
#994470000000
1!
1'
1/
#994480000000
0!
0'
0/
#994490000000
1!
1'
1/
#994500000000
0!
0'
0/
#994510000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#994520000000
0!
0'
0/
#994530000000
1!
1'
1/
#994540000000
0!
0'
0/
#994550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#994560000000
0!
0'
0/
#994570000000
1!
1'
1/
#994580000000
0!
0'
0/
#994590000000
#994600000000
1!
1'
1/
#994610000000
0!
0'
0/
#994620000000
1!
1'
1/
#994630000000
0!
1"
0'
1(
0/
10
#994640000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#994650000000
0!
0'
0/
#994660000000
1!
1'
1/
#994670000000
0!
0'
0/
#994680000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#994690000000
0!
0'
0/
#994700000000
1!
1'
1/
#994710000000
0!
1"
0'
1(
0/
10
#994720000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#994730000000
0!
1$
0'
1+
0/
#994740000000
1!
1'
1/
#994750000000
0!
0'
0/
#994760000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#994770000000
0!
0'
0/
#994780000000
1!
1'
1/
#994790000000
0!
0'
0/
#994800000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#994810000000
0!
0'
0/
#994820000000
1!
1'
1/
#994830000000
0!
0'
0/
#994840000000
1!
1'
1/
#994850000000
0!
0'
0/
#994860000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#994870000000
0!
0'
0/
#994880000000
1!
1'
1/
#994890000000
0!
0'
0/
#994900000000
1!
1'
1/
#994910000000
0!
0'
0/
#994920000000
1!
1'
1/
#994930000000
0!
0'
0/
#994940000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#994950000000
0!
0'
0/
#994960000000
1!
1'
1/
#994970000000
0!
0'
0/
#994980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#994990000000
0!
0'
0/
#995000000000
1!
1'
1/
#995010000000
0!
0'
0/
#995020000000
#995030000000
1!
1'
1/
#995040000000
0!
0'
0/
#995050000000
1!
1'
1/
#995060000000
0!
1"
0'
1(
0/
10
#995070000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#995080000000
0!
0'
0/
#995090000000
1!
1'
1/
#995100000000
0!
0'
0/
#995110000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#995120000000
0!
0'
0/
#995130000000
1!
1'
1/
#995140000000
0!
1"
0'
1(
0/
10
#995150000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#995160000000
0!
1$
0'
1+
0/
#995170000000
1!
1'
1/
#995180000000
0!
0'
0/
#995190000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#995200000000
0!
0'
0/
#995210000000
1!
1'
1/
#995220000000
0!
0'
0/
#995230000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#995240000000
0!
0'
0/
#995250000000
1!
1'
1/
#995260000000
0!
0'
0/
#995270000000
1!
1'
1/
#995280000000
0!
0'
0/
#995290000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#995300000000
0!
0'
0/
#995310000000
1!
1'
1/
#995320000000
0!
0'
0/
#995330000000
1!
1'
1/
#995340000000
0!
0'
0/
#995350000000
1!
1'
1/
#995360000000
0!
0'
0/
#995370000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#995380000000
0!
0'
0/
#995390000000
1!
1'
1/
#995400000000
0!
0'
0/
#995410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#995420000000
0!
0'
0/
#995430000000
1!
1'
1/
#995440000000
0!
0'
0/
#995450000000
#995460000000
1!
1'
1/
#995470000000
0!
0'
0/
#995480000000
1!
1'
1/
#995490000000
0!
1"
0'
1(
0/
10
#995500000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#995510000000
0!
0'
0/
#995520000000
1!
1'
1/
#995530000000
0!
0'
0/
#995540000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#995550000000
0!
0'
0/
#995560000000
1!
1'
1/
#995570000000
0!
1"
0'
1(
0/
10
#995580000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#995590000000
0!
1$
0'
1+
0/
#995600000000
1!
1'
1/
#995610000000
0!
0'
0/
#995620000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#995630000000
0!
0'
0/
#995640000000
1!
1'
1/
#995650000000
0!
0'
0/
#995660000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#995670000000
0!
0'
0/
#995680000000
1!
1'
1/
#995690000000
0!
0'
0/
#995700000000
1!
1'
1/
#995710000000
0!
0'
0/
#995720000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#995730000000
0!
0'
0/
#995740000000
1!
1'
1/
#995750000000
0!
0'
0/
#995760000000
1!
1'
1/
#995770000000
0!
0'
0/
#995780000000
1!
1'
1/
#995790000000
0!
0'
0/
#995800000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#995810000000
0!
0'
0/
#995820000000
1!
1'
1/
#995830000000
0!
0'
0/
#995840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#995850000000
0!
0'
0/
#995860000000
1!
1'
1/
#995870000000
0!
0'
0/
#995880000000
#995890000000
1!
1'
1/
#995900000000
0!
0'
0/
#995910000000
1!
1'
1/
#995920000000
0!
1"
0'
1(
0/
10
#995930000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#995940000000
0!
0'
0/
#995950000000
1!
1'
1/
#995960000000
0!
0'
0/
#995970000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#995980000000
0!
0'
0/
#995990000000
1!
1'
1/
#996000000000
0!
1"
0'
1(
0/
10
#996010000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#996020000000
0!
1$
0'
1+
0/
#996030000000
1!
1'
1/
#996040000000
0!
0'
0/
#996050000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#996060000000
0!
0'
0/
#996070000000
1!
1'
1/
#996080000000
0!
0'
0/
#996090000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#996100000000
0!
0'
0/
#996110000000
1!
1'
1/
#996120000000
0!
0'
0/
#996130000000
1!
1'
1/
#996140000000
0!
0'
0/
#996150000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#996160000000
0!
0'
0/
#996170000000
1!
1'
1/
#996180000000
0!
0'
0/
#996190000000
1!
1'
1/
#996200000000
0!
0'
0/
#996210000000
1!
1'
1/
#996220000000
0!
0'
0/
#996230000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#996240000000
0!
0'
0/
#996250000000
1!
1'
1/
#996260000000
0!
0'
0/
#996270000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#996280000000
0!
0'
0/
#996290000000
1!
1'
1/
#996300000000
0!
0'
0/
#996310000000
#996320000000
1!
1'
1/
#996330000000
0!
0'
0/
#996340000000
1!
1'
1/
#996350000000
0!
1"
0'
1(
0/
10
#996360000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#996370000000
0!
0'
0/
#996380000000
1!
1'
1/
#996390000000
0!
0'
0/
#996400000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#996410000000
0!
0'
0/
#996420000000
1!
1'
1/
#996430000000
0!
1"
0'
1(
0/
10
#996440000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#996450000000
0!
1$
0'
1+
0/
#996460000000
1!
1'
1/
#996470000000
0!
0'
0/
#996480000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#996490000000
0!
0'
0/
#996500000000
1!
1'
1/
#996510000000
0!
0'
0/
#996520000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#996530000000
0!
0'
0/
#996540000000
1!
1'
1/
#996550000000
0!
0'
0/
#996560000000
1!
1'
1/
#996570000000
0!
0'
0/
#996580000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#996590000000
0!
0'
0/
#996600000000
1!
1'
1/
#996610000000
0!
0'
0/
#996620000000
1!
1'
1/
#996630000000
0!
0'
0/
#996640000000
1!
1'
1/
#996650000000
0!
0'
0/
#996660000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#996670000000
0!
0'
0/
#996680000000
1!
1'
1/
#996690000000
0!
0'
0/
#996700000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#996710000000
0!
0'
0/
#996720000000
1!
1'
1/
#996730000000
0!
0'
0/
#996740000000
#996750000000
1!
1'
1/
#996760000000
0!
0'
0/
#996770000000
1!
1'
1/
#996780000000
0!
1"
0'
1(
0/
10
#996790000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#996800000000
0!
0'
0/
#996810000000
1!
1'
1/
#996820000000
0!
0'
0/
#996830000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#996840000000
0!
0'
0/
#996850000000
1!
1'
1/
#996860000000
0!
1"
0'
1(
0/
10
#996870000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#996880000000
0!
1$
0'
1+
0/
#996890000000
1!
1'
1/
#996900000000
0!
0'
0/
#996910000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#996920000000
0!
0'
0/
#996930000000
1!
1'
1/
#996940000000
0!
0'
0/
#996950000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#996960000000
0!
0'
0/
#996970000000
1!
1'
1/
#996980000000
0!
0'
0/
#996990000000
1!
1'
1/
#997000000000
0!
0'
0/
#997010000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#997020000000
0!
0'
0/
#997030000000
1!
1'
1/
#997040000000
0!
0'
0/
#997050000000
1!
1'
1/
#997060000000
0!
0'
0/
#997070000000
1!
1'
1/
#997080000000
0!
0'
0/
#997090000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#997100000000
0!
0'
0/
#997110000000
1!
1'
1/
#997120000000
0!
0'
0/
#997130000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#997140000000
0!
0'
0/
#997150000000
1!
1'
1/
#997160000000
0!
0'
0/
#997170000000
#997180000000
1!
1'
1/
#997190000000
0!
0'
0/
#997200000000
1!
1'
1/
#997210000000
0!
1"
0'
1(
0/
10
#997220000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#997230000000
0!
0'
0/
#997240000000
1!
1'
1/
#997250000000
0!
0'
0/
#997260000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#997270000000
0!
0'
0/
#997280000000
1!
1'
1/
#997290000000
0!
1"
0'
1(
0/
10
#997300000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#997310000000
0!
1$
0'
1+
0/
#997320000000
1!
1'
1/
#997330000000
0!
0'
0/
#997340000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#997350000000
0!
0'
0/
#997360000000
1!
1'
1/
#997370000000
0!
0'
0/
#997380000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#997390000000
0!
0'
0/
#997400000000
1!
1'
1/
#997410000000
0!
0'
0/
#997420000000
1!
1'
1/
#997430000000
0!
0'
0/
#997440000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#997450000000
0!
0'
0/
#997460000000
1!
1'
1/
#997470000000
0!
0'
0/
#997480000000
1!
1'
1/
#997490000000
0!
0'
0/
#997500000000
1!
1'
1/
#997510000000
0!
0'
0/
#997520000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#997530000000
0!
0'
0/
#997540000000
1!
1'
1/
#997550000000
0!
0'
0/
#997560000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#997570000000
0!
0'
0/
#997580000000
1!
1'
1/
#997590000000
0!
0'
0/
#997600000000
#997610000000
1!
1'
1/
#997620000000
0!
0'
0/
#997630000000
1!
1'
1/
#997640000000
0!
1"
0'
1(
0/
10
#997650000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#997660000000
0!
0'
0/
#997670000000
1!
1'
1/
#997680000000
0!
0'
0/
#997690000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#997700000000
0!
0'
0/
#997710000000
1!
1'
1/
#997720000000
0!
1"
0'
1(
0/
10
#997730000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#997740000000
0!
1$
0'
1+
0/
#997750000000
1!
1'
1/
#997760000000
0!
0'
0/
#997770000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#997780000000
0!
0'
0/
#997790000000
1!
1'
1/
#997800000000
0!
0'
0/
#997810000000
1!
1"
b0110000 &
1'
1(
b0110000 )
1-
b0001 .
1/
10
11
12
13
b0110000 4
b0001 5
#997820000000
0!
0'
0/
#997830000000
1!
1'
1/
#997840000000
0!
0'
0/
#997850000000
1!
1'
1/
#997860000000
0!
0'
0/
#997870000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#997880000000
0!
0'
0/
#997890000000
1!
1'
1/
#997900000000
0!
0'
0/
#997910000000
1!
1'
1/
#997920000000
0!
0'
0/
#997930000000
1!
1'
1/
#997940000000
0!
0'
0/
#997950000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#997960000000
0!
0'
0/
#997970000000
1!
1'
1/
#997980000000
0!
0'
0/
#997990000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#998000000000
0!
0'
0/
#998010000000
1!
1'
1/
#998020000000
0!
0'
0/
#998030000000
#998040000000
1!
1'
1/
#998050000000
0!
0'
0/
#998060000000
1!
1'
1/
#998070000000
0!
1"
0'
1(
0/
10
#998080000000
1!
b1111001 &
1'
b1111001 )
1-
b0011 .
1/
11
12
13
b1111001 4
b0011 5
#998090000000
0!
0'
0/
#998100000000
1!
1'
1/
#998110000000
0!
0'
0/
#998120000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#998130000000
0!
0'
0/
#998140000000
1!
1'
1/
#998150000000
0!
1"
0'
1(
0/
10
#998160000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#998170000000
0!
1$
0'
1+
0/
#998180000000
1!
1'
1/
#998190000000
0!
0'
0/
#998200000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#998210000000
0!
0'
0/
#998220000000
1!
1'
1/
#998230000000
0!
0'
0/
#998240000000
1!
1"
b1011011 &
1'
1(
b1011011 )
1-
b0101 .
1/
10
11
12
13
b1011011 4
b0101 5
#998250000000
0!
0'
0/
#998260000000
1!
1'
1/
#998270000000
0!
0'
0/
#998280000000
1!
1'
1/
#998290000000
0!
0'
0/
#998300000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#998310000000
0!
0'
0/
#998320000000
1!
1'
1/
#998330000000
0!
0'
0/
#998340000000
1!
1'
1/
#998350000000
0!
0'
0/
#998360000000
1!
1'
1/
#998370000000
0!
0'
0/
#998380000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#998390000000
0!
0'
0/
#998400000000
1!
1'
1/
#998410000000
0!
0'
0/
#998420000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#998430000000
0!
0'
0/
#998440000000
1!
1'
1/
#998450000000
0!
0'
0/
#998460000000
#998470000000
1!
1'
1/
#998480000000
0!
0'
0/
#998490000000
1!
1'
1/
#998500000000
0!
1"
0'
1(
0/
10
#998510000000
1!
0%
b1111110 &
1'
b1111110 )
0,
1-
b0000 .
1/
11
12
13
b1111110 4
b0000 5
#998520000000
0!
0'
0/
#998530000000
1!
1'
1/
#998540000000
0!
0'
0/
#998550000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#998560000000
0!
0'
0/
#998570000000
1!
1'
1/
#998580000000
0!
1"
0'
1(
0/
10
#998590000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#998600000000
0!
1$
0'
1+
0/
#998610000000
1!
1'
1/
#998620000000
0!
0'
0/
#998630000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#998640000000
0!
0'
0/
#998650000000
1!
1'
1/
#998660000000
0!
0'
0/
#998670000000
1!
1"
b1101101 &
1'
1(
b1101101 )
1-
b0010 .
1/
10
11
12
13
b1101101 4
b0010 5
#998680000000
0!
0'
0/
#998690000000
1!
1'
1/
#998700000000
0!
0'
0/
#998710000000
1!
1'
1/
#998720000000
0!
0'
0/
#998730000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#998740000000
0!
0'
0/
#998750000000
1!
1'
1/
#998760000000
0!
0'
0/
#998770000000
1!
1'
1/
#998780000000
0!
0'
0/
#998790000000
1!
1'
1/
#998800000000
0!
0'
0/
#998810000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#998820000000
0!
0'
0/
#998830000000
1!
1'
1/
#998840000000
0!
0'
0/
#998850000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#998860000000
0!
0'
0/
#998870000000
1!
1'
1/
#998880000000
0!
0'
0/
#998890000000
#998900000000
1!
1'
1/
#998910000000
0!
0'
0/
#998920000000
1!
1'
1/
#998930000000
0!
1"
0'
1(
0/
10
#998940000000
1!
b0110011 &
1'
b0110011 )
1-
b0100 .
1/
11
12
13
b0110011 4
b0100 5
#998950000000
0!
0'
0/
#998960000000
1!
1'
1/
#998970000000
0!
0'
0/
#998980000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#998990000000
0!
0'
0/
#999000000000
1!
1'
1/
#999010000000
0!
1"
0'
1(
0/
10
#999020000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#999030000000
0!
1$
0'
1+
0/
#999040000000
1!
1'
1/
#999050000000
0!
0'
0/
#999060000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#999070000000
0!
0'
0/
#999080000000
1!
1'
1/
#999090000000
0!
0'
0/
#999100000000
1!
1"
1%
b1011111 &
1'
1(
b1011111 )
1,
1-
b0110 .
1/
10
11
12
13
b1011111 4
b0110 5
#999110000000
0!
0'
0/
#999120000000
1!
1'
1/
#999130000000
0!
0'
0/
#999140000000
1!
1'
1/
#999150000000
0!
0'
0/
#999160000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#999170000000
0!
0'
0/
#999180000000
1!
1'
1/
#999190000000
0!
0'
0/
#999200000000
1!
1'
1/
#999210000000
0!
0'
0/
#999220000000
1!
1'
1/
#999230000000
0!
0'
0/
#999240000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#999250000000
0!
0'
0/
#999260000000
1!
1'
1/
#999270000000
0!
0'
0/
#999280000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#999290000000
0!
0'
0/
#999300000000
1!
1'
1/
#999310000000
0!
0'
0/
#999320000000
#999330000000
1!
1'
1/
#999340000000
0!
0'
0/
#999350000000
1!
1'
1/
#999360000000
0!
1"
0'
1(
0/
10
#999370000000
1!
b0110000 &
1'
b0110000 )
1-
b0001 .
1/
11
12
13
b0110000 4
b0001 5
#999380000000
0!
0'
0/
#999390000000
1!
1'
1/
#999400000000
0!
0'
0/
#999410000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#999420000000
0!
0'
0/
#999430000000
1!
1'
1/
#999440000000
0!
1"
0'
1(
0/
10
#999450000000
1!
b1101101 &
1'
b1101101 )
1-
b0010 .
1/
11
12
13
b1101101 4
b0010 5
#999460000000
0!
1$
0'
1+
0/
#999470000000
1!
1'
1/
#999480000000
0!
0'
0/
#999490000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#999500000000
0!
0'
0/
#999510000000
1!
1'
1/
#999520000000
0!
0'
0/
#999530000000
1!
1"
b1111001 &
1'
1(
b1111001 )
1-
b0011 .
1/
10
11
12
13
b1111001 4
b0011 5
#999540000000
0!
0'
0/
#999550000000
1!
1'
1/
#999560000000
0!
0'
0/
#999570000000
1!
1'
1/
#999580000000
0!
0'
0/
#999590000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#999600000000
0!
0'
0/
#999610000000
1!
1'
1/
#999620000000
0!
0'
0/
#999630000000
1!
1'
1/
#999640000000
0!
0'
0/
#999650000000
1!
1'
1/
#999660000000
0!
0'
0/
#999670000000
1!
1"
b0110011 &
1'
1(
b0110011 )
1-
b0100 .
1/
10
11
12
13
b0110011 4
b0100 5
#999680000000
0!
0'
0/
#999690000000
1!
1'
1/
#999700000000
0!
0'
0/
#999710000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#999720000000
0!
0'
0/
#999730000000
1!
1'
1/
#999740000000
0!
0'
0/
#999750000000
#999760000000
1!
1'
1/
#999770000000
0!
0'
0/
#999780000000
1!
1'
1/
#999790000000
0!
1"
0'
1(
0/
10
#999800000000
1!
b1011011 &
1'
b1011011 )
1-
b0101 .
1/
11
12
13
b1011011 4
b0101 5
#999810000000
0!
0'
0/
#999820000000
1!
1'
1/
#999830000000
0!
0'
0/
#999840000000
1!
0"
1'
0(
0-
1/
00
01
02
03
#999850000000
0!
0'
0/
#999860000000
1!
1'
1/
#999870000000
0!
1"
0'
1(
0/
10
#999880000000
1!
1%
b1011111 &
1'
b1011111 )
1,
1-
b0110 .
1/
11
12
13
b1011111 4
b0110 5
#999890000000
0!
1$
0'
1+
0/
#999900000000
1!
1'
1/
#999910000000
0!
0'
0/
#999920000000
1!
0"
0$
1'
0(
0+
0-
1/
00
01
02
03
#999930000000
0!
0'
0/
#999940000000
1!
1'
1/
#999950000000
0!
0'
0/
#999960000000
1!
1"
0%
b1111110 &
1'
1(
b1111110 )
0,
1-
b0000 .
1/
10
11
12
13
b1111110 4
b0000 5
#999970000000
0!
0'
0/
#999980000000
1!
1'
1/
#999990000000
0!
0'
0/
#1000000000000
1!
1'
1/
