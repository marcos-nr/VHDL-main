$date
  Sun May 26 15:16:01 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module math_real $end
$upscope $end
$scope module tb_tx_uart $end
$var reg 1 ! clk $end
$var reg 1 " reset $end
$var reg 1 # send $end
$var reg 1 $ tx $end
$var reg 1 % done $end
$var reg 8 & cadena[7:0] $end
$scope module uut $end
$var reg 1 ' clk $end
$var reg 1 ( reset $end
$var reg 1 ) send $end
$var reg 8 * cadena[7:0] $end
$var reg 1 + tx $end
$var reg 1 , done $end
$comment estado is not handled $end
$var reg 8 - ds[7:0] $end
$var reg 1 . done_aux $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
0"
1#
1$
1%
b01110010 &
0'
0(
1)
b01110010 *
1+
1,
bUUUUUUUU -
1.
#10000000
1!
0$
1'
0+
b01110010 -
#20000000
0!
0'
#30000000
1!
1'
#40000000
0!
0'
#50000000
1!
1'
#60000000
0!
0'
#70000000
1!
1'
#80000000
0!
0'
#90000000
1!
1'
#100000000
0!
0'
#110000000
1!
1'
#120000000
0!
0'
#130000000
1!
1'
#140000000
0!
0'
#150000000
1!
1'
#160000000
0!
0'
#170000000
1!
1'
#180000000
0!
0'
#190000000
1!
1'
#200000000
0!
0'
#210000000
1!
1'
#220000000
0!
0'
#230000000
1!
1'
#240000000
0!
0'
#250000000
1!
1'
#260000000
0!
0'
#270000000
1!
1'
#280000000
0!
0'
#290000000
1!
1'
#300000000
0!
0'
#310000000
1!
1'
#320000000
0!
0'
#330000000
1!
1'
#340000000
0!
0'
#350000000
1!
1'
#360000000
0!
0'
#370000000
1!
1'
#380000000
0!
0'
#390000000
1!
1'
#400000000
0!
0'
#410000000
1!
1'
#420000000
0!
0'
#430000000
1!
1'
#440000000
0!
0'
#450000000
1!
1'
#460000000
0!
0'
#470000000
1!
1'
#480000000
0!
0'
#490000000
1!
1'
#500000000
0!
0'
#510000000
1!
1'
#520000000
0!
0'
#530000000
1!
1'
#540000000
0!
0'
#550000000
1!
1'
#560000000
0!
0'
#570000000
1!
1'
#580000000
0!
0'
#590000000
1!
1'
#600000000
0!
0'
#610000000
1!
1'
#620000000
0!
0'
#630000000
1!
1'
#640000000
0!
0'
#650000000
1!
1'
#660000000
0!
0'
#670000000
1!
1'
#680000000
0!
0'
#690000000
1!
1'
#700000000
0!
0'
#710000000
1!
1'
#720000000
0!
0'
#730000000
1!
1'
#740000000
0!
0'
#750000000
1!
1'
#760000000
0!
0'
#770000000
1!
1'
#780000000
0!
0'
#790000000
1!
1'
#800000000
0!
0'
#810000000
1!
1'
#820000000
0!
0'
#830000000
1!
1'
#840000000
0!
0'
#850000000
1!
1'
#860000000
0!
0'
#870000000
1!
1'
#880000000
0!
0'
#890000000
1!
1'
#900000000
0!
0'
#910000000
1!
1'
#920000000
0!
0'
#930000000
1!
1'
#940000000
0!
0'
#950000000
1!
1'
#960000000
0!
0'
#970000000
1!
1'
#980000000
0!
0'
#990000000
1!
1'
#1000000000
0!
0'
#1010000000
1!
1'
#1020000000
0!
0'
#1030000000
1!
1'
#1040000000
0!
0'
#1050000000
1!
1'
#1060000000
0!
0'
#1070000000
1!
1'
#1080000000
0!
0'
#1090000000
1!
1'
#1100000000
0!
0'
#1110000000
1!
1'
#1120000000
0!
0'
#1130000000
1!
1'
#1140000000
0!
0'
#1150000000
1!
1'
#1160000000
0!
0'
#1170000000
1!
1'
#1180000000
0!
0'
#1190000000
1!
1'
#1200000000
0!
0'
#1210000000
1!
1'
#1220000000
0!
0'
#1230000000
1!
1'
#1240000000
0!
0'
#1250000000
1!
1'
#1260000000
0!
0'
#1270000000
1!
1'
#1280000000
0!
0'
#1290000000
1!
1'
#1300000000
0!
0'
#1310000000
1!
1'
#1320000000
0!
0'
#1330000000
1!
1'
#1340000000
0!
0'
#1350000000
1!
1'
#1360000000
0!
0'
#1370000000
1!
1'
#1380000000
0!
0'
#1390000000
1!
1'
#1400000000
0!
0'
#1410000000
1!
1'
#1420000000
0!
0'
#1430000000
1!
1'
#1440000000
0!
0'
#1450000000
1!
1'
#1460000000
0!
0'
#1470000000
1!
1'
#1480000000
0!
0'
#1490000000
1!
1'
#1500000000
0!
0'
#1510000000
1!
1'
#1520000000
0!
0'
#1530000000
1!
1'
#1540000000
0!
0'
#1550000000
1!
1'
#1560000000
0!
0'
#1570000000
1!
1'
#1580000000
0!
0'
#1590000000
1!
1'
#1600000000
0!
0'
#1610000000
1!
1'
#1620000000
0!
0'
#1630000000
1!
1'
#1640000000
0!
0'
#1650000000
1!
1'
#1660000000
0!
0'
#1670000000
1!
1'
#1680000000
0!
0'
#1690000000
1!
1'
#1700000000
0!
0'
#1710000000
1!
1'
#1720000000
0!
0'
#1730000000
1!
1'
#1740000000
0!
0'
#1750000000
1!
1'
#1760000000
0!
0'
#1770000000
1!
1'
#1780000000
0!
0'
#1790000000
1!
1'
#1800000000
0!
0'
#1810000000
1!
1'
#1820000000
0!
0'
#1830000000
1!
1'
#1840000000
0!
0'
#1850000000
1!
1'
#1860000000
0!
0'
#1870000000
1!
1'
#1880000000
0!
0'
#1890000000
1!
1'
#1900000000
0!
0'
#1910000000
1!
1'
#1920000000
0!
0'
#1930000000
1!
1'
#1940000000
0!
0'
#1950000000
1!
1'
#1960000000
0!
0'
#1970000000
1!
1'
#1980000000
0!
0'
#1990000000
1!
1'
#2000000000
0!
0'
#2010000000
1!
1'
#2020000000
0!
0'
#2030000000
1!
1'
#2040000000
0!
0'
#2050000000
1!
1'
#2060000000
0!
0'
#2070000000
1!
1'
#2080000000
0!
0'
#2090000000
1!
1'
#2100000000
0!
0'
#2110000000
1!
1'
#2120000000
0!
0'
#2130000000
1!
1'
#2140000000
0!
0'
#2150000000
1!
1'
#2160000000
0!
0'
#2170000000
1!
1'
#2180000000
0!
0'
#2190000000
1!
1'
#2200000000
0!
0'
#2210000000
1!
1'
#2220000000
0!
0'
#2230000000
1!
1'
#2240000000
0!
0'
#2250000000
1!
1'
#2260000000
0!
0'
#2270000000
1!
1'
#2280000000
0!
0'
#2290000000
1!
1'
#2300000000
0!
0'
#2310000000
1!
1'
#2320000000
0!
0'
#2330000000
1!
1'
#2340000000
0!
0'
#2350000000
1!
1'
#2360000000
0!
0'
#2370000000
1!
1'
#2380000000
0!
0'
#2390000000
1!
1'
#2400000000
0!
0'
#2410000000
1!
1'
#2420000000
0!
0'
#2430000000
1!
1'
#2440000000
0!
0'
#2450000000
1!
1'
#2460000000
0!
0'
#2470000000
1!
1'
#2480000000
0!
0'
#2490000000
1!
1'
#2500000000
0!
0'
#2510000000
1!
1'
#2520000000
0!
0'
#2530000000
1!
1'
#2540000000
0!
0'
#2550000000
1!
1'
#2560000000
0!
0'
#2570000000
1!
1'
#2580000000
0!
0'
#2590000000
1!
1'
#2600000000
0!
0'
#2610000000
1!
1'
#2620000000
0!
0'
#2630000000
1!
1'
#2640000000
0!
0'
#2650000000
1!
1'
#2660000000
0!
0'
#2670000000
1!
1'
#2680000000
0!
0'
#2690000000
1!
1'
#2700000000
0!
0'
#2710000000
1!
1'
#2720000000
0!
0'
#2730000000
1!
1'
#2740000000
0!
0'
#2750000000
1!
1'
#2760000000
0!
0'
#2770000000
1!
1'
#2780000000
0!
0'
#2790000000
1!
1'
#2800000000
0!
0'
#2810000000
1!
1'
#2820000000
0!
0'
#2830000000
1!
1'
#2840000000
0!
0'
#2850000000
1!
1'
#2860000000
0!
0'
#2870000000
1!
1'
#2880000000
0!
0'
#2890000000
1!
1'
#2900000000
0!
0'
#2910000000
1!
1'
#2920000000
0!
0'
#2930000000
1!
1'
#2940000000
0!
0'
#2950000000
1!
1'
#2960000000
0!
0'
#2970000000
1!
1'
#2980000000
0!
0'
#2990000000
1!
1'
#3000000000
0!
0'
#3010000000
1!
1'
#3020000000
0!
0'
#3030000000
1!
1'
#3040000000
0!
0'
#3050000000
1!
1'
#3060000000
0!
0'
#3070000000
1!
1'
#3080000000
0!
0'
#3090000000
1!
1'
#3100000000
0!
0'
#3110000000
1!
1'
#3120000000
0!
0'
#3130000000
1!
1'
#3140000000
0!
0'
#3150000000
1!
1'
#3160000000
0!
0'
#3170000000
1!
1'
#3180000000
0!
0'
#3190000000
1!
1'
#3200000000
0!
0'
#3210000000
1!
1'
#3220000000
0!
0'
#3230000000
1!
1'
#3240000000
0!
0'
#3250000000
1!
1'
#3260000000
0!
0'
#3270000000
1!
1'
#3280000000
0!
0'
#3290000000
1!
1'
#3300000000
0!
0'
#3310000000
1!
1'
#3320000000
0!
0'
#3330000000
1!
1'
#3340000000
0!
0'
#3350000000
1!
1'
#3360000000
0!
0'
#3370000000
1!
1'
#3380000000
0!
0'
#3390000000
1!
1'
#3400000000
0!
0'
#3410000000
1!
1'
#3420000000
0!
0'
#3430000000
1!
1'
#3440000000
0!
0'
#3450000000
1!
1'
#3460000000
0!
0'
#3470000000
1!
1'
#3480000000
0!
0'
#3490000000
1!
1'
#3500000000
0!
0'
#3510000000
1!
1'
#3520000000
0!
0'
#3530000000
1!
1'
#3540000000
0!
0'
#3550000000
1!
1'
#3560000000
0!
0'
#3570000000
1!
1'
#3580000000
0!
0'
#3590000000
1!
1'
#3600000000
0!
0'
#3610000000
1!
1'
#3620000000
0!
0'
#3630000000
1!
1'
#3640000000
0!
0'
#3650000000
1!
1'
#3660000000
0!
0'
#3670000000
1!
1'
#3680000000
0!
0'
#3690000000
1!
1'
#3700000000
0!
0'
#3710000000
1!
1'
#3720000000
0!
0'
#3730000000
1!
1'
#3740000000
0!
0'
#3750000000
1!
1'
#3760000000
0!
0'
#3770000000
1!
1'
#3780000000
0!
0'
#3790000000
1!
1'
#3800000000
0!
0'
#3810000000
1!
1'
#3820000000
0!
0'
#3830000000
1!
1'
#3840000000
0!
0'
#3850000000
1!
1'
#3860000000
0!
0'
#3870000000
1!
1'
#3880000000
0!
0'
#3890000000
1!
1'
#3900000000
0!
0'
#3910000000
1!
1'
#3920000000
0!
0'
#3930000000
1!
1'
#3940000000
0!
0'
#3950000000
1!
1'
#3960000000
0!
0'
#3970000000
1!
1'
#3980000000
0!
0'
#3990000000
1!
1'
#4000000000
0!
0'
#4010000000
1!
1'
#4020000000
0!
0'
#4030000000
1!
1'
#4040000000
0!
0'
#4050000000
1!
1'
#4060000000
0!
0'
#4070000000
1!
1'
#4080000000
0!
0'
#4090000000
1!
1'
#4100000000
0!
0'
#4110000000
1!
1'
#4120000000
0!
0'
#4130000000
1!
1'
#4140000000
0!
0'
#4150000000
1!
1'
#4160000000
0!
0'
#4170000000
1!
1'
#4180000000
0!
0'
#4190000000
1!
1'
#4200000000
0!
0'
#4210000000
1!
1'
#4220000000
0!
0'
#4230000000
1!
1'
#4240000000
0!
0'
#4250000000
1!
1'
#4260000000
0!
0'
#4270000000
1!
1'
#4280000000
0!
0'
#4290000000
1!
1'
#4300000000
0!
0'
#4310000000
1!
1'
#4320000000
0!
0'
#4330000000
1!
1'
#4340000000
0!
0'
#4350000000
1!
1'
#4360000000
0!
0'
#4370000000
1!
1'
#4380000000
0!
0'
#4390000000
1!
1'
#4400000000
0!
0'
#4410000000
1!
1'
#4420000000
0!
0'
#4430000000
1!
1'
#4440000000
0!
0'
#4450000000
1!
1'
#4460000000
0!
0'
#4470000000
1!
1'
#4480000000
0!
0'
#4490000000
1!
1'
#4500000000
0!
0'
#4510000000
1!
1'
#4520000000
0!
0'
#4530000000
1!
1'
#4540000000
0!
0'
#4550000000
1!
1'
#4560000000
0!
0'
#4570000000
1!
1'
#4580000000
0!
0'
#4590000000
1!
1'
#4600000000
0!
0'
#4610000000
1!
1'
#4620000000
0!
0'
#4630000000
1!
1'
#4640000000
0!
0'
#4650000000
1!
1'
#4660000000
0!
0'
#4670000000
1!
1'
#4680000000
0!
0'
#4690000000
1!
1'
#4700000000
0!
0'
#4710000000
1!
1'
#4720000000
0!
0'
#4730000000
1!
1'
#4740000000
0!
0'
#4750000000
1!
1'
#4760000000
0!
0'
#4770000000
1!
1'
#4780000000
0!
0'
#4790000000
1!
1'
#4800000000
0!
0'
#4810000000
1!
1'
#4820000000
0!
0'
#4830000000
1!
1'
#4840000000
0!
0'
#4850000000
1!
1'
#4860000000
0!
0'
#4870000000
1!
1'
#4880000000
0!
0'
#4890000000
1!
1'
#4900000000
0!
0'
#4910000000
1!
1'
#4920000000
0!
0'
#4930000000
1!
1'
#4940000000
0!
0'
#4950000000
1!
1'
#4960000000
0!
0'
#4970000000
1!
1'
#4980000000
0!
0'
#4990000000
1!
1'
#5000000000
0!
0'
#5010000000
1!
1'
#5020000000
0!
0'
#5030000000
1!
1'
#5040000000
0!
0'
#5050000000
1!
1'
#5060000000
0!
0'
#5070000000
1!
1'
#5080000000
0!
0'
#5090000000
1!
1'
#5100000000
0!
0'
#5110000000
1!
1'
#5120000000
0!
0'
#5130000000
1!
1'
#5140000000
0!
0'
#5150000000
1!
1'
#5160000000
0!
0'
#5170000000
1!
1'
#5180000000
0!
0'
#5190000000
1!
1'
#5200000000
0!
0'
#5210000000
1!
1'
#5220000000
0!
0'
#5230000000
1!
1'
#5240000000
0!
0'
#5250000000
1!
1'
#5260000000
0!
0'
#5270000000
1!
1'
#5280000000
0!
0'
#5290000000
1!
1'
#5300000000
0!
0'
#5310000000
1!
1'
#5320000000
0!
0'
#5330000000
1!
1'
#5340000000
0!
0'
#5350000000
1!
1'
#5360000000
0!
0'
#5370000000
1!
1'
#5380000000
0!
0'
#5390000000
1!
1'
#5400000000
0!
0'
#5410000000
1!
1'
#5420000000
0!
0'
#5430000000
1!
1'
#5440000000
0!
0'
#5450000000
1!
1'
#5460000000
0!
0'
#5470000000
1!
1'
#5480000000
0!
0'
#5490000000
1!
1'
#5500000000
0!
0'
#5510000000
1!
1'
#5520000000
0!
0'
#5530000000
1!
1'
#5540000000
0!
0'
#5550000000
1!
1'
#5560000000
0!
0'
#5570000000
1!
1'
#5580000000
0!
0'
#5590000000
1!
1'
#5600000000
0!
0'
#5610000000
1!
1'
#5620000000
0!
0'
#5630000000
1!
1'
#5640000000
0!
0'
#5650000000
1!
1'
#5660000000
0!
0'
#5670000000
1!
1'
#5680000000
0!
0'
#5690000000
1!
1'
#5700000000
0!
0'
#5710000000
1!
1'
#5720000000
0!
0'
#5730000000
1!
1'
#5740000000
0!
0'
#5750000000
1!
1'
#5760000000
0!
0'
#5770000000
1!
1'
#5780000000
0!
0'
#5790000000
1!
1'
#5800000000
0!
0'
#5810000000
1!
1'
#5820000000
0!
0'
#5830000000
1!
1'
#5840000000
0!
0'
#5850000000
1!
1'
#5860000000
0!
0'
#5870000000
1!
1'
#5880000000
0!
0'
#5890000000
1!
1'
#5900000000
0!
0'
#5910000000
1!
1'
#5920000000
0!
0'
#5930000000
1!
1'
#5940000000
0!
0'
#5950000000
1!
1'
#5960000000
0!
0'
#5970000000
1!
1'
#5980000000
0!
0'
#5990000000
1!
1'
#6000000000
0!
0'
#6010000000
1!
1'
#6020000000
0!
0'
#6030000000
1!
1'
#6040000000
0!
0'
#6050000000
1!
1'
#6060000000
0!
0'
#6070000000
1!
1'
#6080000000
0!
0'
#6090000000
1!
1'
#6100000000
0!
0'
#6110000000
1!
1'
#6120000000
0!
0'
#6130000000
1!
1'
#6140000000
0!
0'
#6150000000
1!
1'
#6160000000
0!
0'
#6170000000
1!
1'
#6180000000
0!
0'
#6190000000
1!
1'
#6200000000
0!
0'
#6210000000
1!
1'
#6220000000
0!
0'
#6230000000
1!
1'
#6240000000
0!
0'
#6250000000
1!
1'
#6260000000
0!
0'
#6270000000
1!
1'
#6280000000
0!
0'
#6290000000
1!
1'
#6300000000
0!
0'
#6310000000
1!
1'
#6320000000
0!
0'
#6330000000
1!
1'
#6340000000
0!
0'
#6350000000
1!
1'
#6360000000
0!
0'
#6370000000
1!
1'
#6380000000
0!
0'
#6390000000
1!
1'
#6400000000
0!
0'
#6410000000
1!
1'
#6420000000
0!
0'
#6430000000
1!
1'
#6440000000
0!
0'
#6450000000
1!
1'
#6460000000
0!
0'
#6470000000
1!
1'
#6480000000
0!
0'
#6490000000
1!
1'
#6500000000
0!
0'
#6510000000
1!
1'
#6520000000
0!
0'
#6530000000
1!
1'
#6540000000
0!
0'
#6550000000
1!
1'
#6560000000
0!
0'
#6570000000
1!
1'
#6580000000
0!
0'
#6590000000
1!
1'
#6600000000
0!
0'
#6610000000
1!
1'
#6620000000
0!
0'
#6630000000
1!
1'
#6640000000
0!
0'
#6650000000
1!
1'
#6660000000
0!
0'
#6670000000
1!
1'
#6680000000
0!
0'
#6690000000
1!
1'
#6700000000
0!
0'
#6710000000
1!
1'
#6720000000
0!
0'
#6730000000
1!
1'
#6740000000
0!
0'
#6750000000
1!
1'
#6760000000
0!
0'
#6770000000
1!
1'
#6780000000
0!
0'
#6790000000
1!
1'
#6800000000
0!
0'
#6810000000
1!
1'
#6820000000
0!
0'
#6830000000
1!
1'
#6840000000
0!
0'
#6850000000
1!
1'
#6860000000
0!
0'
#6870000000
1!
1'
#6880000000
0!
0'
#6890000000
1!
1'
#6900000000
0!
0'
#6910000000
1!
1'
#6920000000
0!
0'
#6930000000
1!
1'
#6940000000
0!
0'
#6950000000
1!
1'
#6960000000
0!
0'
#6970000000
1!
1'
#6980000000
0!
0'
#6990000000
1!
1'
#7000000000
0!
0'
#7010000000
1!
1'
#7020000000
0!
0'
#7030000000
1!
1'
#7040000000
0!
0'
#7050000000
1!
1'
#7060000000
0!
0'
#7070000000
1!
1'
#7080000000
0!
0'
#7090000000
1!
1'
#7100000000
0!
0'
#7110000000
1!
1'
#7120000000
0!
0'
#7130000000
1!
1'
#7140000000
0!
0'
#7150000000
1!
1'
#7160000000
0!
0'
#7170000000
1!
1'
#7180000000
0!
0'
#7190000000
1!
1'
#7200000000
0!
0'
#7210000000
1!
1'
#7220000000
0!
0'
#7230000000
1!
1'
#7240000000
0!
0'
#7250000000
1!
1'
#7260000000
0!
0'
#7270000000
1!
1'
#7280000000
0!
0'
#7290000000
1!
1'
#7300000000
0!
0'
#7310000000
1!
1'
#7320000000
0!
0'
#7330000000
1!
1'
#7340000000
0!
0'
#7350000000
1!
1'
#7360000000
0!
0'
#7370000000
1!
1'
#7380000000
0!
0'
#7390000000
1!
1'
#7400000000
0!
0'
#7410000000
1!
1'
#7420000000
0!
0'
#7430000000
1!
1'
#7440000000
0!
0'
#7450000000
1!
1'
#7460000000
0!
0'
#7470000000
1!
1'
#7480000000
0!
0'
#7490000000
1!
1'
#7500000000
0!
0'
#7510000000
1!
1'
#7520000000
0!
0'
#7530000000
1!
1'
#7540000000
0!
0'
#7550000000
1!
1'
#7560000000
0!
0'
#7570000000
1!
1'
#7580000000
0!
0'
#7590000000
1!
1'
#7600000000
0!
0'
#7610000000
1!
1'
#7620000000
0!
0'
#7630000000
1!
1'
#7640000000
0!
0'
#7650000000
1!
1'
#7660000000
0!
0'
#7670000000
1!
1'
#7680000000
0!
0'
#7690000000
1!
1'
#7700000000
0!
0'
#7710000000
1!
1'
#7720000000
0!
0'
#7730000000
1!
1'
#7740000000
0!
0'
#7750000000
1!
1'
#7760000000
0!
0'
#7770000000
1!
1'
#7780000000
0!
0'
#7790000000
1!
1'
#7800000000
0!
0'
#7810000000
1!
1'
#7820000000
0!
0'
#7830000000
1!
1'
#7840000000
0!
0'
#7850000000
1!
1'
#7860000000
0!
0'
#7870000000
1!
1'
#7880000000
0!
0'
#7890000000
1!
1'
#7900000000
0!
0'
#7910000000
1!
1'
#7920000000
0!
0'
#7930000000
1!
1'
#7940000000
0!
0'
#7950000000
1!
1'
#7960000000
0!
0'
#7970000000
1!
1'
#7980000000
0!
0'
#7990000000
1!
1'
#8000000000
0!
0'
#8010000000
1!
1'
#8020000000
0!
0'
#8030000000
1!
1'
#8040000000
0!
0'
#8050000000
1!
1'
#8060000000
0!
0'
#8070000000
1!
1'
#8080000000
0!
0'
#8090000000
1!
1'
#8100000000
0!
0'
#8110000000
1!
1'
#8120000000
0!
0'
#8130000000
1!
1'
#8140000000
0!
0'
#8150000000
1!
1'
#8160000000
0!
0'
#8170000000
1!
1'
#8180000000
0!
0'
#8190000000
1!
1'
#8200000000
0!
0'
#8210000000
1!
1'
#8220000000
0!
0'
#8230000000
1!
1'
#8240000000
0!
0'
#8250000000
1!
1'
#8260000000
0!
0'
#8270000000
1!
1'
#8280000000
0!
0'
#8290000000
1!
1'
#8300000000
0!
0'
#8310000000
1!
1'
#8320000000
0!
0'
#8330000000
1!
1'
#8340000000
0!
0'
#8350000000
1!
1'
#8360000000
0!
0'
#8370000000
1!
1'
#8380000000
0!
0'
#8390000000
1!
1'
#8400000000
0!
0'
#8410000000
1!
1'
#8420000000
0!
0'
#8430000000
1!
1'
#8440000000
0!
0'
#8450000000
1!
1'
#8460000000
0!
0'
#8470000000
1!
1'
#8480000000
0!
0'
#8490000000
1!
1'
#8500000000
0!
0'
#8510000000
1!
1'
#8520000000
0!
0'
#8530000000
1!
1'
#8540000000
0!
0'
#8550000000
1!
1'
#8560000000
0!
0'
#8570000000
1!
1'
#8580000000
0!
0'
#8590000000
1!
1'
#8600000000
0!
0'
#8610000000
1!
1'
#8620000000
0!
0'
#8630000000
1!
1'
#8640000000
0!
0'
#8650000000
1!
1'
#8660000000
0!
0'
#8670000000
1!
1'
#8680000000
0!
0'
#8690000000
1!
1'
#8700000000
0!
0'
#8710000000
1!
1'
#8720000000
0!
0'
#8730000000
1!
1'
#8740000000
0!
0'
#8750000000
1!
1'
#8760000000
0!
0'
#8770000000
1!
1'
#8780000000
0!
0'
#8790000000
1!
1'
#8800000000
0!
0'
#8810000000
1!
1'
#8820000000
0!
0'
#8830000000
1!
1'
#8840000000
0!
0'
#8850000000
1!
1'
#8860000000
0!
0'
#8870000000
1!
1'
#8880000000
0!
0'
#8890000000
1!
1'
#8900000000
0!
0'
#8910000000
1!
1'
#8920000000
0!
0'
#8930000000
1!
1'
#8940000000
0!
0'
#8950000000
1!
1'
#8960000000
0!
0'
#8970000000
1!
1'
#8980000000
0!
0'
#8990000000
1!
1'
#9000000000
0!
0'
#9010000000
1!
1'
#9020000000
0!
0'
#9030000000
1!
1'
#9040000000
0!
0'
#9050000000
1!
1'
#9060000000
0!
0'
#9070000000
1!
1'
#9080000000
0!
0'
#9090000000
1!
1'
#9100000000
0!
0'
#9110000000
1!
1'
#9120000000
0!
0'
#9130000000
1!
1'
#9140000000
0!
0'
#9150000000
1!
1'
#9160000000
0!
0'
#9170000000
1!
1'
#9180000000
0!
0'
#9190000000
1!
1'
#9200000000
0!
0'
#9210000000
1!
1'
#9220000000
0!
0'
#9230000000
1!
1'
#9240000000
0!
0'
#9250000000
1!
1'
#9260000000
0!
0'
#9270000000
1!
1'
#9280000000
0!
0'
#9290000000
1!
1'
#9300000000
0!
0'
#9310000000
1!
1'
#9320000000
0!
0'
#9330000000
1!
1'
#9340000000
0!
0'
#9350000000
1!
1'
#9360000000
0!
0'
#9370000000
1!
1'
#9380000000
0!
0'
#9390000000
1!
1'
#9400000000
0!
0'
#9410000000
1!
1'
#9420000000
0!
0'
#9430000000
1!
1'
#9440000000
0!
0'
#9450000000
1!
1'
#9460000000
0!
0'
#9470000000
1!
1'
#9480000000
0!
0'
#9490000000
1!
1'
#9500000000
0!
0'
#9510000000
1!
1'
#9520000000
0!
0'
#9530000000
1!
1'
#9540000000
0!
0'
#9550000000
1!
1'
#9560000000
0!
0'
#9570000000
1!
1'
#9580000000
0!
0'
#9590000000
1!
1'
#9600000000
0!
0'
#9610000000
1!
1'
#9620000000
0!
0'
#9630000000
1!
1'
#9640000000
0!
0'
#9650000000
1!
1'
#9660000000
0!
0'
#9670000000
1!
1'
#9680000000
0!
0'
#9690000000
1!
1'
#9700000000
0!
0'
#9710000000
1!
1'
#9720000000
0!
0'
#9730000000
1!
1'
#9740000000
0!
0'
#9750000000
1!
1'
#9760000000
0!
0'
#9770000000
1!
1'
#9780000000
0!
0'
#9790000000
1!
1'
#9800000000
0!
0'
#9810000000
1!
1'
#9820000000
0!
0'
#9830000000
1!
1'
#9840000000
0!
0'
#9850000000
1!
1'
#9860000000
0!
0'
#9870000000
1!
1'
#9880000000
0!
0'
#9890000000
1!
1'
#9900000000
0!
0'
#9910000000
1!
1'
#9920000000
0!
0'
#9930000000
1!
1'
#9940000000
0!
0'
#9950000000
1!
1'
#9960000000
0!
0'
#9970000000
1!
1'
#9980000000
0!
0'
#9990000000
1!
1'
#10000000000
0!
0'
