$date
  Mon Apr 15 19:21:22 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_tp1_3 $end
$var reg 4 ! vot[3:0] $end
$var reg 7 " disp[6:0] $end
$scope module uut $end
$var reg 4 # votos[3:0] $end
$var reg 7 $ display[6:0] $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
b0000 !
b1011110 "
b0000 #
b1011110 $
#10000000
b0001 !
b0001 #
#20000000
b0010 !
b0010 #
#30000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#40000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#50000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#60000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#70000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#80000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#90000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#100000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#110000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#120000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#130000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#140000000
b1110 !
b1110 #
#150000000
b1111 !
b1111 #
#160000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#170000000
b0001 !
b0001 #
#180000000
b0010 !
b0010 #
#190000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#200000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#210000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#220000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#230000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#240000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#250000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#260000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#270000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#280000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#290000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#300000000
b1110 !
b1110 #
#310000000
b1111 !
b1111 #
#320000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#330000000
b0001 !
b0001 #
#340000000
b0010 !
b0010 #
#350000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#360000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#370000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#380000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#390000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#400000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#410000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#420000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#430000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#440000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#450000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#460000000
b1110 !
b1110 #
#470000000
b1111 !
b1111 #
#480000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#490000000
b0001 !
b0001 #
#500000000
b0010 !
b0010 #
#510000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#520000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#530000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#540000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#550000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#560000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#570000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#580000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#590000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#600000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#610000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#620000000
b1110 !
b1110 #
#630000000
b1111 !
b1111 #
#640000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#650000000
b0001 !
b0001 #
#660000000
b0010 !
b0010 #
#670000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#680000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#690000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#700000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#710000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#720000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#730000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#740000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#750000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#760000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#770000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#780000000
b1110 !
b1110 #
#790000000
b1111 !
b1111 #
#800000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#810000000
b0001 !
b0001 #
#820000000
b0010 !
b0010 #
#830000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#840000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#850000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#860000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#870000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#880000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#890000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#900000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#910000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#920000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#930000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#940000000
b1110 !
b1110 #
#950000000
b1111 !
b1111 #
#960000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#970000000
b0001 !
b0001 #
#980000000
b0010 !
b0010 #
#990000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#1000000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#1010000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#1020000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#1030000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#1040000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#1050000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#1060000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#1070000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#1080000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#1090000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#1100000000
b1110 !
b1110 #
#1110000000
b1111 !
b1111 #
#1120000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#1130000000
b0001 !
b0001 #
#1140000000
b0010 !
b0010 #
#1150000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#1160000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#1170000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#1180000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#1190000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#1200000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#1210000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#1220000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#1230000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#1240000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#1250000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#1260000000
b1110 !
b1110 #
#1270000000
b1111 !
b1111 #
#1280000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#1290000000
b0001 !
b0001 #
#1300000000
b0010 !
b0010 #
#1310000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#1320000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#1330000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#1340000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#1350000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#1360000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#1370000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#1380000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#1390000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#1400000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#1410000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#1420000000
b1110 !
b1110 #
#1430000000
b1111 !
b1111 #
#1440000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#1450000000
b0001 !
b0001 #
#1460000000
b0010 !
b0010 #
#1470000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#1480000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#1490000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#1500000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#1510000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#1520000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#1530000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#1540000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#1550000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#1560000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#1570000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#1580000000
b1110 !
b1110 #
#1590000000
b1111 !
b1111 #
#1600000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#1610000000
b0001 !
b0001 #
#1620000000
b0010 !
b0010 #
#1630000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#1640000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#1650000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#1660000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#1670000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#1680000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#1690000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#1700000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#1710000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#1720000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#1730000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#1740000000
b1110 !
b1110 #
#1750000000
b1111 !
b1111 #
#1760000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#1770000000
b0001 !
b0001 #
#1780000000
b0010 !
b0010 #
#1790000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#1800000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#1810000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#1820000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#1830000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#1840000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#1850000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#1860000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#1870000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#1880000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#1890000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#1900000000
b1110 !
b1110 #
#1910000000
b1111 !
b1111 #
#1920000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#1930000000
b0001 !
b0001 #
#1940000000
b0010 !
b0010 #
#1950000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#1960000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#1970000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#1980000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#1990000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#2000000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#2010000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#2020000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#2030000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#2040000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#2050000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#2060000000
b1110 !
b1110 #
#2070000000
b1111 !
b1111 #
#2080000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#2090000000
b0001 !
b0001 #
#2100000000
b0010 !
b0010 #
#2110000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#2120000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#2130000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#2140000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#2150000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#2160000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#2170000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#2180000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#2190000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#2200000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#2210000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#2220000000
b1110 !
b1110 #
#2230000000
b1111 !
b1111 #
#2240000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#2250000000
b0001 !
b0001 #
#2260000000
b0010 !
b0010 #
#2270000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#2280000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#2290000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#2300000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#2310000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#2320000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#2330000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#2340000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#2350000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#2360000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#2370000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#2380000000
b1110 !
b1110 #
#2390000000
b1111 !
b1111 #
#2400000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#2410000000
b0001 !
b0001 #
#2420000000
b0010 !
b0010 #
#2430000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#2440000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#2450000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#2460000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#2470000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#2480000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#2490000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#2500000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#2510000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#2520000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#2530000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#2540000000
b1110 !
b1110 #
#2550000000
b1111 !
b1111 #
#2560000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#2570000000
b0001 !
b0001 #
#2580000000
b0010 !
b0010 #
#2590000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#2600000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#2610000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#2620000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#2630000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#2640000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#2650000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#2660000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#2670000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#2680000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#2690000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#2700000000
b1110 !
b1110 #
#2710000000
b1111 !
b1111 #
#2720000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#2730000000
b0001 !
b0001 #
#2740000000
b0010 !
b0010 #
#2750000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#2760000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#2770000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#2780000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#2790000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#2800000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#2810000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#2820000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#2830000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#2840000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#2850000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#2860000000
b1110 !
b1110 #
#2870000000
b1111 !
b1111 #
#2880000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#2890000000
b0001 !
b0001 #
#2900000000
b0010 !
b0010 #
#2910000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#2920000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#2930000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#2940000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#2950000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#2960000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#2970000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#2980000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#2990000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#3000000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#3010000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#3020000000
b1110 !
b1110 #
#3030000000
b1111 !
b1111 #
#3040000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#3050000000
b0001 !
b0001 #
#3060000000
b0010 !
b0010 #
#3070000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#3080000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#3090000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#3100000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#3110000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#3120000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#3130000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#3140000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#3150000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#3160000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#3170000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#3180000000
b1110 !
b1110 #
#3190000000
b1111 !
b1111 #
#3200000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#3210000000
b0001 !
b0001 #
#3220000000
b0010 !
b0010 #
#3230000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#3240000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#3250000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#3260000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#3270000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#3280000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#3290000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#3300000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#3310000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#3320000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#3330000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#3340000000
b1110 !
b1110 #
#3350000000
b1111 !
b1111 #
#3360000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#3370000000
b0001 !
b0001 #
#3380000000
b0010 !
b0010 #
#3390000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#3400000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#3410000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#3420000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#3430000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#3440000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#3450000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#3460000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#3470000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#3480000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#3490000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#3500000000
b1110 !
b1110 #
#3510000000
b1111 !
b1111 #
#3520000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#3530000000
b0001 !
b0001 #
#3540000000
b0010 !
b0010 #
#3550000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#3560000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#3570000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#3580000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#3590000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#3600000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#3610000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#3620000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#3630000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#3640000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#3650000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#3660000000
b1110 !
b1110 #
#3670000000
b1111 !
b1111 #
#3680000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#3690000000
b0001 !
b0001 #
#3700000000
b0010 !
b0010 #
#3710000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#3720000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#3730000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#3740000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#3750000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#3760000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#3770000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#3780000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#3790000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#3800000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#3810000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#3820000000
b1110 !
b1110 #
#3830000000
b1111 !
b1111 #
#3840000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#3850000000
b0001 !
b0001 #
#3860000000
b0010 !
b0010 #
#3870000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#3880000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#3890000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#3900000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#3910000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#3920000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#3930000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#3940000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#3950000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#3960000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#3970000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#3980000000
b1110 !
b1110 #
#3990000000
b1111 !
b1111 #
#4000000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#4010000000
b0001 !
b0001 #
#4020000000
b0010 !
b0010 #
#4030000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#4040000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#4050000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#4060000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#4070000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#4080000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#4090000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#4100000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#4110000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#4120000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#4130000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#4140000000
b1110 !
b1110 #
#4150000000
b1111 !
b1111 #
#4160000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#4170000000
b0001 !
b0001 #
#4180000000
b0010 !
b0010 #
#4190000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#4200000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#4210000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#4220000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#4230000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#4240000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#4250000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#4260000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#4270000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#4280000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#4290000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#4300000000
b1110 !
b1110 #
#4310000000
b1111 !
b1111 #
#4320000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#4330000000
b0001 !
b0001 #
#4340000000
b0010 !
b0010 #
#4350000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#4360000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#4370000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#4380000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#4390000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#4400000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#4410000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#4420000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#4430000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#4440000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#4450000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#4460000000
b1110 !
b1110 #
#4470000000
b1111 !
b1111 #
#4480000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#4490000000
b0001 !
b0001 #
#4500000000
b0010 !
b0010 #
#4510000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#4520000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#4530000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#4540000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#4550000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#4560000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#4570000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#4580000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#4590000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#4600000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#4610000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#4620000000
b1110 !
b1110 #
#4630000000
b1111 !
b1111 #
#4640000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#4650000000
b0001 !
b0001 #
#4660000000
b0010 !
b0010 #
#4670000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#4680000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#4690000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#4700000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#4710000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#4720000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#4730000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#4740000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#4750000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#4760000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#4770000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#4780000000
b1110 !
b1110 #
#4790000000
b1111 !
b1111 #
#4800000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#4810000000
b0001 !
b0001 #
#4820000000
b0010 !
b0010 #
#4830000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#4840000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#4850000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#4860000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#4870000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#4880000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#4890000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#4900000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#4910000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#4920000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#4930000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#4940000000
b1110 !
b1110 #
#4950000000
b1111 !
b1111 #
#4960000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#4970000000
b0001 !
b0001 #
#4980000000
b0010 !
b0010 #
#4990000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#5000000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#5010000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#5020000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#5030000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#5040000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#5050000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#5060000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#5070000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#5080000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#5090000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#5100000000
b1110 !
b1110 #
#5110000000
b1111 !
b1111 #
#5120000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#5130000000
b0001 !
b0001 #
#5140000000
b0010 !
b0010 #
#5150000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#5160000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#5170000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#5180000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#5190000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#5200000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#5210000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#5220000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#5230000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#5240000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#5250000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#5260000000
b1110 !
b1110 #
#5270000000
b1111 !
b1111 #
#5280000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#5290000000
b0001 !
b0001 #
#5300000000
b0010 !
b0010 #
#5310000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#5320000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#5330000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#5340000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#5350000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#5360000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#5370000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#5380000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#5390000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#5400000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#5410000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#5420000000
b1110 !
b1110 #
#5430000000
b1111 !
b1111 #
#5440000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#5450000000
b0001 !
b0001 #
#5460000000
b0010 !
b0010 #
#5470000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#5480000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#5490000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#5500000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#5510000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#5520000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#5530000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#5540000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#5550000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#5560000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#5570000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#5580000000
b1110 !
b1110 #
#5590000000
b1111 !
b1111 #
#5600000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#5610000000
b0001 !
b0001 #
#5620000000
b0010 !
b0010 #
#5630000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#5640000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#5650000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#5660000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#5670000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#5680000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#5690000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#5700000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#5710000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#5720000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#5730000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#5740000000
b1110 !
b1110 #
#5750000000
b1111 !
b1111 #
#5760000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#5770000000
b0001 !
b0001 #
#5780000000
b0010 !
b0010 #
#5790000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#5800000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#5810000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#5820000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#5830000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#5840000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#5850000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#5860000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#5870000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#5880000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#5890000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#5900000000
b1110 !
b1110 #
#5910000000
b1111 !
b1111 #
#5920000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#5930000000
b0001 !
b0001 #
#5940000000
b0010 !
b0010 #
#5950000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#5960000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#5970000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#5980000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#5990000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#6000000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#6010000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#6020000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#6030000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#6040000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#6050000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#6060000000
b1110 !
b1110 #
#6070000000
b1111 !
b1111 #
#6080000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#6090000000
b0001 !
b0001 #
#6100000000
b0010 !
b0010 #
#6110000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#6120000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#6130000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#6140000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#6150000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#6160000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#6170000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#6180000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#6190000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#6200000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#6210000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#6220000000
b1110 !
b1110 #
#6230000000
b1111 !
b1111 #
#6240000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#6250000000
b0001 !
b0001 #
#6260000000
b0010 !
b0010 #
#6270000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#6280000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#6290000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#6300000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#6310000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#6320000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#6330000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#6340000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#6350000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#6360000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#6370000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#6380000000
b1110 !
b1110 #
#6390000000
b1111 !
b1111 #
#6400000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#6410000000
b0001 !
b0001 #
#6420000000
b0010 !
b0010 #
#6430000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#6440000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#6450000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#6460000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#6470000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#6480000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#6490000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#6500000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#6510000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#6520000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#6530000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#6540000000
b1110 !
b1110 #
#6550000000
b1111 !
b1111 #
#6560000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#6570000000
b0001 !
b0001 #
#6580000000
b0010 !
b0010 #
#6590000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#6600000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#6610000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#6620000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#6630000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#6640000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#6650000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#6660000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#6670000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#6680000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#6690000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#6700000000
b1110 !
b1110 #
#6710000000
b1111 !
b1111 #
#6720000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#6730000000
b0001 !
b0001 #
#6740000000
b0010 !
b0010 #
#6750000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#6760000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#6770000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#6780000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#6790000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#6800000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#6810000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#6820000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#6830000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#6840000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#6850000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#6860000000
b1110 !
b1110 #
#6870000000
b1111 !
b1111 #
#6880000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#6890000000
b0001 !
b0001 #
#6900000000
b0010 !
b0010 #
#6910000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#6920000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#6930000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#6940000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#6950000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#6960000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#6970000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#6980000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#6990000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#7000000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#7010000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#7020000000
b1110 !
b1110 #
#7030000000
b1111 !
b1111 #
#7040000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#7050000000
b0001 !
b0001 #
#7060000000
b0010 !
b0010 #
#7070000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#7080000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#7090000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#7100000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#7110000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#7120000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#7130000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#7140000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#7150000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#7160000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#7170000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#7180000000
b1110 !
b1110 #
#7190000000
b1111 !
b1111 #
#7200000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#7210000000
b0001 !
b0001 #
#7220000000
b0010 !
b0010 #
#7230000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#7240000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#7250000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#7260000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#7270000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#7280000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#7290000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#7300000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#7310000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#7320000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#7330000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#7340000000
b1110 !
b1110 #
#7350000000
b1111 !
b1111 #
#7360000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#7370000000
b0001 !
b0001 #
#7380000000
b0010 !
b0010 #
#7390000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#7400000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#7410000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#7420000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#7430000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#7440000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#7450000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#7460000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#7470000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#7480000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#7490000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#7500000000
b1110 !
b1110 #
#7510000000
b1111 !
b1111 #
#7520000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#7530000000
b0001 !
b0001 #
#7540000000
b0010 !
b0010 #
#7550000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#7560000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#7570000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#7580000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#7590000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#7600000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#7610000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#7620000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#7630000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#7640000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#7650000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#7660000000
b1110 !
b1110 #
#7670000000
b1111 !
b1111 #
#7680000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#7690000000
b0001 !
b0001 #
#7700000000
b0010 !
b0010 #
#7710000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#7720000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#7730000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#7740000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#7750000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#7760000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#7770000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#7780000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#7790000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#7800000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#7810000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#7820000000
b1110 !
b1110 #
#7830000000
b1111 !
b1111 #
#7840000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#7850000000
b0001 !
b0001 #
#7860000000
b0010 !
b0010 #
#7870000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#7880000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#7890000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#7900000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#7910000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#7920000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#7930000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#7940000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#7950000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#7960000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#7970000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#7980000000
b1110 !
b1110 #
#7990000000
b1111 !
b1111 #
#8000000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#8010000000
b0001 !
b0001 #
#8020000000
b0010 !
b0010 #
#8030000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#8040000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#8050000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#8060000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#8070000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#8080000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#8090000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#8100000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#8110000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#8120000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#8130000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#8140000000
b1110 !
b1110 #
#8150000000
b1111 !
b1111 #
#8160000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#8170000000
b0001 !
b0001 #
#8180000000
b0010 !
b0010 #
#8190000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#8200000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#8210000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#8220000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#8230000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#8240000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#8250000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#8260000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#8270000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#8280000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#8290000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#8300000000
b1110 !
b1110 #
#8310000000
b1111 !
b1111 #
#8320000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#8330000000
b0001 !
b0001 #
#8340000000
b0010 !
b0010 #
#8350000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#8360000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#8370000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#8380000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#8390000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#8400000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#8410000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#8420000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#8430000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#8440000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#8450000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#8460000000
b1110 !
b1110 #
#8470000000
b1111 !
b1111 #
#8480000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#8490000000
b0001 !
b0001 #
#8500000000
b0010 !
b0010 #
#8510000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#8520000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#8530000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#8540000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#8550000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#8560000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#8570000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#8580000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#8590000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#8600000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#8610000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#8620000000
b1110 !
b1110 #
#8630000000
b1111 !
b1111 #
#8640000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#8650000000
b0001 !
b0001 #
#8660000000
b0010 !
b0010 #
#8670000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#8680000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#8690000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#8700000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#8710000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#8720000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#8730000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#8740000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#8750000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#8760000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#8770000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#8780000000
b1110 !
b1110 #
#8790000000
b1111 !
b1111 #
#8800000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#8810000000
b0001 !
b0001 #
#8820000000
b0010 !
b0010 #
#8830000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#8840000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#8850000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#8860000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#8870000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#8880000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#8890000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#8900000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#8910000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#8920000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#8930000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#8940000000
b1110 !
b1110 #
#8950000000
b1111 !
b1111 #
#8960000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#8970000000
b0001 !
b0001 #
#8980000000
b0010 !
b0010 #
#8990000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#9000000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#9010000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#9020000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#9030000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#9040000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#9050000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#9060000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#9070000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#9080000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#9090000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#9100000000
b1110 !
b1110 #
#9110000000
b1111 !
b1111 #
#9120000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#9130000000
b0001 !
b0001 #
#9140000000
b0010 !
b0010 #
#9150000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#9160000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#9170000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#9180000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#9190000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#9200000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#9210000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#9220000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#9230000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#9240000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#9250000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#9260000000
b1110 !
b1110 #
#9270000000
b1111 !
b1111 #
#9280000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#9290000000
b0001 !
b0001 #
#9300000000
b0010 !
b0010 #
#9310000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#9320000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#9330000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#9340000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#9350000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#9360000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#9370000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#9380000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#9390000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#9400000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#9410000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#9420000000
b1110 !
b1110 #
#9430000000
b1111 !
b1111 #
#9440000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#9450000000
b0001 !
b0001 #
#9460000000
b0010 !
b0010 #
#9470000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#9480000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#9490000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#9500000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#9510000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#9520000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#9530000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#9540000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#9550000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#9560000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#9570000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#9580000000
b1110 !
b1110 #
#9590000000
b1111 !
b1111 #
#9600000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#9610000000
b0001 !
b0001 #
#9620000000
b0010 !
b0010 #
#9630000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#9640000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#9650000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#9660000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#9670000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#9680000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#9690000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#9700000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#9710000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#9720000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#9730000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#9740000000
b1110 !
b1110 #
#9750000000
b1111 !
b1111 #
#9760000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#9770000000
b0001 !
b0001 #
#9780000000
b0010 !
b0010 #
#9790000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#9800000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#9810000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#9820000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#9830000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#9840000000
b1000 !
b1011110 "
b1000 #
b1011110 $
#9850000000
b1001 !
b1110111 "
b1001 #
b1110111 $
#9860000000
b1010 !
b1011110 "
b1010 #
b1011110 $
#9870000000
b1011 !
b1110111 "
b1011 #
b1110111 $
#9880000000
b1100 !
b1011110 "
b1100 #
b1011110 $
#9890000000
b1101 !
b1110111 "
b1101 #
b1110111 $
#9900000000
b1110 !
b1110 #
#9910000000
b1111 !
b1111 #
#9920000000
b0000 !
b1011110 "
b0000 #
b1011110 $
#9930000000
b0001 !
b0001 #
#9940000000
b0010 !
b0010 #
#9950000000
b0011 !
b1110111 "
b0011 #
b1110111 $
#9960000000
b0100 !
b1011110 "
b0100 #
b1011110 $
#9970000000
b0101 !
b1110111 "
b0101 #
b1110111 $
#9980000000
b0110 !
b1011110 "
b0110 #
b1011110 $
#9990000000
b0111 !
b1110111 "
b0111 #
b1110111 $
#10000000000
b1000 !
b1011110 "
b1000 #
b1011110 $
