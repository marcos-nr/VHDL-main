$date
  Sun May 12 23:26:07 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module textio $end
$upscope $end
$scope module tb_tp3_1 $end
$var integer 32 ! x $end
$var integer 32 " y $end
$var integer 32 # z $end
$scope module uut $end
$var integer 32 $ a $end
$var integer 32 % b $end
$var integer 32 & s $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
b101 !
b110000 "
b11110000 #
b101 $
b110000 %
b11110000 &
#10000000
#60000000
b110 !
b110111 "
b101001010 #
b110 $
b110111 %
b101001010 &
#70000000
#120000000
b101001 !
b110 "
b11110110 #
b101001 $
b110 %
b11110110 &
#130000000
#180000000
b111111 !
b10 "
b1111110 #
b111111 $
b10 %
b1111110 &
#190000000
#240000000
b11111 !
b1001 "
b100010111 #
b11111 $
b1001 %
b100010111 &
#250000000
#300000000
