$date
  Sat May 04 15:45:09 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_prueba $end
$var reg 1 ! clk $end
$var reg 1 " reset $end
$var reg 4 # dig3[3:0] $end
$var reg 4 $ dig2[3:0] $end
$var reg 4 % dig1[3:0] $end
$var reg 4 & dig0[3:0] $end
$var reg 4 ' enable_disp[3:0] $end
$var reg 7 ( segmentos[6:0] $end
$scope module uut $end
$var reg 1 ) clk $end
$var reg 1 * reset $end
$var reg 4 + dig3[3:0] $end
$var reg 4 , dig2[3:0] $end
$var reg 4 - dig1[3:0] $end
$var reg 4 . dig0[3:0] $end
$var reg 4 / enable_disp[3:0] $end
$var reg 7 0 segmentos[6:0] $end
$var reg 1 1 debounced_reset $end
$scope module d $end
$var reg 1 2 clk $end
$var reg 1 3 key $end
$var reg 1 4 debounced_key $end
$var reg 1 5 key_stable $end
$var reg 1 6 last_key $end
$upscope $end
$scope module a $end
$var reg 1 7 clk $end
$var reg 1 8 reset $end
$var reg 4 9 dig3[3:0] $end
$var reg 4 : dig2[3:0] $end
$var reg 4 ; dig1[3:0] $end
$var reg 4 < dig0[3:0] $end
$var reg 4 = enable_disp[3:0] $end
$var reg 7 > segmentos[6:0] $end
$comment state is not handled $end
$var integer 32 ? cuenta $end
$var reg 1 @ debounced_reset $end
$var reg 1 A enable_conta $end
$var reg 4 B bcd[3:0] $end
$scope module a $end
$var reg 1 C clk $end
$var reg 1 D key $end
$var reg 1 E debounced_key $end
$var reg 1 F key_stable $end
$var reg 1 G last_key $end
$upscope $end
$scope module b $end
$var reg 1 H clk $end
$var reg 1 I reset $end
$var reg 1 J enable $end
$var reg 1 K cout $end
$var integer 32 L q $end
$upscope $end
$scope module d $end
$var reg 7 M segmentos[6:0] $end
$var reg 4 N bcd[3:0] $end
$upscope $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
0"
b1000 #
b0110 $
b0100 %
b0010 &
b0001 '
b0111000 (
0)
0*
b1000 +
b0110 ,
b0100 -
b0010 .
b0001 /
b0111000 0
U1
02
03
U4
U5
U6
07
08
b1000 9
b0110 :
b0100 ;
b0010 <
b0001 =
b0111000 >
b0 ?
U@
1A
bUUUU B
0C
0D
UE
UF
UG
0H
UI
1J
UK
b0 L
b0111000 M
bUUUU N
#10000000
1!
1)
01
12
04
05
06
17
0@
1C
0E
0F
0G
1H
0I
0K
#20000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#30000000
1!
1)
12
17
1C
1H
#40000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#50000000
1!
1)
12
17
1C
1H
#60000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#70000000
1!
1)
12
17
1C
1H
1K
#80000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#90000000
1!
1)
12
17
1C
1H
#100000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#110000000
1!
1)
12
17
1C
1H
#120000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#130000000
1!
1)
12
17
1C
1H
#140000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#150000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#160000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#170000000
1!
1)
12
17
1C
1H
#180000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#190000000
1!
1)
12
17
1C
1H
#200000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#210000000
1!
1)
12
17
1C
1H
#220000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#230000000
1!
1)
12
17
1C
1H
1K
#240000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#250000000
1!
1)
12
17
1C
1H
#260000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#270000000
1!
1)
12
17
1C
1H
#280000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#290000000
1!
1)
12
17
1C
1H
#300000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#310000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#320000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#330000000
1!
1)
12
17
1C
1H
#340000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#350000000
1!
1)
12
17
1C
1H
#360000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#370000000
1!
1)
12
17
1C
1H
#380000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#390000000
1!
1)
12
17
1C
1H
1K
#400000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#410000000
1!
1)
12
17
1C
1H
#420000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#430000000
1!
1)
12
17
1C
1H
#440000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#450000000
1!
1)
12
17
1C
1H
#460000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#470000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#480000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#490000000
1!
1)
12
17
1C
1H
#500000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#510000000
1!
1)
12
17
1C
1H
#520000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#530000000
1!
1)
12
17
1C
1H
#540000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#550000000
1!
1)
12
17
1C
1H
1K
#560000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#570000000
1!
1)
12
17
1C
1H
#580000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#590000000
1!
1)
12
17
1C
1H
#600000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#610000000
1!
1)
12
17
1C
1H
#620000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#630000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#640000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#650000000
1!
1)
12
17
1C
1H
#660000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#670000000
1!
1)
12
17
1C
1H
#680000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#690000000
1!
1)
12
17
1C
1H
#700000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#710000000
1!
1)
12
17
1C
1H
1K
#720000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#730000000
1!
1)
12
17
1C
1H
#740000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#750000000
1!
1)
12
17
1C
1H
#760000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#770000000
1!
1)
12
17
1C
1H
#780000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#790000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#800000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#810000000
1!
1)
12
17
1C
1H
#820000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#830000000
1!
1)
12
17
1C
1H
#840000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#850000000
1!
1)
12
17
1C
1H
#860000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#870000000
1!
1)
12
17
1C
1H
1K
#880000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#890000000
1!
1)
12
17
1C
1H
#900000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#910000000
1!
1)
12
17
1C
1H
#920000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#930000000
1!
1)
12
17
1C
1H
#940000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#950000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#960000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#970000000
1!
1)
12
17
1C
1H
#980000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#990000000
1!
1)
12
17
1C
1H
#1000000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#1010000000
1!
1)
12
17
1C
1H
#1020000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#1030000000
1!
1)
12
17
1C
1H
1K
#1040000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#1050000000
1!
1)
12
17
1C
1H
#1060000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#1070000000
1!
1)
12
17
1C
1H
#1080000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#1090000000
1!
1)
12
17
1C
1H
#1100000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#1110000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#1120000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#1130000000
1!
1)
12
17
1C
1H
#1140000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#1150000000
1!
1)
12
17
1C
1H
#1160000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#1170000000
1!
1)
12
17
1C
1H
#1180000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#1190000000
1!
1)
12
17
1C
1H
1K
#1200000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#1210000000
1!
1)
12
17
1C
1H
#1220000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#1230000000
1!
1)
12
17
1C
1H
#1240000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#1250000000
1!
1)
12
17
1C
1H
#1260000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#1270000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#1280000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#1290000000
1!
1)
12
17
1C
1H
#1300000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#1310000000
1!
1)
12
17
1C
1H
#1320000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#1330000000
1!
1)
12
17
1C
1H
#1340000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#1350000000
1!
1)
12
17
1C
1H
1K
#1360000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#1370000000
1!
1)
12
17
1C
1H
#1380000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#1390000000
1!
1)
12
17
1C
1H
#1400000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#1410000000
1!
1)
12
17
1C
1H
#1420000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#1430000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#1440000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#1450000000
1!
1)
12
17
1C
1H
#1460000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#1470000000
1!
1)
12
17
1C
1H
#1480000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#1490000000
1!
1)
12
17
1C
1H
#1500000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#1510000000
1!
1)
12
17
1C
1H
1K
#1520000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#1530000000
1!
1)
12
17
1C
1H
#1540000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#1550000000
1!
1)
12
17
1C
1H
#1560000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#1570000000
1!
1)
12
17
1C
1H
#1580000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#1590000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#1600000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#1610000000
1!
1)
12
17
1C
1H
#1620000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#1630000000
1!
1)
12
17
1C
1H
#1640000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#1650000000
1!
1)
12
17
1C
1H
#1660000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#1670000000
1!
1)
12
17
1C
1H
1K
#1680000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#1690000000
1!
1)
12
17
1C
1H
#1700000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#1710000000
1!
1)
12
17
1C
1H
#1720000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#1730000000
1!
1)
12
17
1C
1H
#1740000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#1750000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#1760000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#1770000000
1!
1)
12
17
1C
1H
#1780000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#1790000000
1!
1)
12
17
1C
1H
#1800000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#1810000000
1!
1)
12
17
1C
1H
#1820000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#1830000000
1!
1)
12
17
1C
1H
1K
#1840000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#1850000000
1!
1)
12
17
1C
1H
#1860000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#1870000000
1!
1)
12
17
1C
1H
#1880000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#1890000000
1!
1)
12
17
1C
1H
#1900000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#1910000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#1920000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#1930000000
1!
1)
12
17
1C
1H
#1940000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#1950000000
1!
1)
12
17
1C
1H
#1960000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#1970000000
1!
1)
12
17
1C
1H
#1980000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#1990000000
1!
1)
12
17
1C
1H
1K
#2000000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#2010000000
1!
1)
12
17
1C
1H
#2020000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#2030000000
1!
1)
12
17
1C
1H
#2040000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#2050000000
1!
1)
12
17
1C
1H
#2060000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#2070000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#2080000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#2090000000
1!
1)
12
17
1C
1H
#2100000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#2110000000
1!
1)
12
17
1C
1H
#2120000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#2130000000
1!
1)
12
17
1C
1H
#2140000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#2150000000
1!
1)
12
17
1C
1H
1K
#2160000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#2170000000
1!
1)
12
17
1C
1H
#2180000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#2190000000
1!
1)
12
17
1C
1H
#2200000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#2210000000
1!
1)
12
17
1C
1H
#2220000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#2230000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#2240000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#2250000000
1!
1)
12
17
1C
1H
#2260000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#2270000000
1!
1)
12
17
1C
1H
#2280000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#2290000000
1!
1)
12
17
1C
1H
#2300000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#2310000000
1!
1)
12
17
1C
1H
1K
#2320000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#2330000000
1!
1)
12
17
1C
1H
#2340000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#2350000000
1!
1)
12
17
1C
1H
#2360000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#2370000000
1!
1)
12
17
1C
1H
#2380000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#2390000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#2400000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#2410000000
1!
1)
12
17
1C
1H
#2420000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#2430000000
1!
1)
12
17
1C
1H
#2440000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#2450000000
1!
1)
12
17
1C
1H
#2460000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#2470000000
1!
1)
12
17
1C
1H
1K
#2480000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#2490000000
1!
1)
12
17
1C
1H
#2500000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#2510000000
1!
1)
12
17
1C
1H
#2520000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#2530000000
1!
1)
12
17
1C
1H
#2540000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#2550000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#2560000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#2570000000
1!
1)
12
17
1C
1H
#2580000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#2590000000
1!
1)
12
17
1C
1H
#2600000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#2610000000
1!
1)
12
17
1C
1H
#2620000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#2630000000
1!
1)
12
17
1C
1H
1K
#2640000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#2650000000
1!
1)
12
17
1C
1H
#2660000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#2670000000
1!
1)
12
17
1C
1H
#2680000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#2690000000
1!
1)
12
17
1C
1H
#2700000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#2710000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#2720000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#2730000000
1!
1)
12
17
1C
1H
#2740000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#2750000000
1!
1)
12
17
1C
1H
#2760000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#2770000000
1!
1)
12
17
1C
1H
#2780000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#2790000000
1!
1)
12
17
1C
1H
1K
#2800000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#2810000000
1!
1)
12
17
1C
1H
#2820000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#2830000000
1!
1)
12
17
1C
1H
#2840000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#2850000000
1!
1)
12
17
1C
1H
#2860000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#2870000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#2880000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#2890000000
1!
1)
12
17
1C
1H
#2900000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#2910000000
1!
1)
12
17
1C
1H
#2920000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#2930000000
1!
1)
12
17
1C
1H
#2940000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#2950000000
1!
1)
12
17
1C
1H
1K
#2960000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#2970000000
1!
1)
12
17
1C
1H
#2980000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#2990000000
1!
1)
12
17
1C
1H
#3000000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#3010000000
1!
1)
12
17
1C
1H
#3020000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#3030000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#3040000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#3050000000
1!
1)
12
17
1C
1H
#3060000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#3070000000
1!
1)
12
17
1C
1H
#3080000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#3090000000
1!
1)
12
17
1C
1H
#3100000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#3110000000
1!
1)
12
17
1C
1H
1K
#3120000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#3130000000
1!
1)
12
17
1C
1H
#3140000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#3150000000
1!
1)
12
17
1C
1H
#3160000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#3170000000
1!
1)
12
17
1C
1H
#3180000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#3190000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#3200000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#3210000000
1!
1)
12
17
1C
1H
#3220000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#3230000000
1!
1)
12
17
1C
1H
#3240000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#3250000000
1!
1)
12
17
1C
1H
#3260000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#3270000000
1!
1)
12
17
1C
1H
1K
#3280000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#3290000000
1!
1)
12
17
1C
1H
#3300000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#3310000000
1!
1)
12
17
1C
1H
#3320000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#3330000000
1!
1)
12
17
1C
1H
#3340000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#3350000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#3360000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#3370000000
1!
1)
12
17
1C
1H
#3380000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#3390000000
1!
1)
12
17
1C
1H
#3400000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#3410000000
1!
1)
12
17
1C
1H
#3420000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#3430000000
1!
1)
12
17
1C
1H
1K
#3440000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#3450000000
1!
1)
12
17
1C
1H
#3460000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#3470000000
1!
1)
12
17
1C
1H
#3480000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#3490000000
1!
1)
12
17
1C
1H
#3500000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#3510000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#3520000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#3530000000
1!
1)
12
17
1C
1H
#3540000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#3550000000
1!
1)
12
17
1C
1H
#3560000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#3570000000
1!
1)
12
17
1C
1H
#3580000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#3590000000
1!
1)
12
17
1C
1H
1K
#3600000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#3610000000
1!
1)
12
17
1C
1H
#3620000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#3630000000
1!
1)
12
17
1C
1H
#3640000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#3650000000
1!
1)
12
17
1C
1H
#3660000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#3670000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#3680000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#3690000000
1!
1)
12
17
1C
1H
#3700000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#3710000000
1!
1)
12
17
1C
1H
#3720000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#3730000000
1!
1)
12
17
1C
1H
#3740000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#3750000000
1!
1)
12
17
1C
1H
1K
#3760000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#3770000000
1!
1)
12
17
1C
1H
#3780000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#3790000000
1!
1)
12
17
1C
1H
#3800000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#3810000000
1!
1)
12
17
1C
1H
#3820000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#3830000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#3840000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#3850000000
1!
1)
12
17
1C
1H
#3860000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#3870000000
1!
1)
12
17
1C
1H
#3880000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#3890000000
1!
1)
12
17
1C
1H
#3900000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#3910000000
1!
1)
12
17
1C
1H
1K
#3920000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#3930000000
1!
1)
12
17
1C
1H
#3940000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#3950000000
1!
1)
12
17
1C
1H
#3960000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#3970000000
1!
1)
12
17
1C
1H
#3980000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#3990000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#4000000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#4010000000
1!
1)
12
17
1C
1H
#4020000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#4030000000
1!
1)
12
17
1C
1H
#4040000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#4050000000
1!
1)
12
17
1C
1H
#4060000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#4070000000
1!
1)
12
17
1C
1H
1K
#4080000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#4090000000
1!
1)
12
17
1C
1H
#4100000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#4110000000
1!
1)
12
17
1C
1H
#4120000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#4130000000
1!
1)
12
17
1C
1H
#4140000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#4150000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#4160000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#4170000000
1!
1)
12
17
1C
1H
#4180000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#4190000000
1!
1)
12
17
1C
1H
#4200000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#4210000000
1!
1)
12
17
1C
1H
#4220000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#4230000000
1!
1)
12
17
1C
1H
1K
#4240000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#4250000000
1!
1)
12
17
1C
1H
#4260000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#4270000000
1!
1)
12
17
1C
1H
#4280000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#4290000000
1!
1)
12
17
1C
1H
#4300000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#4310000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#4320000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#4330000000
1!
1)
12
17
1C
1H
#4340000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#4350000000
1!
1)
12
17
1C
1H
#4360000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#4370000000
1!
1)
12
17
1C
1H
#4380000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#4390000000
1!
1)
12
17
1C
1H
1K
#4400000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#4410000000
1!
1)
12
17
1C
1H
#4420000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#4430000000
1!
1)
12
17
1C
1H
#4440000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#4450000000
1!
1)
12
17
1C
1H
#4460000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#4470000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#4480000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#4490000000
1!
1)
12
17
1C
1H
#4500000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#4510000000
1!
1)
12
17
1C
1H
#4520000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#4530000000
1!
1)
12
17
1C
1H
#4540000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#4550000000
1!
1)
12
17
1C
1H
1K
#4560000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#4570000000
1!
1)
12
17
1C
1H
#4580000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#4590000000
1!
1)
12
17
1C
1H
#4600000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#4610000000
1!
1)
12
17
1C
1H
#4620000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#4630000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#4640000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#4650000000
1!
1)
12
17
1C
1H
#4660000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#4670000000
1!
1)
12
17
1C
1H
#4680000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#4690000000
1!
1)
12
17
1C
1H
#4700000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#4710000000
1!
1)
12
17
1C
1H
1K
#4720000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#4730000000
1!
1)
12
17
1C
1H
#4740000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#4750000000
1!
1)
12
17
1C
1H
#4760000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#4770000000
1!
1)
12
17
1C
1H
#4780000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#4790000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#4800000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#4810000000
1!
1)
12
17
1C
1H
#4820000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#4830000000
1!
1)
12
17
1C
1H
#4840000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#4850000000
1!
1)
12
17
1C
1H
#4860000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#4870000000
1!
1)
12
17
1C
1H
1K
#4880000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#4890000000
1!
1)
12
17
1C
1H
#4900000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#4910000000
1!
1)
12
17
1C
1H
#4920000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#4930000000
1!
1)
12
17
1C
1H
#4940000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#4950000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#4960000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#4970000000
1!
1)
12
17
1C
1H
#4980000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#4990000000
1!
1)
12
17
1C
1H
#5000000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#5010000000
1!
1)
12
17
1C
1H
#5020000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#5030000000
1!
1)
12
17
1C
1H
1K
#5040000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#5050000000
1!
1)
12
17
1C
1H
#5060000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#5070000000
1!
1)
12
17
1C
1H
#5080000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#5090000000
1!
1)
12
17
1C
1H
#5100000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#5110000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#5120000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#5130000000
1!
1)
12
17
1C
1H
#5140000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#5150000000
1!
1)
12
17
1C
1H
#5160000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#5170000000
1!
1)
12
17
1C
1H
#5180000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#5190000000
1!
1)
12
17
1C
1H
1K
#5200000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#5210000000
1!
1)
12
17
1C
1H
#5220000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#5230000000
1!
1)
12
17
1C
1H
#5240000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#5250000000
1!
1)
12
17
1C
1H
#5260000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#5270000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#5280000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#5290000000
1!
1)
12
17
1C
1H
#5300000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#5310000000
1!
1)
12
17
1C
1H
#5320000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#5330000000
1!
1)
12
17
1C
1H
#5340000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#5350000000
1!
1)
12
17
1C
1H
1K
#5360000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#5370000000
1!
1)
12
17
1C
1H
#5380000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#5390000000
1!
1)
12
17
1C
1H
#5400000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#5410000000
1!
1)
12
17
1C
1H
#5420000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#5430000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#5440000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#5450000000
1!
1)
12
17
1C
1H
#5460000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#5470000000
1!
1)
12
17
1C
1H
#5480000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#5490000000
1!
1)
12
17
1C
1H
#5500000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#5510000000
1!
1)
12
17
1C
1H
1K
#5520000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#5530000000
1!
1)
12
17
1C
1H
#5540000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#5550000000
1!
1)
12
17
1C
1H
#5560000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#5570000000
1!
1)
12
17
1C
1H
#5580000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#5590000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#5600000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#5610000000
1!
1)
12
17
1C
1H
#5620000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#5630000000
1!
1)
12
17
1C
1H
#5640000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#5650000000
1!
1)
12
17
1C
1H
#5660000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#5670000000
1!
1)
12
17
1C
1H
1K
#5680000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#5690000000
1!
1)
12
17
1C
1H
#5700000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#5710000000
1!
1)
12
17
1C
1H
#5720000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#5730000000
1!
1)
12
17
1C
1H
#5740000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#5750000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#5760000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#5770000000
1!
1)
12
17
1C
1H
#5780000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#5790000000
1!
1)
12
17
1C
1H
#5800000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#5810000000
1!
1)
12
17
1C
1H
#5820000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#5830000000
1!
1)
12
17
1C
1H
1K
#5840000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#5850000000
1!
1)
12
17
1C
1H
#5860000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#5870000000
1!
1)
12
17
1C
1H
#5880000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#5890000000
1!
1)
12
17
1C
1H
#5900000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#5910000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#5920000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#5930000000
1!
1)
12
17
1C
1H
#5940000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#5950000000
1!
1)
12
17
1C
1H
#5960000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#5970000000
1!
1)
12
17
1C
1H
#5980000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#5990000000
1!
1)
12
17
1C
1H
1K
#6000000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#6010000000
1!
1)
12
17
1C
1H
#6020000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#6030000000
1!
1)
12
17
1C
1H
#6040000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#6050000000
1!
1)
12
17
1C
1H
#6060000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#6070000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#6080000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#6090000000
1!
1)
12
17
1C
1H
#6100000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#6110000000
1!
1)
12
17
1C
1H
#6120000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#6130000000
1!
1)
12
17
1C
1H
#6140000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#6150000000
1!
1)
12
17
1C
1H
1K
#6160000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#6170000000
1!
1)
12
17
1C
1H
#6180000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#6190000000
1!
1)
12
17
1C
1H
#6200000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#6210000000
1!
1)
12
17
1C
1H
#6220000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#6230000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#6240000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#6250000000
1!
1)
12
17
1C
1H
#6260000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#6270000000
1!
1)
12
17
1C
1H
#6280000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#6290000000
1!
1)
12
17
1C
1H
#6300000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#6310000000
1!
1)
12
17
1C
1H
1K
#6320000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#6330000000
1!
1)
12
17
1C
1H
#6340000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#6350000000
1!
1)
12
17
1C
1H
#6360000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#6370000000
1!
1)
12
17
1C
1H
#6380000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#6390000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#6400000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#6410000000
1!
1)
12
17
1C
1H
#6420000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#6430000000
1!
1)
12
17
1C
1H
#6440000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#6450000000
1!
1)
12
17
1C
1H
#6460000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#6470000000
1!
1)
12
17
1C
1H
1K
#6480000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#6490000000
1!
1)
12
17
1C
1H
#6500000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#6510000000
1!
1)
12
17
1C
1H
#6520000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#6530000000
1!
1)
12
17
1C
1H
#6540000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#6550000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#6560000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#6570000000
1!
1)
12
17
1C
1H
#6580000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#6590000000
1!
1)
12
17
1C
1H
#6600000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#6610000000
1!
1)
12
17
1C
1H
#6620000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#6630000000
1!
1)
12
17
1C
1H
1K
#6640000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#6650000000
1!
1)
12
17
1C
1H
#6660000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#6670000000
1!
1)
12
17
1C
1H
#6680000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#6690000000
1!
1)
12
17
1C
1H
#6700000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#6710000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#6720000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#6730000000
1!
1)
12
17
1C
1H
#6740000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#6750000000
1!
1)
12
17
1C
1H
#6760000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#6770000000
1!
1)
12
17
1C
1H
#6780000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#6790000000
1!
1)
12
17
1C
1H
1K
#6800000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#6810000000
1!
1)
12
17
1C
1H
#6820000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#6830000000
1!
1)
12
17
1C
1H
#6840000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#6850000000
1!
1)
12
17
1C
1H
#6860000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#6870000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#6880000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#6890000000
1!
1)
12
17
1C
1H
#6900000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#6910000000
1!
1)
12
17
1C
1H
#6920000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#6930000000
1!
1)
12
17
1C
1H
#6940000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#6950000000
1!
1)
12
17
1C
1H
1K
#6960000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#6970000000
1!
1)
12
17
1C
1H
#6980000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#6990000000
1!
1)
12
17
1C
1H
#7000000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#7010000000
1!
1)
12
17
1C
1H
#7020000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#7030000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#7040000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#7050000000
1!
1)
12
17
1C
1H
#7060000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#7070000000
1!
1)
12
17
1C
1H
#7080000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#7090000000
1!
1)
12
17
1C
1H
#7100000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#7110000000
1!
1)
12
17
1C
1H
1K
#7120000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#7130000000
1!
1)
12
17
1C
1H
#7140000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#7150000000
1!
1)
12
17
1C
1H
#7160000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#7170000000
1!
1)
12
17
1C
1H
#7180000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#7190000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#7200000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#7210000000
1!
1)
12
17
1C
1H
#7220000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#7230000000
1!
1)
12
17
1C
1H
#7240000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#7250000000
1!
1)
12
17
1C
1H
#7260000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#7270000000
1!
1)
12
17
1C
1H
1K
#7280000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#7290000000
1!
1)
12
17
1C
1H
#7300000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#7310000000
1!
1)
12
17
1C
1H
#7320000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#7330000000
1!
1)
12
17
1C
1H
#7340000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#7350000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#7360000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#7370000000
1!
1)
12
17
1C
1H
#7380000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#7390000000
1!
1)
12
17
1C
1H
#7400000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#7410000000
1!
1)
12
17
1C
1H
#7420000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#7430000000
1!
1)
12
17
1C
1H
1K
#7440000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#7450000000
1!
1)
12
17
1C
1H
#7460000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#7470000000
1!
1)
12
17
1C
1H
#7480000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#7490000000
1!
1)
12
17
1C
1H
#7500000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#7510000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#7520000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#7530000000
1!
1)
12
17
1C
1H
#7540000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#7550000000
1!
1)
12
17
1C
1H
#7560000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#7570000000
1!
1)
12
17
1C
1H
#7580000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#7590000000
1!
1)
12
17
1C
1H
1K
#7600000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#7610000000
1!
1)
12
17
1C
1H
#7620000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#7630000000
1!
1)
12
17
1C
1H
#7640000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#7650000000
1!
1)
12
17
1C
1H
#7660000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#7670000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#7680000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#7690000000
1!
1)
12
17
1C
1H
#7700000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#7710000000
1!
1)
12
17
1C
1H
#7720000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#7730000000
1!
1)
12
17
1C
1H
#7740000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#7750000000
1!
1)
12
17
1C
1H
1K
#7760000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#7770000000
1!
1)
12
17
1C
1H
#7780000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#7790000000
1!
1)
12
17
1C
1H
#7800000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#7810000000
1!
1)
12
17
1C
1H
#7820000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#7830000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#7840000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#7850000000
1!
1)
12
17
1C
1H
#7860000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#7870000000
1!
1)
12
17
1C
1H
#7880000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#7890000000
1!
1)
12
17
1C
1H
#7900000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#7910000000
1!
1)
12
17
1C
1H
1K
#7920000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#7930000000
1!
1)
12
17
1C
1H
#7940000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#7950000000
1!
1)
12
17
1C
1H
#7960000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#7970000000
1!
1)
12
17
1C
1H
#7980000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#7990000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#8000000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#8010000000
1!
1)
12
17
1C
1H
#8020000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#8030000000
1!
1)
12
17
1C
1H
#8040000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#8050000000
1!
1)
12
17
1C
1H
#8060000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#8070000000
1!
1)
12
17
1C
1H
1K
#8080000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#8090000000
1!
1)
12
17
1C
1H
#8100000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#8110000000
1!
1)
12
17
1C
1H
#8120000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#8130000000
1!
1)
12
17
1C
1H
#8140000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#8150000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#8160000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#8170000000
1!
1)
12
17
1C
1H
#8180000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#8190000000
1!
1)
12
17
1C
1H
#8200000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#8210000000
1!
1)
12
17
1C
1H
#8220000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#8230000000
1!
1)
12
17
1C
1H
1K
#8240000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#8250000000
1!
1)
12
17
1C
1H
#8260000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#8270000000
1!
1)
12
17
1C
1H
#8280000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#8290000000
1!
1)
12
17
1C
1H
#8300000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#8310000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#8320000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#8330000000
1!
1)
12
17
1C
1H
#8340000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#8350000000
1!
1)
12
17
1C
1H
#8360000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#8370000000
1!
1)
12
17
1C
1H
#8380000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#8390000000
1!
1)
12
17
1C
1H
1K
#8400000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#8410000000
1!
1)
12
17
1C
1H
#8420000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#8430000000
1!
1)
12
17
1C
1H
#8440000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#8450000000
1!
1)
12
17
1C
1H
#8460000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#8470000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#8480000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#8490000000
1!
1)
12
17
1C
1H
#8500000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#8510000000
1!
1)
12
17
1C
1H
#8520000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#8530000000
1!
1)
12
17
1C
1H
#8540000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#8550000000
1!
1)
12
17
1C
1H
1K
#8560000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#8570000000
1!
1)
12
17
1C
1H
#8580000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#8590000000
1!
1)
12
17
1C
1H
#8600000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#8610000000
1!
1)
12
17
1C
1H
#8620000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#8630000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#8640000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#8650000000
1!
1)
12
17
1C
1H
#8660000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#8670000000
1!
1)
12
17
1C
1H
#8680000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#8690000000
1!
1)
12
17
1C
1H
#8700000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#8710000000
1!
1)
12
17
1C
1H
1K
#8720000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#8730000000
1!
1)
12
17
1C
1H
#8740000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#8750000000
1!
1)
12
17
1C
1H
#8760000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#8770000000
1!
1)
12
17
1C
1H
#8780000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#8790000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#8800000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#8810000000
1!
1)
12
17
1C
1H
#8820000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#8830000000
1!
1)
12
17
1C
1H
#8840000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#8850000000
1!
1)
12
17
1C
1H
#8860000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#8870000000
1!
1)
12
17
1C
1H
1K
#8880000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#8890000000
1!
1)
12
17
1C
1H
#8900000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#8910000000
1!
1)
12
17
1C
1H
#8920000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#8930000000
1!
1)
12
17
1C
1H
#8940000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#8950000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#8960000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#8970000000
1!
1)
12
17
1C
1H
#8980000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#8990000000
1!
1)
12
17
1C
1H
#9000000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#9010000000
1!
1)
12
17
1C
1H
#9020000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#9030000000
1!
1)
12
17
1C
1H
1K
#9040000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#9050000000
1!
1)
12
17
1C
1H
#9060000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#9070000000
1!
1)
12
17
1C
1H
#9080000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#9090000000
1!
1)
12
17
1C
1H
#9100000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#9110000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#9120000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#9130000000
1!
1)
12
17
1C
1H
#9140000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#9150000000
1!
1)
12
17
1C
1H
#9160000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#9170000000
1!
1)
12
17
1C
1H
#9180000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#9190000000
1!
1)
12
17
1C
1H
1K
#9200000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#9210000000
1!
1)
12
17
1C
1H
#9220000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#9230000000
1!
1)
12
17
1C
1H
#9240000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#9250000000
1!
1)
12
17
1C
1H
#9260000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#9270000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#9280000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#9290000000
1!
1)
12
17
1C
1H
#9300000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#9310000000
1!
1)
12
17
1C
1H
#9320000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#9330000000
1!
1)
12
17
1C
1H
#9340000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#9350000000
1!
1)
12
17
1C
1H
1K
#9360000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#9370000000
1!
1)
12
17
1C
1H
#9380000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#9390000000
1!
1)
12
17
1C
1H
#9400000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#9410000000
1!
1)
12
17
1C
1H
#9420000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#9430000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
12
17
b1000 =
b0000000 >
b1000 B
1C
1H
0K
b0000000 M
b1000 N
#9440000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#9450000000
1!
1)
12
17
1C
1H
#9460000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#9470000000
1!
1)
12
17
1C
1H
#9480000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#9490000000
1!
1)
12
17
1C
1H
#9500000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#9510000000
1!
1)
12
17
1C
1H
1K
#9520000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#9530000000
1!
1)
12
17
1C
1H
#9540000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#9550000000
1!
1)
12
17
1C
1H
#9560000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#9570000000
1!
1)
12
17
1C
1H
#9580000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#9590000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
12
17
b0001 =
b0010010 >
b0010 B
1C
1H
0K
b0010010 M
b0010 N
#9600000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#9610000000
1!
1)
12
17
1C
1H
#9620000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#9630000000
1!
1)
12
17
1C
1H
#9640000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#9650000000
1!
1)
12
17
1C
1H
#9660000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#9670000000
1!
1)
12
17
1C
1H
1K
#9680000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#9690000000
1!
1)
12
17
1C
1H
#9700000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#9710000000
1!
1)
12
17
1C
1H
#9720000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#9730000000
1!
1)
12
17
1C
1H
#9740000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#9750000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
12
17
b0010 =
b1001100 >
b0100 B
1C
1H
0K
b1001100 M
b0100 N
#9760000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#9770000000
1!
1)
12
17
1C
1H
#9780000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#9790000000
1!
1)
12
17
1C
1H
#9800000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#9810000000
1!
1)
12
17
1C
1H
#9820000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#9830000000
1!
1)
12
17
1C
1H
1K
#9840000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
#9850000000
1!
1)
12
17
1C
1H
#9860000000
0!
0)
02
07
b101 ?
0C
0H
b101 L
#9870000000
1!
1)
12
17
1C
1H
#9880000000
0!
0)
02
07
b110 ?
0C
0H
b110 L
#9890000000
1!
1)
12
17
1C
1H
#9900000000
0!
0)
02
07
b111 ?
0C
0H
b111 L
#9910000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
12
17
b0100 =
b0100000 >
b0110 B
1C
1H
0K
b0100000 M
b0110 N
#9920000000
0!
0)
02
07
b0 ?
0C
0H
b0 L
#9930000000
1!
1)
12
17
1C
1H
#9940000000
0!
0)
02
07
b1 ?
0C
0H
b1 L
#9950000000
1!
1)
12
17
1C
1H
#9960000000
0!
0)
02
07
b10 ?
0C
0H
b10 L
#9970000000
1!
1)
12
17
1C
1H
#9980000000
0!
0)
02
07
b11 ?
0C
0H
b11 L
#9990000000
1!
1)
12
17
1C
1H
1K
#10000000000
0!
0)
02
07
b100 ?
0C
0H
b100 L
