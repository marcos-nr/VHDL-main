$date
  Mon Jun 24 20:07:30 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_pwm $end
$var reg 1 ! clk $end
$var reg 1 " reset $end
$var reg 1 # enable $end
$var reg 1 $ cout $end
$var integer 32 % q $end
$var integer 32 & duty $end
$scope module uud $end
$var reg 1 ' clk $end
$var reg 1 ( reset $end
$var reg 1 ) enable $end
$var reg 1 * cout $end
$var integer 32 + q $end
$var integer 32 , duty $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
1!
0"
1#
1$
b1 %
b10 &
1'
0(
1)
1*
b1 +
b10 ,
#10000000
0!
0'
#20000000
1!
b10 %
1'
b10 +
#30000000
0!
0'
#40000000
1!
b11 %
1'
b11 +
#50000000
0!
0'
#60000000
1!
b100 %
1'
b100 +
#70000000
0!
0'
#80000000
1!
b101 %
1'
b101 +
#90000000
0!
0'
#100000000
1!
0$
b110 %
1'
0*
b110 +
#110000000
0!
0'
#120000000
1!
b111 %
1'
b111 +
#130000000
0!
0'
#140000000
1!
b1000 %
1'
b1000 +
#150000000
0!
0'
#160000000
1!
b1001 %
1'
b1001 +
#170000000
0!
0'
#180000000
1!
b0 %
1'
b0 +
#190000000
0!
0'
#200000000
1!
1$
b1 %
1'
1*
b1 +
#210000000
1"
1(
#220000000
0!
0"
b100 &
0'
0(
b100 ,
#230000000
1!
b10 %
1'
b10 +
#240000000
0!
0'
#250000000
1!
b11 %
1'
b11 +
#260000000
0!
0'
#270000000
1!
b100 %
1'
b100 +
#280000000
0!
0'
#290000000
1!
b101 %
1'
b101 +
#300000000
0!
0'
#310000000
1!
b110 %
1'
b110 +
#320000000
0!
0'
#330000000
1!
b111 %
1'
b111 +
#340000000
0!
0'
#350000000
1!
0$
b1000 %
1'
0*
b1000 +
#360000000
0!
0'
#370000000
1!
b1001 %
1'
b1001 +
#380000000
0!
0'
#390000000
1!
b0 %
1'
b0 +
#400000000
0!
0'
#410000000
1!
1$
b1 %
1'
1*
b1 +
#420000000
0!
0'
#430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#440000000
0!
0'
#450000000
1!
b11 %
1'
b11 +
#460000000
0!
0'
#470000000
1!
b100 %
1'
b100 +
#480000000
0!
0'
#490000000
1!
b101 %
1'
b101 +
#500000000
0!
0'
#510000000
1!
0$
b110 %
1'
0*
b110 +
#520000000
0!
0'
#530000000
1!
b111 %
1'
b111 +
#540000000
0!
0'
#550000000
1!
b1000 %
1'
b1000 +
#560000000
0!
0'
#570000000
1!
b1001 %
1'
b1001 +
#580000000
0!
0'
#590000000
1!
b0 %
1'
b0 +
#600000000
0!
0'
#610000000
1!
1$
b1 %
1'
1*
b1 +
#620000000
0!
0'
#630000000
1!
b10 %
1'
b10 +
#640000000
1"
1(
#650000000
0!
0"
b100 &
0'
0(
b100 ,
#660000000
1!
b11 %
1'
b11 +
#670000000
0!
0'
#680000000
1!
b100 %
1'
b100 +
#690000000
0!
0'
#700000000
1!
b101 %
1'
b101 +
#710000000
0!
0'
#720000000
1!
b110 %
1'
b110 +
#730000000
0!
0'
#740000000
1!
b111 %
1'
b111 +
#750000000
0!
0'
#760000000
1!
0$
b1000 %
1'
0*
b1000 +
#770000000
0!
0'
#780000000
1!
b1001 %
1'
b1001 +
#790000000
0!
0'
#800000000
1!
b0 %
1'
b0 +
#810000000
0!
0'
#820000000
1!
1$
b1 %
1'
1*
b1 +
#830000000
0!
0'
#840000000
1!
b10 %
1'
b10 +
#850000000
0!
0'
#860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#870000000
0!
0'
#880000000
1!
b100 %
1'
b100 +
#890000000
0!
0'
#900000000
1!
b101 %
1'
b101 +
#910000000
0!
0'
#920000000
1!
0$
b110 %
1'
0*
b110 +
#930000000
0!
0'
#940000000
1!
b111 %
1'
b111 +
#950000000
0!
0'
#960000000
1!
b1000 %
1'
b1000 +
#970000000
0!
0'
#980000000
1!
b1001 %
1'
b1001 +
#990000000
0!
0'
#1000000000
1!
b0 %
1'
b0 +
#1010000000
0!
0'
#1020000000
1!
1$
b1 %
1'
1*
b1 +
#1030000000
0!
0'
#1040000000
1!
b10 %
1'
b10 +
#1050000000
0!
0'
#1060000000
1!
b11 %
1'
b11 +
#1070000000
1"
1(
#1080000000
0!
0"
b100 &
0'
0(
b100 ,
#1090000000
1!
b100 %
1'
b100 +
#1100000000
0!
0'
#1110000000
1!
b101 %
1'
b101 +
#1120000000
0!
0'
#1130000000
1!
b110 %
1'
b110 +
#1140000000
0!
0'
#1150000000
1!
b111 %
1'
b111 +
#1160000000
0!
0'
#1170000000
1!
0$
b1000 %
1'
0*
b1000 +
#1180000000
0!
0'
#1190000000
1!
b1001 %
1'
b1001 +
#1200000000
0!
0'
#1210000000
1!
b0 %
1'
b0 +
#1220000000
0!
0'
#1230000000
1!
1$
b1 %
1'
1*
b1 +
#1240000000
0!
0'
#1250000000
1!
b10 %
1'
b10 +
#1260000000
0!
0'
#1270000000
1!
b11 %
1'
b11 +
#1280000000
0!
0'
#1290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#1300000000
0!
0'
#1310000000
1!
b101 %
1'
b101 +
#1320000000
0!
0'
#1330000000
1!
0$
b110 %
1'
0*
b110 +
#1340000000
0!
0'
#1350000000
1!
b111 %
1'
b111 +
#1360000000
0!
0'
#1370000000
1!
b1000 %
1'
b1000 +
#1380000000
0!
0'
#1390000000
1!
b1001 %
1'
b1001 +
#1400000000
0!
0'
#1410000000
1!
b0 %
1'
b0 +
#1420000000
0!
0'
#1430000000
1!
1$
b1 %
1'
1*
b1 +
#1440000000
0!
0'
#1450000000
1!
b10 %
1'
b10 +
#1460000000
0!
0'
#1470000000
1!
b11 %
1'
b11 +
#1480000000
0!
0'
#1490000000
1!
b100 %
1'
b100 +
#1500000000
1"
1(
#1510000000
0!
0"
b100 &
0'
0(
b100 ,
#1520000000
1!
b101 %
1'
b101 +
#1530000000
0!
0'
#1540000000
1!
b110 %
1'
b110 +
#1550000000
0!
0'
#1560000000
1!
b111 %
1'
b111 +
#1570000000
0!
0'
#1580000000
1!
0$
b1000 %
1'
0*
b1000 +
#1590000000
0!
0'
#1600000000
1!
b1001 %
1'
b1001 +
#1610000000
0!
0'
#1620000000
1!
b0 %
1'
b0 +
#1630000000
0!
0'
#1640000000
1!
1$
b1 %
1'
1*
b1 +
#1650000000
0!
0'
#1660000000
1!
b10 %
1'
b10 +
#1670000000
0!
0'
#1680000000
1!
b11 %
1'
b11 +
#1690000000
0!
0'
#1700000000
1!
b100 %
1'
b100 +
#1710000000
0!
0'
#1720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#1730000000
0!
0'
#1740000000
1!
0$
b110 %
1'
0*
b110 +
#1750000000
0!
0'
#1760000000
1!
b111 %
1'
b111 +
#1770000000
0!
0'
#1780000000
1!
b1000 %
1'
b1000 +
#1790000000
0!
0'
#1800000000
1!
b1001 %
1'
b1001 +
#1810000000
0!
0'
#1820000000
1!
b0 %
1'
b0 +
#1830000000
0!
0'
#1840000000
1!
1$
b1 %
1'
1*
b1 +
#1850000000
0!
0'
#1860000000
1!
b10 %
1'
b10 +
#1870000000
0!
0'
#1880000000
1!
b11 %
1'
b11 +
#1890000000
0!
0'
#1900000000
1!
b100 %
1'
b100 +
#1910000000
0!
0'
#1920000000
1!
b101 %
1'
b101 +
#1930000000
1"
1(
#1940000000
0!
0"
b100 &
0'
0(
b100 ,
#1950000000
1!
b110 %
1'
b110 +
#1960000000
0!
0'
#1970000000
1!
b111 %
1'
b111 +
#1980000000
0!
0'
#1990000000
1!
0$
b1000 %
1'
0*
b1000 +
#2000000000
0!
0'
#2010000000
1!
b1001 %
1'
b1001 +
#2020000000
0!
0'
#2030000000
1!
b0 %
1'
b0 +
#2040000000
0!
0'
#2050000000
1!
1$
b1 %
1'
1*
b1 +
#2060000000
0!
0'
#2070000000
1!
b10 %
1'
b10 +
#2080000000
0!
0'
#2090000000
1!
b11 %
1'
b11 +
#2100000000
0!
0'
#2110000000
1!
b100 %
1'
b100 +
#2120000000
0!
0'
#2130000000
1!
b101 %
1'
b101 +
#2140000000
0!
0'
#2150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#2160000000
0!
0'
#2170000000
1!
b111 %
1'
b111 +
#2180000000
0!
0'
#2190000000
1!
b1000 %
1'
b1000 +
#2200000000
0!
0'
#2210000000
1!
b1001 %
1'
b1001 +
#2220000000
0!
0'
#2230000000
1!
b0 %
1'
b0 +
#2240000000
0!
0'
#2250000000
1!
1$
b1 %
1'
1*
b1 +
#2260000000
0!
0'
#2270000000
1!
b10 %
1'
b10 +
#2280000000
0!
0'
#2290000000
1!
b11 %
1'
b11 +
#2300000000
0!
0'
#2310000000
1!
b100 %
1'
b100 +
#2320000000
0!
0'
#2330000000
1!
b101 %
1'
b101 +
#2340000000
0!
0'
#2350000000
1!
0$
b110 %
1'
0*
b110 +
#2360000000
1"
1(
#2370000000
0!
0"
b100 &
0'
0(
b100 ,
#2380000000
1!
1$
b111 %
1'
1*
b111 +
#2390000000
0!
0'
#2400000000
1!
0$
b1000 %
1'
0*
b1000 +
#2410000000
0!
0'
#2420000000
1!
b1001 %
1'
b1001 +
#2430000000
0!
0'
#2440000000
1!
b0 %
1'
b0 +
#2450000000
0!
0'
#2460000000
1!
1$
b1 %
1'
1*
b1 +
#2470000000
0!
0'
#2480000000
1!
b10 %
1'
b10 +
#2490000000
0!
0'
#2500000000
1!
b11 %
1'
b11 +
#2510000000
0!
0'
#2520000000
1!
b100 %
1'
b100 +
#2530000000
0!
0'
#2540000000
1!
b101 %
1'
b101 +
#2550000000
0!
0'
#2560000000
1!
b110 %
1'
b110 +
#2570000000
0!
0'
#2580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#2590000000
0!
0'
#2600000000
1!
b1000 %
1'
b1000 +
#2610000000
0!
0'
#2620000000
1!
b1001 %
1'
b1001 +
#2630000000
0!
0'
#2640000000
1!
b0 %
1'
b0 +
#2650000000
0!
0'
#2660000000
1!
1$
b1 %
1'
1*
b1 +
#2670000000
0!
0'
#2680000000
1!
b10 %
1'
b10 +
#2690000000
0!
0'
#2700000000
1!
b11 %
1'
b11 +
#2710000000
0!
0'
#2720000000
1!
b100 %
1'
b100 +
#2730000000
0!
0'
#2740000000
1!
b101 %
1'
b101 +
#2750000000
0!
0'
#2760000000
1!
0$
b110 %
1'
0*
b110 +
#2770000000
0!
0'
#2780000000
1!
b111 %
1'
b111 +
#2790000000
1"
1(
#2800000000
0!
0"
b100 &
0'
0(
b100 ,
#2810000000
1!
b1000 %
1'
b1000 +
#2820000000
0!
0'
#2830000000
1!
b1001 %
1'
b1001 +
#2840000000
0!
0'
#2850000000
1!
b0 %
1'
b0 +
#2860000000
0!
0'
#2870000000
1!
1$
b1 %
1'
1*
b1 +
#2880000000
0!
0'
#2890000000
1!
b10 %
1'
b10 +
#2900000000
0!
0'
#2910000000
1!
b11 %
1'
b11 +
#2920000000
0!
0'
#2930000000
1!
b100 %
1'
b100 +
#2940000000
0!
0'
#2950000000
1!
b101 %
1'
b101 +
#2960000000
0!
0'
#2970000000
1!
b110 %
1'
b110 +
#2980000000
0!
0'
#2990000000
1!
b111 %
1'
b111 +
#3000000000
0!
0'
#3010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#3020000000
0!
0'
#3030000000
1!
b1001 %
1'
b1001 +
#3040000000
0!
0'
#3050000000
1!
b0 %
1'
b0 +
#3060000000
0!
0'
#3070000000
1!
1$
b1 %
1'
1*
b1 +
#3080000000
0!
0'
#3090000000
1!
b10 %
1'
b10 +
#3100000000
0!
0'
#3110000000
1!
b11 %
1'
b11 +
#3120000000
0!
0'
#3130000000
1!
b100 %
1'
b100 +
#3140000000
0!
0'
#3150000000
1!
b101 %
1'
b101 +
#3160000000
0!
0'
#3170000000
1!
0$
b110 %
1'
0*
b110 +
#3180000000
0!
0'
#3190000000
1!
b111 %
1'
b111 +
#3200000000
0!
0'
#3210000000
1!
b1000 %
1'
b1000 +
#3220000000
1"
1(
#3230000000
0!
0"
b100 &
0'
0(
b100 ,
#3240000000
1!
b1001 %
1'
b1001 +
#3250000000
0!
0'
#3260000000
1!
b0 %
1'
b0 +
#3270000000
0!
0'
#3280000000
1!
1$
b1 %
1'
1*
b1 +
#3290000000
0!
0'
#3300000000
1!
b10 %
1'
b10 +
#3310000000
0!
0'
#3320000000
1!
b11 %
1'
b11 +
#3330000000
0!
0'
#3340000000
1!
b100 %
1'
b100 +
#3350000000
0!
0'
#3360000000
1!
b101 %
1'
b101 +
#3370000000
0!
0'
#3380000000
1!
b110 %
1'
b110 +
#3390000000
0!
0'
#3400000000
1!
b111 %
1'
b111 +
#3410000000
0!
0'
#3420000000
1!
0$
b1000 %
1'
0*
b1000 +
#3430000000
0!
0'
#3440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#3450000000
0!
0'
#3460000000
1!
b0 %
1'
b0 +
#3470000000
0!
0'
#3480000000
1!
1$
b1 %
1'
1*
b1 +
#3490000000
0!
0'
#3500000000
1!
b10 %
1'
b10 +
#3510000000
0!
0'
#3520000000
1!
b11 %
1'
b11 +
#3530000000
0!
0'
#3540000000
1!
b100 %
1'
b100 +
#3550000000
0!
0'
#3560000000
1!
b101 %
1'
b101 +
#3570000000
0!
0'
#3580000000
1!
0$
b110 %
1'
0*
b110 +
#3590000000
0!
0'
#3600000000
1!
b111 %
1'
b111 +
#3610000000
0!
0'
#3620000000
1!
b1000 %
1'
b1000 +
#3630000000
0!
0'
#3640000000
1!
b1001 %
1'
b1001 +
#3650000000
1"
1(
#3660000000
0!
0"
b100 &
0'
0(
b100 ,
#3670000000
1!
b0 %
1'
b0 +
#3680000000
0!
0'
#3690000000
1!
1$
b1 %
1'
1*
b1 +
#3700000000
0!
0'
#3710000000
1!
b10 %
1'
b10 +
#3720000000
0!
0'
#3730000000
1!
b11 %
1'
b11 +
#3740000000
0!
0'
#3750000000
1!
b100 %
1'
b100 +
#3760000000
0!
0'
#3770000000
1!
b101 %
1'
b101 +
#3780000000
0!
0'
#3790000000
1!
b110 %
1'
b110 +
#3800000000
0!
0'
#3810000000
1!
b111 %
1'
b111 +
#3820000000
0!
0'
#3830000000
1!
0$
b1000 %
1'
0*
b1000 +
#3840000000
0!
0'
#3850000000
1!
b1001 %
1'
b1001 +
#3860000000
0!
0'
#3870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#3880000000
0!
0'
#3890000000
1!
1$
b1 %
1'
1*
b1 +
#3900000000
0!
0'
#3910000000
1!
b10 %
1'
b10 +
#3920000000
0!
0'
#3930000000
1!
b11 %
1'
b11 +
#3940000000
0!
0'
#3950000000
1!
b100 %
1'
b100 +
#3960000000
0!
0'
#3970000000
1!
b101 %
1'
b101 +
#3980000000
0!
0'
#3990000000
1!
0$
b110 %
1'
0*
b110 +
#4000000000
0!
0'
#4010000000
1!
b111 %
1'
b111 +
#4020000000
0!
0'
#4030000000
1!
b1000 %
1'
b1000 +
#4040000000
0!
0'
#4050000000
1!
b1001 %
1'
b1001 +
#4060000000
0!
0'
#4070000000
1!
b0 %
1'
b0 +
#4080000000
1"
1(
#4090000000
0!
0"
b100 &
0'
0(
b100 ,
#4100000000
1!
1$
b1 %
1'
1*
b1 +
#4110000000
0!
0'
#4120000000
1!
b10 %
1'
b10 +
#4130000000
0!
0'
#4140000000
1!
b11 %
1'
b11 +
#4150000000
0!
0'
#4160000000
1!
b100 %
1'
b100 +
#4170000000
0!
0'
#4180000000
1!
b101 %
1'
b101 +
#4190000000
0!
0'
#4200000000
1!
b110 %
1'
b110 +
#4210000000
0!
0'
#4220000000
1!
b111 %
1'
b111 +
#4230000000
0!
0'
#4240000000
1!
0$
b1000 %
1'
0*
b1000 +
#4250000000
0!
0'
#4260000000
1!
b1001 %
1'
b1001 +
#4270000000
0!
0'
#4280000000
1!
b0 %
1'
b0 +
#4290000000
0!
0'
#4300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#4310000000
0!
0'
#4320000000
1!
b10 %
1'
b10 +
#4330000000
0!
0'
#4340000000
1!
b11 %
1'
b11 +
#4350000000
0!
0'
#4360000000
1!
b100 %
1'
b100 +
#4370000000
0!
0'
#4380000000
1!
b101 %
1'
b101 +
#4390000000
0!
0'
#4400000000
1!
0$
b110 %
1'
0*
b110 +
#4410000000
0!
0'
#4420000000
1!
b111 %
1'
b111 +
#4430000000
0!
0'
#4440000000
1!
b1000 %
1'
b1000 +
#4450000000
0!
0'
#4460000000
1!
b1001 %
1'
b1001 +
#4470000000
0!
0'
#4480000000
1!
b0 %
1'
b0 +
#4490000000
0!
0'
#4500000000
1!
1$
b1 %
1'
1*
b1 +
#4510000000
1"
1(
#4520000000
0!
0"
b100 &
0'
0(
b100 ,
#4530000000
1!
b10 %
1'
b10 +
#4540000000
0!
0'
#4550000000
1!
b11 %
1'
b11 +
#4560000000
0!
0'
#4570000000
1!
b100 %
1'
b100 +
#4580000000
0!
0'
#4590000000
1!
b101 %
1'
b101 +
#4600000000
0!
0'
#4610000000
1!
b110 %
1'
b110 +
#4620000000
0!
0'
#4630000000
1!
b111 %
1'
b111 +
#4640000000
0!
0'
#4650000000
1!
0$
b1000 %
1'
0*
b1000 +
#4660000000
0!
0'
#4670000000
1!
b1001 %
1'
b1001 +
#4680000000
0!
0'
#4690000000
1!
b0 %
1'
b0 +
#4700000000
0!
0'
#4710000000
1!
1$
b1 %
1'
1*
b1 +
#4720000000
0!
0'
#4730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#4740000000
0!
0'
#4750000000
1!
b11 %
1'
b11 +
#4760000000
0!
0'
#4770000000
1!
b100 %
1'
b100 +
#4780000000
0!
0'
#4790000000
1!
b101 %
1'
b101 +
#4800000000
0!
0'
#4810000000
1!
0$
b110 %
1'
0*
b110 +
#4820000000
0!
0'
#4830000000
1!
b111 %
1'
b111 +
#4840000000
0!
0'
#4850000000
1!
b1000 %
1'
b1000 +
#4860000000
0!
0'
#4870000000
1!
b1001 %
1'
b1001 +
#4880000000
0!
0'
#4890000000
1!
b0 %
1'
b0 +
#4900000000
0!
0'
#4910000000
1!
1$
b1 %
1'
1*
b1 +
#4920000000
0!
0'
#4930000000
1!
b10 %
1'
b10 +
#4940000000
1"
1(
#4950000000
0!
0"
b100 &
0'
0(
b100 ,
#4960000000
1!
b11 %
1'
b11 +
#4970000000
0!
0'
#4980000000
1!
b100 %
1'
b100 +
#4990000000
0!
0'
#5000000000
1!
b101 %
1'
b101 +
#5010000000
0!
0'
#5020000000
1!
b110 %
1'
b110 +
#5030000000
0!
0'
#5040000000
1!
b111 %
1'
b111 +
#5050000000
0!
0'
#5060000000
1!
0$
b1000 %
1'
0*
b1000 +
#5070000000
0!
0'
#5080000000
1!
b1001 %
1'
b1001 +
#5090000000
0!
0'
#5100000000
1!
b0 %
1'
b0 +
#5110000000
0!
0'
#5120000000
1!
1$
b1 %
1'
1*
b1 +
#5130000000
0!
0'
#5140000000
1!
b10 %
1'
b10 +
#5150000000
0!
0'
#5160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#5170000000
0!
0'
#5180000000
1!
b100 %
1'
b100 +
#5190000000
0!
0'
#5200000000
1!
b101 %
1'
b101 +
#5210000000
0!
0'
#5220000000
1!
0$
b110 %
1'
0*
b110 +
#5230000000
0!
0'
#5240000000
1!
b111 %
1'
b111 +
#5250000000
0!
0'
#5260000000
1!
b1000 %
1'
b1000 +
#5270000000
0!
0'
#5280000000
1!
b1001 %
1'
b1001 +
#5290000000
0!
0'
#5300000000
1!
b0 %
1'
b0 +
#5310000000
0!
0'
#5320000000
1!
1$
b1 %
1'
1*
b1 +
#5330000000
0!
0'
#5340000000
1!
b10 %
1'
b10 +
#5350000000
0!
0'
#5360000000
1!
b11 %
1'
b11 +
#5370000000
1"
1(
#5380000000
0!
0"
b100 &
0'
0(
b100 ,
#5390000000
1!
b100 %
1'
b100 +
#5400000000
0!
0'
#5410000000
1!
b101 %
1'
b101 +
#5420000000
0!
0'
#5430000000
1!
b110 %
1'
b110 +
#5440000000
0!
0'
#5450000000
1!
b111 %
1'
b111 +
#5460000000
0!
0'
#5470000000
1!
0$
b1000 %
1'
0*
b1000 +
#5480000000
0!
0'
#5490000000
1!
b1001 %
1'
b1001 +
#5500000000
0!
0'
#5510000000
1!
b0 %
1'
b0 +
#5520000000
0!
0'
#5530000000
1!
1$
b1 %
1'
1*
b1 +
#5540000000
0!
0'
#5550000000
1!
b10 %
1'
b10 +
#5560000000
0!
0'
#5570000000
1!
b11 %
1'
b11 +
#5580000000
0!
0'
#5590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#5600000000
0!
0'
#5610000000
1!
b101 %
1'
b101 +
#5620000000
0!
0'
#5630000000
1!
0$
b110 %
1'
0*
b110 +
#5640000000
0!
0'
#5650000000
1!
b111 %
1'
b111 +
#5660000000
0!
0'
#5670000000
1!
b1000 %
1'
b1000 +
#5680000000
0!
0'
#5690000000
1!
b1001 %
1'
b1001 +
#5700000000
0!
0'
#5710000000
1!
b0 %
1'
b0 +
#5720000000
0!
0'
#5730000000
1!
1$
b1 %
1'
1*
b1 +
#5740000000
0!
0'
#5750000000
1!
b10 %
1'
b10 +
#5760000000
0!
0'
#5770000000
1!
b11 %
1'
b11 +
#5780000000
0!
0'
#5790000000
1!
b100 %
1'
b100 +
#5800000000
1"
1(
#5810000000
0!
0"
b100 &
0'
0(
b100 ,
#5820000000
1!
b101 %
1'
b101 +
#5830000000
0!
0'
#5840000000
1!
b110 %
1'
b110 +
#5850000000
0!
0'
#5860000000
1!
b111 %
1'
b111 +
#5870000000
0!
0'
#5880000000
1!
0$
b1000 %
1'
0*
b1000 +
#5890000000
0!
0'
#5900000000
1!
b1001 %
1'
b1001 +
#5910000000
0!
0'
#5920000000
1!
b0 %
1'
b0 +
#5930000000
0!
0'
#5940000000
1!
1$
b1 %
1'
1*
b1 +
#5950000000
0!
0'
#5960000000
1!
b10 %
1'
b10 +
#5970000000
0!
0'
#5980000000
1!
b11 %
1'
b11 +
#5990000000
0!
0'
#6000000000
1!
b100 %
1'
b100 +
#6010000000
0!
0'
#6020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#6030000000
0!
0'
#6040000000
1!
0$
b110 %
1'
0*
b110 +
#6050000000
0!
0'
#6060000000
1!
b111 %
1'
b111 +
#6070000000
0!
0'
#6080000000
1!
b1000 %
1'
b1000 +
#6090000000
0!
0'
#6100000000
1!
b1001 %
1'
b1001 +
#6110000000
0!
0'
#6120000000
1!
b0 %
1'
b0 +
#6130000000
0!
0'
#6140000000
1!
1$
b1 %
1'
1*
b1 +
#6150000000
0!
0'
#6160000000
1!
b10 %
1'
b10 +
#6170000000
0!
0'
#6180000000
1!
b11 %
1'
b11 +
#6190000000
0!
0'
#6200000000
1!
b100 %
1'
b100 +
#6210000000
0!
0'
#6220000000
1!
b101 %
1'
b101 +
#6230000000
1"
1(
#6240000000
0!
0"
b100 &
0'
0(
b100 ,
#6250000000
1!
b110 %
1'
b110 +
#6260000000
0!
0'
#6270000000
1!
b111 %
1'
b111 +
#6280000000
0!
0'
#6290000000
1!
0$
b1000 %
1'
0*
b1000 +
#6300000000
0!
0'
#6310000000
1!
b1001 %
1'
b1001 +
#6320000000
0!
0'
#6330000000
1!
b0 %
1'
b0 +
#6340000000
0!
0'
#6350000000
1!
1$
b1 %
1'
1*
b1 +
#6360000000
0!
0'
#6370000000
1!
b10 %
1'
b10 +
#6380000000
0!
0'
#6390000000
1!
b11 %
1'
b11 +
#6400000000
0!
0'
#6410000000
1!
b100 %
1'
b100 +
#6420000000
0!
0'
#6430000000
1!
b101 %
1'
b101 +
#6440000000
0!
0'
#6450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#6460000000
0!
0'
#6470000000
1!
b111 %
1'
b111 +
#6480000000
0!
0'
#6490000000
1!
b1000 %
1'
b1000 +
#6500000000
0!
0'
#6510000000
1!
b1001 %
1'
b1001 +
#6520000000
0!
0'
#6530000000
1!
b0 %
1'
b0 +
#6540000000
0!
0'
#6550000000
1!
1$
b1 %
1'
1*
b1 +
#6560000000
0!
0'
#6570000000
1!
b10 %
1'
b10 +
#6580000000
0!
0'
#6590000000
1!
b11 %
1'
b11 +
#6600000000
0!
0'
#6610000000
1!
b100 %
1'
b100 +
#6620000000
0!
0'
#6630000000
1!
b101 %
1'
b101 +
#6640000000
0!
0'
#6650000000
1!
0$
b110 %
1'
0*
b110 +
#6660000000
1"
1(
#6670000000
0!
0"
b100 &
0'
0(
b100 ,
#6680000000
1!
1$
b111 %
1'
1*
b111 +
#6690000000
0!
0'
#6700000000
1!
0$
b1000 %
1'
0*
b1000 +
#6710000000
0!
0'
#6720000000
1!
b1001 %
1'
b1001 +
#6730000000
0!
0'
#6740000000
1!
b0 %
1'
b0 +
#6750000000
0!
0'
#6760000000
1!
1$
b1 %
1'
1*
b1 +
#6770000000
0!
0'
#6780000000
1!
b10 %
1'
b10 +
#6790000000
0!
0'
#6800000000
1!
b11 %
1'
b11 +
#6810000000
0!
0'
#6820000000
1!
b100 %
1'
b100 +
#6830000000
0!
0'
#6840000000
1!
b101 %
1'
b101 +
#6850000000
0!
0'
#6860000000
1!
b110 %
1'
b110 +
#6870000000
0!
0'
#6880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#6890000000
0!
0'
#6900000000
1!
b1000 %
1'
b1000 +
#6910000000
0!
0'
#6920000000
1!
b1001 %
1'
b1001 +
#6930000000
0!
0'
#6940000000
1!
b0 %
1'
b0 +
#6950000000
0!
0'
#6960000000
1!
1$
b1 %
1'
1*
b1 +
#6970000000
0!
0'
#6980000000
1!
b10 %
1'
b10 +
#6990000000
0!
0'
#7000000000
1!
b11 %
1'
b11 +
#7010000000
0!
0'
#7020000000
1!
b100 %
1'
b100 +
#7030000000
0!
0'
#7040000000
1!
b101 %
1'
b101 +
#7050000000
0!
0'
#7060000000
1!
0$
b110 %
1'
0*
b110 +
#7070000000
0!
0'
#7080000000
1!
b111 %
1'
b111 +
#7090000000
1"
1(
#7100000000
0!
0"
b100 &
0'
0(
b100 ,
#7110000000
1!
b1000 %
1'
b1000 +
#7120000000
0!
0'
#7130000000
1!
b1001 %
1'
b1001 +
#7140000000
0!
0'
#7150000000
1!
b0 %
1'
b0 +
#7160000000
0!
0'
#7170000000
1!
1$
b1 %
1'
1*
b1 +
#7180000000
0!
0'
#7190000000
1!
b10 %
1'
b10 +
#7200000000
0!
0'
#7210000000
1!
b11 %
1'
b11 +
#7220000000
0!
0'
#7230000000
1!
b100 %
1'
b100 +
#7240000000
0!
0'
#7250000000
1!
b101 %
1'
b101 +
#7260000000
0!
0'
#7270000000
1!
b110 %
1'
b110 +
#7280000000
0!
0'
#7290000000
1!
b111 %
1'
b111 +
#7300000000
0!
0'
#7310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#7320000000
0!
0'
#7330000000
1!
b1001 %
1'
b1001 +
#7340000000
0!
0'
#7350000000
1!
b0 %
1'
b0 +
#7360000000
0!
0'
#7370000000
1!
1$
b1 %
1'
1*
b1 +
#7380000000
0!
0'
#7390000000
1!
b10 %
1'
b10 +
#7400000000
0!
0'
#7410000000
1!
b11 %
1'
b11 +
#7420000000
0!
0'
#7430000000
1!
b100 %
1'
b100 +
#7440000000
0!
0'
#7450000000
1!
b101 %
1'
b101 +
#7460000000
0!
0'
#7470000000
1!
0$
b110 %
1'
0*
b110 +
#7480000000
0!
0'
#7490000000
1!
b111 %
1'
b111 +
#7500000000
0!
0'
#7510000000
1!
b1000 %
1'
b1000 +
#7520000000
1"
1(
#7530000000
0!
0"
b100 &
0'
0(
b100 ,
#7540000000
1!
b1001 %
1'
b1001 +
#7550000000
0!
0'
#7560000000
1!
b0 %
1'
b0 +
#7570000000
0!
0'
#7580000000
1!
1$
b1 %
1'
1*
b1 +
#7590000000
0!
0'
#7600000000
1!
b10 %
1'
b10 +
#7610000000
0!
0'
#7620000000
1!
b11 %
1'
b11 +
#7630000000
0!
0'
#7640000000
1!
b100 %
1'
b100 +
#7650000000
0!
0'
#7660000000
1!
b101 %
1'
b101 +
#7670000000
0!
0'
#7680000000
1!
b110 %
1'
b110 +
#7690000000
0!
0'
#7700000000
1!
b111 %
1'
b111 +
#7710000000
0!
0'
#7720000000
1!
0$
b1000 %
1'
0*
b1000 +
#7730000000
0!
0'
#7740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#7750000000
0!
0'
#7760000000
1!
b0 %
1'
b0 +
#7770000000
0!
0'
#7780000000
1!
1$
b1 %
1'
1*
b1 +
#7790000000
0!
0'
#7800000000
1!
b10 %
1'
b10 +
#7810000000
0!
0'
#7820000000
1!
b11 %
1'
b11 +
#7830000000
0!
0'
#7840000000
1!
b100 %
1'
b100 +
#7850000000
0!
0'
#7860000000
1!
b101 %
1'
b101 +
#7870000000
0!
0'
#7880000000
1!
0$
b110 %
1'
0*
b110 +
#7890000000
0!
0'
#7900000000
1!
b111 %
1'
b111 +
#7910000000
0!
0'
#7920000000
1!
b1000 %
1'
b1000 +
#7930000000
0!
0'
#7940000000
1!
b1001 %
1'
b1001 +
#7950000000
1"
1(
#7960000000
0!
0"
b100 &
0'
0(
b100 ,
#7970000000
1!
b0 %
1'
b0 +
#7980000000
0!
0'
#7990000000
1!
1$
b1 %
1'
1*
b1 +
#8000000000
0!
0'
#8010000000
1!
b10 %
1'
b10 +
#8020000000
0!
0'
#8030000000
1!
b11 %
1'
b11 +
#8040000000
0!
0'
#8050000000
1!
b100 %
1'
b100 +
#8060000000
0!
0'
#8070000000
1!
b101 %
1'
b101 +
#8080000000
0!
0'
#8090000000
1!
b110 %
1'
b110 +
#8100000000
0!
0'
#8110000000
1!
b111 %
1'
b111 +
#8120000000
0!
0'
#8130000000
1!
0$
b1000 %
1'
0*
b1000 +
#8140000000
0!
0'
#8150000000
1!
b1001 %
1'
b1001 +
#8160000000
0!
0'
#8170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#8180000000
0!
0'
#8190000000
1!
1$
b1 %
1'
1*
b1 +
#8200000000
0!
0'
#8210000000
1!
b10 %
1'
b10 +
#8220000000
0!
0'
#8230000000
1!
b11 %
1'
b11 +
#8240000000
0!
0'
#8250000000
1!
b100 %
1'
b100 +
#8260000000
0!
0'
#8270000000
1!
b101 %
1'
b101 +
#8280000000
0!
0'
#8290000000
1!
0$
b110 %
1'
0*
b110 +
#8300000000
0!
0'
#8310000000
1!
b111 %
1'
b111 +
#8320000000
0!
0'
#8330000000
1!
b1000 %
1'
b1000 +
#8340000000
0!
0'
#8350000000
1!
b1001 %
1'
b1001 +
#8360000000
0!
0'
#8370000000
1!
b0 %
1'
b0 +
#8380000000
1"
1(
#8390000000
0!
0"
b100 &
0'
0(
b100 ,
#8400000000
1!
1$
b1 %
1'
1*
b1 +
#8410000000
0!
0'
#8420000000
1!
b10 %
1'
b10 +
#8430000000
0!
0'
#8440000000
1!
b11 %
1'
b11 +
#8450000000
0!
0'
#8460000000
1!
b100 %
1'
b100 +
#8470000000
0!
0'
#8480000000
1!
b101 %
1'
b101 +
#8490000000
0!
0'
#8500000000
1!
b110 %
1'
b110 +
#8510000000
0!
0'
#8520000000
1!
b111 %
1'
b111 +
#8530000000
0!
0'
#8540000000
1!
0$
b1000 %
1'
0*
b1000 +
#8550000000
0!
0'
#8560000000
1!
b1001 %
1'
b1001 +
#8570000000
0!
0'
#8580000000
1!
b0 %
1'
b0 +
#8590000000
0!
0'
#8600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#8610000000
0!
0'
#8620000000
1!
b10 %
1'
b10 +
#8630000000
0!
0'
#8640000000
1!
b11 %
1'
b11 +
#8650000000
0!
0'
#8660000000
1!
b100 %
1'
b100 +
#8670000000
0!
0'
#8680000000
1!
b101 %
1'
b101 +
#8690000000
0!
0'
#8700000000
1!
0$
b110 %
1'
0*
b110 +
#8710000000
0!
0'
#8720000000
1!
b111 %
1'
b111 +
#8730000000
0!
0'
#8740000000
1!
b1000 %
1'
b1000 +
#8750000000
0!
0'
#8760000000
1!
b1001 %
1'
b1001 +
#8770000000
0!
0'
#8780000000
1!
b0 %
1'
b0 +
#8790000000
0!
0'
#8800000000
1!
1$
b1 %
1'
1*
b1 +
#8810000000
1"
1(
#8820000000
0!
0"
b100 &
0'
0(
b100 ,
#8830000000
1!
b10 %
1'
b10 +
#8840000000
0!
0'
#8850000000
1!
b11 %
1'
b11 +
#8860000000
0!
0'
#8870000000
1!
b100 %
1'
b100 +
#8880000000
0!
0'
#8890000000
1!
b101 %
1'
b101 +
#8900000000
0!
0'
#8910000000
1!
b110 %
1'
b110 +
#8920000000
0!
0'
#8930000000
1!
b111 %
1'
b111 +
#8940000000
0!
0'
#8950000000
1!
0$
b1000 %
1'
0*
b1000 +
#8960000000
0!
0'
#8970000000
1!
b1001 %
1'
b1001 +
#8980000000
0!
0'
#8990000000
1!
b0 %
1'
b0 +
#9000000000
0!
0'
#9010000000
1!
1$
b1 %
1'
1*
b1 +
#9020000000
0!
0'
#9030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#9040000000
0!
0'
#9050000000
1!
b11 %
1'
b11 +
#9060000000
0!
0'
#9070000000
1!
b100 %
1'
b100 +
#9080000000
0!
0'
#9090000000
1!
b101 %
1'
b101 +
#9100000000
0!
0'
#9110000000
1!
0$
b110 %
1'
0*
b110 +
#9120000000
0!
0'
#9130000000
1!
b111 %
1'
b111 +
#9140000000
0!
0'
#9150000000
1!
b1000 %
1'
b1000 +
#9160000000
0!
0'
#9170000000
1!
b1001 %
1'
b1001 +
#9180000000
0!
0'
#9190000000
1!
b0 %
1'
b0 +
#9200000000
0!
0'
#9210000000
1!
1$
b1 %
1'
1*
b1 +
#9220000000
0!
0'
#9230000000
1!
b10 %
1'
b10 +
#9240000000
1"
1(
#9250000000
0!
0"
b100 &
0'
0(
b100 ,
#9260000000
1!
b11 %
1'
b11 +
#9270000000
0!
0'
#9280000000
1!
b100 %
1'
b100 +
#9290000000
0!
0'
#9300000000
1!
b101 %
1'
b101 +
#9310000000
0!
0'
#9320000000
1!
b110 %
1'
b110 +
#9330000000
0!
0'
#9340000000
1!
b111 %
1'
b111 +
#9350000000
0!
0'
#9360000000
1!
0$
b1000 %
1'
0*
b1000 +
#9370000000
0!
0'
#9380000000
1!
b1001 %
1'
b1001 +
#9390000000
0!
0'
#9400000000
1!
b0 %
1'
b0 +
#9410000000
0!
0'
#9420000000
1!
1$
b1 %
1'
1*
b1 +
#9430000000
0!
0'
#9440000000
1!
b10 %
1'
b10 +
#9450000000
0!
0'
#9460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#9470000000
0!
0'
#9480000000
1!
b100 %
1'
b100 +
#9490000000
0!
0'
#9500000000
1!
b101 %
1'
b101 +
#9510000000
0!
0'
#9520000000
1!
0$
b110 %
1'
0*
b110 +
#9530000000
0!
0'
#9540000000
1!
b111 %
1'
b111 +
#9550000000
0!
0'
#9560000000
1!
b1000 %
1'
b1000 +
#9570000000
0!
0'
#9580000000
1!
b1001 %
1'
b1001 +
#9590000000
0!
0'
#9600000000
1!
b0 %
1'
b0 +
#9610000000
0!
0'
#9620000000
1!
1$
b1 %
1'
1*
b1 +
#9630000000
0!
0'
#9640000000
1!
b10 %
1'
b10 +
#9650000000
0!
0'
#9660000000
1!
b11 %
1'
b11 +
#9670000000
1"
1(
#9680000000
0!
0"
b100 &
0'
0(
b100 ,
#9690000000
1!
b100 %
1'
b100 +
#9700000000
0!
0'
#9710000000
1!
b101 %
1'
b101 +
#9720000000
0!
0'
#9730000000
1!
b110 %
1'
b110 +
#9740000000
0!
0'
#9750000000
1!
b111 %
1'
b111 +
#9760000000
0!
0'
#9770000000
1!
0$
b1000 %
1'
0*
b1000 +
#9780000000
0!
0'
#9790000000
1!
b1001 %
1'
b1001 +
#9800000000
0!
0'
#9810000000
1!
b0 %
1'
b0 +
#9820000000
0!
0'
#9830000000
1!
1$
b1 %
1'
1*
b1 +
#9840000000
0!
0'
#9850000000
1!
b10 %
1'
b10 +
#9860000000
0!
0'
#9870000000
1!
b11 %
1'
b11 +
#9880000000
0!
0'
#9890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#9900000000
0!
0'
#9910000000
1!
b101 %
1'
b101 +
#9920000000
0!
0'
#9930000000
1!
0$
b110 %
1'
0*
b110 +
#9940000000
0!
0'
#9950000000
1!
b111 %
1'
b111 +
#9960000000
0!
0'
#9970000000
1!
b1000 %
1'
b1000 +
#9980000000
0!
0'
#9990000000
1!
b1001 %
1'
b1001 +
#10000000000
0!
0'
#10010000000
1!
b0 %
1'
b0 +
#10020000000
0!
0'
#10030000000
1!
1$
b1 %
1'
1*
b1 +
#10040000000
0!
0'
#10050000000
1!
b10 %
1'
b10 +
#10060000000
0!
0'
#10070000000
1!
b11 %
1'
b11 +
#10080000000
0!
0'
#10090000000
1!
b100 %
1'
b100 +
#10100000000
1"
1(
#10110000000
0!
0"
b100 &
0'
0(
b100 ,
#10120000000
1!
b101 %
1'
b101 +
#10130000000
0!
0'
#10140000000
1!
b110 %
1'
b110 +
#10150000000
0!
0'
#10160000000
1!
b111 %
1'
b111 +
#10170000000
0!
0'
#10180000000
1!
0$
b1000 %
1'
0*
b1000 +
#10190000000
0!
0'
#10200000000
1!
b1001 %
1'
b1001 +
#10210000000
0!
0'
#10220000000
1!
b0 %
1'
b0 +
#10230000000
0!
0'
#10240000000
1!
1$
b1 %
1'
1*
b1 +
#10250000000
0!
0'
#10260000000
1!
b10 %
1'
b10 +
#10270000000
0!
0'
#10280000000
1!
b11 %
1'
b11 +
#10290000000
0!
0'
#10300000000
1!
b100 %
1'
b100 +
#10310000000
0!
0'
#10320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#10330000000
0!
0'
#10340000000
1!
0$
b110 %
1'
0*
b110 +
#10350000000
0!
0'
#10360000000
1!
b111 %
1'
b111 +
#10370000000
0!
0'
#10380000000
1!
b1000 %
1'
b1000 +
#10390000000
0!
0'
#10400000000
1!
b1001 %
1'
b1001 +
#10410000000
0!
0'
#10420000000
1!
b0 %
1'
b0 +
#10430000000
0!
0'
#10440000000
1!
1$
b1 %
1'
1*
b1 +
#10450000000
0!
0'
#10460000000
1!
b10 %
1'
b10 +
#10470000000
0!
0'
#10480000000
1!
b11 %
1'
b11 +
#10490000000
0!
0'
#10500000000
1!
b100 %
1'
b100 +
#10510000000
0!
0'
#10520000000
1!
b101 %
1'
b101 +
#10530000000
1"
1(
#10540000000
0!
0"
b100 &
0'
0(
b100 ,
#10550000000
1!
b110 %
1'
b110 +
#10560000000
0!
0'
#10570000000
1!
b111 %
1'
b111 +
#10580000000
0!
0'
#10590000000
1!
0$
b1000 %
1'
0*
b1000 +
#10600000000
0!
0'
#10610000000
1!
b1001 %
1'
b1001 +
#10620000000
0!
0'
#10630000000
1!
b0 %
1'
b0 +
#10640000000
0!
0'
#10650000000
1!
1$
b1 %
1'
1*
b1 +
#10660000000
0!
0'
#10670000000
1!
b10 %
1'
b10 +
#10680000000
0!
0'
#10690000000
1!
b11 %
1'
b11 +
#10700000000
0!
0'
#10710000000
1!
b100 %
1'
b100 +
#10720000000
0!
0'
#10730000000
1!
b101 %
1'
b101 +
#10740000000
0!
0'
#10750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#10760000000
0!
0'
#10770000000
1!
b111 %
1'
b111 +
#10780000000
0!
0'
#10790000000
1!
b1000 %
1'
b1000 +
#10800000000
0!
0'
#10810000000
1!
b1001 %
1'
b1001 +
#10820000000
0!
0'
#10830000000
1!
b0 %
1'
b0 +
#10840000000
0!
0'
#10850000000
1!
1$
b1 %
1'
1*
b1 +
#10860000000
0!
0'
#10870000000
1!
b10 %
1'
b10 +
#10880000000
0!
0'
#10890000000
1!
b11 %
1'
b11 +
#10900000000
0!
0'
#10910000000
1!
b100 %
1'
b100 +
#10920000000
0!
0'
#10930000000
1!
b101 %
1'
b101 +
#10940000000
0!
0'
#10950000000
1!
0$
b110 %
1'
0*
b110 +
#10960000000
1"
1(
#10970000000
0!
0"
b100 &
0'
0(
b100 ,
#10980000000
1!
1$
b111 %
1'
1*
b111 +
#10990000000
0!
0'
#11000000000
1!
0$
b1000 %
1'
0*
b1000 +
#11010000000
0!
0'
#11020000000
1!
b1001 %
1'
b1001 +
#11030000000
0!
0'
#11040000000
1!
b0 %
1'
b0 +
#11050000000
0!
0'
#11060000000
1!
1$
b1 %
1'
1*
b1 +
#11070000000
0!
0'
#11080000000
1!
b10 %
1'
b10 +
#11090000000
0!
0'
#11100000000
1!
b11 %
1'
b11 +
#11110000000
0!
0'
#11120000000
1!
b100 %
1'
b100 +
#11130000000
0!
0'
#11140000000
1!
b101 %
1'
b101 +
#11150000000
0!
0'
#11160000000
1!
b110 %
1'
b110 +
#11170000000
0!
0'
#11180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#11190000000
0!
0'
#11200000000
1!
b1000 %
1'
b1000 +
#11210000000
0!
0'
#11220000000
1!
b1001 %
1'
b1001 +
#11230000000
0!
0'
#11240000000
1!
b0 %
1'
b0 +
#11250000000
0!
0'
#11260000000
1!
1$
b1 %
1'
1*
b1 +
#11270000000
0!
0'
#11280000000
1!
b10 %
1'
b10 +
#11290000000
0!
0'
#11300000000
1!
b11 %
1'
b11 +
#11310000000
0!
0'
#11320000000
1!
b100 %
1'
b100 +
#11330000000
0!
0'
#11340000000
1!
b101 %
1'
b101 +
#11350000000
0!
0'
#11360000000
1!
0$
b110 %
1'
0*
b110 +
#11370000000
0!
0'
#11380000000
1!
b111 %
1'
b111 +
#11390000000
1"
1(
#11400000000
0!
0"
b100 &
0'
0(
b100 ,
#11410000000
1!
b1000 %
1'
b1000 +
#11420000000
0!
0'
#11430000000
1!
b1001 %
1'
b1001 +
#11440000000
0!
0'
#11450000000
1!
b0 %
1'
b0 +
#11460000000
0!
0'
#11470000000
1!
1$
b1 %
1'
1*
b1 +
#11480000000
0!
0'
#11490000000
1!
b10 %
1'
b10 +
#11500000000
0!
0'
#11510000000
1!
b11 %
1'
b11 +
#11520000000
0!
0'
#11530000000
1!
b100 %
1'
b100 +
#11540000000
0!
0'
#11550000000
1!
b101 %
1'
b101 +
#11560000000
0!
0'
#11570000000
1!
b110 %
1'
b110 +
#11580000000
0!
0'
#11590000000
1!
b111 %
1'
b111 +
#11600000000
0!
0'
#11610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#11620000000
0!
0'
#11630000000
1!
b1001 %
1'
b1001 +
#11640000000
0!
0'
#11650000000
1!
b0 %
1'
b0 +
#11660000000
0!
0'
#11670000000
1!
1$
b1 %
1'
1*
b1 +
#11680000000
0!
0'
#11690000000
1!
b10 %
1'
b10 +
#11700000000
0!
0'
#11710000000
1!
b11 %
1'
b11 +
#11720000000
0!
0'
#11730000000
1!
b100 %
1'
b100 +
#11740000000
0!
0'
#11750000000
1!
b101 %
1'
b101 +
#11760000000
0!
0'
#11770000000
1!
0$
b110 %
1'
0*
b110 +
#11780000000
0!
0'
#11790000000
1!
b111 %
1'
b111 +
#11800000000
0!
0'
#11810000000
1!
b1000 %
1'
b1000 +
#11820000000
1"
1(
#11830000000
0!
0"
b100 &
0'
0(
b100 ,
#11840000000
1!
b1001 %
1'
b1001 +
#11850000000
0!
0'
#11860000000
1!
b0 %
1'
b0 +
#11870000000
0!
0'
#11880000000
1!
1$
b1 %
1'
1*
b1 +
#11890000000
0!
0'
#11900000000
1!
b10 %
1'
b10 +
#11910000000
0!
0'
#11920000000
1!
b11 %
1'
b11 +
#11930000000
0!
0'
#11940000000
1!
b100 %
1'
b100 +
#11950000000
0!
0'
#11960000000
1!
b101 %
1'
b101 +
#11970000000
0!
0'
#11980000000
1!
b110 %
1'
b110 +
#11990000000
0!
0'
#12000000000
1!
b111 %
1'
b111 +
#12010000000
0!
0'
#12020000000
1!
0$
b1000 %
1'
0*
b1000 +
#12030000000
0!
0'
#12040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#12050000000
0!
0'
#12060000000
1!
b0 %
1'
b0 +
#12070000000
0!
0'
#12080000000
1!
1$
b1 %
1'
1*
b1 +
#12090000000
0!
0'
#12100000000
1!
b10 %
1'
b10 +
#12110000000
0!
0'
#12120000000
1!
b11 %
1'
b11 +
#12130000000
0!
0'
#12140000000
1!
b100 %
1'
b100 +
#12150000000
0!
0'
#12160000000
1!
b101 %
1'
b101 +
#12170000000
0!
0'
#12180000000
1!
0$
b110 %
1'
0*
b110 +
#12190000000
0!
0'
#12200000000
1!
b111 %
1'
b111 +
#12210000000
0!
0'
#12220000000
1!
b1000 %
1'
b1000 +
#12230000000
0!
0'
#12240000000
1!
b1001 %
1'
b1001 +
#12250000000
1"
1(
#12260000000
0!
0"
b100 &
0'
0(
b100 ,
#12270000000
1!
b0 %
1'
b0 +
#12280000000
0!
0'
#12290000000
1!
1$
b1 %
1'
1*
b1 +
#12300000000
0!
0'
#12310000000
1!
b10 %
1'
b10 +
#12320000000
0!
0'
#12330000000
1!
b11 %
1'
b11 +
#12340000000
0!
0'
#12350000000
1!
b100 %
1'
b100 +
#12360000000
0!
0'
#12370000000
1!
b101 %
1'
b101 +
#12380000000
0!
0'
#12390000000
1!
b110 %
1'
b110 +
#12400000000
0!
0'
#12410000000
1!
b111 %
1'
b111 +
#12420000000
0!
0'
#12430000000
1!
0$
b1000 %
1'
0*
b1000 +
#12440000000
0!
0'
#12450000000
1!
b1001 %
1'
b1001 +
#12460000000
0!
0'
#12470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#12480000000
0!
0'
#12490000000
1!
1$
b1 %
1'
1*
b1 +
#12500000000
0!
0'
#12510000000
1!
b10 %
1'
b10 +
#12520000000
0!
0'
#12530000000
1!
b11 %
1'
b11 +
#12540000000
0!
0'
#12550000000
1!
b100 %
1'
b100 +
#12560000000
0!
0'
#12570000000
1!
b101 %
1'
b101 +
#12580000000
0!
0'
#12590000000
1!
0$
b110 %
1'
0*
b110 +
#12600000000
0!
0'
#12610000000
1!
b111 %
1'
b111 +
#12620000000
0!
0'
#12630000000
1!
b1000 %
1'
b1000 +
#12640000000
0!
0'
#12650000000
1!
b1001 %
1'
b1001 +
#12660000000
0!
0'
#12670000000
1!
b0 %
1'
b0 +
#12680000000
1"
1(
#12690000000
0!
0"
b100 &
0'
0(
b100 ,
#12700000000
1!
1$
b1 %
1'
1*
b1 +
#12710000000
0!
0'
#12720000000
1!
b10 %
1'
b10 +
#12730000000
0!
0'
#12740000000
1!
b11 %
1'
b11 +
#12750000000
0!
0'
#12760000000
1!
b100 %
1'
b100 +
#12770000000
0!
0'
#12780000000
1!
b101 %
1'
b101 +
#12790000000
0!
0'
#12800000000
1!
b110 %
1'
b110 +
#12810000000
0!
0'
#12820000000
1!
b111 %
1'
b111 +
#12830000000
0!
0'
#12840000000
1!
0$
b1000 %
1'
0*
b1000 +
#12850000000
0!
0'
#12860000000
1!
b1001 %
1'
b1001 +
#12870000000
0!
0'
#12880000000
1!
b0 %
1'
b0 +
#12890000000
0!
0'
#12900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#12910000000
0!
0'
#12920000000
1!
b10 %
1'
b10 +
#12930000000
0!
0'
#12940000000
1!
b11 %
1'
b11 +
#12950000000
0!
0'
#12960000000
1!
b100 %
1'
b100 +
#12970000000
0!
0'
#12980000000
1!
b101 %
1'
b101 +
#12990000000
0!
0'
#13000000000
1!
0$
b110 %
1'
0*
b110 +
#13010000000
0!
0'
#13020000000
1!
b111 %
1'
b111 +
#13030000000
0!
0'
#13040000000
1!
b1000 %
1'
b1000 +
#13050000000
0!
0'
#13060000000
1!
b1001 %
1'
b1001 +
#13070000000
0!
0'
#13080000000
1!
b0 %
1'
b0 +
#13090000000
0!
0'
#13100000000
1!
1$
b1 %
1'
1*
b1 +
#13110000000
1"
1(
#13120000000
0!
0"
b100 &
0'
0(
b100 ,
#13130000000
1!
b10 %
1'
b10 +
#13140000000
0!
0'
#13150000000
1!
b11 %
1'
b11 +
#13160000000
0!
0'
#13170000000
1!
b100 %
1'
b100 +
#13180000000
0!
0'
#13190000000
1!
b101 %
1'
b101 +
#13200000000
0!
0'
#13210000000
1!
b110 %
1'
b110 +
#13220000000
0!
0'
#13230000000
1!
b111 %
1'
b111 +
#13240000000
0!
0'
#13250000000
1!
0$
b1000 %
1'
0*
b1000 +
#13260000000
0!
0'
#13270000000
1!
b1001 %
1'
b1001 +
#13280000000
0!
0'
#13290000000
1!
b0 %
1'
b0 +
#13300000000
0!
0'
#13310000000
1!
1$
b1 %
1'
1*
b1 +
#13320000000
0!
0'
#13330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#13340000000
0!
0'
#13350000000
1!
b11 %
1'
b11 +
#13360000000
0!
0'
#13370000000
1!
b100 %
1'
b100 +
#13380000000
0!
0'
#13390000000
1!
b101 %
1'
b101 +
#13400000000
0!
0'
#13410000000
1!
0$
b110 %
1'
0*
b110 +
#13420000000
0!
0'
#13430000000
1!
b111 %
1'
b111 +
#13440000000
0!
0'
#13450000000
1!
b1000 %
1'
b1000 +
#13460000000
0!
0'
#13470000000
1!
b1001 %
1'
b1001 +
#13480000000
0!
0'
#13490000000
1!
b0 %
1'
b0 +
#13500000000
0!
0'
#13510000000
1!
1$
b1 %
1'
1*
b1 +
#13520000000
0!
0'
#13530000000
1!
b10 %
1'
b10 +
#13540000000
1"
1(
#13550000000
0!
0"
b100 &
0'
0(
b100 ,
#13560000000
1!
b11 %
1'
b11 +
#13570000000
0!
0'
#13580000000
1!
b100 %
1'
b100 +
#13590000000
0!
0'
#13600000000
1!
b101 %
1'
b101 +
#13610000000
0!
0'
#13620000000
1!
b110 %
1'
b110 +
#13630000000
0!
0'
#13640000000
1!
b111 %
1'
b111 +
#13650000000
0!
0'
#13660000000
1!
0$
b1000 %
1'
0*
b1000 +
#13670000000
0!
0'
#13680000000
1!
b1001 %
1'
b1001 +
#13690000000
0!
0'
#13700000000
1!
b0 %
1'
b0 +
#13710000000
0!
0'
#13720000000
1!
1$
b1 %
1'
1*
b1 +
#13730000000
0!
0'
#13740000000
1!
b10 %
1'
b10 +
#13750000000
0!
0'
#13760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#13770000000
0!
0'
#13780000000
1!
b100 %
1'
b100 +
#13790000000
0!
0'
#13800000000
1!
b101 %
1'
b101 +
#13810000000
0!
0'
#13820000000
1!
0$
b110 %
1'
0*
b110 +
#13830000000
0!
0'
#13840000000
1!
b111 %
1'
b111 +
#13850000000
0!
0'
#13860000000
1!
b1000 %
1'
b1000 +
#13870000000
0!
0'
#13880000000
1!
b1001 %
1'
b1001 +
#13890000000
0!
0'
#13900000000
1!
b0 %
1'
b0 +
#13910000000
0!
0'
#13920000000
1!
1$
b1 %
1'
1*
b1 +
#13930000000
0!
0'
#13940000000
1!
b10 %
1'
b10 +
#13950000000
0!
0'
#13960000000
1!
b11 %
1'
b11 +
#13970000000
1"
1(
#13980000000
0!
0"
b100 &
0'
0(
b100 ,
#13990000000
1!
b100 %
1'
b100 +
#14000000000
0!
0'
#14010000000
1!
b101 %
1'
b101 +
#14020000000
0!
0'
#14030000000
1!
b110 %
1'
b110 +
#14040000000
0!
0'
#14050000000
1!
b111 %
1'
b111 +
#14060000000
0!
0'
#14070000000
1!
0$
b1000 %
1'
0*
b1000 +
#14080000000
0!
0'
#14090000000
1!
b1001 %
1'
b1001 +
#14100000000
0!
0'
#14110000000
1!
b0 %
1'
b0 +
#14120000000
0!
0'
#14130000000
1!
1$
b1 %
1'
1*
b1 +
#14140000000
0!
0'
#14150000000
1!
b10 %
1'
b10 +
#14160000000
0!
0'
#14170000000
1!
b11 %
1'
b11 +
#14180000000
0!
0'
#14190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#14200000000
0!
0'
#14210000000
1!
b101 %
1'
b101 +
#14220000000
0!
0'
#14230000000
1!
0$
b110 %
1'
0*
b110 +
#14240000000
0!
0'
#14250000000
1!
b111 %
1'
b111 +
#14260000000
0!
0'
#14270000000
1!
b1000 %
1'
b1000 +
#14280000000
0!
0'
#14290000000
1!
b1001 %
1'
b1001 +
#14300000000
0!
0'
#14310000000
1!
b0 %
1'
b0 +
#14320000000
0!
0'
#14330000000
1!
1$
b1 %
1'
1*
b1 +
#14340000000
0!
0'
#14350000000
1!
b10 %
1'
b10 +
#14360000000
0!
0'
#14370000000
1!
b11 %
1'
b11 +
#14380000000
0!
0'
#14390000000
1!
b100 %
1'
b100 +
#14400000000
1"
1(
#14410000000
0!
0"
b100 &
0'
0(
b100 ,
#14420000000
1!
b101 %
1'
b101 +
#14430000000
0!
0'
#14440000000
1!
b110 %
1'
b110 +
#14450000000
0!
0'
#14460000000
1!
b111 %
1'
b111 +
#14470000000
0!
0'
#14480000000
1!
0$
b1000 %
1'
0*
b1000 +
#14490000000
0!
0'
#14500000000
1!
b1001 %
1'
b1001 +
#14510000000
0!
0'
#14520000000
1!
b0 %
1'
b0 +
#14530000000
0!
0'
#14540000000
1!
1$
b1 %
1'
1*
b1 +
#14550000000
0!
0'
#14560000000
1!
b10 %
1'
b10 +
#14570000000
0!
0'
#14580000000
1!
b11 %
1'
b11 +
#14590000000
0!
0'
#14600000000
1!
b100 %
1'
b100 +
#14610000000
0!
0'
#14620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#14630000000
0!
0'
#14640000000
1!
0$
b110 %
1'
0*
b110 +
#14650000000
0!
0'
#14660000000
1!
b111 %
1'
b111 +
#14670000000
0!
0'
#14680000000
1!
b1000 %
1'
b1000 +
#14690000000
0!
0'
#14700000000
1!
b1001 %
1'
b1001 +
#14710000000
0!
0'
#14720000000
1!
b0 %
1'
b0 +
#14730000000
0!
0'
#14740000000
1!
1$
b1 %
1'
1*
b1 +
#14750000000
0!
0'
#14760000000
1!
b10 %
1'
b10 +
#14770000000
0!
0'
#14780000000
1!
b11 %
1'
b11 +
#14790000000
0!
0'
#14800000000
1!
b100 %
1'
b100 +
#14810000000
0!
0'
#14820000000
1!
b101 %
1'
b101 +
#14830000000
1"
1(
#14840000000
0!
0"
b100 &
0'
0(
b100 ,
#14850000000
1!
b110 %
1'
b110 +
#14860000000
0!
0'
#14870000000
1!
b111 %
1'
b111 +
#14880000000
0!
0'
#14890000000
1!
0$
b1000 %
1'
0*
b1000 +
#14900000000
0!
0'
#14910000000
1!
b1001 %
1'
b1001 +
#14920000000
0!
0'
#14930000000
1!
b0 %
1'
b0 +
#14940000000
0!
0'
#14950000000
1!
1$
b1 %
1'
1*
b1 +
#14960000000
0!
0'
#14970000000
1!
b10 %
1'
b10 +
#14980000000
0!
0'
#14990000000
1!
b11 %
1'
b11 +
#15000000000
0!
0'
#15010000000
1!
b100 %
1'
b100 +
#15020000000
0!
0'
#15030000000
1!
b101 %
1'
b101 +
#15040000000
0!
0'
#15050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#15060000000
0!
0'
#15070000000
1!
b111 %
1'
b111 +
#15080000000
0!
0'
#15090000000
1!
b1000 %
1'
b1000 +
#15100000000
0!
0'
#15110000000
1!
b1001 %
1'
b1001 +
#15120000000
0!
0'
#15130000000
1!
b0 %
1'
b0 +
#15140000000
0!
0'
#15150000000
1!
1$
b1 %
1'
1*
b1 +
#15160000000
0!
0'
#15170000000
1!
b10 %
1'
b10 +
#15180000000
0!
0'
#15190000000
1!
b11 %
1'
b11 +
#15200000000
0!
0'
#15210000000
1!
b100 %
1'
b100 +
#15220000000
0!
0'
#15230000000
1!
b101 %
1'
b101 +
#15240000000
0!
0'
#15250000000
1!
0$
b110 %
1'
0*
b110 +
#15260000000
1"
1(
#15270000000
0!
0"
b100 &
0'
0(
b100 ,
#15280000000
1!
1$
b111 %
1'
1*
b111 +
#15290000000
0!
0'
#15300000000
1!
0$
b1000 %
1'
0*
b1000 +
#15310000000
0!
0'
#15320000000
1!
b1001 %
1'
b1001 +
#15330000000
0!
0'
#15340000000
1!
b0 %
1'
b0 +
#15350000000
0!
0'
#15360000000
1!
1$
b1 %
1'
1*
b1 +
#15370000000
0!
0'
#15380000000
1!
b10 %
1'
b10 +
#15390000000
0!
0'
#15400000000
1!
b11 %
1'
b11 +
#15410000000
0!
0'
#15420000000
1!
b100 %
1'
b100 +
#15430000000
0!
0'
#15440000000
1!
b101 %
1'
b101 +
#15450000000
0!
0'
#15460000000
1!
b110 %
1'
b110 +
#15470000000
0!
0'
#15480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#15490000000
0!
0'
#15500000000
1!
b1000 %
1'
b1000 +
#15510000000
0!
0'
#15520000000
1!
b1001 %
1'
b1001 +
#15530000000
0!
0'
#15540000000
1!
b0 %
1'
b0 +
#15550000000
0!
0'
#15560000000
1!
1$
b1 %
1'
1*
b1 +
#15570000000
0!
0'
#15580000000
1!
b10 %
1'
b10 +
#15590000000
0!
0'
#15600000000
1!
b11 %
1'
b11 +
#15610000000
0!
0'
#15620000000
1!
b100 %
1'
b100 +
#15630000000
0!
0'
#15640000000
1!
b101 %
1'
b101 +
#15650000000
0!
0'
#15660000000
1!
0$
b110 %
1'
0*
b110 +
#15670000000
0!
0'
#15680000000
1!
b111 %
1'
b111 +
#15690000000
1"
1(
#15700000000
0!
0"
b100 &
0'
0(
b100 ,
#15710000000
1!
b1000 %
1'
b1000 +
#15720000000
0!
0'
#15730000000
1!
b1001 %
1'
b1001 +
#15740000000
0!
0'
#15750000000
1!
b0 %
1'
b0 +
#15760000000
0!
0'
#15770000000
1!
1$
b1 %
1'
1*
b1 +
#15780000000
0!
0'
#15790000000
1!
b10 %
1'
b10 +
#15800000000
0!
0'
#15810000000
1!
b11 %
1'
b11 +
#15820000000
0!
0'
#15830000000
1!
b100 %
1'
b100 +
#15840000000
0!
0'
#15850000000
1!
b101 %
1'
b101 +
#15860000000
0!
0'
#15870000000
1!
b110 %
1'
b110 +
#15880000000
0!
0'
#15890000000
1!
b111 %
1'
b111 +
#15900000000
0!
0'
#15910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#15920000000
0!
0'
#15930000000
1!
b1001 %
1'
b1001 +
#15940000000
0!
0'
#15950000000
1!
b0 %
1'
b0 +
#15960000000
0!
0'
#15970000000
1!
1$
b1 %
1'
1*
b1 +
#15980000000
0!
0'
#15990000000
1!
b10 %
1'
b10 +
#16000000000
0!
0'
#16010000000
1!
b11 %
1'
b11 +
#16020000000
0!
0'
#16030000000
1!
b100 %
1'
b100 +
#16040000000
0!
0'
#16050000000
1!
b101 %
1'
b101 +
#16060000000
0!
0'
#16070000000
1!
0$
b110 %
1'
0*
b110 +
#16080000000
0!
0'
#16090000000
1!
b111 %
1'
b111 +
#16100000000
0!
0'
#16110000000
1!
b1000 %
1'
b1000 +
#16120000000
1"
1(
#16130000000
0!
0"
b100 &
0'
0(
b100 ,
#16140000000
1!
b1001 %
1'
b1001 +
#16150000000
0!
0'
#16160000000
1!
b0 %
1'
b0 +
#16170000000
0!
0'
#16180000000
1!
1$
b1 %
1'
1*
b1 +
#16190000000
0!
0'
#16200000000
1!
b10 %
1'
b10 +
#16210000000
0!
0'
#16220000000
1!
b11 %
1'
b11 +
#16230000000
0!
0'
#16240000000
1!
b100 %
1'
b100 +
#16250000000
0!
0'
#16260000000
1!
b101 %
1'
b101 +
#16270000000
0!
0'
#16280000000
1!
b110 %
1'
b110 +
#16290000000
0!
0'
#16300000000
1!
b111 %
1'
b111 +
#16310000000
0!
0'
#16320000000
1!
0$
b1000 %
1'
0*
b1000 +
#16330000000
0!
0'
#16340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#16350000000
0!
0'
#16360000000
1!
b0 %
1'
b0 +
#16370000000
0!
0'
#16380000000
1!
1$
b1 %
1'
1*
b1 +
#16390000000
0!
0'
#16400000000
1!
b10 %
1'
b10 +
#16410000000
0!
0'
#16420000000
1!
b11 %
1'
b11 +
#16430000000
0!
0'
#16440000000
1!
b100 %
1'
b100 +
#16450000000
0!
0'
#16460000000
1!
b101 %
1'
b101 +
#16470000000
0!
0'
#16480000000
1!
0$
b110 %
1'
0*
b110 +
#16490000000
0!
0'
#16500000000
1!
b111 %
1'
b111 +
#16510000000
0!
0'
#16520000000
1!
b1000 %
1'
b1000 +
#16530000000
0!
0'
#16540000000
1!
b1001 %
1'
b1001 +
#16550000000
1"
1(
#16560000000
0!
0"
b100 &
0'
0(
b100 ,
#16570000000
1!
b0 %
1'
b0 +
#16580000000
0!
0'
#16590000000
1!
1$
b1 %
1'
1*
b1 +
#16600000000
0!
0'
#16610000000
1!
b10 %
1'
b10 +
#16620000000
0!
0'
#16630000000
1!
b11 %
1'
b11 +
#16640000000
0!
0'
#16650000000
1!
b100 %
1'
b100 +
#16660000000
0!
0'
#16670000000
1!
b101 %
1'
b101 +
#16680000000
0!
0'
#16690000000
1!
b110 %
1'
b110 +
#16700000000
0!
0'
#16710000000
1!
b111 %
1'
b111 +
#16720000000
0!
0'
#16730000000
1!
0$
b1000 %
1'
0*
b1000 +
#16740000000
0!
0'
#16750000000
1!
b1001 %
1'
b1001 +
#16760000000
0!
0'
#16770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#16780000000
0!
0'
#16790000000
1!
1$
b1 %
1'
1*
b1 +
#16800000000
0!
0'
#16810000000
1!
b10 %
1'
b10 +
#16820000000
0!
0'
#16830000000
1!
b11 %
1'
b11 +
#16840000000
0!
0'
#16850000000
1!
b100 %
1'
b100 +
#16860000000
0!
0'
#16870000000
1!
b101 %
1'
b101 +
#16880000000
0!
0'
#16890000000
1!
0$
b110 %
1'
0*
b110 +
#16900000000
0!
0'
#16910000000
1!
b111 %
1'
b111 +
#16920000000
0!
0'
#16930000000
1!
b1000 %
1'
b1000 +
#16940000000
0!
0'
#16950000000
1!
b1001 %
1'
b1001 +
#16960000000
0!
0'
#16970000000
1!
b0 %
1'
b0 +
#16980000000
1"
1(
#16990000000
0!
0"
b100 &
0'
0(
b100 ,
#17000000000
1!
1$
b1 %
1'
1*
b1 +
#17010000000
0!
0'
#17020000000
1!
b10 %
1'
b10 +
#17030000000
0!
0'
#17040000000
1!
b11 %
1'
b11 +
#17050000000
0!
0'
#17060000000
1!
b100 %
1'
b100 +
#17070000000
0!
0'
#17080000000
1!
b101 %
1'
b101 +
#17090000000
0!
0'
#17100000000
1!
b110 %
1'
b110 +
#17110000000
0!
0'
#17120000000
1!
b111 %
1'
b111 +
#17130000000
0!
0'
#17140000000
1!
0$
b1000 %
1'
0*
b1000 +
#17150000000
0!
0'
#17160000000
1!
b1001 %
1'
b1001 +
#17170000000
0!
0'
#17180000000
1!
b0 %
1'
b0 +
#17190000000
0!
0'
#17200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#17210000000
0!
0'
#17220000000
1!
b10 %
1'
b10 +
#17230000000
0!
0'
#17240000000
1!
b11 %
1'
b11 +
#17250000000
0!
0'
#17260000000
1!
b100 %
1'
b100 +
#17270000000
0!
0'
#17280000000
1!
b101 %
1'
b101 +
#17290000000
0!
0'
#17300000000
1!
0$
b110 %
1'
0*
b110 +
#17310000000
0!
0'
#17320000000
1!
b111 %
1'
b111 +
#17330000000
0!
0'
#17340000000
1!
b1000 %
1'
b1000 +
#17350000000
0!
0'
#17360000000
1!
b1001 %
1'
b1001 +
#17370000000
0!
0'
#17380000000
1!
b0 %
1'
b0 +
#17390000000
0!
0'
#17400000000
1!
1$
b1 %
1'
1*
b1 +
#17410000000
1"
1(
#17420000000
0!
0"
b100 &
0'
0(
b100 ,
#17430000000
1!
b10 %
1'
b10 +
#17440000000
0!
0'
#17450000000
1!
b11 %
1'
b11 +
#17460000000
0!
0'
#17470000000
1!
b100 %
1'
b100 +
#17480000000
0!
0'
#17490000000
1!
b101 %
1'
b101 +
#17500000000
0!
0'
#17510000000
1!
b110 %
1'
b110 +
#17520000000
0!
0'
#17530000000
1!
b111 %
1'
b111 +
#17540000000
0!
0'
#17550000000
1!
0$
b1000 %
1'
0*
b1000 +
#17560000000
0!
0'
#17570000000
1!
b1001 %
1'
b1001 +
#17580000000
0!
0'
#17590000000
1!
b0 %
1'
b0 +
#17600000000
0!
0'
#17610000000
1!
1$
b1 %
1'
1*
b1 +
#17620000000
0!
0'
#17630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#17640000000
0!
0'
#17650000000
1!
b11 %
1'
b11 +
#17660000000
0!
0'
#17670000000
1!
b100 %
1'
b100 +
#17680000000
0!
0'
#17690000000
1!
b101 %
1'
b101 +
#17700000000
0!
0'
#17710000000
1!
0$
b110 %
1'
0*
b110 +
#17720000000
0!
0'
#17730000000
1!
b111 %
1'
b111 +
#17740000000
0!
0'
#17750000000
1!
b1000 %
1'
b1000 +
#17760000000
0!
0'
#17770000000
1!
b1001 %
1'
b1001 +
#17780000000
0!
0'
#17790000000
1!
b0 %
1'
b0 +
#17800000000
0!
0'
#17810000000
1!
1$
b1 %
1'
1*
b1 +
#17820000000
0!
0'
#17830000000
1!
b10 %
1'
b10 +
#17840000000
1"
1(
#17850000000
0!
0"
b100 &
0'
0(
b100 ,
#17860000000
1!
b11 %
1'
b11 +
#17870000000
0!
0'
#17880000000
1!
b100 %
1'
b100 +
#17890000000
0!
0'
#17900000000
1!
b101 %
1'
b101 +
#17910000000
0!
0'
#17920000000
1!
b110 %
1'
b110 +
#17930000000
0!
0'
#17940000000
1!
b111 %
1'
b111 +
#17950000000
0!
0'
#17960000000
1!
0$
b1000 %
1'
0*
b1000 +
#17970000000
0!
0'
#17980000000
1!
b1001 %
1'
b1001 +
#17990000000
0!
0'
#18000000000
1!
b0 %
1'
b0 +
#18010000000
0!
0'
#18020000000
1!
1$
b1 %
1'
1*
b1 +
#18030000000
0!
0'
#18040000000
1!
b10 %
1'
b10 +
#18050000000
0!
0'
#18060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#18070000000
0!
0'
#18080000000
1!
b100 %
1'
b100 +
#18090000000
0!
0'
#18100000000
1!
b101 %
1'
b101 +
#18110000000
0!
0'
#18120000000
1!
0$
b110 %
1'
0*
b110 +
#18130000000
0!
0'
#18140000000
1!
b111 %
1'
b111 +
#18150000000
0!
0'
#18160000000
1!
b1000 %
1'
b1000 +
#18170000000
0!
0'
#18180000000
1!
b1001 %
1'
b1001 +
#18190000000
0!
0'
#18200000000
1!
b0 %
1'
b0 +
#18210000000
0!
0'
#18220000000
1!
1$
b1 %
1'
1*
b1 +
#18230000000
0!
0'
#18240000000
1!
b10 %
1'
b10 +
#18250000000
0!
0'
#18260000000
1!
b11 %
1'
b11 +
#18270000000
1"
1(
#18280000000
0!
0"
b100 &
0'
0(
b100 ,
#18290000000
1!
b100 %
1'
b100 +
#18300000000
0!
0'
#18310000000
1!
b101 %
1'
b101 +
#18320000000
0!
0'
#18330000000
1!
b110 %
1'
b110 +
#18340000000
0!
0'
#18350000000
1!
b111 %
1'
b111 +
#18360000000
0!
0'
#18370000000
1!
0$
b1000 %
1'
0*
b1000 +
#18380000000
0!
0'
#18390000000
1!
b1001 %
1'
b1001 +
#18400000000
0!
0'
#18410000000
1!
b0 %
1'
b0 +
#18420000000
0!
0'
#18430000000
1!
1$
b1 %
1'
1*
b1 +
#18440000000
0!
0'
#18450000000
1!
b10 %
1'
b10 +
#18460000000
0!
0'
#18470000000
1!
b11 %
1'
b11 +
#18480000000
0!
0'
#18490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#18500000000
0!
0'
#18510000000
1!
b101 %
1'
b101 +
#18520000000
0!
0'
#18530000000
1!
0$
b110 %
1'
0*
b110 +
#18540000000
0!
0'
#18550000000
1!
b111 %
1'
b111 +
#18560000000
0!
0'
#18570000000
1!
b1000 %
1'
b1000 +
#18580000000
0!
0'
#18590000000
1!
b1001 %
1'
b1001 +
#18600000000
0!
0'
#18610000000
1!
b0 %
1'
b0 +
#18620000000
0!
0'
#18630000000
1!
1$
b1 %
1'
1*
b1 +
#18640000000
0!
0'
#18650000000
1!
b10 %
1'
b10 +
#18660000000
0!
0'
#18670000000
1!
b11 %
1'
b11 +
#18680000000
0!
0'
#18690000000
1!
b100 %
1'
b100 +
#18700000000
1"
1(
#18710000000
0!
0"
b100 &
0'
0(
b100 ,
#18720000000
1!
b101 %
1'
b101 +
#18730000000
0!
0'
#18740000000
1!
b110 %
1'
b110 +
#18750000000
0!
0'
#18760000000
1!
b111 %
1'
b111 +
#18770000000
0!
0'
#18780000000
1!
0$
b1000 %
1'
0*
b1000 +
#18790000000
0!
0'
#18800000000
1!
b1001 %
1'
b1001 +
#18810000000
0!
0'
#18820000000
1!
b0 %
1'
b0 +
#18830000000
0!
0'
#18840000000
1!
1$
b1 %
1'
1*
b1 +
#18850000000
0!
0'
#18860000000
1!
b10 %
1'
b10 +
#18870000000
0!
0'
#18880000000
1!
b11 %
1'
b11 +
#18890000000
0!
0'
#18900000000
1!
b100 %
1'
b100 +
#18910000000
0!
0'
#18920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#18930000000
0!
0'
#18940000000
1!
0$
b110 %
1'
0*
b110 +
#18950000000
0!
0'
#18960000000
1!
b111 %
1'
b111 +
#18970000000
0!
0'
#18980000000
1!
b1000 %
1'
b1000 +
#18990000000
0!
0'
#19000000000
1!
b1001 %
1'
b1001 +
#19010000000
0!
0'
#19020000000
1!
b0 %
1'
b0 +
#19030000000
0!
0'
#19040000000
1!
1$
b1 %
1'
1*
b1 +
#19050000000
0!
0'
#19060000000
1!
b10 %
1'
b10 +
#19070000000
0!
0'
#19080000000
1!
b11 %
1'
b11 +
#19090000000
0!
0'
#19100000000
1!
b100 %
1'
b100 +
#19110000000
0!
0'
#19120000000
1!
b101 %
1'
b101 +
#19130000000
1"
1(
#19140000000
0!
0"
b100 &
0'
0(
b100 ,
#19150000000
1!
b110 %
1'
b110 +
#19160000000
0!
0'
#19170000000
1!
b111 %
1'
b111 +
#19180000000
0!
0'
#19190000000
1!
0$
b1000 %
1'
0*
b1000 +
#19200000000
0!
0'
#19210000000
1!
b1001 %
1'
b1001 +
#19220000000
0!
0'
#19230000000
1!
b0 %
1'
b0 +
#19240000000
0!
0'
#19250000000
1!
1$
b1 %
1'
1*
b1 +
#19260000000
0!
0'
#19270000000
1!
b10 %
1'
b10 +
#19280000000
0!
0'
#19290000000
1!
b11 %
1'
b11 +
#19300000000
0!
0'
#19310000000
1!
b100 %
1'
b100 +
#19320000000
0!
0'
#19330000000
1!
b101 %
1'
b101 +
#19340000000
0!
0'
#19350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#19360000000
0!
0'
#19370000000
1!
b111 %
1'
b111 +
#19380000000
0!
0'
#19390000000
1!
b1000 %
1'
b1000 +
#19400000000
0!
0'
#19410000000
1!
b1001 %
1'
b1001 +
#19420000000
0!
0'
#19430000000
1!
b0 %
1'
b0 +
#19440000000
0!
0'
#19450000000
1!
1$
b1 %
1'
1*
b1 +
#19460000000
0!
0'
#19470000000
1!
b10 %
1'
b10 +
#19480000000
0!
0'
#19490000000
1!
b11 %
1'
b11 +
#19500000000
0!
0'
#19510000000
1!
b100 %
1'
b100 +
#19520000000
0!
0'
#19530000000
1!
b101 %
1'
b101 +
#19540000000
0!
0'
#19550000000
1!
0$
b110 %
1'
0*
b110 +
#19560000000
1"
1(
#19570000000
0!
0"
b100 &
0'
0(
b100 ,
#19580000000
1!
1$
b111 %
1'
1*
b111 +
#19590000000
0!
0'
#19600000000
1!
0$
b1000 %
1'
0*
b1000 +
#19610000000
0!
0'
#19620000000
1!
b1001 %
1'
b1001 +
#19630000000
0!
0'
#19640000000
1!
b0 %
1'
b0 +
#19650000000
0!
0'
#19660000000
1!
1$
b1 %
1'
1*
b1 +
#19670000000
0!
0'
#19680000000
1!
b10 %
1'
b10 +
#19690000000
0!
0'
#19700000000
1!
b11 %
1'
b11 +
#19710000000
0!
0'
#19720000000
1!
b100 %
1'
b100 +
#19730000000
0!
0'
#19740000000
1!
b101 %
1'
b101 +
#19750000000
0!
0'
#19760000000
1!
b110 %
1'
b110 +
#19770000000
0!
0'
#19780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#19790000000
0!
0'
#19800000000
1!
b1000 %
1'
b1000 +
#19810000000
0!
0'
#19820000000
1!
b1001 %
1'
b1001 +
#19830000000
0!
0'
#19840000000
1!
b0 %
1'
b0 +
#19850000000
0!
0'
#19860000000
1!
1$
b1 %
1'
1*
b1 +
#19870000000
0!
0'
#19880000000
1!
b10 %
1'
b10 +
#19890000000
0!
0'
#19900000000
1!
b11 %
1'
b11 +
#19910000000
0!
0'
#19920000000
1!
b100 %
1'
b100 +
#19930000000
0!
0'
#19940000000
1!
b101 %
1'
b101 +
#19950000000
0!
0'
#19960000000
1!
0$
b110 %
1'
0*
b110 +
#19970000000
0!
0'
#19980000000
1!
b111 %
1'
b111 +
#19990000000
1"
1(
#20000000000
0!
0"
b100 &
0'
0(
b100 ,
#20010000000
1!
b1000 %
1'
b1000 +
#20020000000
0!
0'
#20030000000
1!
b1001 %
1'
b1001 +
#20040000000
0!
0'
#20050000000
1!
b0 %
1'
b0 +
#20060000000
0!
0'
#20070000000
1!
1$
b1 %
1'
1*
b1 +
#20080000000
0!
0'
#20090000000
1!
b10 %
1'
b10 +
#20100000000
0!
0'
#20110000000
1!
b11 %
1'
b11 +
#20120000000
0!
0'
#20130000000
1!
b100 %
1'
b100 +
#20140000000
0!
0'
#20150000000
1!
b101 %
1'
b101 +
#20160000000
0!
0'
#20170000000
1!
b110 %
1'
b110 +
#20180000000
0!
0'
#20190000000
1!
b111 %
1'
b111 +
#20200000000
0!
0'
#20210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#20220000000
0!
0'
#20230000000
1!
b1001 %
1'
b1001 +
#20240000000
0!
0'
#20250000000
1!
b0 %
1'
b0 +
#20260000000
0!
0'
#20270000000
1!
1$
b1 %
1'
1*
b1 +
#20280000000
0!
0'
#20290000000
1!
b10 %
1'
b10 +
#20300000000
0!
0'
#20310000000
1!
b11 %
1'
b11 +
#20320000000
0!
0'
#20330000000
1!
b100 %
1'
b100 +
#20340000000
0!
0'
#20350000000
1!
b101 %
1'
b101 +
#20360000000
0!
0'
#20370000000
1!
0$
b110 %
1'
0*
b110 +
#20380000000
0!
0'
#20390000000
1!
b111 %
1'
b111 +
#20400000000
0!
0'
#20410000000
1!
b1000 %
1'
b1000 +
#20420000000
1"
1(
#20430000000
0!
0"
b100 &
0'
0(
b100 ,
#20440000000
1!
b1001 %
1'
b1001 +
#20450000000
0!
0'
#20460000000
1!
b0 %
1'
b0 +
#20470000000
0!
0'
#20480000000
1!
1$
b1 %
1'
1*
b1 +
#20490000000
0!
0'
#20500000000
1!
b10 %
1'
b10 +
#20510000000
0!
0'
#20520000000
1!
b11 %
1'
b11 +
#20530000000
0!
0'
#20540000000
1!
b100 %
1'
b100 +
#20550000000
0!
0'
#20560000000
1!
b101 %
1'
b101 +
#20570000000
0!
0'
#20580000000
1!
b110 %
1'
b110 +
#20590000000
0!
0'
#20600000000
1!
b111 %
1'
b111 +
#20610000000
0!
0'
#20620000000
1!
0$
b1000 %
1'
0*
b1000 +
#20630000000
0!
0'
#20640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#20650000000
0!
0'
#20660000000
1!
b0 %
1'
b0 +
#20670000000
0!
0'
#20680000000
1!
1$
b1 %
1'
1*
b1 +
#20690000000
0!
0'
#20700000000
1!
b10 %
1'
b10 +
#20710000000
0!
0'
#20720000000
1!
b11 %
1'
b11 +
#20730000000
0!
0'
#20740000000
1!
b100 %
1'
b100 +
#20750000000
0!
0'
#20760000000
1!
b101 %
1'
b101 +
#20770000000
0!
0'
#20780000000
1!
0$
b110 %
1'
0*
b110 +
#20790000000
0!
0'
#20800000000
1!
b111 %
1'
b111 +
#20810000000
0!
0'
#20820000000
1!
b1000 %
1'
b1000 +
#20830000000
0!
0'
#20840000000
1!
b1001 %
1'
b1001 +
#20850000000
1"
1(
#20860000000
0!
0"
b100 &
0'
0(
b100 ,
#20870000000
1!
b0 %
1'
b0 +
#20880000000
0!
0'
#20890000000
1!
1$
b1 %
1'
1*
b1 +
#20900000000
0!
0'
#20910000000
1!
b10 %
1'
b10 +
#20920000000
0!
0'
#20930000000
1!
b11 %
1'
b11 +
#20940000000
0!
0'
#20950000000
1!
b100 %
1'
b100 +
#20960000000
0!
0'
#20970000000
1!
b101 %
1'
b101 +
#20980000000
0!
0'
#20990000000
1!
b110 %
1'
b110 +
#21000000000
0!
0'
#21010000000
1!
b111 %
1'
b111 +
#21020000000
0!
0'
#21030000000
1!
0$
b1000 %
1'
0*
b1000 +
#21040000000
0!
0'
#21050000000
1!
b1001 %
1'
b1001 +
#21060000000
0!
0'
#21070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#21080000000
0!
0'
#21090000000
1!
1$
b1 %
1'
1*
b1 +
#21100000000
0!
0'
#21110000000
1!
b10 %
1'
b10 +
#21120000000
0!
0'
#21130000000
1!
b11 %
1'
b11 +
#21140000000
0!
0'
#21150000000
1!
b100 %
1'
b100 +
#21160000000
0!
0'
#21170000000
1!
b101 %
1'
b101 +
#21180000000
0!
0'
#21190000000
1!
0$
b110 %
1'
0*
b110 +
#21200000000
0!
0'
#21210000000
1!
b111 %
1'
b111 +
#21220000000
0!
0'
#21230000000
1!
b1000 %
1'
b1000 +
#21240000000
0!
0'
#21250000000
1!
b1001 %
1'
b1001 +
#21260000000
0!
0'
#21270000000
1!
b0 %
1'
b0 +
#21280000000
1"
1(
#21290000000
0!
0"
b100 &
0'
0(
b100 ,
#21300000000
1!
1$
b1 %
1'
1*
b1 +
#21310000000
0!
0'
#21320000000
1!
b10 %
1'
b10 +
#21330000000
0!
0'
#21340000000
1!
b11 %
1'
b11 +
#21350000000
0!
0'
#21360000000
1!
b100 %
1'
b100 +
#21370000000
0!
0'
#21380000000
1!
b101 %
1'
b101 +
#21390000000
0!
0'
#21400000000
1!
b110 %
1'
b110 +
#21410000000
0!
0'
#21420000000
1!
b111 %
1'
b111 +
#21430000000
0!
0'
#21440000000
1!
0$
b1000 %
1'
0*
b1000 +
#21450000000
0!
0'
#21460000000
1!
b1001 %
1'
b1001 +
#21470000000
0!
0'
#21480000000
1!
b0 %
1'
b0 +
#21490000000
0!
0'
#21500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#21510000000
0!
0'
#21520000000
1!
b10 %
1'
b10 +
#21530000000
0!
0'
#21540000000
1!
b11 %
1'
b11 +
#21550000000
0!
0'
#21560000000
1!
b100 %
1'
b100 +
#21570000000
0!
0'
#21580000000
1!
b101 %
1'
b101 +
#21590000000
0!
0'
#21600000000
1!
0$
b110 %
1'
0*
b110 +
#21610000000
0!
0'
#21620000000
1!
b111 %
1'
b111 +
#21630000000
0!
0'
#21640000000
1!
b1000 %
1'
b1000 +
#21650000000
0!
0'
#21660000000
1!
b1001 %
1'
b1001 +
#21670000000
0!
0'
#21680000000
1!
b0 %
1'
b0 +
#21690000000
0!
0'
#21700000000
1!
1$
b1 %
1'
1*
b1 +
#21710000000
1"
1(
#21720000000
0!
0"
b100 &
0'
0(
b100 ,
#21730000000
1!
b10 %
1'
b10 +
#21740000000
0!
0'
#21750000000
1!
b11 %
1'
b11 +
#21760000000
0!
0'
#21770000000
1!
b100 %
1'
b100 +
#21780000000
0!
0'
#21790000000
1!
b101 %
1'
b101 +
#21800000000
0!
0'
#21810000000
1!
b110 %
1'
b110 +
#21820000000
0!
0'
#21830000000
1!
b111 %
1'
b111 +
#21840000000
0!
0'
#21850000000
1!
0$
b1000 %
1'
0*
b1000 +
#21860000000
0!
0'
#21870000000
1!
b1001 %
1'
b1001 +
#21880000000
0!
0'
#21890000000
1!
b0 %
1'
b0 +
#21900000000
0!
0'
#21910000000
1!
1$
b1 %
1'
1*
b1 +
#21920000000
0!
0'
#21930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#21940000000
0!
0'
#21950000000
1!
b11 %
1'
b11 +
#21960000000
0!
0'
#21970000000
1!
b100 %
1'
b100 +
#21980000000
0!
0'
#21990000000
1!
b101 %
1'
b101 +
#22000000000
0!
0'
#22010000000
1!
0$
b110 %
1'
0*
b110 +
#22020000000
0!
0'
#22030000000
1!
b111 %
1'
b111 +
#22040000000
0!
0'
#22050000000
1!
b1000 %
1'
b1000 +
#22060000000
0!
0'
#22070000000
1!
b1001 %
1'
b1001 +
#22080000000
0!
0'
#22090000000
1!
b0 %
1'
b0 +
#22100000000
0!
0'
#22110000000
1!
1$
b1 %
1'
1*
b1 +
#22120000000
0!
0'
#22130000000
1!
b10 %
1'
b10 +
#22140000000
1"
1(
#22150000000
0!
0"
b100 &
0'
0(
b100 ,
#22160000000
1!
b11 %
1'
b11 +
#22170000000
0!
0'
#22180000000
1!
b100 %
1'
b100 +
#22190000000
0!
0'
#22200000000
1!
b101 %
1'
b101 +
#22210000000
0!
0'
#22220000000
1!
b110 %
1'
b110 +
#22230000000
0!
0'
#22240000000
1!
b111 %
1'
b111 +
#22250000000
0!
0'
#22260000000
1!
0$
b1000 %
1'
0*
b1000 +
#22270000000
0!
0'
#22280000000
1!
b1001 %
1'
b1001 +
#22290000000
0!
0'
#22300000000
1!
b0 %
1'
b0 +
#22310000000
0!
0'
#22320000000
1!
1$
b1 %
1'
1*
b1 +
#22330000000
0!
0'
#22340000000
1!
b10 %
1'
b10 +
#22350000000
0!
0'
#22360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#22370000000
0!
0'
#22380000000
1!
b100 %
1'
b100 +
#22390000000
0!
0'
#22400000000
1!
b101 %
1'
b101 +
#22410000000
0!
0'
#22420000000
1!
0$
b110 %
1'
0*
b110 +
#22430000000
0!
0'
#22440000000
1!
b111 %
1'
b111 +
#22450000000
0!
0'
#22460000000
1!
b1000 %
1'
b1000 +
#22470000000
0!
0'
#22480000000
1!
b1001 %
1'
b1001 +
#22490000000
0!
0'
#22500000000
1!
b0 %
1'
b0 +
#22510000000
0!
0'
#22520000000
1!
1$
b1 %
1'
1*
b1 +
#22530000000
0!
0'
#22540000000
1!
b10 %
1'
b10 +
#22550000000
0!
0'
#22560000000
1!
b11 %
1'
b11 +
#22570000000
1"
1(
#22580000000
0!
0"
b100 &
0'
0(
b100 ,
#22590000000
1!
b100 %
1'
b100 +
#22600000000
0!
0'
#22610000000
1!
b101 %
1'
b101 +
#22620000000
0!
0'
#22630000000
1!
b110 %
1'
b110 +
#22640000000
0!
0'
#22650000000
1!
b111 %
1'
b111 +
#22660000000
0!
0'
#22670000000
1!
0$
b1000 %
1'
0*
b1000 +
#22680000000
0!
0'
#22690000000
1!
b1001 %
1'
b1001 +
#22700000000
0!
0'
#22710000000
1!
b0 %
1'
b0 +
#22720000000
0!
0'
#22730000000
1!
1$
b1 %
1'
1*
b1 +
#22740000000
0!
0'
#22750000000
1!
b10 %
1'
b10 +
#22760000000
0!
0'
#22770000000
1!
b11 %
1'
b11 +
#22780000000
0!
0'
#22790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#22800000000
0!
0'
#22810000000
1!
b101 %
1'
b101 +
#22820000000
0!
0'
#22830000000
1!
0$
b110 %
1'
0*
b110 +
#22840000000
0!
0'
#22850000000
1!
b111 %
1'
b111 +
#22860000000
0!
0'
#22870000000
1!
b1000 %
1'
b1000 +
#22880000000
0!
0'
#22890000000
1!
b1001 %
1'
b1001 +
#22900000000
0!
0'
#22910000000
1!
b0 %
1'
b0 +
#22920000000
0!
0'
#22930000000
1!
1$
b1 %
1'
1*
b1 +
#22940000000
0!
0'
#22950000000
1!
b10 %
1'
b10 +
#22960000000
0!
0'
#22970000000
1!
b11 %
1'
b11 +
#22980000000
0!
0'
#22990000000
1!
b100 %
1'
b100 +
#23000000000
1"
1(
#23010000000
0!
0"
b100 &
0'
0(
b100 ,
#23020000000
1!
b101 %
1'
b101 +
#23030000000
0!
0'
#23040000000
1!
b110 %
1'
b110 +
#23050000000
0!
0'
#23060000000
1!
b111 %
1'
b111 +
#23070000000
0!
0'
#23080000000
1!
0$
b1000 %
1'
0*
b1000 +
#23090000000
0!
0'
#23100000000
1!
b1001 %
1'
b1001 +
#23110000000
0!
0'
#23120000000
1!
b0 %
1'
b0 +
#23130000000
0!
0'
#23140000000
1!
1$
b1 %
1'
1*
b1 +
#23150000000
0!
0'
#23160000000
1!
b10 %
1'
b10 +
#23170000000
0!
0'
#23180000000
1!
b11 %
1'
b11 +
#23190000000
0!
0'
#23200000000
1!
b100 %
1'
b100 +
#23210000000
0!
0'
#23220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#23230000000
0!
0'
#23240000000
1!
0$
b110 %
1'
0*
b110 +
#23250000000
0!
0'
#23260000000
1!
b111 %
1'
b111 +
#23270000000
0!
0'
#23280000000
1!
b1000 %
1'
b1000 +
#23290000000
0!
0'
#23300000000
1!
b1001 %
1'
b1001 +
#23310000000
0!
0'
#23320000000
1!
b0 %
1'
b0 +
#23330000000
0!
0'
#23340000000
1!
1$
b1 %
1'
1*
b1 +
#23350000000
0!
0'
#23360000000
1!
b10 %
1'
b10 +
#23370000000
0!
0'
#23380000000
1!
b11 %
1'
b11 +
#23390000000
0!
0'
#23400000000
1!
b100 %
1'
b100 +
#23410000000
0!
0'
#23420000000
1!
b101 %
1'
b101 +
#23430000000
1"
1(
#23440000000
0!
0"
b100 &
0'
0(
b100 ,
#23450000000
1!
b110 %
1'
b110 +
#23460000000
0!
0'
#23470000000
1!
b111 %
1'
b111 +
#23480000000
0!
0'
#23490000000
1!
0$
b1000 %
1'
0*
b1000 +
#23500000000
0!
0'
#23510000000
1!
b1001 %
1'
b1001 +
#23520000000
0!
0'
#23530000000
1!
b0 %
1'
b0 +
#23540000000
0!
0'
#23550000000
1!
1$
b1 %
1'
1*
b1 +
#23560000000
0!
0'
#23570000000
1!
b10 %
1'
b10 +
#23580000000
0!
0'
#23590000000
1!
b11 %
1'
b11 +
#23600000000
0!
0'
#23610000000
1!
b100 %
1'
b100 +
#23620000000
0!
0'
#23630000000
1!
b101 %
1'
b101 +
#23640000000
0!
0'
#23650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#23660000000
0!
0'
#23670000000
1!
b111 %
1'
b111 +
#23680000000
0!
0'
#23690000000
1!
b1000 %
1'
b1000 +
#23700000000
0!
0'
#23710000000
1!
b1001 %
1'
b1001 +
#23720000000
0!
0'
#23730000000
1!
b0 %
1'
b0 +
#23740000000
0!
0'
#23750000000
1!
1$
b1 %
1'
1*
b1 +
#23760000000
0!
0'
#23770000000
1!
b10 %
1'
b10 +
#23780000000
0!
0'
#23790000000
1!
b11 %
1'
b11 +
#23800000000
0!
0'
#23810000000
1!
b100 %
1'
b100 +
#23820000000
0!
0'
#23830000000
1!
b101 %
1'
b101 +
#23840000000
0!
0'
#23850000000
1!
0$
b110 %
1'
0*
b110 +
#23860000000
1"
1(
#23870000000
0!
0"
b100 &
0'
0(
b100 ,
#23880000000
1!
1$
b111 %
1'
1*
b111 +
#23890000000
0!
0'
#23900000000
1!
0$
b1000 %
1'
0*
b1000 +
#23910000000
0!
0'
#23920000000
1!
b1001 %
1'
b1001 +
#23930000000
0!
0'
#23940000000
1!
b0 %
1'
b0 +
#23950000000
0!
0'
#23960000000
1!
1$
b1 %
1'
1*
b1 +
#23970000000
0!
0'
#23980000000
1!
b10 %
1'
b10 +
#23990000000
0!
0'
#24000000000
1!
b11 %
1'
b11 +
#24010000000
0!
0'
#24020000000
1!
b100 %
1'
b100 +
#24030000000
0!
0'
#24040000000
1!
b101 %
1'
b101 +
#24050000000
0!
0'
#24060000000
1!
b110 %
1'
b110 +
#24070000000
0!
0'
#24080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#24090000000
0!
0'
#24100000000
1!
b1000 %
1'
b1000 +
#24110000000
0!
0'
#24120000000
1!
b1001 %
1'
b1001 +
#24130000000
0!
0'
#24140000000
1!
b0 %
1'
b0 +
#24150000000
0!
0'
#24160000000
1!
1$
b1 %
1'
1*
b1 +
#24170000000
0!
0'
#24180000000
1!
b10 %
1'
b10 +
#24190000000
0!
0'
#24200000000
1!
b11 %
1'
b11 +
#24210000000
0!
0'
#24220000000
1!
b100 %
1'
b100 +
#24230000000
0!
0'
#24240000000
1!
b101 %
1'
b101 +
#24250000000
0!
0'
#24260000000
1!
0$
b110 %
1'
0*
b110 +
#24270000000
0!
0'
#24280000000
1!
b111 %
1'
b111 +
#24290000000
1"
1(
#24300000000
0!
0"
b100 &
0'
0(
b100 ,
#24310000000
1!
b1000 %
1'
b1000 +
#24320000000
0!
0'
#24330000000
1!
b1001 %
1'
b1001 +
#24340000000
0!
0'
#24350000000
1!
b0 %
1'
b0 +
#24360000000
0!
0'
#24370000000
1!
1$
b1 %
1'
1*
b1 +
#24380000000
0!
0'
#24390000000
1!
b10 %
1'
b10 +
#24400000000
0!
0'
#24410000000
1!
b11 %
1'
b11 +
#24420000000
0!
0'
#24430000000
1!
b100 %
1'
b100 +
#24440000000
0!
0'
#24450000000
1!
b101 %
1'
b101 +
#24460000000
0!
0'
#24470000000
1!
b110 %
1'
b110 +
#24480000000
0!
0'
#24490000000
1!
b111 %
1'
b111 +
#24500000000
0!
0'
#24510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#24520000000
0!
0'
#24530000000
1!
b1001 %
1'
b1001 +
#24540000000
0!
0'
#24550000000
1!
b0 %
1'
b0 +
#24560000000
0!
0'
#24570000000
1!
1$
b1 %
1'
1*
b1 +
#24580000000
0!
0'
#24590000000
1!
b10 %
1'
b10 +
#24600000000
0!
0'
#24610000000
1!
b11 %
1'
b11 +
#24620000000
0!
0'
#24630000000
1!
b100 %
1'
b100 +
#24640000000
0!
0'
#24650000000
1!
b101 %
1'
b101 +
#24660000000
0!
0'
#24670000000
1!
0$
b110 %
1'
0*
b110 +
#24680000000
0!
0'
#24690000000
1!
b111 %
1'
b111 +
#24700000000
0!
0'
#24710000000
1!
b1000 %
1'
b1000 +
#24720000000
1"
1(
#24730000000
0!
0"
b100 &
0'
0(
b100 ,
#24740000000
1!
b1001 %
1'
b1001 +
#24750000000
0!
0'
#24760000000
1!
b0 %
1'
b0 +
#24770000000
0!
0'
#24780000000
1!
1$
b1 %
1'
1*
b1 +
#24790000000
0!
0'
#24800000000
1!
b10 %
1'
b10 +
#24810000000
0!
0'
#24820000000
1!
b11 %
1'
b11 +
#24830000000
0!
0'
#24840000000
1!
b100 %
1'
b100 +
#24850000000
0!
0'
#24860000000
1!
b101 %
1'
b101 +
#24870000000
0!
0'
#24880000000
1!
b110 %
1'
b110 +
#24890000000
0!
0'
#24900000000
1!
b111 %
1'
b111 +
#24910000000
0!
0'
#24920000000
1!
0$
b1000 %
1'
0*
b1000 +
#24930000000
0!
0'
#24940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#24950000000
0!
0'
#24960000000
1!
b0 %
1'
b0 +
#24970000000
0!
0'
#24980000000
1!
1$
b1 %
1'
1*
b1 +
#24990000000
0!
0'
#25000000000
1!
b10 %
1'
b10 +
#25010000000
0!
0'
#25020000000
1!
b11 %
1'
b11 +
#25030000000
0!
0'
#25040000000
1!
b100 %
1'
b100 +
#25050000000
0!
0'
#25060000000
1!
b101 %
1'
b101 +
#25070000000
0!
0'
#25080000000
1!
0$
b110 %
1'
0*
b110 +
#25090000000
0!
0'
#25100000000
1!
b111 %
1'
b111 +
#25110000000
0!
0'
#25120000000
1!
b1000 %
1'
b1000 +
#25130000000
0!
0'
#25140000000
1!
b1001 %
1'
b1001 +
#25150000000
1"
1(
#25160000000
0!
0"
b100 &
0'
0(
b100 ,
#25170000000
1!
b0 %
1'
b0 +
#25180000000
0!
0'
#25190000000
1!
1$
b1 %
1'
1*
b1 +
#25200000000
0!
0'
#25210000000
1!
b10 %
1'
b10 +
#25220000000
0!
0'
#25230000000
1!
b11 %
1'
b11 +
#25240000000
0!
0'
#25250000000
1!
b100 %
1'
b100 +
#25260000000
0!
0'
#25270000000
1!
b101 %
1'
b101 +
#25280000000
0!
0'
#25290000000
1!
b110 %
1'
b110 +
#25300000000
0!
0'
#25310000000
1!
b111 %
1'
b111 +
#25320000000
0!
0'
#25330000000
1!
0$
b1000 %
1'
0*
b1000 +
#25340000000
0!
0'
#25350000000
1!
b1001 %
1'
b1001 +
#25360000000
0!
0'
#25370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#25380000000
0!
0'
#25390000000
1!
1$
b1 %
1'
1*
b1 +
#25400000000
0!
0'
#25410000000
1!
b10 %
1'
b10 +
#25420000000
0!
0'
#25430000000
1!
b11 %
1'
b11 +
#25440000000
0!
0'
#25450000000
1!
b100 %
1'
b100 +
#25460000000
0!
0'
#25470000000
1!
b101 %
1'
b101 +
#25480000000
0!
0'
#25490000000
1!
0$
b110 %
1'
0*
b110 +
#25500000000
0!
0'
#25510000000
1!
b111 %
1'
b111 +
#25520000000
0!
0'
#25530000000
1!
b1000 %
1'
b1000 +
#25540000000
0!
0'
#25550000000
1!
b1001 %
1'
b1001 +
#25560000000
0!
0'
#25570000000
1!
b0 %
1'
b0 +
#25580000000
1"
1(
#25590000000
0!
0"
b100 &
0'
0(
b100 ,
#25600000000
1!
1$
b1 %
1'
1*
b1 +
#25610000000
0!
0'
#25620000000
1!
b10 %
1'
b10 +
#25630000000
0!
0'
#25640000000
1!
b11 %
1'
b11 +
#25650000000
0!
0'
#25660000000
1!
b100 %
1'
b100 +
#25670000000
0!
0'
#25680000000
1!
b101 %
1'
b101 +
#25690000000
0!
0'
#25700000000
1!
b110 %
1'
b110 +
#25710000000
0!
0'
#25720000000
1!
b111 %
1'
b111 +
#25730000000
0!
0'
#25740000000
1!
0$
b1000 %
1'
0*
b1000 +
#25750000000
0!
0'
#25760000000
1!
b1001 %
1'
b1001 +
#25770000000
0!
0'
#25780000000
1!
b0 %
1'
b0 +
#25790000000
0!
0'
#25800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#25810000000
0!
0'
#25820000000
1!
b10 %
1'
b10 +
#25830000000
0!
0'
#25840000000
1!
b11 %
1'
b11 +
#25850000000
0!
0'
#25860000000
1!
b100 %
1'
b100 +
#25870000000
0!
0'
#25880000000
1!
b101 %
1'
b101 +
#25890000000
0!
0'
#25900000000
1!
0$
b110 %
1'
0*
b110 +
#25910000000
0!
0'
#25920000000
1!
b111 %
1'
b111 +
#25930000000
0!
0'
#25940000000
1!
b1000 %
1'
b1000 +
#25950000000
0!
0'
#25960000000
1!
b1001 %
1'
b1001 +
#25970000000
0!
0'
#25980000000
1!
b0 %
1'
b0 +
#25990000000
0!
0'
#26000000000
1!
1$
b1 %
1'
1*
b1 +
#26010000000
1"
1(
#26020000000
0!
0"
b100 &
0'
0(
b100 ,
#26030000000
1!
b10 %
1'
b10 +
#26040000000
0!
0'
#26050000000
1!
b11 %
1'
b11 +
#26060000000
0!
0'
#26070000000
1!
b100 %
1'
b100 +
#26080000000
0!
0'
#26090000000
1!
b101 %
1'
b101 +
#26100000000
0!
0'
#26110000000
1!
b110 %
1'
b110 +
#26120000000
0!
0'
#26130000000
1!
b111 %
1'
b111 +
#26140000000
0!
0'
#26150000000
1!
0$
b1000 %
1'
0*
b1000 +
#26160000000
0!
0'
#26170000000
1!
b1001 %
1'
b1001 +
#26180000000
0!
0'
#26190000000
1!
b0 %
1'
b0 +
#26200000000
0!
0'
#26210000000
1!
1$
b1 %
1'
1*
b1 +
#26220000000
0!
0'
#26230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#26240000000
0!
0'
#26250000000
1!
b11 %
1'
b11 +
#26260000000
0!
0'
#26270000000
1!
b100 %
1'
b100 +
#26280000000
0!
0'
#26290000000
1!
b101 %
1'
b101 +
#26300000000
0!
0'
#26310000000
1!
0$
b110 %
1'
0*
b110 +
#26320000000
0!
0'
#26330000000
1!
b111 %
1'
b111 +
#26340000000
0!
0'
#26350000000
1!
b1000 %
1'
b1000 +
#26360000000
0!
0'
#26370000000
1!
b1001 %
1'
b1001 +
#26380000000
0!
0'
#26390000000
1!
b0 %
1'
b0 +
#26400000000
0!
0'
#26410000000
1!
1$
b1 %
1'
1*
b1 +
#26420000000
0!
0'
#26430000000
1!
b10 %
1'
b10 +
#26440000000
1"
1(
#26450000000
0!
0"
b100 &
0'
0(
b100 ,
#26460000000
1!
b11 %
1'
b11 +
#26470000000
0!
0'
#26480000000
1!
b100 %
1'
b100 +
#26490000000
0!
0'
#26500000000
1!
b101 %
1'
b101 +
#26510000000
0!
0'
#26520000000
1!
b110 %
1'
b110 +
#26530000000
0!
0'
#26540000000
1!
b111 %
1'
b111 +
#26550000000
0!
0'
#26560000000
1!
0$
b1000 %
1'
0*
b1000 +
#26570000000
0!
0'
#26580000000
1!
b1001 %
1'
b1001 +
#26590000000
0!
0'
#26600000000
1!
b0 %
1'
b0 +
#26610000000
0!
0'
#26620000000
1!
1$
b1 %
1'
1*
b1 +
#26630000000
0!
0'
#26640000000
1!
b10 %
1'
b10 +
#26650000000
0!
0'
#26660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#26670000000
0!
0'
#26680000000
1!
b100 %
1'
b100 +
#26690000000
0!
0'
#26700000000
1!
b101 %
1'
b101 +
#26710000000
0!
0'
#26720000000
1!
0$
b110 %
1'
0*
b110 +
#26730000000
0!
0'
#26740000000
1!
b111 %
1'
b111 +
#26750000000
0!
0'
#26760000000
1!
b1000 %
1'
b1000 +
#26770000000
0!
0'
#26780000000
1!
b1001 %
1'
b1001 +
#26790000000
0!
0'
#26800000000
1!
b0 %
1'
b0 +
#26810000000
0!
0'
#26820000000
1!
1$
b1 %
1'
1*
b1 +
#26830000000
0!
0'
#26840000000
1!
b10 %
1'
b10 +
#26850000000
0!
0'
#26860000000
1!
b11 %
1'
b11 +
#26870000000
1"
1(
#26880000000
0!
0"
b100 &
0'
0(
b100 ,
#26890000000
1!
b100 %
1'
b100 +
#26900000000
0!
0'
#26910000000
1!
b101 %
1'
b101 +
#26920000000
0!
0'
#26930000000
1!
b110 %
1'
b110 +
#26940000000
0!
0'
#26950000000
1!
b111 %
1'
b111 +
#26960000000
0!
0'
#26970000000
1!
0$
b1000 %
1'
0*
b1000 +
#26980000000
0!
0'
#26990000000
1!
b1001 %
1'
b1001 +
#27000000000
0!
0'
#27010000000
1!
b0 %
1'
b0 +
#27020000000
0!
0'
#27030000000
1!
1$
b1 %
1'
1*
b1 +
#27040000000
0!
0'
#27050000000
1!
b10 %
1'
b10 +
#27060000000
0!
0'
#27070000000
1!
b11 %
1'
b11 +
#27080000000
0!
0'
#27090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#27100000000
0!
0'
#27110000000
1!
b101 %
1'
b101 +
#27120000000
0!
0'
#27130000000
1!
0$
b110 %
1'
0*
b110 +
#27140000000
0!
0'
#27150000000
1!
b111 %
1'
b111 +
#27160000000
0!
0'
#27170000000
1!
b1000 %
1'
b1000 +
#27180000000
0!
0'
#27190000000
1!
b1001 %
1'
b1001 +
#27200000000
0!
0'
#27210000000
1!
b0 %
1'
b0 +
#27220000000
0!
0'
#27230000000
1!
1$
b1 %
1'
1*
b1 +
#27240000000
0!
0'
#27250000000
1!
b10 %
1'
b10 +
#27260000000
0!
0'
#27270000000
1!
b11 %
1'
b11 +
#27280000000
0!
0'
#27290000000
1!
b100 %
1'
b100 +
#27300000000
1"
1(
#27310000000
0!
0"
b100 &
0'
0(
b100 ,
#27320000000
1!
b101 %
1'
b101 +
#27330000000
0!
0'
#27340000000
1!
b110 %
1'
b110 +
#27350000000
0!
0'
#27360000000
1!
b111 %
1'
b111 +
#27370000000
0!
0'
#27380000000
1!
0$
b1000 %
1'
0*
b1000 +
#27390000000
0!
0'
#27400000000
1!
b1001 %
1'
b1001 +
#27410000000
0!
0'
#27420000000
1!
b0 %
1'
b0 +
#27430000000
0!
0'
#27440000000
1!
1$
b1 %
1'
1*
b1 +
#27450000000
0!
0'
#27460000000
1!
b10 %
1'
b10 +
#27470000000
0!
0'
#27480000000
1!
b11 %
1'
b11 +
#27490000000
0!
0'
#27500000000
1!
b100 %
1'
b100 +
#27510000000
0!
0'
#27520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#27530000000
0!
0'
#27540000000
1!
0$
b110 %
1'
0*
b110 +
#27550000000
0!
0'
#27560000000
1!
b111 %
1'
b111 +
#27570000000
0!
0'
#27580000000
1!
b1000 %
1'
b1000 +
#27590000000
0!
0'
#27600000000
1!
b1001 %
1'
b1001 +
#27610000000
0!
0'
#27620000000
1!
b0 %
1'
b0 +
#27630000000
0!
0'
#27640000000
1!
1$
b1 %
1'
1*
b1 +
#27650000000
0!
0'
#27660000000
1!
b10 %
1'
b10 +
#27670000000
0!
0'
#27680000000
1!
b11 %
1'
b11 +
#27690000000
0!
0'
#27700000000
1!
b100 %
1'
b100 +
#27710000000
0!
0'
#27720000000
1!
b101 %
1'
b101 +
#27730000000
1"
1(
#27740000000
0!
0"
b100 &
0'
0(
b100 ,
#27750000000
1!
b110 %
1'
b110 +
#27760000000
0!
0'
#27770000000
1!
b111 %
1'
b111 +
#27780000000
0!
0'
#27790000000
1!
0$
b1000 %
1'
0*
b1000 +
#27800000000
0!
0'
#27810000000
1!
b1001 %
1'
b1001 +
#27820000000
0!
0'
#27830000000
1!
b0 %
1'
b0 +
#27840000000
0!
0'
#27850000000
1!
1$
b1 %
1'
1*
b1 +
#27860000000
0!
0'
#27870000000
1!
b10 %
1'
b10 +
#27880000000
0!
0'
#27890000000
1!
b11 %
1'
b11 +
#27900000000
0!
0'
#27910000000
1!
b100 %
1'
b100 +
#27920000000
0!
0'
#27930000000
1!
b101 %
1'
b101 +
#27940000000
0!
0'
#27950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#27960000000
0!
0'
#27970000000
1!
b111 %
1'
b111 +
#27980000000
0!
0'
#27990000000
1!
b1000 %
1'
b1000 +
#28000000000
0!
0'
#28010000000
1!
b1001 %
1'
b1001 +
#28020000000
0!
0'
#28030000000
1!
b0 %
1'
b0 +
#28040000000
0!
0'
#28050000000
1!
1$
b1 %
1'
1*
b1 +
#28060000000
0!
0'
#28070000000
1!
b10 %
1'
b10 +
#28080000000
0!
0'
#28090000000
1!
b11 %
1'
b11 +
#28100000000
0!
0'
#28110000000
1!
b100 %
1'
b100 +
#28120000000
0!
0'
#28130000000
1!
b101 %
1'
b101 +
#28140000000
0!
0'
#28150000000
1!
0$
b110 %
1'
0*
b110 +
#28160000000
1"
1(
#28170000000
0!
0"
b100 &
0'
0(
b100 ,
#28180000000
1!
1$
b111 %
1'
1*
b111 +
#28190000000
0!
0'
#28200000000
1!
0$
b1000 %
1'
0*
b1000 +
#28210000000
0!
0'
#28220000000
1!
b1001 %
1'
b1001 +
#28230000000
0!
0'
#28240000000
1!
b0 %
1'
b0 +
#28250000000
0!
0'
#28260000000
1!
1$
b1 %
1'
1*
b1 +
#28270000000
0!
0'
#28280000000
1!
b10 %
1'
b10 +
#28290000000
0!
0'
#28300000000
1!
b11 %
1'
b11 +
#28310000000
0!
0'
#28320000000
1!
b100 %
1'
b100 +
#28330000000
0!
0'
#28340000000
1!
b101 %
1'
b101 +
#28350000000
0!
0'
#28360000000
1!
b110 %
1'
b110 +
#28370000000
0!
0'
#28380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#28390000000
0!
0'
#28400000000
1!
b1000 %
1'
b1000 +
#28410000000
0!
0'
#28420000000
1!
b1001 %
1'
b1001 +
#28430000000
0!
0'
#28440000000
1!
b0 %
1'
b0 +
#28450000000
0!
0'
#28460000000
1!
1$
b1 %
1'
1*
b1 +
#28470000000
0!
0'
#28480000000
1!
b10 %
1'
b10 +
#28490000000
0!
0'
#28500000000
1!
b11 %
1'
b11 +
#28510000000
0!
0'
#28520000000
1!
b100 %
1'
b100 +
#28530000000
0!
0'
#28540000000
1!
b101 %
1'
b101 +
#28550000000
0!
0'
#28560000000
1!
0$
b110 %
1'
0*
b110 +
#28570000000
0!
0'
#28580000000
1!
b111 %
1'
b111 +
#28590000000
1"
1(
#28600000000
0!
0"
b100 &
0'
0(
b100 ,
#28610000000
1!
b1000 %
1'
b1000 +
#28620000000
0!
0'
#28630000000
1!
b1001 %
1'
b1001 +
#28640000000
0!
0'
#28650000000
1!
b0 %
1'
b0 +
#28660000000
0!
0'
#28670000000
1!
1$
b1 %
1'
1*
b1 +
#28680000000
0!
0'
#28690000000
1!
b10 %
1'
b10 +
#28700000000
0!
0'
#28710000000
1!
b11 %
1'
b11 +
#28720000000
0!
0'
#28730000000
1!
b100 %
1'
b100 +
#28740000000
0!
0'
#28750000000
1!
b101 %
1'
b101 +
#28760000000
0!
0'
#28770000000
1!
b110 %
1'
b110 +
#28780000000
0!
0'
#28790000000
1!
b111 %
1'
b111 +
#28800000000
0!
0'
#28810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#28820000000
0!
0'
#28830000000
1!
b1001 %
1'
b1001 +
#28840000000
0!
0'
#28850000000
1!
b0 %
1'
b0 +
#28860000000
0!
0'
#28870000000
1!
1$
b1 %
1'
1*
b1 +
#28880000000
0!
0'
#28890000000
1!
b10 %
1'
b10 +
#28900000000
0!
0'
#28910000000
1!
b11 %
1'
b11 +
#28920000000
0!
0'
#28930000000
1!
b100 %
1'
b100 +
#28940000000
0!
0'
#28950000000
1!
b101 %
1'
b101 +
#28960000000
0!
0'
#28970000000
1!
0$
b110 %
1'
0*
b110 +
#28980000000
0!
0'
#28990000000
1!
b111 %
1'
b111 +
#29000000000
0!
0'
#29010000000
1!
b1000 %
1'
b1000 +
#29020000000
1"
1(
#29030000000
0!
0"
b100 &
0'
0(
b100 ,
#29040000000
1!
b1001 %
1'
b1001 +
#29050000000
0!
0'
#29060000000
1!
b0 %
1'
b0 +
#29070000000
0!
0'
#29080000000
1!
1$
b1 %
1'
1*
b1 +
#29090000000
0!
0'
#29100000000
1!
b10 %
1'
b10 +
#29110000000
0!
0'
#29120000000
1!
b11 %
1'
b11 +
#29130000000
0!
0'
#29140000000
1!
b100 %
1'
b100 +
#29150000000
0!
0'
#29160000000
1!
b101 %
1'
b101 +
#29170000000
0!
0'
#29180000000
1!
b110 %
1'
b110 +
#29190000000
0!
0'
#29200000000
1!
b111 %
1'
b111 +
#29210000000
0!
0'
#29220000000
1!
0$
b1000 %
1'
0*
b1000 +
#29230000000
0!
0'
#29240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#29250000000
0!
0'
#29260000000
1!
b0 %
1'
b0 +
#29270000000
0!
0'
#29280000000
1!
1$
b1 %
1'
1*
b1 +
#29290000000
0!
0'
#29300000000
1!
b10 %
1'
b10 +
#29310000000
0!
0'
#29320000000
1!
b11 %
1'
b11 +
#29330000000
0!
0'
#29340000000
1!
b100 %
1'
b100 +
#29350000000
0!
0'
#29360000000
1!
b101 %
1'
b101 +
#29370000000
0!
0'
#29380000000
1!
0$
b110 %
1'
0*
b110 +
#29390000000
0!
0'
#29400000000
1!
b111 %
1'
b111 +
#29410000000
0!
0'
#29420000000
1!
b1000 %
1'
b1000 +
#29430000000
0!
0'
#29440000000
1!
b1001 %
1'
b1001 +
#29450000000
1"
1(
#29460000000
0!
0"
b100 &
0'
0(
b100 ,
#29470000000
1!
b0 %
1'
b0 +
#29480000000
0!
0'
#29490000000
1!
1$
b1 %
1'
1*
b1 +
#29500000000
0!
0'
#29510000000
1!
b10 %
1'
b10 +
#29520000000
0!
0'
#29530000000
1!
b11 %
1'
b11 +
#29540000000
0!
0'
#29550000000
1!
b100 %
1'
b100 +
#29560000000
0!
0'
#29570000000
1!
b101 %
1'
b101 +
#29580000000
0!
0'
#29590000000
1!
b110 %
1'
b110 +
#29600000000
0!
0'
#29610000000
1!
b111 %
1'
b111 +
#29620000000
0!
0'
#29630000000
1!
0$
b1000 %
1'
0*
b1000 +
#29640000000
0!
0'
#29650000000
1!
b1001 %
1'
b1001 +
#29660000000
0!
0'
#29670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#29680000000
0!
0'
#29690000000
1!
1$
b1 %
1'
1*
b1 +
#29700000000
0!
0'
#29710000000
1!
b10 %
1'
b10 +
#29720000000
0!
0'
#29730000000
1!
b11 %
1'
b11 +
#29740000000
0!
0'
#29750000000
1!
b100 %
1'
b100 +
#29760000000
0!
0'
#29770000000
1!
b101 %
1'
b101 +
#29780000000
0!
0'
#29790000000
1!
0$
b110 %
1'
0*
b110 +
#29800000000
0!
0'
#29810000000
1!
b111 %
1'
b111 +
#29820000000
0!
0'
#29830000000
1!
b1000 %
1'
b1000 +
#29840000000
0!
0'
#29850000000
1!
b1001 %
1'
b1001 +
#29860000000
0!
0'
#29870000000
1!
b0 %
1'
b0 +
#29880000000
1"
1(
#29890000000
0!
0"
b100 &
0'
0(
b100 ,
#29900000000
1!
1$
b1 %
1'
1*
b1 +
#29910000000
0!
0'
#29920000000
1!
b10 %
1'
b10 +
#29930000000
0!
0'
#29940000000
1!
b11 %
1'
b11 +
#29950000000
0!
0'
#29960000000
1!
b100 %
1'
b100 +
#29970000000
0!
0'
#29980000000
1!
b101 %
1'
b101 +
#29990000000
0!
0'
#30000000000
1!
b110 %
1'
b110 +
#30010000000
0!
0'
#30020000000
1!
b111 %
1'
b111 +
#30030000000
0!
0'
#30040000000
1!
0$
b1000 %
1'
0*
b1000 +
#30050000000
0!
0'
#30060000000
1!
b1001 %
1'
b1001 +
#30070000000
0!
0'
#30080000000
1!
b0 %
1'
b0 +
#30090000000
0!
0'
#30100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#30110000000
0!
0'
#30120000000
1!
b10 %
1'
b10 +
#30130000000
0!
0'
#30140000000
1!
b11 %
1'
b11 +
#30150000000
0!
0'
#30160000000
1!
b100 %
1'
b100 +
#30170000000
0!
0'
#30180000000
1!
b101 %
1'
b101 +
#30190000000
0!
0'
#30200000000
1!
0$
b110 %
1'
0*
b110 +
#30210000000
0!
0'
#30220000000
1!
b111 %
1'
b111 +
#30230000000
0!
0'
#30240000000
1!
b1000 %
1'
b1000 +
#30250000000
0!
0'
#30260000000
1!
b1001 %
1'
b1001 +
#30270000000
0!
0'
#30280000000
1!
b0 %
1'
b0 +
#30290000000
0!
0'
#30300000000
1!
1$
b1 %
1'
1*
b1 +
#30310000000
1"
1(
#30320000000
0!
0"
b100 &
0'
0(
b100 ,
#30330000000
1!
b10 %
1'
b10 +
#30340000000
0!
0'
#30350000000
1!
b11 %
1'
b11 +
#30360000000
0!
0'
#30370000000
1!
b100 %
1'
b100 +
#30380000000
0!
0'
#30390000000
1!
b101 %
1'
b101 +
#30400000000
0!
0'
#30410000000
1!
b110 %
1'
b110 +
#30420000000
0!
0'
#30430000000
1!
b111 %
1'
b111 +
#30440000000
0!
0'
#30450000000
1!
0$
b1000 %
1'
0*
b1000 +
#30460000000
0!
0'
#30470000000
1!
b1001 %
1'
b1001 +
#30480000000
0!
0'
#30490000000
1!
b0 %
1'
b0 +
#30500000000
0!
0'
#30510000000
1!
1$
b1 %
1'
1*
b1 +
#30520000000
0!
0'
#30530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#30540000000
0!
0'
#30550000000
1!
b11 %
1'
b11 +
#30560000000
0!
0'
#30570000000
1!
b100 %
1'
b100 +
#30580000000
0!
0'
#30590000000
1!
b101 %
1'
b101 +
#30600000000
0!
0'
#30610000000
1!
0$
b110 %
1'
0*
b110 +
#30620000000
0!
0'
#30630000000
1!
b111 %
1'
b111 +
#30640000000
0!
0'
#30650000000
1!
b1000 %
1'
b1000 +
#30660000000
0!
0'
#30670000000
1!
b1001 %
1'
b1001 +
#30680000000
0!
0'
#30690000000
1!
b0 %
1'
b0 +
#30700000000
0!
0'
#30710000000
1!
1$
b1 %
1'
1*
b1 +
#30720000000
0!
0'
#30730000000
1!
b10 %
1'
b10 +
#30740000000
1"
1(
#30750000000
0!
0"
b100 &
0'
0(
b100 ,
#30760000000
1!
b11 %
1'
b11 +
#30770000000
0!
0'
#30780000000
1!
b100 %
1'
b100 +
#30790000000
0!
0'
#30800000000
1!
b101 %
1'
b101 +
#30810000000
0!
0'
#30820000000
1!
b110 %
1'
b110 +
#30830000000
0!
0'
#30840000000
1!
b111 %
1'
b111 +
#30850000000
0!
0'
#30860000000
1!
0$
b1000 %
1'
0*
b1000 +
#30870000000
0!
0'
#30880000000
1!
b1001 %
1'
b1001 +
#30890000000
0!
0'
#30900000000
1!
b0 %
1'
b0 +
#30910000000
0!
0'
#30920000000
1!
1$
b1 %
1'
1*
b1 +
#30930000000
0!
0'
#30940000000
1!
b10 %
1'
b10 +
#30950000000
0!
0'
#30960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#30970000000
0!
0'
#30980000000
1!
b100 %
1'
b100 +
#30990000000
0!
0'
#31000000000
1!
b101 %
1'
b101 +
#31010000000
0!
0'
#31020000000
1!
0$
b110 %
1'
0*
b110 +
#31030000000
0!
0'
#31040000000
1!
b111 %
1'
b111 +
#31050000000
0!
0'
#31060000000
1!
b1000 %
1'
b1000 +
#31070000000
0!
0'
#31080000000
1!
b1001 %
1'
b1001 +
#31090000000
0!
0'
#31100000000
1!
b0 %
1'
b0 +
#31110000000
0!
0'
#31120000000
1!
1$
b1 %
1'
1*
b1 +
#31130000000
0!
0'
#31140000000
1!
b10 %
1'
b10 +
#31150000000
0!
0'
#31160000000
1!
b11 %
1'
b11 +
#31170000000
1"
1(
#31180000000
0!
0"
b100 &
0'
0(
b100 ,
#31190000000
1!
b100 %
1'
b100 +
#31200000000
0!
0'
#31210000000
1!
b101 %
1'
b101 +
#31220000000
0!
0'
#31230000000
1!
b110 %
1'
b110 +
#31240000000
0!
0'
#31250000000
1!
b111 %
1'
b111 +
#31260000000
0!
0'
#31270000000
1!
0$
b1000 %
1'
0*
b1000 +
#31280000000
0!
0'
#31290000000
1!
b1001 %
1'
b1001 +
#31300000000
0!
0'
#31310000000
1!
b0 %
1'
b0 +
#31320000000
0!
0'
#31330000000
1!
1$
b1 %
1'
1*
b1 +
#31340000000
0!
0'
#31350000000
1!
b10 %
1'
b10 +
#31360000000
0!
0'
#31370000000
1!
b11 %
1'
b11 +
#31380000000
0!
0'
#31390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#31400000000
0!
0'
#31410000000
1!
b101 %
1'
b101 +
#31420000000
0!
0'
#31430000000
1!
0$
b110 %
1'
0*
b110 +
#31440000000
0!
0'
#31450000000
1!
b111 %
1'
b111 +
#31460000000
0!
0'
#31470000000
1!
b1000 %
1'
b1000 +
#31480000000
0!
0'
#31490000000
1!
b1001 %
1'
b1001 +
#31500000000
0!
0'
#31510000000
1!
b0 %
1'
b0 +
#31520000000
0!
0'
#31530000000
1!
1$
b1 %
1'
1*
b1 +
#31540000000
0!
0'
#31550000000
1!
b10 %
1'
b10 +
#31560000000
0!
0'
#31570000000
1!
b11 %
1'
b11 +
#31580000000
0!
0'
#31590000000
1!
b100 %
1'
b100 +
#31600000000
1"
1(
#31610000000
0!
0"
b100 &
0'
0(
b100 ,
#31620000000
1!
b101 %
1'
b101 +
#31630000000
0!
0'
#31640000000
1!
b110 %
1'
b110 +
#31650000000
0!
0'
#31660000000
1!
b111 %
1'
b111 +
#31670000000
0!
0'
#31680000000
1!
0$
b1000 %
1'
0*
b1000 +
#31690000000
0!
0'
#31700000000
1!
b1001 %
1'
b1001 +
#31710000000
0!
0'
#31720000000
1!
b0 %
1'
b0 +
#31730000000
0!
0'
#31740000000
1!
1$
b1 %
1'
1*
b1 +
#31750000000
0!
0'
#31760000000
1!
b10 %
1'
b10 +
#31770000000
0!
0'
#31780000000
1!
b11 %
1'
b11 +
#31790000000
0!
0'
#31800000000
1!
b100 %
1'
b100 +
#31810000000
0!
0'
#31820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#31830000000
0!
0'
#31840000000
1!
0$
b110 %
1'
0*
b110 +
#31850000000
0!
0'
#31860000000
1!
b111 %
1'
b111 +
#31870000000
0!
0'
#31880000000
1!
b1000 %
1'
b1000 +
#31890000000
0!
0'
#31900000000
1!
b1001 %
1'
b1001 +
#31910000000
0!
0'
#31920000000
1!
b0 %
1'
b0 +
#31930000000
0!
0'
#31940000000
1!
1$
b1 %
1'
1*
b1 +
#31950000000
0!
0'
#31960000000
1!
b10 %
1'
b10 +
#31970000000
0!
0'
#31980000000
1!
b11 %
1'
b11 +
#31990000000
0!
0'
#32000000000
1!
b100 %
1'
b100 +
#32010000000
0!
0'
#32020000000
1!
b101 %
1'
b101 +
#32030000000
1"
1(
#32040000000
0!
0"
b100 &
0'
0(
b100 ,
#32050000000
1!
b110 %
1'
b110 +
#32060000000
0!
0'
#32070000000
1!
b111 %
1'
b111 +
#32080000000
0!
0'
#32090000000
1!
0$
b1000 %
1'
0*
b1000 +
#32100000000
0!
0'
#32110000000
1!
b1001 %
1'
b1001 +
#32120000000
0!
0'
#32130000000
1!
b0 %
1'
b0 +
#32140000000
0!
0'
#32150000000
1!
1$
b1 %
1'
1*
b1 +
#32160000000
0!
0'
#32170000000
1!
b10 %
1'
b10 +
#32180000000
0!
0'
#32190000000
1!
b11 %
1'
b11 +
#32200000000
0!
0'
#32210000000
1!
b100 %
1'
b100 +
#32220000000
0!
0'
#32230000000
1!
b101 %
1'
b101 +
#32240000000
0!
0'
#32250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#32260000000
0!
0'
#32270000000
1!
b111 %
1'
b111 +
#32280000000
0!
0'
#32290000000
1!
b1000 %
1'
b1000 +
#32300000000
0!
0'
#32310000000
1!
b1001 %
1'
b1001 +
#32320000000
0!
0'
#32330000000
1!
b0 %
1'
b0 +
#32340000000
0!
0'
#32350000000
1!
1$
b1 %
1'
1*
b1 +
#32360000000
0!
0'
#32370000000
1!
b10 %
1'
b10 +
#32380000000
0!
0'
#32390000000
1!
b11 %
1'
b11 +
#32400000000
0!
0'
#32410000000
1!
b100 %
1'
b100 +
#32420000000
0!
0'
#32430000000
1!
b101 %
1'
b101 +
#32440000000
0!
0'
#32450000000
1!
0$
b110 %
1'
0*
b110 +
#32460000000
1"
1(
#32470000000
0!
0"
b100 &
0'
0(
b100 ,
#32480000000
1!
1$
b111 %
1'
1*
b111 +
#32490000000
0!
0'
#32500000000
1!
0$
b1000 %
1'
0*
b1000 +
#32510000000
0!
0'
#32520000000
1!
b1001 %
1'
b1001 +
#32530000000
0!
0'
#32540000000
1!
b0 %
1'
b0 +
#32550000000
0!
0'
#32560000000
1!
1$
b1 %
1'
1*
b1 +
#32570000000
0!
0'
#32580000000
1!
b10 %
1'
b10 +
#32590000000
0!
0'
#32600000000
1!
b11 %
1'
b11 +
#32610000000
0!
0'
#32620000000
1!
b100 %
1'
b100 +
#32630000000
0!
0'
#32640000000
1!
b101 %
1'
b101 +
#32650000000
0!
0'
#32660000000
1!
b110 %
1'
b110 +
#32670000000
0!
0'
#32680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#32690000000
0!
0'
#32700000000
1!
b1000 %
1'
b1000 +
#32710000000
0!
0'
#32720000000
1!
b1001 %
1'
b1001 +
#32730000000
0!
0'
#32740000000
1!
b0 %
1'
b0 +
#32750000000
0!
0'
#32760000000
1!
1$
b1 %
1'
1*
b1 +
#32770000000
0!
0'
#32780000000
1!
b10 %
1'
b10 +
#32790000000
0!
0'
#32800000000
1!
b11 %
1'
b11 +
#32810000000
0!
0'
#32820000000
1!
b100 %
1'
b100 +
#32830000000
0!
0'
#32840000000
1!
b101 %
1'
b101 +
#32850000000
0!
0'
#32860000000
1!
0$
b110 %
1'
0*
b110 +
#32870000000
0!
0'
#32880000000
1!
b111 %
1'
b111 +
#32890000000
1"
1(
#32900000000
0!
0"
b100 &
0'
0(
b100 ,
#32910000000
1!
b1000 %
1'
b1000 +
#32920000000
0!
0'
#32930000000
1!
b1001 %
1'
b1001 +
#32940000000
0!
0'
#32950000000
1!
b0 %
1'
b0 +
#32960000000
0!
0'
#32970000000
1!
1$
b1 %
1'
1*
b1 +
#32980000000
0!
0'
#32990000000
1!
b10 %
1'
b10 +
#33000000000
0!
0'
#33010000000
1!
b11 %
1'
b11 +
#33020000000
0!
0'
#33030000000
1!
b100 %
1'
b100 +
#33040000000
0!
0'
#33050000000
1!
b101 %
1'
b101 +
#33060000000
0!
0'
#33070000000
1!
b110 %
1'
b110 +
#33080000000
0!
0'
#33090000000
1!
b111 %
1'
b111 +
#33100000000
0!
0'
#33110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#33120000000
0!
0'
#33130000000
1!
b1001 %
1'
b1001 +
#33140000000
0!
0'
#33150000000
1!
b0 %
1'
b0 +
#33160000000
0!
0'
#33170000000
1!
1$
b1 %
1'
1*
b1 +
#33180000000
0!
0'
#33190000000
1!
b10 %
1'
b10 +
#33200000000
0!
0'
#33210000000
1!
b11 %
1'
b11 +
#33220000000
0!
0'
#33230000000
1!
b100 %
1'
b100 +
#33240000000
0!
0'
#33250000000
1!
b101 %
1'
b101 +
#33260000000
0!
0'
#33270000000
1!
0$
b110 %
1'
0*
b110 +
#33280000000
0!
0'
#33290000000
1!
b111 %
1'
b111 +
#33300000000
0!
0'
#33310000000
1!
b1000 %
1'
b1000 +
#33320000000
1"
1(
#33330000000
0!
0"
b100 &
0'
0(
b100 ,
#33340000000
1!
b1001 %
1'
b1001 +
#33350000000
0!
0'
#33360000000
1!
b0 %
1'
b0 +
#33370000000
0!
0'
#33380000000
1!
1$
b1 %
1'
1*
b1 +
#33390000000
0!
0'
#33400000000
1!
b10 %
1'
b10 +
#33410000000
0!
0'
#33420000000
1!
b11 %
1'
b11 +
#33430000000
0!
0'
#33440000000
1!
b100 %
1'
b100 +
#33450000000
0!
0'
#33460000000
1!
b101 %
1'
b101 +
#33470000000
0!
0'
#33480000000
1!
b110 %
1'
b110 +
#33490000000
0!
0'
#33500000000
1!
b111 %
1'
b111 +
#33510000000
0!
0'
#33520000000
1!
0$
b1000 %
1'
0*
b1000 +
#33530000000
0!
0'
#33540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#33550000000
0!
0'
#33560000000
1!
b0 %
1'
b0 +
#33570000000
0!
0'
#33580000000
1!
1$
b1 %
1'
1*
b1 +
#33590000000
0!
0'
#33600000000
1!
b10 %
1'
b10 +
#33610000000
0!
0'
#33620000000
1!
b11 %
1'
b11 +
#33630000000
0!
0'
#33640000000
1!
b100 %
1'
b100 +
#33650000000
0!
0'
#33660000000
1!
b101 %
1'
b101 +
#33670000000
0!
0'
#33680000000
1!
0$
b110 %
1'
0*
b110 +
#33690000000
0!
0'
#33700000000
1!
b111 %
1'
b111 +
#33710000000
0!
0'
#33720000000
1!
b1000 %
1'
b1000 +
#33730000000
0!
0'
#33740000000
1!
b1001 %
1'
b1001 +
#33750000000
1"
1(
#33760000000
0!
0"
b100 &
0'
0(
b100 ,
#33770000000
1!
b0 %
1'
b0 +
#33780000000
0!
0'
#33790000000
1!
1$
b1 %
1'
1*
b1 +
#33800000000
0!
0'
#33810000000
1!
b10 %
1'
b10 +
#33820000000
0!
0'
#33830000000
1!
b11 %
1'
b11 +
#33840000000
0!
0'
#33850000000
1!
b100 %
1'
b100 +
#33860000000
0!
0'
#33870000000
1!
b101 %
1'
b101 +
#33880000000
0!
0'
#33890000000
1!
b110 %
1'
b110 +
#33900000000
0!
0'
#33910000000
1!
b111 %
1'
b111 +
#33920000000
0!
0'
#33930000000
1!
0$
b1000 %
1'
0*
b1000 +
#33940000000
0!
0'
#33950000000
1!
b1001 %
1'
b1001 +
#33960000000
0!
0'
#33970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#33980000000
0!
0'
#33990000000
1!
1$
b1 %
1'
1*
b1 +
#34000000000
0!
0'
#34010000000
1!
b10 %
1'
b10 +
#34020000000
0!
0'
#34030000000
1!
b11 %
1'
b11 +
#34040000000
0!
0'
#34050000000
1!
b100 %
1'
b100 +
#34060000000
0!
0'
#34070000000
1!
b101 %
1'
b101 +
#34080000000
0!
0'
#34090000000
1!
0$
b110 %
1'
0*
b110 +
#34100000000
0!
0'
#34110000000
1!
b111 %
1'
b111 +
#34120000000
0!
0'
#34130000000
1!
b1000 %
1'
b1000 +
#34140000000
0!
0'
#34150000000
1!
b1001 %
1'
b1001 +
#34160000000
0!
0'
#34170000000
1!
b0 %
1'
b0 +
#34180000000
1"
1(
#34190000000
0!
0"
b100 &
0'
0(
b100 ,
#34200000000
1!
1$
b1 %
1'
1*
b1 +
#34210000000
0!
0'
#34220000000
1!
b10 %
1'
b10 +
#34230000000
0!
0'
#34240000000
1!
b11 %
1'
b11 +
#34250000000
0!
0'
#34260000000
1!
b100 %
1'
b100 +
#34270000000
0!
0'
#34280000000
1!
b101 %
1'
b101 +
#34290000000
0!
0'
#34300000000
1!
b110 %
1'
b110 +
#34310000000
0!
0'
#34320000000
1!
b111 %
1'
b111 +
#34330000000
0!
0'
#34340000000
1!
0$
b1000 %
1'
0*
b1000 +
#34350000000
0!
0'
#34360000000
1!
b1001 %
1'
b1001 +
#34370000000
0!
0'
#34380000000
1!
b0 %
1'
b0 +
#34390000000
0!
0'
#34400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#34410000000
0!
0'
#34420000000
1!
b10 %
1'
b10 +
#34430000000
0!
0'
#34440000000
1!
b11 %
1'
b11 +
#34450000000
0!
0'
#34460000000
1!
b100 %
1'
b100 +
#34470000000
0!
0'
#34480000000
1!
b101 %
1'
b101 +
#34490000000
0!
0'
#34500000000
1!
0$
b110 %
1'
0*
b110 +
#34510000000
0!
0'
#34520000000
1!
b111 %
1'
b111 +
#34530000000
0!
0'
#34540000000
1!
b1000 %
1'
b1000 +
#34550000000
0!
0'
#34560000000
1!
b1001 %
1'
b1001 +
#34570000000
0!
0'
#34580000000
1!
b0 %
1'
b0 +
#34590000000
0!
0'
#34600000000
1!
1$
b1 %
1'
1*
b1 +
#34610000000
1"
1(
#34620000000
0!
0"
b100 &
0'
0(
b100 ,
#34630000000
1!
b10 %
1'
b10 +
#34640000000
0!
0'
#34650000000
1!
b11 %
1'
b11 +
#34660000000
0!
0'
#34670000000
1!
b100 %
1'
b100 +
#34680000000
0!
0'
#34690000000
1!
b101 %
1'
b101 +
#34700000000
0!
0'
#34710000000
1!
b110 %
1'
b110 +
#34720000000
0!
0'
#34730000000
1!
b111 %
1'
b111 +
#34740000000
0!
0'
#34750000000
1!
0$
b1000 %
1'
0*
b1000 +
#34760000000
0!
0'
#34770000000
1!
b1001 %
1'
b1001 +
#34780000000
0!
0'
#34790000000
1!
b0 %
1'
b0 +
#34800000000
0!
0'
#34810000000
1!
1$
b1 %
1'
1*
b1 +
#34820000000
0!
0'
#34830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#34840000000
0!
0'
#34850000000
1!
b11 %
1'
b11 +
#34860000000
0!
0'
#34870000000
1!
b100 %
1'
b100 +
#34880000000
0!
0'
#34890000000
1!
b101 %
1'
b101 +
#34900000000
0!
0'
#34910000000
1!
0$
b110 %
1'
0*
b110 +
#34920000000
0!
0'
#34930000000
1!
b111 %
1'
b111 +
#34940000000
0!
0'
#34950000000
1!
b1000 %
1'
b1000 +
#34960000000
0!
0'
#34970000000
1!
b1001 %
1'
b1001 +
#34980000000
0!
0'
#34990000000
1!
b0 %
1'
b0 +
#35000000000
0!
0'
#35010000000
1!
1$
b1 %
1'
1*
b1 +
#35020000000
0!
0'
#35030000000
1!
b10 %
1'
b10 +
#35040000000
1"
1(
#35050000000
0!
0"
b100 &
0'
0(
b100 ,
#35060000000
1!
b11 %
1'
b11 +
#35070000000
0!
0'
#35080000000
1!
b100 %
1'
b100 +
#35090000000
0!
0'
#35100000000
1!
b101 %
1'
b101 +
#35110000000
0!
0'
#35120000000
1!
b110 %
1'
b110 +
#35130000000
0!
0'
#35140000000
1!
b111 %
1'
b111 +
#35150000000
0!
0'
#35160000000
1!
0$
b1000 %
1'
0*
b1000 +
#35170000000
0!
0'
#35180000000
1!
b1001 %
1'
b1001 +
#35190000000
0!
0'
#35200000000
1!
b0 %
1'
b0 +
#35210000000
0!
0'
#35220000000
1!
1$
b1 %
1'
1*
b1 +
#35230000000
0!
0'
#35240000000
1!
b10 %
1'
b10 +
#35250000000
0!
0'
#35260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#35270000000
0!
0'
#35280000000
1!
b100 %
1'
b100 +
#35290000000
0!
0'
#35300000000
1!
b101 %
1'
b101 +
#35310000000
0!
0'
#35320000000
1!
0$
b110 %
1'
0*
b110 +
#35330000000
0!
0'
#35340000000
1!
b111 %
1'
b111 +
#35350000000
0!
0'
#35360000000
1!
b1000 %
1'
b1000 +
#35370000000
0!
0'
#35380000000
1!
b1001 %
1'
b1001 +
#35390000000
0!
0'
#35400000000
1!
b0 %
1'
b0 +
#35410000000
0!
0'
#35420000000
1!
1$
b1 %
1'
1*
b1 +
#35430000000
0!
0'
#35440000000
1!
b10 %
1'
b10 +
#35450000000
0!
0'
#35460000000
1!
b11 %
1'
b11 +
#35470000000
1"
1(
#35480000000
0!
0"
b100 &
0'
0(
b100 ,
#35490000000
1!
b100 %
1'
b100 +
#35500000000
0!
0'
#35510000000
1!
b101 %
1'
b101 +
#35520000000
0!
0'
#35530000000
1!
b110 %
1'
b110 +
#35540000000
0!
0'
#35550000000
1!
b111 %
1'
b111 +
#35560000000
0!
0'
#35570000000
1!
0$
b1000 %
1'
0*
b1000 +
#35580000000
0!
0'
#35590000000
1!
b1001 %
1'
b1001 +
#35600000000
0!
0'
#35610000000
1!
b0 %
1'
b0 +
#35620000000
0!
0'
#35630000000
1!
1$
b1 %
1'
1*
b1 +
#35640000000
0!
0'
#35650000000
1!
b10 %
1'
b10 +
#35660000000
0!
0'
#35670000000
1!
b11 %
1'
b11 +
#35680000000
0!
0'
#35690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#35700000000
0!
0'
#35710000000
1!
b101 %
1'
b101 +
#35720000000
0!
0'
#35730000000
1!
0$
b110 %
1'
0*
b110 +
#35740000000
0!
0'
#35750000000
1!
b111 %
1'
b111 +
#35760000000
0!
0'
#35770000000
1!
b1000 %
1'
b1000 +
#35780000000
0!
0'
#35790000000
1!
b1001 %
1'
b1001 +
#35800000000
0!
0'
#35810000000
1!
b0 %
1'
b0 +
#35820000000
0!
0'
#35830000000
1!
1$
b1 %
1'
1*
b1 +
#35840000000
0!
0'
#35850000000
1!
b10 %
1'
b10 +
#35860000000
0!
0'
#35870000000
1!
b11 %
1'
b11 +
#35880000000
0!
0'
#35890000000
1!
b100 %
1'
b100 +
#35900000000
1"
1(
#35910000000
0!
0"
b100 &
0'
0(
b100 ,
#35920000000
1!
b101 %
1'
b101 +
#35930000000
0!
0'
#35940000000
1!
b110 %
1'
b110 +
#35950000000
0!
0'
#35960000000
1!
b111 %
1'
b111 +
#35970000000
0!
0'
#35980000000
1!
0$
b1000 %
1'
0*
b1000 +
#35990000000
0!
0'
#36000000000
1!
b1001 %
1'
b1001 +
#36010000000
0!
0'
#36020000000
1!
b0 %
1'
b0 +
#36030000000
0!
0'
#36040000000
1!
1$
b1 %
1'
1*
b1 +
#36050000000
0!
0'
#36060000000
1!
b10 %
1'
b10 +
#36070000000
0!
0'
#36080000000
1!
b11 %
1'
b11 +
#36090000000
0!
0'
#36100000000
1!
b100 %
1'
b100 +
#36110000000
0!
0'
#36120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#36130000000
0!
0'
#36140000000
1!
0$
b110 %
1'
0*
b110 +
#36150000000
0!
0'
#36160000000
1!
b111 %
1'
b111 +
#36170000000
0!
0'
#36180000000
1!
b1000 %
1'
b1000 +
#36190000000
0!
0'
#36200000000
1!
b1001 %
1'
b1001 +
#36210000000
0!
0'
#36220000000
1!
b0 %
1'
b0 +
#36230000000
0!
0'
#36240000000
1!
1$
b1 %
1'
1*
b1 +
#36250000000
0!
0'
#36260000000
1!
b10 %
1'
b10 +
#36270000000
0!
0'
#36280000000
1!
b11 %
1'
b11 +
#36290000000
0!
0'
#36300000000
1!
b100 %
1'
b100 +
#36310000000
0!
0'
#36320000000
1!
b101 %
1'
b101 +
#36330000000
1"
1(
#36340000000
0!
0"
b100 &
0'
0(
b100 ,
#36350000000
1!
b110 %
1'
b110 +
#36360000000
0!
0'
#36370000000
1!
b111 %
1'
b111 +
#36380000000
0!
0'
#36390000000
1!
0$
b1000 %
1'
0*
b1000 +
#36400000000
0!
0'
#36410000000
1!
b1001 %
1'
b1001 +
#36420000000
0!
0'
#36430000000
1!
b0 %
1'
b0 +
#36440000000
0!
0'
#36450000000
1!
1$
b1 %
1'
1*
b1 +
#36460000000
0!
0'
#36470000000
1!
b10 %
1'
b10 +
#36480000000
0!
0'
#36490000000
1!
b11 %
1'
b11 +
#36500000000
0!
0'
#36510000000
1!
b100 %
1'
b100 +
#36520000000
0!
0'
#36530000000
1!
b101 %
1'
b101 +
#36540000000
0!
0'
#36550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#36560000000
0!
0'
#36570000000
1!
b111 %
1'
b111 +
#36580000000
0!
0'
#36590000000
1!
b1000 %
1'
b1000 +
#36600000000
0!
0'
#36610000000
1!
b1001 %
1'
b1001 +
#36620000000
0!
0'
#36630000000
1!
b0 %
1'
b0 +
#36640000000
0!
0'
#36650000000
1!
1$
b1 %
1'
1*
b1 +
#36660000000
0!
0'
#36670000000
1!
b10 %
1'
b10 +
#36680000000
0!
0'
#36690000000
1!
b11 %
1'
b11 +
#36700000000
0!
0'
#36710000000
1!
b100 %
1'
b100 +
#36720000000
0!
0'
#36730000000
1!
b101 %
1'
b101 +
#36740000000
0!
0'
#36750000000
1!
0$
b110 %
1'
0*
b110 +
#36760000000
1"
1(
#36770000000
0!
0"
b100 &
0'
0(
b100 ,
#36780000000
1!
1$
b111 %
1'
1*
b111 +
#36790000000
0!
0'
#36800000000
1!
0$
b1000 %
1'
0*
b1000 +
#36810000000
0!
0'
#36820000000
1!
b1001 %
1'
b1001 +
#36830000000
0!
0'
#36840000000
1!
b0 %
1'
b0 +
#36850000000
0!
0'
#36860000000
1!
1$
b1 %
1'
1*
b1 +
#36870000000
0!
0'
#36880000000
1!
b10 %
1'
b10 +
#36890000000
0!
0'
#36900000000
1!
b11 %
1'
b11 +
#36910000000
0!
0'
#36920000000
1!
b100 %
1'
b100 +
#36930000000
0!
0'
#36940000000
1!
b101 %
1'
b101 +
#36950000000
0!
0'
#36960000000
1!
b110 %
1'
b110 +
#36970000000
0!
0'
#36980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#36990000000
0!
0'
#37000000000
1!
b1000 %
1'
b1000 +
#37010000000
0!
0'
#37020000000
1!
b1001 %
1'
b1001 +
#37030000000
0!
0'
#37040000000
1!
b0 %
1'
b0 +
#37050000000
0!
0'
#37060000000
1!
1$
b1 %
1'
1*
b1 +
#37070000000
0!
0'
#37080000000
1!
b10 %
1'
b10 +
#37090000000
0!
0'
#37100000000
1!
b11 %
1'
b11 +
#37110000000
0!
0'
#37120000000
1!
b100 %
1'
b100 +
#37130000000
0!
0'
#37140000000
1!
b101 %
1'
b101 +
#37150000000
0!
0'
#37160000000
1!
0$
b110 %
1'
0*
b110 +
#37170000000
0!
0'
#37180000000
1!
b111 %
1'
b111 +
#37190000000
1"
1(
#37200000000
0!
0"
b100 &
0'
0(
b100 ,
#37210000000
1!
b1000 %
1'
b1000 +
#37220000000
0!
0'
#37230000000
1!
b1001 %
1'
b1001 +
#37240000000
0!
0'
#37250000000
1!
b0 %
1'
b0 +
#37260000000
0!
0'
#37270000000
1!
1$
b1 %
1'
1*
b1 +
#37280000000
0!
0'
#37290000000
1!
b10 %
1'
b10 +
#37300000000
0!
0'
#37310000000
1!
b11 %
1'
b11 +
#37320000000
0!
0'
#37330000000
1!
b100 %
1'
b100 +
#37340000000
0!
0'
#37350000000
1!
b101 %
1'
b101 +
#37360000000
0!
0'
#37370000000
1!
b110 %
1'
b110 +
#37380000000
0!
0'
#37390000000
1!
b111 %
1'
b111 +
#37400000000
0!
0'
#37410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#37420000000
0!
0'
#37430000000
1!
b1001 %
1'
b1001 +
#37440000000
0!
0'
#37450000000
1!
b0 %
1'
b0 +
#37460000000
0!
0'
#37470000000
1!
1$
b1 %
1'
1*
b1 +
#37480000000
0!
0'
#37490000000
1!
b10 %
1'
b10 +
#37500000000
0!
0'
#37510000000
1!
b11 %
1'
b11 +
#37520000000
0!
0'
#37530000000
1!
b100 %
1'
b100 +
#37540000000
0!
0'
#37550000000
1!
b101 %
1'
b101 +
#37560000000
0!
0'
#37570000000
1!
0$
b110 %
1'
0*
b110 +
#37580000000
0!
0'
#37590000000
1!
b111 %
1'
b111 +
#37600000000
0!
0'
#37610000000
1!
b1000 %
1'
b1000 +
#37620000000
1"
1(
#37630000000
0!
0"
b100 &
0'
0(
b100 ,
#37640000000
1!
b1001 %
1'
b1001 +
#37650000000
0!
0'
#37660000000
1!
b0 %
1'
b0 +
#37670000000
0!
0'
#37680000000
1!
1$
b1 %
1'
1*
b1 +
#37690000000
0!
0'
#37700000000
1!
b10 %
1'
b10 +
#37710000000
0!
0'
#37720000000
1!
b11 %
1'
b11 +
#37730000000
0!
0'
#37740000000
1!
b100 %
1'
b100 +
#37750000000
0!
0'
#37760000000
1!
b101 %
1'
b101 +
#37770000000
0!
0'
#37780000000
1!
b110 %
1'
b110 +
#37790000000
0!
0'
#37800000000
1!
b111 %
1'
b111 +
#37810000000
0!
0'
#37820000000
1!
0$
b1000 %
1'
0*
b1000 +
#37830000000
0!
0'
#37840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#37850000000
0!
0'
#37860000000
1!
b0 %
1'
b0 +
#37870000000
0!
0'
#37880000000
1!
1$
b1 %
1'
1*
b1 +
#37890000000
0!
0'
#37900000000
1!
b10 %
1'
b10 +
#37910000000
0!
0'
#37920000000
1!
b11 %
1'
b11 +
#37930000000
0!
0'
#37940000000
1!
b100 %
1'
b100 +
#37950000000
0!
0'
#37960000000
1!
b101 %
1'
b101 +
#37970000000
0!
0'
#37980000000
1!
0$
b110 %
1'
0*
b110 +
#37990000000
0!
0'
#38000000000
1!
b111 %
1'
b111 +
#38010000000
0!
0'
#38020000000
1!
b1000 %
1'
b1000 +
#38030000000
0!
0'
#38040000000
1!
b1001 %
1'
b1001 +
#38050000000
1"
1(
#38060000000
0!
0"
b100 &
0'
0(
b100 ,
#38070000000
1!
b0 %
1'
b0 +
#38080000000
0!
0'
#38090000000
1!
1$
b1 %
1'
1*
b1 +
#38100000000
0!
0'
#38110000000
1!
b10 %
1'
b10 +
#38120000000
0!
0'
#38130000000
1!
b11 %
1'
b11 +
#38140000000
0!
0'
#38150000000
1!
b100 %
1'
b100 +
#38160000000
0!
0'
#38170000000
1!
b101 %
1'
b101 +
#38180000000
0!
0'
#38190000000
1!
b110 %
1'
b110 +
#38200000000
0!
0'
#38210000000
1!
b111 %
1'
b111 +
#38220000000
0!
0'
#38230000000
1!
0$
b1000 %
1'
0*
b1000 +
#38240000000
0!
0'
#38250000000
1!
b1001 %
1'
b1001 +
#38260000000
0!
0'
#38270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#38280000000
0!
0'
#38290000000
1!
1$
b1 %
1'
1*
b1 +
#38300000000
0!
0'
#38310000000
1!
b10 %
1'
b10 +
#38320000000
0!
0'
#38330000000
1!
b11 %
1'
b11 +
#38340000000
0!
0'
#38350000000
1!
b100 %
1'
b100 +
#38360000000
0!
0'
#38370000000
1!
b101 %
1'
b101 +
#38380000000
0!
0'
#38390000000
1!
0$
b110 %
1'
0*
b110 +
#38400000000
0!
0'
#38410000000
1!
b111 %
1'
b111 +
#38420000000
0!
0'
#38430000000
1!
b1000 %
1'
b1000 +
#38440000000
0!
0'
#38450000000
1!
b1001 %
1'
b1001 +
#38460000000
0!
0'
#38470000000
1!
b0 %
1'
b0 +
#38480000000
1"
1(
#38490000000
0!
0"
b100 &
0'
0(
b100 ,
#38500000000
1!
1$
b1 %
1'
1*
b1 +
#38510000000
0!
0'
#38520000000
1!
b10 %
1'
b10 +
#38530000000
0!
0'
#38540000000
1!
b11 %
1'
b11 +
#38550000000
0!
0'
#38560000000
1!
b100 %
1'
b100 +
#38570000000
0!
0'
#38580000000
1!
b101 %
1'
b101 +
#38590000000
0!
0'
#38600000000
1!
b110 %
1'
b110 +
#38610000000
0!
0'
#38620000000
1!
b111 %
1'
b111 +
#38630000000
0!
0'
#38640000000
1!
0$
b1000 %
1'
0*
b1000 +
#38650000000
0!
0'
#38660000000
1!
b1001 %
1'
b1001 +
#38670000000
0!
0'
#38680000000
1!
b0 %
1'
b0 +
#38690000000
0!
0'
#38700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#38710000000
0!
0'
#38720000000
1!
b10 %
1'
b10 +
#38730000000
0!
0'
#38740000000
1!
b11 %
1'
b11 +
#38750000000
0!
0'
#38760000000
1!
b100 %
1'
b100 +
#38770000000
0!
0'
#38780000000
1!
b101 %
1'
b101 +
#38790000000
0!
0'
#38800000000
1!
0$
b110 %
1'
0*
b110 +
#38810000000
0!
0'
#38820000000
1!
b111 %
1'
b111 +
#38830000000
0!
0'
#38840000000
1!
b1000 %
1'
b1000 +
#38850000000
0!
0'
#38860000000
1!
b1001 %
1'
b1001 +
#38870000000
0!
0'
#38880000000
1!
b0 %
1'
b0 +
#38890000000
0!
0'
#38900000000
1!
1$
b1 %
1'
1*
b1 +
#38910000000
1"
1(
#38920000000
0!
0"
b100 &
0'
0(
b100 ,
#38930000000
1!
b10 %
1'
b10 +
#38940000000
0!
0'
#38950000000
1!
b11 %
1'
b11 +
#38960000000
0!
0'
#38970000000
1!
b100 %
1'
b100 +
#38980000000
0!
0'
#38990000000
1!
b101 %
1'
b101 +
#39000000000
0!
0'
#39010000000
1!
b110 %
1'
b110 +
#39020000000
0!
0'
#39030000000
1!
b111 %
1'
b111 +
#39040000000
0!
0'
#39050000000
1!
0$
b1000 %
1'
0*
b1000 +
#39060000000
0!
0'
#39070000000
1!
b1001 %
1'
b1001 +
#39080000000
0!
0'
#39090000000
1!
b0 %
1'
b0 +
#39100000000
0!
0'
#39110000000
1!
1$
b1 %
1'
1*
b1 +
#39120000000
0!
0'
#39130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#39140000000
0!
0'
#39150000000
1!
b11 %
1'
b11 +
#39160000000
0!
0'
#39170000000
1!
b100 %
1'
b100 +
#39180000000
0!
0'
#39190000000
1!
b101 %
1'
b101 +
#39200000000
0!
0'
#39210000000
1!
0$
b110 %
1'
0*
b110 +
#39220000000
0!
0'
#39230000000
1!
b111 %
1'
b111 +
#39240000000
0!
0'
#39250000000
1!
b1000 %
1'
b1000 +
#39260000000
0!
0'
#39270000000
1!
b1001 %
1'
b1001 +
#39280000000
0!
0'
#39290000000
1!
b0 %
1'
b0 +
#39300000000
0!
0'
#39310000000
1!
1$
b1 %
1'
1*
b1 +
#39320000000
0!
0'
#39330000000
1!
b10 %
1'
b10 +
#39340000000
1"
1(
#39350000000
0!
0"
b100 &
0'
0(
b100 ,
#39360000000
1!
b11 %
1'
b11 +
#39370000000
0!
0'
#39380000000
1!
b100 %
1'
b100 +
#39390000000
0!
0'
#39400000000
1!
b101 %
1'
b101 +
#39410000000
0!
0'
#39420000000
1!
b110 %
1'
b110 +
#39430000000
0!
0'
#39440000000
1!
b111 %
1'
b111 +
#39450000000
0!
0'
#39460000000
1!
0$
b1000 %
1'
0*
b1000 +
#39470000000
0!
0'
#39480000000
1!
b1001 %
1'
b1001 +
#39490000000
0!
0'
#39500000000
1!
b0 %
1'
b0 +
#39510000000
0!
0'
#39520000000
1!
1$
b1 %
1'
1*
b1 +
#39530000000
0!
0'
#39540000000
1!
b10 %
1'
b10 +
#39550000000
0!
0'
#39560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#39570000000
0!
0'
#39580000000
1!
b100 %
1'
b100 +
#39590000000
0!
0'
#39600000000
1!
b101 %
1'
b101 +
#39610000000
0!
0'
#39620000000
1!
0$
b110 %
1'
0*
b110 +
#39630000000
0!
0'
#39640000000
1!
b111 %
1'
b111 +
#39650000000
0!
0'
#39660000000
1!
b1000 %
1'
b1000 +
#39670000000
0!
0'
#39680000000
1!
b1001 %
1'
b1001 +
#39690000000
0!
0'
#39700000000
1!
b0 %
1'
b0 +
#39710000000
0!
0'
#39720000000
1!
1$
b1 %
1'
1*
b1 +
#39730000000
0!
0'
#39740000000
1!
b10 %
1'
b10 +
#39750000000
0!
0'
#39760000000
1!
b11 %
1'
b11 +
#39770000000
1"
1(
#39780000000
0!
0"
b100 &
0'
0(
b100 ,
#39790000000
1!
b100 %
1'
b100 +
#39800000000
0!
0'
#39810000000
1!
b101 %
1'
b101 +
#39820000000
0!
0'
#39830000000
1!
b110 %
1'
b110 +
#39840000000
0!
0'
#39850000000
1!
b111 %
1'
b111 +
#39860000000
0!
0'
#39870000000
1!
0$
b1000 %
1'
0*
b1000 +
#39880000000
0!
0'
#39890000000
1!
b1001 %
1'
b1001 +
#39900000000
0!
0'
#39910000000
1!
b0 %
1'
b0 +
#39920000000
0!
0'
#39930000000
1!
1$
b1 %
1'
1*
b1 +
#39940000000
0!
0'
#39950000000
1!
b10 %
1'
b10 +
#39960000000
0!
0'
#39970000000
1!
b11 %
1'
b11 +
#39980000000
0!
0'
#39990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#40000000000
0!
0'
#40010000000
1!
b101 %
1'
b101 +
#40020000000
0!
0'
#40030000000
1!
0$
b110 %
1'
0*
b110 +
#40040000000
0!
0'
#40050000000
1!
b111 %
1'
b111 +
#40060000000
0!
0'
#40070000000
1!
b1000 %
1'
b1000 +
#40080000000
0!
0'
#40090000000
1!
b1001 %
1'
b1001 +
#40100000000
0!
0'
#40110000000
1!
b0 %
1'
b0 +
#40120000000
0!
0'
#40130000000
1!
1$
b1 %
1'
1*
b1 +
#40140000000
0!
0'
#40150000000
1!
b10 %
1'
b10 +
#40160000000
0!
0'
#40170000000
1!
b11 %
1'
b11 +
#40180000000
0!
0'
#40190000000
1!
b100 %
1'
b100 +
#40200000000
1"
1(
#40210000000
0!
0"
b100 &
0'
0(
b100 ,
#40220000000
1!
b101 %
1'
b101 +
#40230000000
0!
0'
#40240000000
1!
b110 %
1'
b110 +
#40250000000
0!
0'
#40260000000
1!
b111 %
1'
b111 +
#40270000000
0!
0'
#40280000000
1!
0$
b1000 %
1'
0*
b1000 +
#40290000000
0!
0'
#40300000000
1!
b1001 %
1'
b1001 +
#40310000000
0!
0'
#40320000000
1!
b0 %
1'
b0 +
#40330000000
0!
0'
#40340000000
1!
1$
b1 %
1'
1*
b1 +
#40350000000
0!
0'
#40360000000
1!
b10 %
1'
b10 +
#40370000000
0!
0'
#40380000000
1!
b11 %
1'
b11 +
#40390000000
0!
0'
#40400000000
1!
b100 %
1'
b100 +
#40410000000
0!
0'
#40420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#40430000000
0!
0'
#40440000000
1!
0$
b110 %
1'
0*
b110 +
#40450000000
0!
0'
#40460000000
1!
b111 %
1'
b111 +
#40470000000
0!
0'
#40480000000
1!
b1000 %
1'
b1000 +
#40490000000
0!
0'
#40500000000
1!
b1001 %
1'
b1001 +
#40510000000
0!
0'
#40520000000
1!
b0 %
1'
b0 +
#40530000000
0!
0'
#40540000000
1!
1$
b1 %
1'
1*
b1 +
#40550000000
0!
0'
#40560000000
1!
b10 %
1'
b10 +
#40570000000
0!
0'
#40580000000
1!
b11 %
1'
b11 +
#40590000000
0!
0'
#40600000000
1!
b100 %
1'
b100 +
#40610000000
0!
0'
#40620000000
1!
b101 %
1'
b101 +
#40630000000
1"
1(
#40640000000
0!
0"
b100 &
0'
0(
b100 ,
#40650000000
1!
b110 %
1'
b110 +
#40660000000
0!
0'
#40670000000
1!
b111 %
1'
b111 +
#40680000000
0!
0'
#40690000000
1!
0$
b1000 %
1'
0*
b1000 +
#40700000000
0!
0'
#40710000000
1!
b1001 %
1'
b1001 +
#40720000000
0!
0'
#40730000000
1!
b0 %
1'
b0 +
#40740000000
0!
0'
#40750000000
1!
1$
b1 %
1'
1*
b1 +
#40760000000
0!
0'
#40770000000
1!
b10 %
1'
b10 +
#40780000000
0!
0'
#40790000000
1!
b11 %
1'
b11 +
#40800000000
0!
0'
#40810000000
1!
b100 %
1'
b100 +
#40820000000
0!
0'
#40830000000
1!
b101 %
1'
b101 +
#40840000000
0!
0'
#40850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#40860000000
0!
0'
#40870000000
1!
b111 %
1'
b111 +
#40880000000
0!
0'
#40890000000
1!
b1000 %
1'
b1000 +
#40900000000
0!
0'
#40910000000
1!
b1001 %
1'
b1001 +
#40920000000
0!
0'
#40930000000
1!
b0 %
1'
b0 +
#40940000000
0!
0'
#40950000000
1!
1$
b1 %
1'
1*
b1 +
#40960000000
0!
0'
#40970000000
1!
b10 %
1'
b10 +
#40980000000
0!
0'
#40990000000
1!
b11 %
1'
b11 +
#41000000000
0!
0'
#41010000000
1!
b100 %
1'
b100 +
#41020000000
0!
0'
#41030000000
1!
b101 %
1'
b101 +
#41040000000
0!
0'
#41050000000
1!
0$
b110 %
1'
0*
b110 +
#41060000000
1"
1(
#41070000000
0!
0"
b100 &
0'
0(
b100 ,
#41080000000
1!
1$
b111 %
1'
1*
b111 +
#41090000000
0!
0'
#41100000000
1!
0$
b1000 %
1'
0*
b1000 +
#41110000000
0!
0'
#41120000000
1!
b1001 %
1'
b1001 +
#41130000000
0!
0'
#41140000000
1!
b0 %
1'
b0 +
#41150000000
0!
0'
#41160000000
1!
1$
b1 %
1'
1*
b1 +
#41170000000
0!
0'
#41180000000
1!
b10 %
1'
b10 +
#41190000000
0!
0'
#41200000000
1!
b11 %
1'
b11 +
#41210000000
0!
0'
#41220000000
1!
b100 %
1'
b100 +
#41230000000
0!
0'
#41240000000
1!
b101 %
1'
b101 +
#41250000000
0!
0'
#41260000000
1!
b110 %
1'
b110 +
#41270000000
0!
0'
#41280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#41290000000
0!
0'
#41300000000
1!
b1000 %
1'
b1000 +
#41310000000
0!
0'
#41320000000
1!
b1001 %
1'
b1001 +
#41330000000
0!
0'
#41340000000
1!
b0 %
1'
b0 +
#41350000000
0!
0'
#41360000000
1!
1$
b1 %
1'
1*
b1 +
#41370000000
0!
0'
#41380000000
1!
b10 %
1'
b10 +
#41390000000
0!
0'
#41400000000
1!
b11 %
1'
b11 +
#41410000000
0!
0'
#41420000000
1!
b100 %
1'
b100 +
#41430000000
0!
0'
#41440000000
1!
b101 %
1'
b101 +
#41450000000
0!
0'
#41460000000
1!
0$
b110 %
1'
0*
b110 +
#41470000000
0!
0'
#41480000000
1!
b111 %
1'
b111 +
#41490000000
1"
1(
#41500000000
0!
0"
b100 &
0'
0(
b100 ,
#41510000000
1!
b1000 %
1'
b1000 +
#41520000000
0!
0'
#41530000000
1!
b1001 %
1'
b1001 +
#41540000000
0!
0'
#41550000000
1!
b0 %
1'
b0 +
#41560000000
0!
0'
#41570000000
1!
1$
b1 %
1'
1*
b1 +
#41580000000
0!
0'
#41590000000
1!
b10 %
1'
b10 +
#41600000000
0!
0'
#41610000000
1!
b11 %
1'
b11 +
#41620000000
0!
0'
#41630000000
1!
b100 %
1'
b100 +
#41640000000
0!
0'
#41650000000
1!
b101 %
1'
b101 +
#41660000000
0!
0'
#41670000000
1!
b110 %
1'
b110 +
#41680000000
0!
0'
#41690000000
1!
b111 %
1'
b111 +
#41700000000
0!
0'
#41710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#41720000000
0!
0'
#41730000000
1!
b1001 %
1'
b1001 +
#41740000000
0!
0'
#41750000000
1!
b0 %
1'
b0 +
#41760000000
0!
0'
#41770000000
1!
1$
b1 %
1'
1*
b1 +
#41780000000
0!
0'
#41790000000
1!
b10 %
1'
b10 +
#41800000000
0!
0'
#41810000000
1!
b11 %
1'
b11 +
#41820000000
0!
0'
#41830000000
1!
b100 %
1'
b100 +
#41840000000
0!
0'
#41850000000
1!
b101 %
1'
b101 +
#41860000000
0!
0'
#41870000000
1!
0$
b110 %
1'
0*
b110 +
#41880000000
0!
0'
#41890000000
1!
b111 %
1'
b111 +
#41900000000
0!
0'
#41910000000
1!
b1000 %
1'
b1000 +
#41920000000
1"
1(
#41930000000
0!
0"
b100 &
0'
0(
b100 ,
#41940000000
1!
b1001 %
1'
b1001 +
#41950000000
0!
0'
#41960000000
1!
b0 %
1'
b0 +
#41970000000
0!
0'
#41980000000
1!
1$
b1 %
1'
1*
b1 +
#41990000000
0!
0'
#42000000000
1!
b10 %
1'
b10 +
#42010000000
0!
0'
#42020000000
1!
b11 %
1'
b11 +
#42030000000
0!
0'
#42040000000
1!
b100 %
1'
b100 +
#42050000000
0!
0'
#42060000000
1!
b101 %
1'
b101 +
#42070000000
0!
0'
#42080000000
1!
b110 %
1'
b110 +
#42090000000
0!
0'
#42100000000
1!
b111 %
1'
b111 +
#42110000000
0!
0'
#42120000000
1!
0$
b1000 %
1'
0*
b1000 +
#42130000000
0!
0'
#42140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#42150000000
0!
0'
#42160000000
1!
b0 %
1'
b0 +
#42170000000
0!
0'
#42180000000
1!
1$
b1 %
1'
1*
b1 +
#42190000000
0!
0'
#42200000000
1!
b10 %
1'
b10 +
#42210000000
0!
0'
#42220000000
1!
b11 %
1'
b11 +
#42230000000
0!
0'
#42240000000
1!
b100 %
1'
b100 +
#42250000000
0!
0'
#42260000000
1!
b101 %
1'
b101 +
#42270000000
0!
0'
#42280000000
1!
0$
b110 %
1'
0*
b110 +
#42290000000
0!
0'
#42300000000
1!
b111 %
1'
b111 +
#42310000000
0!
0'
#42320000000
1!
b1000 %
1'
b1000 +
#42330000000
0!
0'
#42340000000
1!
b1001 %
1'
b1001 +
#42350000000
1"
1(
#42360000000
0!
0"
b100 &
0'
0(
b100 ,
#42370000000
1!
b0 %
1'
b0 +
#42380000000
0!
0'
#42390000000
1!
1$
b1 %
1'
1*
b1 +
#42400000000
0!
0'
#42410000000
1!
b10 %
1'
b10 +
#42420000000
0!
0'
#42430000000
1!
b11 %
1'
b11 +
#42440000000
0!
0'
#42450000000
1!
b100 %
1'
b100 +
#42460000000
0!
0'
#42470000000
1!
b101 %
1'
b101 +
#42480000000
0!
0'
#42490000000
1!
b110 %
1'
b110 +
#42500000000
0!
0'
#42510000000
1!
b111 %
1'
b111 +
#42520000000
0!
0'
#42530000000
1!
0$
b1000 %
1'
0*
b1000 +
#42540000000
0!
0'
#42550000000
1!
b1001 %
1'
b1001 +
#42560000000
0!
0'
#42570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#42580000000
0!
0'
#42590000000
1!
1$
b1 %
1'
1*
b1 +
#42600000000
0!
0'
#42610000000
1!
b10 %
1'
b10 +
#42620000000
0!
0'
#42630000000
1!
b11 %
1'
b11 +
#42640000000
0!
0'
#42650000000
1!
b100 %
1'
b100 +
#42660000000
0!
0'
#42670000000
1!
b101 %
1'
b101 +
#42680000000
0!
0'
#42690000000
1!
0$
b110 %
1'
0*
b110 +
#42700000000
0!
0'
#42710000000
1!
b111 %
1'
b111 +
#42720000000
0!
0'
#42730000000
1!
b1000 %
1'
b1000 +
#42740000000
0!
0'
#42750000000
1!
b1001 %
1'
b1001 +
#42760000000
0!
0'
#42770000000
1!
b0 %
1'
b0 +
#42780000000
1"
1(
#42790000000
0!
0"
b100 &
0'
0(
b100 ,
#42800000000
1!
1$
b1 %
1'
1*
b1 +
#42810000000
0!
0'
#42820000000
1!
b10 %
1'
b10 +
#42830000000
0!
0'
#42840000000
1!
b11 %
1'
b11 +
#42850000000
0!
0'
#42860000000
1!
b100 %
1'
b100 +
#42870000000
0!
0'
#42880000000
1!
b101 %
1'
b101 +
#42890000000
0!
0'
#42900000000
1!
b110 %
1'
b110 +
#42910000000
0!
0'
#42920000000
1!
b111 %
1'
b111 +
#42930000000
0!
0'
#42940000000
1!
0$
b1000 %
1'
0*
b1000 +
#42950000000
0!
0'
#42960000000
1!
b1001 %
1'
b1001 +
#42970000000
0!
0'
#42980000000
1!
b0 %
1'
b0 +
#42990000000
0!
0'
#43000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#43010000000
0!
0'
#43020000000
1!
b10 %
1'
b10 +
#43030000000
0!
0'
#43040000000
1!
b11 %
1'
b11 +
#43050000000
0!
0'
#43060000000
1!
b100 %
1'
b100 +
#43070000000
0!
0'
#43080000000
1!
b101 %
1'
b101 +
#43090000000
0!
0'
#43100000000
1!
0$
b110 %
1'
0*
b110 +
#43110000000
0!
0'
#43120000000
1!
b111 %
1'
b111 +
#43130000000
0!
0'
#43140000000
1!
b1000 %
1'
b1000 +
#43150000000
0!
0'
#43160000000
1!
b1001 %
1'
b1001 +
#43170000000
0!
0'
#43180000000
1!
b0 %
1'
b0 +
#43190000000
0!
0'
#43200000000
1!
1$
b1 %
1'
1*
b1 +
#43210000000
1"
1(
#43220000000
0!
0"
b100 &
0'
0(
b100 ,
#43230000000
1!
b10 %
1'
b10 +
#43240000000
0!
0'
#43250000000
1!
b11 %
1'
b11 +
#43260000000
0!
0'
#43270000000
1!
b100 %
1'
b100 +
#43280000000
0!
0'
#43290000000
1!
b101 %
1'
b101 +
#43300000000
0!
0'
#43310000000
1!
b110 %
1'
b110 +
#43320000000
0!
0'
#43330000000
1!
b111 %
1'
b111 +
#43340000000
0!
0'
#43350000000
1!
0$
b1000 %
1'
0*
b1000 +
#43360000000
0!
0'
#43370000000
1!
b1001 %
1'
b1001 +
#43380000000
0!
0'
#43390000000
1!
b0 %
1'
b0 +
#43400000000
0!
0'
#43410000000
1!
1$
b1 %
1'
1*
b1 +
#43420000000
0!
0'
#43430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#43440000000
0!
0'
#43450000000
1!
b11 %
1'
b11 +
#43460000000
0!
0'
#43470000000
1!
b100 %
1'
b100 +
#43480000000
0!
0'
#43490000000
1!
b101 %
1'
b101 +
#43500000000
0!
0'
#43510000000
1!
0$
b110 %
1'
0*
b110 +
#43520000000
0!
0'
#43530000000
1!
b111 %
1'
b111 +
#43540000000
0!
0'
#43550000000
1!
b1000 %
1'
b1000 +
#43560000000
0!
0'
#43570000000
1!
b1001 %
1'
b1001 +
#43580000000
0!
0'
#43590000000
1!
b0 %
1'
b0 +
#43600000000
0!
0'
#43610000000
1!
1$
b1 %
1'
1*
b1 +
#43620000000
0!
0'
#43630000000
1!
b10 %
1'
b10 +
#43640000000
1"
1(
#43650000000
0!
0"
b100 &
0'
0(
b100 ,
#43660000000
1!
b11 %
1'
b11 +
#43670000000
0!
0'
#43680000000
1!
b100 %
1'
b100 +
#43690000000
0!
0'
#43700000000
1!
b101 %
1'
b101 +
#43710000000
0!
0'
#43720000000
1!
b110 %
1'
b110 +
#43730000000
0!
0'
#43740000000
1!
b111 %
1'
b111 +
#43750000000
0!
0'
#43760000000
1!
0$
b1000 %
1'
0*
b1000 +
#43770000000
0!
0'
#43780000000
1!
b1001 %
1'
b1001 +
#43790000000
0!
0'
#43800000000
1!
b0 %
1'
b0 +
#43810000000
0!
0'
#43820000000
1!
1$
b1 %
1'
1*
b1 +
#43830000000
0!
0'
#43840000000
1!
b10 %
1'
b10 +
#43850000000
0!
0'
#43860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#43870000000
0!
0'
#43880000000
1!
b100 %
1'
b100 +
#43890000000
0!
0'
#43900000000
1!
b101 %
1'
b101 +
#43910000000
0!
0'
#43920000000
1!
0$
b110 %
1'
0*
b110 +
#43930000000
0!
0'
#43940000000
1!
b111 %
1'
b111 +
#43950000000
0!
0'
#43960000000
1!
b1000 %
1'
b1000 +
#43970000000
0!
0'
#43980000000
1!
b1001 %
1'
b1001 +
#43990000000
0!
0'
#44000000000
1!
b0 %
1'
b0 +
#44010000000
0!
0'
#44020000000
1!
1$
b1 %
1'
1*
b1 +
#44030000000
0!
0'
#44040000000
1!
b10 %
1'
b10 +
#44050000000
0!
0'
#44060000000
1!
b11 %
1'
b11 +
#44070000000
1"
1(
#44080000000
0!
0"
b100 &
0'
0(
b100 ,
#44090000000
1!
b100 %
1'
b100 +
#44100000000
0!
0'
#44110000000
1!
b101 %
1'
b101 +
#44120000000
0!
0'
#44130000000
1!
b110 %
1'
b110 +
#44140000000
0!
0'
#44150000000
1!
b111 %
1'
b111 +
#44160000000
0!
0'
#44170000000
1!
0$
b1000 %
1'
0*
b1000 +
#44180000000
0!
0'
#44190000000
1!
b1001 %
1'
b1001 +
#44200000000
0!
0'
#44210000000
1!
b0 %
1'
b0 +
#44220000000
0!
0'
#44230000000
1!
1$
b1 %
1'
1*
b1 +
#44240000000
0!
0'
#44250000000
1!
b10 %
1'
b10 +
#44260000000
0!
0'
#44270000000
1!
b11 %
1'
b11 +
#44280000000
0!
0'
#44290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#44300000000
0!
0'
#44310000000
1!
b101 %
1'
b101 +
#44320000000
0!
0'
#44330000000
1!
0$
b110 %
1'
0*
b110 +
#44340000000
0!
0'
#44350000000
1!
b111 %
1'
b111 +
#44360000000
0!
0'
#44370000000
1!
b1000 %
1'
b1000 +
#44380000000
0!
0'
#44390000000
1!
b1001 %
1'
b1001 +
#44400000000
0!
0'
#44410000000
1!
b0 %
1'
b0 +
#44420000000
0!
0'
#44430000000
1!
1$
b1 %
1'
1*
b1 +
#44440000000
0!
0'
#44450000000
1!
b10 %
1'
b10 +
#44460000000
0!
0'
#44470000000
1!
b11 %
1'
b11 +
#44480000000
0!
0'
#44490000000
1!
b100 %
1'
b100 +
#44500000000
1"
1(
#44510000000
0!
0"
b100 &
0'
0(
b100 ,
#44520000000
1!
b101 %
1'
b101 +
#44530000000
0!
0'
#44540000000
1!
b110 %
1'
b110 +
#44550000000
0!
0'
#44560000000
1!
b111 %
1'
b111 +
#44570000000
0!
0'
#44580000000
1!
0$
b1000 %
1'
0*
b1000 +
#44590000000
0!
0'
#44600000000
1!
b1001 %
1'
b1001 +
#44610000000
0!
0'
#44620000000
1!
b0 %
1'
b0 +
#44630000000
0!
0'
#44640000000
1!
1$
b1 %
1'
1*
b1 +
#44650000000
0!
0'
#44660000000
1!
b10 %
1'
b10 +
#44670000000
0!
0'
#44680000000
1!
b11 %
1'
b11 +
#44690000000
0!
0'
#44700000000
1!
b100 %
1'
b100 +
#44710000000
0!
0'
#44720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#44730000000
0!
0'
#44740000000
1!
0$
b110 %
1'
0*
b110 +
#44750000000
0!
0'
#44760000000
1!
b111 %
1'
b111 +
#44770000000
0!
0'
#44780000000
1!
b1000 %
1'
b1000 +
#44790000000
0!
0'
#44800000000
1!
b1001 %
1'
b1001 +
#44810000000
0!
0'
#44820000000
1!
b0 %
1'
b0 +
#44830000000
0!
0'
#44840000000
1!
1$
b1 %
1'
1*
b1 +
#44850000000
0!
0'
#44860000000
1!
b10 %
1'
b10 +
#44870000000
0!
0'
#44880000000
1!
b11 %
1'
b11 +
#44890000000
0!
0'
#44900000000
1!
b100 %
1'
b100 +
#44910000000
0!
0'
#44920000000
1!
b101 %
1'
b101 +
#44930000000
1"
1(
#44940000000
0!
0"
b100 &
0'
0(
b100 ,
#44950000000
1!
b110 %
1'
b110 +
#44960000000
0!
0'
#44970000000
1!
b111 %
1'
b111 +
#44980000000
0!
0'
#44990000000
1!
0$
b1000 %
1'
0*
b1000 +
#45000000000
0!
0'
#45010000000
1!
b1001 %
1'
b1001 +
#45020000000
0!
0'
#45030000000
1!
b0 %
1'
b0 +
#45040000000
0!
0'
#45050000000
1!
1$
b1 %
1'
1*
b1 +
#45060000000
0!
0'
#45070000000
1!
b10 %
1'
b10 +
#45080000000
0!
0'
#45090000000
1!
b11 %
1'
b11 +
#45100000000
0!
0'
#45110000000
1!
b100 %
1'
b100 +
#45120000000
0!
0'
#45130000000
1!
b101 %
1'
b101 +
#45140000000
0!
0'
#45150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#45160000000
0!
0'
#45170000000
1!
b111 %
1'
b111 +
#45180000000
0!
0'
#45190000000
1!
b1000 %
1'
b1000 +
#45200000000
0!
0'
#45210000000
1!
b1001 %
1'
b1001 +
#45220000000
0!
0'
#45230000000
1!
b0 %
1'
b0 +
#45240000000
0!
0'
#45250000000
1!
1$
b1 %
1'
1*
b1 +
#45260000000
0!
0'
#45270000000
1!
b10 %
1'
b10 +
#45280000000
0!
0'
#45290000000
1!
b11 %
1'
b11 +
#45300000000
0!
0'
#45310000000
1!
b100 %
1'
b100 +
#45320000000
0!
0'
#45330000000
1!
b101 %
1'
b101 +
#45340000000
0!
0'
#45350000000
1!
0$
b110 %
1'
0*
b110 +
#45360000000
1"
1(
#45370000000
0!
0"
b100 &
0'
0(
b100 ,
#45380000000
1!
1$
b111 %
1'
1*
b111 +
#45390000000
0!
0'
#45400000000
1!
0$
b1000 %
1'
0*
b1000 +
#45410000000
0!
0'
#45420000000
1!
b1001 %
1'
b1001 +
#45430000000
0!
0'
#45440000000
1!
b0 %
1'
b0 +
#45450000000
0!
0'
#45460000000
1!
1$
b1 %
1'
1*
b1 +
#45470000000
0!
0'
#45480000000
1!
b10 %
1'
b10 +
#45490000000
0!
0'
#45500000000
1!
b11 %
1'
b11 +
#45510000000
0!
0'
#45520000000
1!
b100 %
1'
b100 +
#45530000000
0!
0'
#45540000000
1!
b101 %
1'
b101 +
#45550000000
0!
0'
#45560000000
1!
b110 %
1'
b110 +
#45570000000
0!
0'
#45580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#45590000000
0!
0'
#45600000000
1!
b1000 %
1'
b1000 +
#45610000000
0!
0'
#45620000000
1!
b1001 %
1'
b1001 +
#45630000000
0!
0'
#45640000000
1!
b0 %
1'
b0 +
#45650000000
0!
0'
#45660000000
1!
1$
b1 %
1'
1*
b1 +
#45670000000
0!
0'
#45680000000
1!
b10 %
1'
b10 +
#45690000000
0!
0'
#45700000000
1!
b11 %
1'
b11 +
#45710000000
0!
0'
#45720000000
1!
b100 %
1'
b100 +
#45730000000
0!
0'
#45740000000
1!
b101 %
1'
b101 +
#45750000000
0!
0'
#45760000000
1!
0$
b110 %
1'
0*
b110 +
#45770000000
0!
0'
#45780000000
1!
b111 %
1'
b111 +
#45790000000
1"
1(
#45800000000
0!
0"
b100 &
0'
0(
b100 ,
#45810000000
1!
b1000 %
1'
b1000 +
#45820000000
0!
0'
#45830000000
1!
b1001 %
1'
b1001 +
#45840000000
0!
0'
#45850000000
1!
b0 %
1'
b0 +
#45860000000
0!
0'
#45870000000
1!
1$
b1 %
1'
1*
b1 +
#45880000000
0!
0'
#45890000000
1!
b10 %
1'
b10 +
#45900000000
0!
0'
#45910000000
1!
b11 %
1'
b11 +
#45920000000
0!
0'
#45930000000
1!
b100 %
1'
b100 +
#45940000000
0!
0'
#45950000000
1!
b101 %
1'
b101 +
#45960000000
0!
0'
#45970000000
1!
b110 %
1'
b110 +
#45980000000
0!
0'
#45990000000
1!
b111 %
1'
b111 +
#46000000000
0!
0'
#46010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#46020000000
0!
0'
#46030000000
1!
b1001 %
1'
b1001 +
#46040000000
0!
0'
#46050000000
1!
b0 %
1'
b0 +
#46060000000
0!
0'
#46070000000
1!
1$
b1 %
1'
1*
b1 +
#46080000000
0!
0'
#46090000000
1!
b10 %
1'
b10 +
#46100000000
0!
0'
#46110000000
1!
b11 %
1'
b11 +
#46120000000
0!
0'
#46130000000
1!
b100 %
1'
b100 +
#46140000000
0!
0'
#46150000000
1!
b101 %
1'
b101 +
#46160000000
0!
0'
#46170000000
1!
0$
b110 %
1'
0*
b110 +
#46180000000
0!
0'
#46190000000
1!
b111 %
1'
b111 +
#46200000000
0!
0'
#46210000000
1!
b1000 %
1'
b1000 +
#46220000000
1"
1(
#46230000000
0!
0"
b100 &
0'
0(
b100 ,
#46240000000
1!
b1001 %
1'
b1001 +
#46250000000
0!
0'
#46260000000
1!
b0 %
1'
b0 +
#46270000000
0!
0'
#46280000000
1!
1$
b1 %
1'
1*
b1 +
#46290000000
0!
0'
#46300000000
1!
b10 %
1'
b10 +
#46310000000
0!
0'
#46320000000
1!
b11 %
1'
b11 +
#46330000000
0!
0'
#46340000000
1!
b100 %
1'
b100 +
#46350000000
0!
0'
#46360000000
1!
b101 %
1'
b101 +
#46370000000
0!
0'
#46380000000
1!
b110 %
1'
b110 +
#46390000000
0!
0'
#46400000000
1!
b111 %
1'
b111 +
#46410000000
0!
0'
#46420000000
1!
0$
b1000 %
1'
0*
b1000 +
#46430000000
0!
0'
#46440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#46450000000
0!
0'
#46460000000
1!
b0 %
1'
b0 +
#46470000000
0!
0'
#46480000000
1!
1$
b1 %
1'
1*
b1 +
#46490000000
0!
0'
#46500000000
1!
b10 %
1'
b10 +
#46510000000
0!
0'
#46520000000
1!
b11 %
1'
b11 +
#46530000000
0!
0'
#46540000000
1!
b100 %
1'
b100 +
#46550000000
0!
0'
#46560000000
1!
b101 %
1'
b101 +
#46570000000
0!
0'
#46580000000
1!
0$
b110 %
1'
0*
b110 +
#46590000000
0!
0'
#46600000000
1!
b111 %
1'
b111 +
#46610000000
0!
0'
#46620000000
1!
b1000 %
1'
b1000 +
#46630000000
0!
0'
#46640000000
1!
b1001 %
1'
b1001 +
#46650000000
1"
1(
#46660000000
0!
0"
b100 &
0'
0(
b100 ,
#46670000000
1!
b0 %
1'
b0 +
#46680000000
0!
0'
#46690000000
1!
1$
b1 %
1'
1*
b1 +
#46700000000
0!
0'
#46710000000
1!
b10 %
1'
b10 +
#46720000000
0!
0'
#46730000000
1!
b11 %
1'
b11 +
#46740000000
0!
0'
#46750000000
1!
b100 %
1'
b100 +
#46760000000
0!
0'
#46770000000
1!
b101 %
1'
b101 +
#46780000000
0!
0'
#46790000000
1!
b110 %
1'
b110 +
#46800000000
0!
0'
#46810000000
1!
b111 %
1'
b111 +
#46820000000
0!
0'
#46830000000
1!
0$
b1000 %
1'
0*
b1000 +
#46840000000
0!
0'
#46850000000
1!
b1001 %
1'
b1001 +
#46860000000
0!
0'
#46870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#46880000000
0!
0'
#46890000000
1!
1$
b1 %
1'
1*
b1 +
#46900000000
0!
0'
#46910000000
1!
b10 %
1'
b10 +
#46920000000
0!
0'
#46930000000
1!
b11 %
1'
b11 +
#46940000000
0!
0'
#46950000000
1!
b100 %
1'
b100 +
#46960000000
0!
0'
#46970000000
1!
b101 %
1'
b101 +
#46980000000
0!
0'
#46990000000
1!
0$
b110 %
1'
0*
b110 +
#47000000000
0!
0'
#47010000000
1!
b111 %
1'
b111 +
#47020000000
0!
0'
#47030000000
1!
b1000 %
1'
b1000 +
#47040000000
0!
0'
#47050000000
1!
b1001 %
1'
b1001 +
#47060000000
0!
0'
#47070000000
1!
b0 %
1'
b0 +
#47080000000
1"
1(
#47090000000
0!
0"
b100 &
0'
0(
b100 ,
#47100000000
1!
1$
b1 %
1'
1*
b1 +
#47110000000
0!
0'
#47120000000
1!
b10 %
1'
b10 +
#47130000000
0!
0'
#47140000000
1!
b11 %
1'
b11 +
#47150000000
0!
0'
#47160000000
1!
b100 %
1'
b100 +
#47170000000
0!
0'
#47180000000
1!
b101 %
1'
b101 +
#47190000000
0!
0'
#47200000000
1!
b110 %
1'
b110 +
#47210000000
0!
0'
#47220000000
1!
b111 %
1'
b111 +
#47230000000
0!
0'
#47240000000
1!
0$
b1000 %
1'
0*
b1000 +
#47250000000
0!
0'
#47260000000
1!
b1001 %
1'
b1001 +
#47270000000
0!
0'
#47280000000
1!
b0 %
1'
b0 +
#47290000000
0!
0'
#47300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#47310000000
0!
0'
#47320000000
1!
b10 %
1'
b10 +
#47330000000
0!
0'
#47340000000
1!
b11 %
1'
b11 +
#47350000000
0!
0'
#47360000000
1!
b100 %
1'
b100 +
#47370000000
0!
0'
#47380000000
1!
b101 %
1'
b101 +
#47390000000
0!
0'
#47400000000
1!
0$
b110 %
1'
0*
b110 +
#47410000000
0!
0'
#47420000000
1!
b111 %
1'
b111 +
#47430000000
0!
0'
#47440000000
1!
b1000 %
1'
b1000 +
#47450000000
0!
0'
#47460000000
1!
b1001 %
1'
b1001 +
#47470000000
0!
0'
#47480000000
1!
b0 %
1'
b0 +
#47490000000
0!
0'
#47500000000
1!
1$
b1 %
1'
1*
b1 +
#47510000000
1"
1(
#47520000000
0!
0"
b100 &
0'
0(
b100 ,
#47530000000
1!
b10 %
1'
b10 +
#47540000000
0!
0'
#47550000000
1!
b11 %
1'
b11 +
#47560000000
0!
0'
#47570000000
1!
b100 %
1'
b100 +
#47580000000
0!
0'
#47590000000
1!
b101 %
1'
b101 +
#47600000000
0!
0'
#47610000000
1!
b110 %
1'
b110 +
#47620000000
0!
0'
#47630000000
1!
b111 %
1'
b111 +
#47640000000
0!
0'
#47650000000
1!
0$
b1000 %
1'
0*
b1000 +
#47660000000
0!
0'
#47670000000
1!
b1001 %
1'
b1001 +
#47680000000
0!
0'
#47690000000
1!
b0 %
1'
b0 +
#47700000000
0!
0'
#47710000000
1!
1$
b1 %
1'
1*
b1 +
#47720000000
0!
0'
#47730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#47740000000
0!
0'
#47750000000
1!
b11 %
1'
b11 +
#47760000000
0!
0'
#47770000000
1!
b100 %
1'
b100 +
#47780000000
0!
0'
#47790000000
1!
b101 %
1'
b101 +
#47800000000
0!
0'
#47810000000
1!
0$
b110 %
1'
0*
b110 +
#47820000000
0!
0'
#47830000000
1!
b111 %
1'
b111 +
#47840000000
0!
0'
#47850000000
1!
b1000 %
1'
b1000 +
#47860000000
0!
0'
#47870000000
1!
b1001 %
1'
b1001 +
#47880000000
0!
0'
#47890000000
1!
b0 %
1'
b0 +
#47900000000
0!
0'
#47910000000
1!
1$
b1 %
1'
1*
b1 +
#47920000000
0!
0'
#47930000000
1!
b10 %
1'
b10 +
#47940000000
1"
1(
#47950000000
0!
0"
b100 &
0'
0(
b100 ,
#47960000000
1!
b11 %
1'
b11 +
#47970000000
0!
0'
#47980000000
1!
b100 %
1'
b100 +
#47990000000
0!
0'
#48000000000
1!
b101 %
1'
b101 +
#48010000000
0!
0'
#48020000000
1!
b110 %
1'
b110 +
#48030000000
0!
0'
#48040000000
1!
b111 %
1'
b111 +
#48050000000
0!
0'
#48060000000
1!
0$
b1000 %
1'
0*
b1000 +
#48070000000
0!
0'
#48080000000
1!
b1001 %
1'
b1001 +
#48090000000
0!
0'
#48100000000
1!
b0 %
1'
b0 +
#48110000000
0!
0'
#48120000000
1!
1$
b1 %
1'
1*
b1 +
#48130000000
0!
0'
#48140000000
1!
b10 %
1'
b10 +
#48150000000
0!
0'
#48160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#48170000000
0!
0'
#48180000000
1!
b100 %
1'
b100 +
#48190000000
0!
0'
#48200000000
1!
b101 %
1'
b101 +
#48210000000
0!
0'
#48220000000
1!
0$
b110 %
1'
0*
b110 +
#48230000000
0!
0'
#48240000000
1!
b111 %
1'
b111 +
#48250000000
0!
0'
#48260000000
1!
b1000 %
1'
b1000 +
#48270000000
0!
0'
#48280000000
1!
b1001 %
1'
b1001 +
#48290000000
0!
0'
#48300000000
1!
b0 %
1'
b0 +
#48310000000
0!
0'
#48320000000
1!
1$
b1 %
1'
1*
b1 +
#48330000000
0!
0'
#48340000000
1!
b10 %
1'
b10 +
#48350000000
0!
0'
#48360000000
1!
b11 %
1'
b11 +
#48370000000
1"
1(
#48380000000
0!
0"
b100 &
0'
0(
b100 ,
#48390000000
1!
b100 %
1'
b100 +
#48400000000
0!
0'
#48410000000
1!
b101 %
1'
b101 +
#48420000000
0!
0'
#48430000000
1!
b110 %
1'
b110 +
#48440000000
0!
0'
#48450000000
1!
b111 %
1'
b111 +
#48460000000
0!
0'
#48470000000
1!
0$
b1000 %
1'
0*
b1000 +
#48480000000
0!
0'
#48490000000
1!
b1001 %
1'
b1001 +
#48500000000
0!
0'
#48510000000
1!
b0 %
1'
b0 +
#48520000000
0!
0'
#48530000000
1!
1$
b1 %
1'
1*
b1 +
#48540000000
0!
0'
#48550000000
1!
b10 %
1'
b10 +
#48560000000
0!
0'
#48570000000
1!
b11 %
1'
b11 +
#48580000000
0!
0'
#48590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#48600000000
0!
0'
#48610000000
1!
b101 %
1'
b101 +
#48620000000
0!
0'
#48630000000
1!
0$
b110 %
1'
0*
b110 +
#48640000000
0!
0'
#48650000000
1!
b111 %
1'
b111 +
#48660000000
0!
0'
#48670000000
1!
b1000 %
1'
b1000 +
#48680000000
0!
0'
#48690000000
1!
b1001 %
1'
b1001 +
#48700000000
0!
0'
#48710000000
1!
b0 %
1'
b0 +
#48720000000
0!
0'
#48730000000
1!
1$
b1 %
1'
1*
b1 +
#48740000000
0!
0'
#48750000000
1!
b10 %
1'
b10 +
#48760000000
0!
0'
#48770000000
1!
b11 %
1'
b11 +
#48780000000
0!
0'
#48790000000
1!
b100 %
1'
b100 +
#48800000000
1"
1(
#48810000000
0!
0"
b100 &
0'
0(
b100 ,
#48820000000
1!
b101 %
1'
b101 +
#48830000000
0!
0'
#48840000000
1!
b110 %
1'
b110 +
#48850000000
0!
0'
#48860000000
1!
b111 %
1'
b111 +
#48870000000
0!
0'
#48880000000
1!
0$
b1000 %
1'
0*
b1000 +
#48890000000
0!
0'
#48900000000
1!
b1001 %
1'
b1001 +
#48910000000
0!
0'
#48920000000
1!
b0 %
1'
b0 +
#48930000000
0!
0'
#48940000000
1!
1$
b1 %
1'
1*
b1 +
#48950000000
0!
0'
#48960000000
1!
b10 %
1'
b10 +
#48970000000
0!
0'
#48980000000
1!
b11 %
1'
b11 +
#48990000000
0!
0'
#49000000000
1!
b100 %
1'
b100 +
#49010000000
0!
0'
#49020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#49030000000
0!
0'
#49040000000
1!
0$
b110 %
1'
0*
b110 +
#49050000000
0!
0'
#49060000000
1!
b111 %
1'
b111 +
#49070000000
0!
0'
#49080000000
1!
b1000 %
1'
b1000 +
#49090000000
0!
0'
#49100000000
1!
b1001 %
1'
b1001 +
#49110000000
0!
0'
#49120000000
1!
b0 %
1'
b0 +
#49130000000
0!
0'
#49140000000
1!
1$
b1 %
1'
1*
b1 +
#49150000000
0!
0'
#49160000000
1!
b10 %
1'
b10 +
#49170000000
0!
0'
#49180000000
1!
b11 %
1'
b11 +
#49190000000
0!
0'
#49200000000
1!
b100 %
1'
b100 +
#49210000000
0!
0'
#49220000000
1!
b101 %
1'
b101 +
#49230000000
1"
1(
#49240000000
0!
0"
b100 &
0'
0(
b100 ,
#49250000000
1!
b110 %
1'
b110 +
#49260000000
0!
0'
#49270000000
1!
b111 %
1'
b111 +
#49280000000
0!
0'
#49290000000
1!
0$
b1000 %
1'
0*
b1000 +
#49300000000
0!
0'
#49310000000
1!
b1001 %
1'
b1001 +
#49320000000
0!
0'
#49330000000
1!
b0 %
1'
b0 +
#49340000000
0!
0'
#49350000000
1!
1$
b1 %
1'
1*
b1 +
#49360000000
0!
0'
#49370000000
1!
b10 %
1'
b10 +
#49380000000
0!
0'
#49390000000
1!
b11 %
1'
b11 +
#49400000000
0!
0'
#49410000000
1!
b100 %
1'
b100 +
#49420000000
0!
0'
#49430000000
1!
b101 %
1'
b101 +
#49440000000
0!
0'
#49450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#49460000000
0!
0'
#49470000000
1!
b111 %
1'
b111 +
#49480000000
0!
0'
#49490000000
1!
b1000 %
1'
b1000 +
#49500000000
0!
0'
#49510000000
1!
b1001 %
1'
b1001 +
#49520000000
0!
0'
#49530000000
1!
b0 %
1'
b0 +
#49540000000
0!
0'
#49550000000
1!
1$
b1 %
1'
1*
b1 +
#49560000000
0!
0'
#49570000000
1!
b10 %
1'
b10 +
#49580000000
0!
0'
#49590000000
1!
b11 %
1'
b11 +
#49600000000
0!
0'
#49610000000
1!
b100 %
1'
b100 +
#49620000000
0!
0'
#49630000000
1!
b101 %
1'
b101 +
#49640000000
0!
0'
#49650000000
1!
0$
b110 %
1'
0*
b110 +
#49660000000
1"
1(
#49670000000
0!
0"
b100 &
0'
0(
b100 ,
#49680000000
1!
1$
b111 %
1'
1*
b111 +
#49690000000
0!
0'
#49700000000
1!
0$
b1000 %
1'
0*
b1000 +
#49710000000
0!
0'
#49720000000
1!
b1001 %
1'
b1001 +
#49730000000
0!
0'
#49740000000
1!
b0 %
1'
b0 +
#49750000000
0!
0'
#49760000000
1!
1$
b1 %
1'
1*
b1 +
#49770000000
0!
0'
#49780000000
1!
b10 %
1'
b10 +
#49790000000
0!
0'
#49800000000
1!
b11 %
1'
b11 +
#49810000000
0!
0'
#49820000000
1!
b100 %
1'
b100 +
#49830000000
0!
0'
#49840000000
1!
b101 %
1'
b101 +
#49850000000
0!
0'
#49860000000
1!
b110 %
1'
b110 +
#49870000000
0!
0'
#49880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#49890000000
0!
0'
#49900000000
1!
b1000 %
1'
b1000 +
#49910000000
0!
0'
#49920000000
1!
b1001 %
1'
b1001 +
#49930000000
0!
0'
#49940000000
1!
b0 %
1'
b0 +
#49950000000
0!
0'
#49960000000
1!
1$
b1 %
1'
1*
b1 +
#49970000000
0!
0'
#49980000000
1!
b10 %
1'
b10 +
#49990000000
0!
0'
#50000000000
1!
b11 %
1'
b11 +
#50010000000
0!
0'
#50020000000
1!
b100 %
1'
b100 +
#50030000000
0!
0'
#50040000000
1!
b101 %
1'
b101 +
#50050000000
0!
0'
#50060000000
1!
0$
b110 %
1'
0*
b110 +
#50070000000
0!
0'
#50080000000
1!
b111 %
1'
b111 +
#50090000000
1"
1(
#50100000000
0!
0"
b100 &
0'
0(
b100 ,
#50110000000
1!
b1000 %
1'
b1000 +
#50120000000
0!
0'
#50130000000
1!
b1001 %
1'
b1001 +
#50140000000
0!
0'
#50150000000
1!
b0 %
1'
b0 +
#50160000000
0!
0'
#50170000000
1!
1$
b1 %
1'
1*
b1 +
#50180000000
0!
0'
#50190000000
1!
b10 %
1'
b10 +
#50200000000
0!
0'
#50210000000
1!
b11 %
1'
b11 +
#50220000000
0!
0'
#50230000000
1!
b100 %
1'
b100 +
#50240000000
0!
0'
#50250000000
1!
b101 %
1'
b101 +
#50260000000
0!
0'
#50270000000
1!
b110 %
1'
b110 +
#50280000000
0!
0'
#50290000000
1!
b111 %
1'
b111 +
#50300000000
0!
0'
#50310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#50320000000
0!
0'
#50330000000
1!
b1001 %
1'
b1001 +
#50340000000
0!
0'
#50350000000
1!
b0 %
1'
b0 +
#50360000000
0!
0'
#50370000000
1!
1$
b1 %
1'
1*
b1 +
#50380000000
0!
0'
#50390000000
1!
b10 %
1'
b10 +
#50400000000
0!
0'
#50410000000
1!
b11 %
1'
b11 +
#50420000000
0!
0'
#50430000000
1!
b100 %
1'
b100 +
#50440000000
0!
0'
#50450000000
1!
b101 %
1'
b101 +
#50460000000
0!
0'
#50470000000
1!
0$
b110 %
1'
0*
b110 +
#50480000000
0!
0'
#50490000000
1!
b111 %
1'
b111 +
#50500000000
0!
0'
#50510000000
1!
b1000 %
1'
b1000 +
#50520000000
1"
1(
#50530000000
0!
0"
b100 &
0'
0(
b100 ,
#50540000000
1!
b1001 %
1'
b1001 +
#50550000000
0!
0'
#50560000000
1!
b0 %
1'
b0 +
#50570000000
0!
0'
#50580000000
1!
1$
b1 %
1'
1*
b1 +
#50590000000
0!
0'
#50600000000
1!
b10 %
1'
b10 +
#50610000000
0!
0'
#50620000000
1!
b11 %
1'
b11 +
#50630000000
0!
0'
#50640000000
1!
b100 %
1'
b100 +
#50650000000
0!
0'
#50660000000
1!
b101 %
1'
b101 +
#50670000000
0!
0'
#50680000000
1!
b110 %
1'
b110 +
#50690000000
0!
0'
#50700000000
1!
b111 %
1'
b111 +
#50710000000
0!
0'
#50720000000
1!
0$
b1000 %
1'
0*
b1000 +
#50730000000
0!
0'
#50740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#50750000000
0!
0'
#50760000000
1!
b0 %
1'
b0 +
#50770000000
0!
0'
#50780000000
1!
1$
b1 %
1'
1*
b1 +
#50790000000
0!
0'
#50800000000
1!
b10 %
1'
b10 +
#50810000000
0!
0'
#50820000000
1!
b11 %
1'
b11 +
#50830000000
0!
0'
#50840000000
1!
b100 %
1'
b100 +
#50850000000
0!
0'
#50860000000
1!
b101 %
1'
b101 +
#50870000000
0!
0'
#50880000000
1!
0$
b110 %
1'
0*
b110 +
#50890000000
0!
0'
#50900000000
1!
b111 %
1'
b111 +
#50910000000
0!
0'
#50920000000
1!
b1000 %
1'
b1000 +
#50930000000
0!
0'
#50940000000
1!
b1001 %
1'
b1001 +
#50950000000
1"
1(
#50960000000
0!
0"
b100 &
0'
0(
b100 ,
#50970000000
1!
b0 %
1'
b0 +
#50980000000
0!
0'
#50990000000
1!
1$
b1 %
1'
1*
b1 +
#51000000000
0!
0'
#51010000000
1!
b10 %
1'
b10 +
#51020000000
0!
0'
#51030000000
1!
b11 %
1'
b11 +
#51040000000
0!
0'
#51050000000
1!
b100 %
1'
b100 +
#51060000000
0!
0'
#51070000000
1!
b101 %
1'
b101 +
#51080000000
0!
0'
#51090000000
1!
b110 %
1'
b110 +
#51100000000
0!
0'
#51110000000
1!
b111 %
1'
b111 +
#51120000000
0!
0'
#51130000000
1!
0$
b1000 %
1'
0*
b1000 +
#51140000000
0!
0'
#51150000000
1!
b1001 %
1'
b1001 +
#51160000000
0!
0'
#51170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#51180000000
0!
0'
#51190000000
1!
1$
b1 %
1'
1*
b1 +
#51200000000
0!
0'
#51210000000
1!
b10 %
1'
b10 +
#51220000000
0!
0'
#51230000000
1!
b11 %
1'
b11 +
#51240000000
0!
0'
#51250000000
1!
b100 %
1'
b100 +
#51260000000
0!
0'
#51270000000
1!
b101 %
1'
b101 +
#51280000000
0!
0'
#51290000000
1!
0$
b110 %
1'
0*
b110 +
#51300000000
0!
0'
#51310000000
1!
b111 %
1'
b111 +
#51320000000
0!
0'
#51330000000
1!
b1000 %
1'
b1000 +
#51340000000
0!
0'
#51350000000
1!
b1001 %
1'
b1001 +
#51360000000
0!
0'
#51370000000
1!
b0 %
1'
b0 +
#51380000000
1"
1(
#51390000000
0!
0"
b100 &
0'
0(
b100 ,
#51400000000
1!
1$
b1 %
1'
1*
b1 +
#51410000000
0!
0'
#51420000000
1!
b10 %
1'
b10 +
#51430000000
0!
0'
#51440000000
1!
b11 %
1'
b11 +
#51450000000
0!
0'
#51460000000
1!
b100 %
1'
b100 +
#51470000000
0!
0'
#51480000000
1!
b101 %
1'
b101 +
#51490000000
0!
0'
#51500000000
1!
b110 %
1'
b110 +
#51510000000
0!
0'
#51520000000
1!
b111 %
1'
b111 +
#51530000000
0!
0'
#51540000000
1!
0$
b1000 %
1'
0*
b1000 +
#51550000000
0!
0'
#51560000000
1!
b1001 %
1'
b1001 +
#51570000000
0!
0'
#51580000000
1!
b0 %
1'
b0 +
#51590000000
0!
0'
#51600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#51610000000
0!
0'
#51620000000
1!
b10 %
1'
b10 +
#51630000000
0!
0'
#51640000000
1!
b11 %
1'
b11 +
#51650000000
0!
0'
#51660000000
1!
b100 %
1'
b100 +
#51670000000
0!
0'
#51680000000
1!
b101 %
1'
b101 +
#51690000000
0!
0'
#51700000000
1!
0$
b110 %
1'
0*
b110 +
#51710000000
0!
0'
#51720000000
1!
b111 %
1'
b111 +
#51730000000
0!
0'
#51740000000
1!
b1000 %
1'
b1000 +
#51750000000
0!
0'
#51760000000
1!
b1001 %
1'
b1001 +
#51770000000
0!
0'
#51780000000
1!
b0 %
1'
b0 +
#51790000000
0!
0'
#51800000000
1!
1$
b1 %
1'
1*
b1 +
#51810000000
1"
1(
#51820000000
0!
0"
b100 &
0'
0(
b100 ,
#51830000000
1!
b10 %
1'
b10 +
#51840000000
0!
0'
#51850000000
1!
b11 %
1'
b11 +
#51860000000
0!
0'
#51870000000
1!
b100 %
1'
b100 +
#51880000000
0!
0'
#51890000000
1!
b101 %
1'
b101 +
#51900000000
0!
0'
#51910000000
1!
b110 %
1'
b110 +
#51920000000
0!
0'
#51930000000
1!
b111 %
1'
b111 +
#51940000000
0!
0'
#51950000000
1!
0$
b1000 %
1'
0*
b1000 +
#51960000000
0!
0'
#51970000000
1!
b1001 %
1'
b1001 +
#51980000000
0!
0'
#51990000000
1!
b0 %
1'
b0 +
#52000000000
0!
0'
#52010000000
1!
1$
b1 %
1'
1*
b1 +
#52020000000
0!
0'
#52030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#52040000000
0!
0'
#52050000000
1!
b11 %
1'
b11 +
#52060000000
0!
0'
#52070000000
1!
b100 %
1'
b100 +
#52080000000
0!
0'
#52090000000
1!
b101 %
1'
b101 +
#52100000000
0!
0'
#52110000000
1!
0$
b110 %
1'
0*
b110 +
#52120000000
0!
0'
#52130000000
1!
b111 %
1'
b111 +
#52140000000
0!
0'
#52150000000
1!
b1000 %
1'
b1000 +
#52160000000
0!
0'
#52170000000
1!
b1001 %
1'
b1001 +
#52180000000
0!
0'
#52190000000
1!
b0 %
1'
b0 +
#52200000000
0!
0'
#52210000000
1!
1$
b1 %
1'
1*
b1 +
#52220000000
0!
0'
#52230000000
1!
b10 %
1'
b10 +
#52240000000
1"
1(
#52250000000
0!
0"
b100 &
0'
0(
b100 ,
#52260000000
1!
b11 %
1'
b11 +
#52270000000
0!
0'
#52280000000
1!
b100 %
1'
b100 +
#52290000000
0!
0'
#52300000000
1!
b101 %
1'
b101 +
#52310000000
0!
0'
#52320000000
1!
b110 %
1'
b110 +
#52330000000
0!
0'
#52340000000
1!
b111 %
1'
b111 +
#52350000000
0!
0'
#52360000000
1!
0$
b1000 %
1'
0*
b1000 +
#52370000000
0!
0'
#52380000000
1!
b1001 %
1'
b1001 +
#52390000000
0!
0'
#52400000000
1!
b0 %
1'
b0 +
#52410000000
0!
0'
#52420000000
1!
1$
b1 %
1'
1*
b1 +
#52430000000
0!
0'
#52440000000
1!
b10 %
1'
b10 +
#52450000000
0!
0'
#52460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#52470000000
0!
0'
#52480000000
1!
b100 %
1'
b100 +
#52490000000
0!
0'
#52500000000
1!
b101 %
1'
b101 +
#52510000000
0!
0'
#52520000000
1!
0$
b110 %
1'
0*
b110 +
#52530000000
0!
0'
#52540000000
1!
b111 %
1'
b111 +
#52550000000
0!
0'
#52560000000
1!
b1000 %
1'
b1000 +
#52570000000
0!
0'
#52580000000
1!
b1001 %
1'
b1001 +
#52590000000
0!
0'
#52600000000
1!
b0 %
1'
b0 +
#52610000000
0!
0'
#52620000000
1!
1$
b1 %
1'
1*
b1 +
#52630000000
0!
0'
#52640000000
1!
b10 %
1'
b10 +
#52650000000
0!
0'
#52660000000
1!
b11 %
1'
b11 +
#52670000000
1"
1(
#52680000000
0!
0"
b100 &
0'
0(
b100 ,
#52690000000
1!
b100 %
1'
b100 +
#52700000000
0!
0'
#52710000000
1!
b101 %
1'
b101 +
#52720000000
0!
0'
#52730000000
1!
b110 %
1'
b110 +
#52740000000
0!
0'
#52750000000
1!
b111 %
1'
b111 +
#52760000000
0!
0'
#52770000000
1!
0$
b1000 %
1'
0*
b1000 +
#52780000000
0!
0'
#52790000000
1!
b1001 %
1'
b1001 +
#52800000000
0!
0'
#52810000000
1!
b0 %
1'
b0 +
#52820000000
0!
0'
#52830000000
1!
1$
b1 %
1'
1*
b1 +
#52840000000
0!
0'
#52850000000
1!
b10 %
1'
b10 +
#52860000000
0!
0'
#52870000000
1!
b11 %
1'
b11 +
#52880000000
0!
0'
#52890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#52900000000
0!
0'
#52910000000
1!
b101 %
1'
b101 +
#52920000000
0!
0'
#52930000000
1!
0$
b110 %
1'
0*
b110 +
#52940000000
0!
0'
#52950000000
1!
b111 %
1'
b111 +
#52960000000
0!
0'
#52970000000
1!
b1000 %
1'
b1000 +
#52980000000
0!
0'
#52990000000
1!
b1001 %
1'
b1001 +
#53000000000
0!
0'
#53010000000
1!
b0 %
1'
b0 +
#53020000000
0!
0'
#53030000000
1!
1$
b1 %
1'
1*
b1 +
#53040000000
0!
0'
#53050000000
1!
b10 %
1'
b10 +
#53060000000
0!
0'
#53070000000
1!
b11 %
1'
b11 +
#53080000000
0!
0'
#53090000000
1!
b100 %
1'
b100 +
#53100000000
1"
1(
#53110000000
0!
0"
b100 &
0'
0(
b100 ,
#53120000000
1!
b101 %
1'
b101 +
#53130000000
0!
0'
#53140000000
1!
b110 %
1'
b110 +
#53150000000
0!
0'
#53160000000
1!
b111 %
1'
b111 +
#53170000000
0!
0'
#53180000000
1!
0$
b1000 %
1'
0*
b1000 +
#53190000000
0!
0'
#53200000000
1!
b1001 %
1'
b1001 +
#53210000000
0!
0'
#53220000000
1!
b0 %
1'
b0 +
#53230000000
0!
0'
#53240000000
1!
1$
b1 %
1'
1*
b1 +
#53250000000
0!
0'
#53260000000
1!
b10 %
1'
b10 +
#53270000000
0!
0'
#53280000000
1!
b11 %
1'
b11 +
#53290000000
0!
0'
#53300000000
1!
b100 %
1'
b100 +
#53310000000
0!
0'
#53320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#53330000000
0!
0'
#53340000000
1!
0$
b110 %
1'
0*
b110 +
#53350000000
0!
0'
#53360000000
1!
b111 %
1'
b111 +
#53370000000
0!
0'
#53380000000
1!
b1000 %
1'
b1000 +
#53390000000
0!
0'
#53400000000
1!
b1001 %
1'
b1001 +
#53410000000
0!
0'
#53420000000
1!
b0 %
1'
b0 +
#53430000000
0!
0'
#53440000000
1!
1$
b1 %
1'
1*
b1 +
#53450000000
0!
0'
#53460000000
1!
b10 %
1'
b10 +
#53470000000
0!
0'
#53480000000
1!
b11 %
1'
b11 +
#53490000000
0!
0'
#53500000000
1!
b100 %
1'
b100 +
#53510000000
0!
0'
#53520000000
1!
b101 %
1'
b101 +
#53530000000
1"
1(
#53540000000
0!
0"
b100 &
0'
0(
b100 ,
#53550000000
1!
b110 %
1'
b110 +
#53560000000
0!
0'
#53570000000
1!
b111 %
1'
b111 +
#53580000000
0!
0'
#53590000000
1!
0$
b1000 %
1'
0*
b1000 +
#53600000000
0!
0'
#53610000000
1!
b1001 %
1'
b1001 +
#53620000000
0!
0'
#53630000000
1!
b0 %
1'
b0 +
#53640000000
0!
0'
#53650000000
1!
1$
b1 %
1'
1*
b1 +
#53660000000
0!
0'
#53670000000
1!
b10 %
1'
b10 +
#53680000000
0!
0'
#53690000000
1!
b11 %
1'
b11 +
#53700000000
0!
0'
#53710000000
1!
b100 %
1'
b100 +
#53720000000
0!
0'
#53730000000
1!
b101 %
1'
b101 +
#53740000000
0!
0'
#53750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#53760000000
0!
0'
#53770000000
1!
b111 %
1'
b111 +
#53780000000
0!
0'
#53790000000
1!
b1000 %
1'
b1000 +
#53800000000
0!
0'
#53810000000
1!
b1001 %
1'
b1001 +
#53820000000
0!
0'
#53830000000
1!
b0 %
1'
b0 +
#53840000000
0!
0'
#53850000000
1!
1$
b1 %
1'
1*
b1 +
#53860000000
0!
0'
#53870000000
1!
b10 %
1'
b10 +
#53880000000
0!
0'
#53890000000
1!
b11 %
1'
b11 +
#53900000000
0!
0'
#53910000000
1!
b100 %
1'
b100 +
#53920000000
0!
0'
#53930000000
1!
b101 %
1'
b101 +
#53940000000
0!
0'
#53950000000
1!
0$
b110 %
1'
0*
b110 +
#53960000000
1"
1(
#53970000000
0!
0"
b100 &
0'
0(
b100 ,
#53980000000
1!
1$
b111 %
1'
1*
b111 +
#53990000000
0!
0'
#54000000000
1!
0$
b1000 %
1'
0*
b1000 +
#54010000000
0!
0'
#54020000000
1!
b1001 %
1'
b1001 +
#54030000000
0!
0'
#54040000000
1!
b0 %
1'
b0 +
#54050000000
0!
0'
#54060000000
1!
1$
b1 %
1'
1*
b1 +
#54070000000
0!
0'
#54080000000
1!
b10 %
1'
b10 +
#54090000000
0!
0'
#54100000000
1!
b11 %
1'
b11 +
#54110000000
0!
0'
#54120000000
1!
b100 %
1'
b100 +
#54130000000
0!
0'
#54140000000
1!
b101 %
1'
b101 +
#54150000000
0!
0'
#54160000000
1!
b110 %
1'
b110 +
#54170000000
0!
0'
#54180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#54190000000
0!
0'
#54200000000
1!
b1000 %
1'
b1000 +
#54210000000
0!
0'
#54220000000
1!
b1001 %
1'
b1001 +
#54230000000
0!
0'
#54240000000
1!
b0 %
1'
b0 +
#54250000000
0!
0'
#54260000000
1!
1$
b1 %
1'
1*
b1 +
#54270000000
0!
0'
#54280000000
1!
b10 %
1'
b10 +
#54290000000
0!
0'
#54300000000
1!
b11 %
1'
b11 +
#54310000000
0!
0'
#54320000000
1!
b100 %
1'
b100 +
#54330000000
0!
0'
#54340000000
1!
b101 %
1'
b101 +
#54350000000
0!
0'
#54360000000
1!
0$
b110 %
1'
0*
b110 +
#54370000000
0!
0'
#54380000000
1!
b111 %
1'
b111 +
#54390000000
1"
1(
#54400000000
0!
0"
b100 &
0'
0(
b100 ,
#54410000000
1!
b1000 %
1'
b1000 +
#54420000000
0!
0'
#54430000000
1!
b1001 %
1'
b1001 +
#54440000000
0!
0'
#54450000000
1!
b0 %
1'
b0 +
#54460000000
0!
0'
#54470000000
1!
1$
b1 %
1'
1*
b1 +
#54480000000
0!
0'
#54490000000
1!
b10 %
1'
b10 +
#54500000000
0!
0'
#54510000000
1!
b11 %
1'
b11 +
#54520000000
0!
0'
#54530000000
1!
b100 %
1'
b100 +
#54540000000
0!
0'
#54550000000
1!
b101 %
1'
b101 +
#54560000000
0!
0'
#54570000000
1!
b110 %
1'
b110 +
#54580000000
0!
0'
#54590000000
1!
b111 %
1'
b111 +
#54600000000
0!
0'
#54610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#54620000000
0!
0'
#54630000000
1!
b1001 %
1'
b1001 +
#54640000000
0!
0'
#54650000000
1!
b0 %
1'
b0 +
#54660000000
0!
0'
#54670000000
1!
1$
b1 %
1'
1*
b1 +
#54680000000
0!
0'
#54690000000
1!
b10 %
1'
b10 +
#54700000000
0!
0'
#54710000000
1!
b11 %
1'
b11 +
#54720000000
0!
0'
#54730000000
1!
b100 %
1'
b100 +
#54740000000
0!
0'
#54750000000
1!
b101 %
1'
b101 +
#54760000000
0!
0'
#54770000000
1!
0$
b110 %
1'
0*
b110 +
#54780000000
0!
0'
#54790000000
1!
b111 %
1'
b111 +
#54800000000
0!
0'
#54810000000
1!
b1000 %
1'
b1000 +
#54820000000
1"
1(
#54830000000
0!
0"
b100 &
0'
0(
b100 ,
#54840000000
1!
b1001 %
1'
b1001 +
#54850000000
0!
0'
#54860000000
1!
b0 %
1'
b0 +
#54870000000
0!
0'
#54880000000
1!
1$
b1 %
1'
1*
b1 +
#54890000000
0!
0'
#54900000000
1!
b10 %
1'
b10 +
#54910000000
0!
0'
#54920000000
1!
b11 %
1'
b11 +
#54930000000
0!
0'
#54940000000
1!
b100 %
1'
b100 +
#54950000000
0!
0'
#54960000000
1!
b101 %
1'
b101 +
#54970000000
0!
0'
#54980000000
1!
b110 %
1'
b110 +
#54990000000
0!
0'
#55000000000
1!
b111 %
1'
b111 +
#55010000000
0!
0'
#55020000000
1!
0$
b1000 %
1'
0*
b1000 +
#55030000000
0!
0'
#55040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#55050000000
0!
0'
#55060000000
1!
b0 %
1'
b0 +
#55070000000
0!
0'
#55080000000
1!
1$
b1 %
1'
1*
b1 +
#55090000000
0!
0'
#55100000000
1!
b10 %
1'
b10 +
#55110000000
0!
0'
#55120000000
1!
b11 %
1'
b11 +
#55130000000
0!
0'
#55140000000
1!
b100 %
1'
b100 +
#55150000000
0!
0'
#55160000000
1!
b101 %
1'
b101 +
#55170000000
0!
0'
#55180000000
1!
0$
b110 %
1'
0*
b110 +
#55190000000
0!
0'
#55200000000
1!
b111 %
1'
b111 +
#55210000000
0!
0'
#55220000000
1!
b1000 %
1'
b1000 +
#55230000000
0!
0'
#55240000000
1!
b1001 %
1'
b1001 +
#55250000000
1"
1(
#55260000000
0!
0"
b100 &
0'
0(
b100 ,
#55270000000
1!
b0 %
1'
b0 +
#55280000000
0!
0'
#55290000000
1!
1$
b1 %
1'
1*
b1 +
#55300000000
0!
0'
#55310000000
1!
b10 %
1'
b10 +
#55320000000
0!
0'
#55330000000
1!
b11 %
1'
b11 +
#55340000000
0!
0'
#55350000000
1!
b100 %
1'
b100 +
#55360000000
0!
0'
#55370000000
1!
b101 %
1'
b101 +
#55380000000
0!
0'
#55390000000
1!
b110 %
1'
b110 +
#55400000000
0!
0'
#55410000000
1!
b111 %
1'
b111 +
#55420000000
0!
0'
#55430000000
1!
0$
b1000 %
1'
0*
b1000 +
#55440000000
0!
0'
#55450000000
1!
b1001 %
1'
b1001 +
#55460000000
0!
0'
#55470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#55480000000
0!
0'
#55490000000
1!
1$
b1 %
1'
1*
b1 +
#55500000000
0!
0'
#55510000000
1!
b10 %
1'
b10 +
#55520000000
0!
0'
#55530000000
1!
b11 %
1'
b11 +
#55540000000
0!
0'
#55550000000
1!
b100 %
1'
b100 +
#55560000000
0!
0'
#55570000000
1!
b101 %
1'
b101 +
#55580000000
0!
0'
#55590000000
1!
0$
b110 %
1'
0*
b110 +
#55600000000
0!
0'
#55610000000
1!
b111 %
1'
b111 +
#55620000000
0!
0'
#55630000000
1!
b1000 %
1'
b1000 +
#55640000000
0!
0'
#55650000000
1!
b1001 %
1'
b1001 +
#55660000000
0!
0'
#55670000000
1!
b0 %
1'
b0 +
#55680000000
1"
1(
#55690000000
0!
0"
b100 &
0'
0(
b100 ,
#55700000000
1!
1$
b1 %
1'
1*
b1 +
#55710000000
0!
0'
#55720000000
1!
b10 %
1'
b10 +
#55730000000
0!
0'
#55740000000
1!
b11 %
1'
b11 +
#55750000000
0!
0'
#55760000000
1!
b100 %
1'
b100 +
#55770000000
0!
0'
#55780000000
1!
b101 %
1'
b101 +
#55790000000
0!
0'
#55800000000
1!
b110 %
1'
b110 +
#55810000000
0!
0'
#55820000000
1!
b111 %
1'
b111 +
#55830000000
0!
0'
#55840000000
1!
0$
b1000 %
1'
0*
b1000 +
#55850000000
0!
0'
#55860000000
1!
b1001 %
1'
b1001 +
#55870000000
0!
0'
#55880000000
1!
b0 %
1'
b0 +
#55890000000
0!
0'
#55900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#55910000000
0!
0'
#55920000000
1!
b10 %
1'
b10 +
#55930000000
0!
0'
#55940000000
1!
b11 %
1'
b11 +
#55950000000
0!
0'
#55960000000
1!
b100 %
1'
b100 +
#55970000000
0!
0'
#55980000000
1!
b101 %
1'
b101 +
#55990000000
0!
0'
#56000000000
1!
0$
b110 %
1'
0*
b110 +
#56010000000
0!
0'
#56020000000
1!
b111 %
1'
b111 +
#56030000000
0!
0'
#56040000000
1!
b1000 %
1'
b1000 +
#56050000000
0!
0'
#56060000000
1!
b1001 %
1'
b1001 +
#56070000000
0!
0'
#56080000000
1!
b0 %
1'
b0 +
#56090000000
0!
0'
#56100000000
1!
1$
b1 %
1'
1*
b1 +
#56110000000
1"
1(
#56120000000
0!
0"
b100 &
0'
0(
b100 ,
#56130000000
1!
b10 %
1'
b10 +
#56140000000
0!
0'
#56150000000
1!
b11 %
1'
b11 +
#56160000000
0!
0'
#56170000000
1!
b100 %
1'
b100 +
#56180000000
0!
0'
#56190000000
1!
b101 %
1'
b101 +
#56200000000
0!
0'
#56210000000
1!
b110 %
1'
b110 +
#56220000000
0!
0'
#56230000000
1!
b111 %
1'
b111 +
#56240000000
0!
0'
#56250000000
1!
0$
b1000 %
1'
0*
b1000 +
#56260000000
0!
0'
#56270000000
1!
b1001 %
1'
b1001 +
#56280000000
0!
0'
#56290000000
1!
b0 %
1'
b0 +
#56300000000
0!
0'
#56310000000
1!
1$
b1 %
1'
1*
b1 +
#56320000000
0!
0'
#56330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#56340000000
0!
0'
#56350000000
1!
b11 %
1'
b11 +
#56360000000
0!
0'
#56370000000
1!
b100 %
1'
b100 +
#56380000000
0!
0'
#56390000000
1!
b101 %
1'
b101 +
#56400000000
0!
0'
#56410000000
1!
0$
b110 %
1'
0*
b110 +
#56420000000
0!
0'
#56430000000
1!
b111 %
1'
b111 +
#56440000000
0!
0'
#56450000000
1!
b1000 %
1'
b1000 +
#56460000000
0!
0'
#56470000000
1!
b1001 %
1'
b1001 +
#56480000000
0!
0'
#56490000000
1!
b0 %
1'
b0 +
#56500000000
0!
0'
#56510000000
1!
1$
b1 %
1'
1*
b1 +
#56520000000
0!
0'
#56530000000
1!
b10 %
1'
b10 +
#56540000000
1"
1(
#56550000000
0!
0"
b100 &
0'
0(
b100 ,
#56560000000
1!
b11 %
1'
b11 +
#56570000000
0!
0'
#56580000000
1!
b100 %
1'
b100 +
#56590000000
0!
0'
#56600000000
1!
b101 %
1'
b101 +
#56610000000
0!
0'
#56620000000
1!
b110 %
1'
b110 +
#56630000000
0!
0'
#56640000000
1!
b111 %
1'
b111 +
#56650000000
0!
0'
#56660000000
1!
0$
b1000 %
1'
0*
b1000 +
#56670000000
0!
0'
#56680000000
1!
b1001 %
1'
b1001 +
#56690000000
0!
0'
#56700000000
1!
b0 %
1'
b0 +
#56710000000
0!
0'
#56720000000
1!
1$
b1 %
1'
1*
b1 +
#56730000000
0!
0'
#56740000000
1!
b10 %
1'
b10 +
#56750000000
0!
0'
#56760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#56770000000
0!
0'
#56780000000
1!
b100 %
1'
b100 +
#56790000000
0!
0'
#56800000000
1!
b101 %
1'
b101 +
#56810000000
0!
0'
#56820000000
1!
0$
b110 %
1'
0*
b110 +
#56830000000
0!
0'
#56840000000
1!
b111 %
1'
b111 +
#56850000000
0!
0'
#56860000000
1!
b1000 %
1'
b1000 +
#56870000000
0!
0'
#56880000000
1!
b1001 %
1'
b1001 +
#56890000000
0!
0'
#56900000000
1!
b0 %
1'
b0 +
#56910000000
0!
0'
#56920000000
1!
1$
b1 %
1'
1*
b1 +
#56930000000
0!
0'
#56940000000
1!
b10 %
1'
b10 +
#56950000000
0!
0'
#56960000000
1!
b11 %
1'
b11 +
#56970000000
1"
1(
#56980000000
0!
0"
b100 &
0'
0(
b100 ,
#56990000000
1!
b100 %
1'
b100 +
#57000000000
0!
0'
#57010000000
1!
b101 %
1'
b101 +
#57020000000
0!
0'
#57030000000
1!
b110 %
1'
b110 +
#57040000000
0!
0'
#57050000000
1!
b111 %
1'
b111 +
#57060000000
0!
0'
#57070000000
1!
0$
b1000 %
1'
0*
b1000 +
#57080000000
0!
0'
#57090000000
1!
b1001 %
1'
b1001 +
#57100000000
0!
0'
#57110000000
1!
b0 %
1'
b0 +
#57120000000
0!
0'
#57130000000
1!
1$
b1 %
1'
1*
b1 +
#57140000000
0!
0'
#57150000000
1!
b10 %
1'
b10 +
#57160000000
0!
0'
#57170000000
1!
b11 %
1'
b11 +
#57180000000
0!
0'
#57190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#57200000000
0!
0'
#57210000000
1!
b101 %
1'
b101 +
#57220000000
0!
0'
#57230000000
1!
0$
b110 %
1'
0*
b110 +
#57240000000
0!
0'
#57250000000
1!
b111 %
1'
b111 +
#57260000000
0!
0'
#57270000000
1!
b1000 %
1'
b1000 +
#57280000000
0!
0'
#57290000000
1!
b1001 %
1'
b1001 +
#57300000000
0!
0'
#57310000000
1!
b0 %
1'
b0 +
#57320000000
0!
0'
#57330000000
1!
1$
b1 %
1'
1*
b1 +
#57340000000
0!
0'
#57350000000
1!
b10 %
1'
b10 +
#57360000000
0!
0'
#57370000000
1!
b11 %
1'
b11 +
#57380000000
0!
0'
#57390000000
1!
b100 %
1'
b100 +
#57400000000
1"
1(
#57410000000
0!
0"
b100 &
0'
0(
b100 ,
#57420000000
1!
b101 %
1'
b101 +
#57430000000
0!
0'
#57440000000
1!
b110 %
1'
b110 +
#57450000000
0!
0'
#57460000000
1!
b111 %
1'
b111 +
#57470000000
0!
0'
#57480000000
1!
0$
b1000 %
1'
0*
b1000 +
#57490000000
0!
0'
#57500000000
1!
b1001 %
1'
b1001 +
#57510000000
0!
0'
#57520000000
1!
b0 %
1'
b0 +
#57530000000
0!
0'
#57540000000
1!
1$
b1 %
1'
1*
b1 +
#57550000000
0!
0'
#57560000000
1!
b10 %
1'
b10 +
#57570000000
0!
0'
#57580000000
1!
b11 %
1'
b11 +
#57590000000
0!
0'
#57600000000
1!
b100 %
1'
b100 +
#57610000000
0!
0'
#57620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#57630000000
0!
0'
#57640000000
1!
0$
b110 %
1'
0*
b110 +
#57650000000
0!
0'
#57660000000
1!
b111 %
1'
b111 +
#57670000000
0!
0'
#57680000000
1!
b1000 %
1'
b1000 +
#57690000000
0!
0'
#57700000000
1!
b1001 %
1'
b1001 +
#57710000000
0!
0'
#57720000000
1!
b0 %
1'
b0 +
#57730000000
0!
0'
#57740000000
1!
1$
b1 %
1'
1*
b1 +
#57750000000
0!
0'
#57760000000
1!
b10 %
1'
b10 +
#57770000000
0!
0'
#57780000000
1!
b11 %
1'
b11 +
#57790000000
0!
0'
#57800000000
1!
b100 %
1'
b100 +
#57810000000
0!
0'
#57820000000
1!
b101 %
1'
b101 +
#57830000000
1"
1(
#57840000000
0!
0"
b100 &
0'
0(
b100 ,
#57850000000
1!
b110 %
1'
b110 +
#57860000000
0!
0'
#57870000000
1!
b111 %
1'
b111 +
#57880000000
0!
0'
#57890000000
1!
0$
b1000 %
1'
0*
b1000 +
#57900000000
0!
0'
#57910000000
1!
b1001 %
1'
b1001 +
#57920000000
0!
0'
#57930000000
1!
b0 %
1'
b0 +
#57940000000
0!
0'
#57950000000
1!
1$
b1 %
1'
1*
b1 +
#57960000000
0!
0'
#57970000000
1!
b10 %
1'
b10 +
#57980000000
0!
0'
#57990000000
1!
b11 %
1'
b11 +
#58000000000
0!
0'
#58010000000
1!
b100 %
1'
b100 +
#58020000000
0!
0'
#58030000000
1!
b101 %
1'
b101 +
#58040000000
0!
0'
#58050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#58060000000
0!
0'
#58070000000
1!
b111 %
1'
b111 +
#58080000000
0!
0'
#58090000000
1!
b1000 %
1'
b1000 +
#58100000000
0!
0'
#58110000000
1!
b1001 %
1'
b1001 +
#58120000000
0!
0'
#58130000000
1!
b0 %
1'
b0 +
#58140000000
0!
0'
#58150000000
1!
1$
b1 %
1'
1*
b1 +
#58160000000
0!
0'
#58170000000
1!
b10 %
1'
b10 +
#58180000000
0!
0'
#58190000000
1!
b11 %
1'
b11 +
#58200000000
0!
0'
#58210000000
1!
b100 %
1'
b100 +
#58220000000
0!
0'
#58230000000
1!
b101 %
1'
b101 +
#58240000000
0!
0'
#58250000000
1!
0$
b110 %
1'
0*
b110 +
#58260000000
1"
1(
#58270000000
0!
0"
b100 &
0'
0(
b100 ,
#58280000000
1!
1$
b111 %
1'
1*
b111 +
#58290000000
0!
0'
#58300000000
1!
0$
b1000 %
1'
0*
b1000 +
#58310000000
0!
0'
#58320000000
1!
b1001 %
1'
b1001 +
#58330000000
0!
0'
#58340000000
1!
b0 %
1'
b0 +
#58350000000
0!
0'
#58360000000
1!
1$
b1 %
1'
1*
b1 +
#58370000000
0!
0'
#58380000000
1!
b10 %
1'
b10 +
#58390000000
0!
0'
#58400000000
1!
b11 %
1'
b11 +
#58410000000
0!
0'
#58420000000
1!
b100 %
1'
b100 +
#58430000000
0!
0'
#58440000000
1!
b101 %
1'
b101 +
#58450000000
0!
0'
#58460000000
1!
b110 %
1'
b110 +
#58470000000
0!
0'
#58480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#58490000000
0!
0'
#58500000000
1!
b1000 %
1'
b1000 +
#58510000000
0!
0'
#58520000000
1!
b1001 %
1'
b1001 +
#58530000000
0!
0'
#58540000000
1!
b0 %
1'
b0 +
#58550000000
0!
0'
#58560000000
1!
1$
b1 %
1'
1*
b1 +
#58570000000
0!
0'
#58580000000
1!
b10 %
1'
b10 +
#58590000000
0!
0'
#58600000000
1!
b11 %
1'
b11 +
#58610000000
0!
0'
#58620000000
1!
b100 %
1'
b100 +
#58630000000
0!
0'
#58640000000
1!
b101 %
1'
b101 +
#58650000000
0!
0'
#58660000000
1!
0$
b110 %
1'
0*
b110 +
#58670000000
0!
0'
#58680000000
1!
b111 %
1'
b111 +
#58690000000
1"
1(
#58700000000
0!
0"
b100 &
0'
0(
b100 ,
#58710000000
1!
b1000 %
1'
b1000 +
#58720000000
0!
0'
#58730000000
1!
b1001 %
1'
b1001 +
#58740000000
0!
0'
#58750000000
1!
b0 %
1'
b0 +
#58760000000
0!
0'
#58770000000
1!
1$
b1 %
1'
1*
b1 +
#58780000000
0!
0'
#58790000000
1!
b10 %
1'
b10 +
#58800000000
0!
0'
#58810000000
1!
b11 %
1'
b11 +
#58820000000
0!
0'
#58830000000
1!
b100 %
1'
b100 +
#58840000000
0!
0'
#58850000000
1!
b101 %
1'
b101 +
#58860000000
0!
0'
#58870000000
1!
b110 %
1'
b110 +
#58880000000
0!
0'
#58890000000
1!
b111 %
1'
b111 +
#58900000000
0!
0'
#58910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#58920000000
0!
0'
#58930000000
1!
b1001 %
1'
b1001 +
#58940000000
0!
0'
#58950000000
1!
b0 %
1'
b0 +
#58960000000
0!
0'
#58970000000
1!
1$
b1 %
1'
1*
b1 +
#58980000000
0!
0'
#58990000000
1!
b10 %
1'
b10 +
#59000000000
0!
0'
#59010000000
1!
b11 %
1'
b11 +
#59020000000
0!
0'
#59030000000
1!
b100 %
1'
b100 +
#59040000000
0!
0'
#59050000000
1!
b101 %
1'
b101 +
#59060000000
0!
0'
#59070000000
1!
0$
b110 %
1'
0*
b110 +
#59080000000
0!
0'
#59090000000
1!
b111 %
1'
b111 +
#59100000000
0!
0'
#59110000000
1!
b1000 %
1'
b1000 +
#59120000000
1"
1(
#59130000000
0!
0"
b100 &
0'
0(
b100 ,
#59140000000
1!
b1001 %
1'
b1001 +
#59150000000
0!
0'
#59160000000
1!
b0 %
1'
b0 +
#59170000000
0!
0'
#59180000000
1!
1$
b1 %
1'
1*
b1 +
#59190000000
0!
0'
#59200000000
1!
b10 %
1'
b10 +
#59210000000
0!
0'
#59220000000
1!
b11 %
1'
b11 +
#59230000000
0!
0'
#59240000000
1!
b100 %
1'
b100 +
#59250000000
0!
0'
#59260000000
1!
b101 %
1'
b101 +
#59270000000
0!
0'
#59280000000
1!
b110 %
1'
b110 +
#59290000000
0!
0'
#59300000000
1!
b111 %
1'
b111 +
#59310000000
0!
0'
#59320000000
1!
0$
b1000 %
1'
0*
b1000 +
#59330000000
0!
0'
#59340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#59350000000
0!
0'
#59360000000
1!
b0 %
1'
b0 +
#59370000000
0!
0'
#59380000000
1!
1$
b1 %
1'
1*
b1 +
#59390000000
0!
0'
#59400000000
1!
b10 %
1'
b10 +
#59410000000
0!
0'
#59420000000
1!
b11 %
1'
b11 +
#59430000000
0!
0'
#59440000000
1!
b100 %
1'
b100 +
#59450000000
0!
0'
#59460000000
1!
b101 %
1'
b101 +
#59470000000
0!
0'
#59480000000
1!
0$
b110 %
1'
0*
b110 +
#59490000000
0!
0'
#59500000000
1!
b111 %
1'
b111 +
#59510000000
0!
0'
#59520000000
1!
b1000 %
1'
b1000 +
#59530000000
0!
0'
#59540000000
1!
b1001 %
1'
b1001 +
#59550000000
1"
1(
#59560000000
0!
0"
b100 &
0'
0(
b100 ,
#59570000000
1!
b0 %
1'
b0 +
#59580000000
0!
0'
#59590000000
1!
1$
b1 %
1'
1*
b1 +
#59600000000
0!
0'
#59610000000
1!
b10 %
1'
b10 +
#59620000000
0!
0'
#59630000000
1!
b11 %
1'
b11 +
#59640000000
0!
0'
#59650000000
1!
b100 %
1'
b100 +
#59660000000
0!
0'
#59670000000
1!
b101 %
1'
b101 +
#59680000000
0!
0'
#59690000000
1!
b110 %
1'
b110 +
#59700000000
0!
0'
#59710000000
1!
b111 %
1'
b111 +
#59720000000
0!
0'
#59730000000
1!
0$
b1000 %
1'
0*
b1000 +
#59740000000
0!
0'
#59750000000
1!
b1001 %
1'
b1001 +
#59760000000
0!
0'
#59770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#59780000000
0!
0'
#59790000000
1!
1$
b1 %
1'
1*
b1 +
#59800000000
0!
0'
#59810000000
1!
b10 %
1'
b10 +
#59820000000
0!
0'
#59830000000
1!
b11 %
1'
b11 +
#59840000000
0!
0'
#59850000000
1!
b100 %
1'
b100 +
#59860000000
0!
0'
#59870000000
1!
b101 %
1'
b101 +
#59880000000
0!
0'
#59890000000
1!
0$
b110 %
1'
0*
b110 +
#59900000000
0!
0'
#59910000000
1!
b111 %
1'
b111 +
#59920000000
0!
0'
#59930000000
1!
b1000 %
1'
b1000 +
#59940000000
0!
0'
#59950000000
1!
b1001 %
1'
b1001 +
#59960000000
0!
0'
#59970000000
1!
b0 %
1'
b0 +
#59980000000
1"
1(
#59990000000
0!
0"
b100 &
0'
0(
b100 ,
#60000000000
1!
1$
b1 %
1'
1*
b1 +
#60010000000
0!
0'
#60020000000
1!
b10 %
1'
b10 +
#60030000000
0!
0'
#60040000000
1!
b11 %
1'
b11 +
#60050000000
0!
0'
#60060000000
1!
b100 %
1'
b100 +
#60070000000
0!
0'
#60080000000
1!
b101 %
1'
b101 +
#60090000000
0!
0'
#60100000000
1!
b110 %
1'
b110 +
#60110000000
0!
0'
#60120000000
1!
b111 %
1'
b111 +
#60130000000
0!
0'
#60140000000
1!
0$
b1000 %
1'
0*
b1000 +
#60150000000
0!
0'
#60160000000
1!
b1001 %
1'
b1001 +
#60170000000
0!
0'
#60180000000
1!
b0 %
1'
b0 +
#60190000000
0!
0'
#60200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#60210000000
0!
0'
#60220000000
1!
b10 %
1'
b10 +
#60230000000
0!
0'
#60240000000
1!
b11 %
1'
b11 +
#60250000000
0!
0'
#60260000000
1!
b100 %
1'
b100 +
#60270000000
0!
0'
#60280000000
1!
b101 %
1'
b101 +
#60290000000
0!
0'
#60300000000
1!
0$
b110 %
1'
0*
b110 +
#60310000000
0!
0'
#60320000000
1!
b111 %
1'
b111 +
#60330000000
0!
0'
#60340000000
1!
b1000 %
1'
b1000 +
#60350000000
0!
0'
#60360000000
1!
b1001 %
1'
b1001 +
#60370000000
0!
0'
#60380000000
1!
b0 %
1'
b0 +
#60390000000
0!
0'
#60400000000
1!
1$
b1 %
1'
1*
b1 +
#60410000000
1"
1(
#60420000000
0!
0"
b100 &
0'
0(
b100 ,
#60430000000
1!
b10 %
1'
b10 +
#60440000000
0!
0'
#60450000000
1!
b11 %
1'
b11 +
#60460000000
0!
0'
#60470000000
1!
b100 %
1'
b100 +
#60480000000
0!
0'
#60490000000
1!
b101 %
1'
b101 +
#60500000000
0!
0'
#60510000000
1!
b110 %
1'
b110 +
#60520000000
0!
0'
#60530000000
1!
b111 %
1'
b111 +
#60540000000
0!
0'
#60550000000
1!
0$
b1000 %
1'
0*
b1000 +
#60560000000
0!
0'
#60570000000
1!
b1001 %
1'
b1001 +
#60580000000
0!
0'
#60590000000
1!
b0 %
1'
b0 +
#60600000000
0!
0'
#60610000000
1!
1$
b1 %
1'
1*
b1 +
#60620000000
0!
0'
#60630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#60640000000
0!
0'
#60650000000
1!
b11 %
1'
b11 +
#60660000000
0!
0'
#60670000000
1!
b100 %
1'
b100 +
#60680000000
0!
0'
#60690000000
1!
b101 %
1'
b101 +
#60700000000
0!
0'
#60710000000
1!
0$
b110 %
1'
0*
b110 +
#60720000000
0!
0'
#60730000000
1!
b111 %
1'
b111 +
#60740000000
0!
0'
#60750000000
1!
b1000 %
1'
b1000 +
#60760000000
0!
0'
#60770000000
1!
b1001 %
1'
b1001 +
#60780000000
0!
0'
#60790000000
1!
b0 %
1'
b0 +
#60800000000
0!
0'
#60810000000
1!
1$
b1 %
1'
1*
b1 +
#60820000000
0!
0'
#60830000000
1!
b10 %
1'
b10 +
#60840000000
1"
1(
#60850000000
0!
0"
b100 &
0'
0(
b100 ,
#60860000000
1!
b11 %
1'
b11 +
#60870000000
0!
0'
#60880000000
1!
b100 %
1'
b100 +
#60890000000
0!
0'
#60900000000
1!
b101 %
1'
b101 +
#60910000000
0!
0'
#60920000000
1!
b110 %
1'
b110 +
#60930000000
0!
0'
#60940000000
1!
b111 %
1'
b111 +
#60950000000
0!
0'
#60960000000
1!
0$
b1000 %
1'
0*
b1000 +
#60970000000
0!
0'
#60980000000
1!
b1001 %
1'
b1001 +
#60990000000
0!
0'
#61000000000
1!
b0 %
1'
b0 +
#61010000000
0!
0'
#61020000000
1!
1$
b1 %
1'
1*
b1 +
#61030000000
0!
0'
#61040000000
1!
b10 %
1'
b10 +
#61050000000
0!
0'
#61060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#61070000000
0!
0'
#61080000000
1!
b100 %
1'
b100 +
#61090000000
0!
0'
#61100000000
1!
b101 %
1'
b101 +
#61110000000
0!
0'
#61120000000
1!
0$
b110 %
1'
0*
b110 +
#61130000000
0!
0'
#61140000000
1!
b111 %
1'
b111 +
#61150000000
0!
0'
#61160000000
1!
b1000 %
1'
b1000 +
#61170000000
0!
0'
#61180000000
1!
b1001 %
1'
b1001 +
#61190000000
0!
0'
#61200000000
1!
b0 %
1'
b0 +
#61210000000
0!
0'
#61220000000
1!
1$
b1 %
1'
1*
b1 +
#61230000000
0!
0'
#61240000000
1!
b10 %
1'
b10 +
#61250000000
0!
0'
#61260000000
1!
b11 %
1'
b11 +
#61270000000
1"
1(
#61280000000
0!
0"
b100 &
0'
0(
b100 ,
#61290000000
1!
b100 %
1'
b100 +
#61300000000
0!
0'
#61310000000
1!
b101 %
1'
b101 +
#61320000000
0!
0'
#61330000000
1!
b110 %
1'
b110 +
#61340000000
0!
0'
#61350000000
1!
b111 %
1'
b111 +
#61360000000
0!
0'
#61370000000
1!
0$
b1000 %
1'
0*
b1000 +
#61380000000
0!
0'
#61390000000
1!
b1001 %
1'
b1001 +
#61400000000
0!
0'
#61410000000
1!
b0 %
1'
b0 +
#61420000000
0!
0'
#61430000000
1!
1$
b1 %
1'
1*
b1 +
#61440000000
0!
0'
#61450000000
1!
b10 %
1'
b10 +
#61460000000
0!
0'
#61470000000
1!
b11 %
1'
b11 +
#61480000000
0!
0'
#61490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#61500000000
0!
0'
#61510000000
1!
b101 %
1'
b101 +
#61520000000
0!
0'
#61530000000
1!
0$
b110 %
1'
0*
b110 +
#61540000000
0!
0'
#61550000000
1!
b111 %
1'
b111 +
#61560000000
0!
0'
#61570000000
1!
b1000 %
1'
b1000 +
#61580000000
0!
0'
#61590000000
1!
b1001 %
1'
b1001 +
#61600000000
0!
0'
#61610000000
1!
b0 %
1'
b0 +
#61620000000
0!
0'
#61630000000
1!
1$
b1 %
1'
1*
b1 +
#61640000000
0!
0'
#61650000000
1!
b10 %
1'
b10 +
#61660000000
0!
0'
#61670000000
1!
b11 %
1'
b11 +
#61680000000
0!
0'
#61690000000
1!
b100 %
1'
b100 +
#61700000000
1"
1(
#61710000000
0!
0"
b100 &
0'
0(
b100 ,
#61720000000
1!
b101 %
1'
b101 +
#61730000000
0!
0'
#61740000000
1!
b110 %
1'
b110 +
#61750000000
0!
0'
#61760000000
1!
b111 %
1'
b111 +
#61770000000
0!
0'
#61780000000
1!
0$
b1000 %
1'
0*
b1000 +
#61790000000
0!
0'
#61800000000
1!
b1001 %
1'
b1001 +
#61810000000
0!
0'
#61820000000
1!
b0 %
1'
b0 +
#61830000000
0!
0'
#61840000000
1!
1$
b1 %
1'
1*
b1 +
#61850000000
0!
0'
#61860000000
1!
b10 %
1'
b10 +
#61870000000
0!
0'
#61880000000
1!
b11 %
1'
b11 +
#61890000000
0!
0'
#61900000000
1!
b100 %
1'
b100 +
#61910000000
0!
0'
#61920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#61930000000
0!
0'
#61940000000
1!
0$
b110 %
1'
0*
b110 +
#61950000000
0!
0'
#61960000000
1!
b111 %
1'
b111 +
#61970000000
0!
0'
#61980000000
1!
b1000 %
1'
b1000 +
#61990000000
0!
0'
#62000000000
1!
b1001 %
1'
b1001 +
#62010000000
0!
0'
#62020000000
1!
b0 %
1'
b0 +
#62030000000
0!
0'
#62040000000
1!
1$
b1 %
1'
1*
b1 +
#62050000000
0!
0'
#62060000000
1!
b10 %
1'
b10 +
#62070000000
0!
0'
#62080000000
1!
b11 %
1'
b11 +
#62090000000
0!
0'
#62100000000
1!
b100 %
1'
b100 +
#62110000000
0!
0'
#62120000000
1!
b101 %
1'
b101 +
#62130000000
1"
1(
#62140000000
0!
0"
b100 &
0'
0(
b100 ,
#62150000000
1!
b110 %
1'
b110 +
#62160000000
0!
0'
#62170000000
1!
b111 %
1'
b111 +
#62180000000
0!
0'
#62190000000
1!
0$
b1000 %
1'
0*
b1000 +
#62200000000
0!
0'
#62210000000
1!
b1001 %
1'
b1001 +
#62220000000
0!
0'
#62230000000
1!
b0 %
1'
b0 +
#62240000000
0!
0'
#62250000000
1!
1$
b1 %
1'
1*
b1 +
#62260000000
0!
0'
#62270000000
1!
b10 %
1'
b10 +
#62280000000
0!
0'
#62290000000
1!
b11 %
1'
b11 +
#62300000000
0!
0'
#62310000000
1!
b100 %
1'
b100 +
#62320000000
0!
0'
#62330000000
1!
b101 %
1'
b101 +
#62340000000
0!
0'
#62350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#62360000000
0!
0'
#62370000000
1!
b111 %
1'
b111 +
#62380000000
0!
0'
#62390000000
1!
b1000 %
1'
b1000 +
#62400000000
0!
0'
#62410000000
1!
b1001 %
1'
b1001 +
#62420000000
0!
0'
#62430000000
1!
b0 %
1'
b0 +
#62440000000
0!
0'
#62450000000
1!
1$
b1 %
1'
1*
b1 +
#62460000000
0!
0'
#62470000000
1!
b10 %
1'
b10 +
#62480000000
0!
0'
#62490000000
1!
b11 %
1'
b11 +
#62500000000
0!
0'
#62510000000
1!
b100 %
1'
b100 +
#62520000000
0!
0'
#62530000000
1!
b101 %
1'
b101 +
#62540000000
0!
0'
#62550000000
1!
0$
b110 %
1'
0*
b110 +
#62560000000
1"
1(
#62570000000
0!
0"
b100 &
0'
0(
b100 ,
#62580000000
1!
1$
b111 %
1'
1*
b111 +
#62590000000
0!
0'
#62600000000
1!
0$
b1000 %
1'
0*
b1000 +
#62610000000
0!
0'
#62620000000
1!
b1001 %
1'
b1001 +
#62630000000
0!
0'
#62640000000
1!
b0 %
1'
b0 +
#62650000000
0!
0'
#62660000000
1!
1$
b1 %
1'
1*
b1 +
#62670000000
0!
0'
#62680000000
1!
b10 %
1'
b10 +
#62690000000
0!
0'
#62700000000
1!
b11 %
1'
b11 +
#62710000000
0!
0'
#62720000000
1!
b100 %
1'
b100 +
#62730000000
0!
0'
#62740000000
1!
b101 %
1'
b101 +
#62750000000
0!
0'
#62760000000
1!
b110 %
1'
b110 +
#62770000000
0!
0'
#62780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#62790000000
0!
0'
#62800000000
1!
b1000 %
1'
b1000 +
#62810000000
0!
0'
#62820000000
1!
b1001 %
1'
b1001 +
#62830000000
0!
0'
#62840000000
1!
b0 %
1'
b0 +
#62850000000
0!
0'
#62860000000
1!
1$
b1 %
1'
1*
b1 +
#62870000000
0!
0'
#62880000000
1!
b10 %
1'
b10 +
#62890000000
0!
0'
#62900000000
1!
b11 %
1'
b11 +
#62910000000
0!
0'
#62920000000
1!
b100 %
1'
b100 +
#62930000000
0!
0'
#62940000000
1!
b101 %
1'
b101 +
#62950000000
0!
0'
#62960000000
1!
0$
b110 %
1'
0*
b110 +
#62970000000
0!
0'
#62980000000
1!
b111 %
1'
b111 +
#62990000000
1"
1(
#63000000000
0!
0"
b100 &
0'
0(
b100 ,
#63010000000
1!
b1000 %
1'
b1000 +
#63020000000
0!
0'
#63030000000
1!
b1001 %
1'
b1001 +
#63040000000
0!
0'
#63050000000
1!
b0 %
1'
b0 +
#63060000000
0!
0'
#63070000000
1!
1$
b1 %
1'
1*
b1 +
#63080000000
0!
0'
#63090000000
1!
b10 %
1'
b10 +
#63100000000
0!
0'
#63110000000
1!
b11 %
1'
b11 +
#63120000000
0!
0'
#63130000000
1!
b100 %
1'
b100 +
#63140000000
0!
0'
#63150000000
1!
b101 %
1'
b101 +
#63160000000
0!
0'
#63170000000
1!
b110 %
1'
b110 +
#63180000000
0!
0'
#63190000000
1!
b111 %
1'
b111 +
#63200000000
0!
0'
#63210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#63220000000
0!
0'
#63230000000
1!
b1001 %
1'
b1001 +
#63240000000
0!
0'
#63250000000
1!
b0 %
1'
b0 +
#63260000000
0!
0'
#63270000000
1!
1$
b1 %
1'
1*
b1 +
#63280000000
0!
0'
#63290000000
1!
b10 %
1'
b10 +
#63300000000
0!
0'
#63310000000
1!
b11 %
1'
b11 +
#63320000000
0!
0'
#63330000000
1!
b100 %
1'
b100 +
#63340000000
0!
0'
#63350000000
1!
b101 %
1'
b101 +
#63360000000
0!
0'
#63370000000
1!
0$
b110 %
1'
0*
b110 +
#63380000000
0!
0'
#63390000000
1!
b111 %
1'
b111 +
#63400000000
0!
0'
#63410000000
1!
b1000 %
1'
b1000 +
#63420000000
1"
1(
#63430000000
0!
0"
b100 &
0'
0(
b100 ,
#63440000000
1!
b1001 %
1'
b1001 +
#63450000000
0!
0'
#63460000000
1!
b0 %
1'
b0 +
#63470000000
0!
0'
#63480000000
1!
1$
b1 %
1'
1*
b1 +
#63490000000
0!
0'
#63500000000
1!
b10 %
1'
b10 +
#63510000000
0!
0'
#63520000000
1!
b11 %
1'
b11 +
#63530000000
0!
0'
#63540000000
1!
b100 %
1'
b100 +
#63550000000
0!
0'
#63560000000
1!
b101 %
1'
b101 +
#63570000000
0!
0'
#63580000000
1!
b110 %
1'
b110 +
#63590000000
0!
0'
#63600000000
1!
b111 %
1'
b111 +
#63610000000
0!
0'
#63620000000
1!
0$
b1000 %
1'
0*
b1000 +
#63630000000
0!
0'
#63640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#63650000000
0!
0'
#63660000000
1!
b0 %
1'
b0 +
#63670000000
0!
0'
#63680000000
1!
1$
b1 %
1'
1*
b1 +
#63690000000
0!
0'
#63700000000
1!
b10 %
1'
b10 +
#63710000000
0!
0'
#63720000000
1!
b11 %
1'
b11 +
#63730000000
0!
0'
#63740000000
1!
b100 %
1'
b100 +
#63750000000
0!
0'
#63760000000
1!
b101 %
1'
b101 +
#63770000000
0!
0'
#63780000000
1!
0$
b110 %
1'
0*
b110 +
#63790000000
0!
0'
#63800000000
1!
b111 %
1'
b111 +
#63810000000
0!
0'
#63820000000
1!
b1000 %
1'
b1000 +
#63830000000
0!
0'
#63840000000
1!
b1001 %
1'
b1001 +
#63850000000
1"
1(
#63860000000
0!
0"
b100 &
0'
0(
b100 ,
#63870000000
1!
b0 %
1'
b0 +
#63880000000
0!
0'
#63890000000
1!
1$
b1 %
1'
1*
b1 +
#63900000000
0!
0'
#63910000000
1!
b10 %
1'
b10 +
#63920000000
0!
0'
#63930000000
1!
b11 %
1'
b11 +
#63940000000
0!
0'
#63950000000
1!
b100 %
1'
b100 +
#63960000000
0!
0'
#63970000000
1!
b101 %
1'
b101 +
#63980000000
0!
0'
#63990000000
1!
b110 %
1'
b110 +
#64000000000
0!
0'
#64010000000
1!
b111 %
1'
b111 +
#64020000000
0!
0'
#64030000000
1!
0$
b1000 %
1'
0*
b1000 +
#64040000000
0!
0'
#64050000000
1!
b1001 %
1'
b1001 +
#64060000000
0!
0'
#64070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#64080000000
0!
0'
#64090000000
1!
1$
b1 %
1'
1*
b1 +
#64100000000
0!
0'
#64110000000
1!
b10 %
1'
b10 +
#64120000000
0!
0'
#64130000000
1!
b11 %
1'
b11 +
#64140000000
0!
0'
#64150000000
1!
b100 %
1'
b100 +
#64160000000
0!
0'
#64170000000
1!
b101 %
1'
b101 +
#64180000000
0!
0'
#64190000000
1!
0$
b110 %
1'
0*
b110 +
#64200000000
0!
0'
#64210000000
1!
b111 %
1'
b111 +
#64220000000
0!
0'
#64230000000
1!
b1000 %
1'
b1000 +
#64240000000
0!
0'
#64250000000
1!
b1001 %
1'
b1001 +
#64260000000
0!
0'
#64270000000
1!
b0 %
1'
b0 +
#64280000000
1"
1(
#64290000000
0!
0"
b100 &
0'
0(
b100 ,
#64300000000
1!
1$
b1 %
1'
1*
b1 +
#64310000000
0!
0'
#64320000000
1!
b10 %
1'
b10 +
#64330000000
0!
0'
#64340000000
1!
b11 %
1'
b11 +
#64350000000
0!
0'
#64360000000
1!
b100 %
1'
b100 +
#64370000000
0!
0'
#64380000000
1!
b101 %
1'
b101 +
#64390000000
0!
0'
#64400000000
1!
b110 %
1'
b110 +
#64410000000
0!
0'
#64420000000
1!
b111 %
1'
b111 +
#64430000000
0!
0'
#64440000000
1!
0$
b1000 %
1'
0*
b1000 +
#64450000000
0!
0'
#64460000000
1!
b1001 %
1'
b1001 +
#64470000000
0!
0'
#64480000000
1!
b0 %
1'
b0 +
#64490000000
0!
0'
#64500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#64510000000
0!
0'
#64520000000
1!
b10 %
1'
b10 +
#64530000000
0!
0'
#64540000000
1!
b11 %
1'
b11 +
#64550000000
0!
0'
#64560000000
1!
b100 %
1'
b100 +
#64570000000
0!
0'
#64580000000
1!
b101 %
1'
b101 +
#64590000000
0!
0'
#64600000000
1!
0$
b110 %
1'
0*
b110 +
#64610000000
0!
0'
#64620000000
1!
b111 %
1'
b111 +
#64630000000
0!
0'
#64640000000
1!
b1000 %
1'
b1000 +
#64650000000
0!
0'
#64660000000
1!
b1001 %
1'
b1001 +
#64670000000
0!
0'
#64680000000
1!
b0 %
1'
b0 +
#64690000000
0!
0'
#64700000000
1!
1$
b1 %
1'
1*
b1 +
#64710000000
1"
1(
#64720000000
0!
0"
b100 &
0'
0(
b100 ,
#64730000000
1!
b10 %
1'
b10 +
#64740000000
0!
0'
#64750000000
1!
b11 %
1'
b11 +
#64760000000
0!
0'
#64770000000
1!
b100 %
1'
b100 +
#64780000000
0!
0'
#64790000000
1!
b101 %
1'
b101 +
#64800000000
0!
0'
#64810000000
1!
b110 %
1'
b110 +
#64820000000
0!
0'
#64830000000
1!
b111 %
1'
b111 +
#64840000000
0!
0'
#64850000000
1!
0$
b1000 %
1'
0*
b1000 +
#64860000000
0!
0'
#64870000000
1!
b1001 %
1'
b1001 +
#64880000000
0!
0'
#64890000000
1!
b0 %
1'
b0 +
#64900000000
0!
0'
#64910000000
1!
1$
b1 %
1'
1*
b1 +
#64920000000
0!
0'
#64930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#64940000000
0!
0'
#64950000000
1!
b11 %
1'
b11 +
#64960000000
0!
0'
#64970000000
1!
b100 %
1'
b100 +
#64980000000
0!
0'
#64990000000
1!
b101 %
1'
b101 +
#65000000000
0!
0'
#65010000000
1!
0$
b110 %
1'
0*
b110 +
#65020000000
0!
0'
#65030000000
1!
b111 %
1'
b111 +
#65040000000
0!
0'
#65050000000
1!
b1000 %
1'
b1000 +
#65060000000
0!
0'
#65070000000
1!
b1001 %
1'
b1001 +
#65080000000
0!
0'
#65090000000
1!
b0 %
1'
b0 +
#65100000000
0!
0'
#65110000000
1!
1$
b1 %
1'
1*
b1 +
#65120000000
0!
0'
#65130000000
1!
b10 %
1'
b10 +
#65140000000
1"
1(
#65150000000
0!
0"
b100 &
0'
0(
b100 ,
#65160000000
1!
b11 %
1'
b11 +
#65170000000
0!
0'
#65180000000
1!
b100 %
1'
b100 +
#65190000000
0!
0'
#65200000000
1!
b101 %
1'
b101 +
#65210000000
0!
0'
#65220000000
1!
b110 %
1'
b110 +
#65230000000
0!
0'
#65240000000
1!
b111 %
1'
b111 +
#65250000000
0!
0'
#65260000000
1!
0$
b1000 %
1'
0*
b1000 +
#65270000000
0!
0'
#65280000000
1!
b1001 %
1'
b1001 +
#65290000000
0!
0'
#65300000000
1!
b0 %
1'
b0 +
#65310000000
0!
0'
#65320000000
1!
1$
b1 %
1'
1*
b1 +
#65330000000
0!
0'
#65340000000
1!
b10 %
1'
b10 +
#65350000000
0!
0'
#65360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#65370000000
0!
0'
#65380000000
1!
b100 %
1'
b100 +
#65390000000
0!
0'
#65400000000
1!
b101 %
1'
b101 +
#65410000000
0!
0'
#65420000000
1!
0$
b110 %
1'
0*
b110 +
#65430000000
0!
0'
#65440000000
1!
b111 %
1'
b111 +
#65450000000
0!
0'
#65460000000
1!
b1000 %
1'
b1000 +
#65470000000
0!
0'
#65480000000
1!
b1001 %
1'
b1001 +
#65490000000
0!
0'
#65500000000
1!
b0 %
1'
b0 +
#65510000000
0!
0'
#65520000000
1!
1$
b1 %
1'
1*
b1 +
#65530000000
0!
0'
#65540000000
1!
b10 %
1'
b10 +
#65550000000
0!
0'
#65560000000
1!
b11 %
1'
b11 +
#65570000000
1"
1(
#65580000000
0!
0"
b100 &
0'
0(
b100 ,
#65590000000
1!
b100 %
1'
b100 +
#65600000000
0!
0'
#65610000000
1!
b101 %
1'
b101 +
#65620000000
0!
0'
#65630000000
1!
b110 %
1'
b110 +
#65640000000
0!
0'
#65650000000
1!
b111 %
1'
b111 +
#65660000000
0!
0'
#65670000000
1!
0$
b1000 %
1'
0*
b1000 +
#65680000000
0!
0'
#65690000000
1!
b1001 %
1'
b1001 +
#65700000000
0!
0'
#65710000000
1!
b0 %
1'
b0 +
#65720000000
0!
0'
#65730000000
1!
1$
b1 %
1'
1*
b1 +
#65740000000
0!
0'
#65750000000
1!
b10 %
1'
b10 +
#65760000000
0!
0'
#65770000000
1!
b11 %
1'
b11 +
#65780000000
0!
0'
#65790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#65800000000
0!
0'
#65810000000
1!
b101 %
1'
b101 +
#65820000000
0!
0'
#65830000000
1!
0$
b110 %
1'
0*
b110 +
#65840000000
0!
0'
#65850000000
1!
b111 %
1'
b111 +
#65860000000
0!
0'
#65870000000
1!
b1000 %
1'
b1000 +
#65880000000
0!
0'
#65890000000
1!
b1001 %
1'
b1001 +
#65900000000
0!
0'
#65910000000
1!
b0 %
1'
b0 +
#65920000000
0!
0'
#65930000000
1!
1$
b1 %
1'
1*
b1 +
#65940000000
0!
0'
#65950000000
1!
b10 %
1'
b10 +
#65960000000
0!
0'
#65970000000
1!
b11 %
1'
b11 +
#65980000000
0!
0'
#65990000000
1!
b100 %
1'
b100 +
#66000000000
1"
1(
#66010000000
0!
0"
b100 &
0'
0(
b100 ,
#66020000000
1!
b101 %
1'
b101 +
#66030000000
0!
0'
#66040000000
1!
b110 %
1'
b110 +
#66050000000
0!
0'
#66060000000
1!
b111 %
1'
b111 +
#66070000000
0!
0'
#66080000000
1!
0$
b1000 %
1'
0*
b1000 +
#66090000000
0!
0'
#66100000000
1!
b1001 %
1'
b1001 +
#66110000000
0!
0'
#66120000000
1!
b0 %
1'
b0 +
#66130000000
0!
0'
#66140000000
1!
1$
b1 %
1'
1*
b1 +
#66150000000
0!
0'
#66160000000
1!
b10 %
1'
b10 +
#66170000000
0!
0'
#66180000000
1!
b11 %
1'
b11 +
#66190000000
0!
0'
#66200000000
1!
b100 %
1'
b100 +
#66210000000
0!
0'
#66220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#66230000000
0!
0'
#66240000000
1!
0$
b110 %
1'
0*
b110 +
#66250000000
0!
0'
#66260000000
1!
b111 %
1'
b111 +
#66270000000
0!
0'
#66280000000
1!
b1000 %
1'
b1000 +
#66290000000
0!
0'
#66300000000
1!
b1001 %
1'
b1001 +
#66310000000
0!
0'
#66320000000
1!
b0 %
1'
b0 +
#66330000000
0!
0'
#66340000000
1!
1$
b1 %
1'
1*
b1 +
#66350000000
0!
0'
#66360000000
1!
b10 %
1'
b10 +
#66370000000
0!
0'
#66380000000
1!
b11 %
1'
b11 +
#66390000000
0!
0'
#66400000000
1!
b100 %
1'
b100 +
#66410000000
0!
0'
#66420000000
1!
b101 %
1'
b101 +
#66430000000
1"
1(
#66440000000
0!
0"
b100 &
0'
0(
b100 ,
#66450000000
1!
b110 %
1'
b110 +
#66460000000
0!
0'
#66470000000
1!
b111 %
1'
b111 +
#66480000000
0!
0'
#66490000000
1!
0$
b1000 %
1'
0*
b1000 +
#66500000000
0!
0'
#66510000000
1!
b1001 %
1'
b1001 +
#66520000000
0!
0'
#66530000000
1!
b0 %
1'
b0 +
#66540000000
0!
0'
#66550000000
1!
1$
b1 %
1'
1*
b1 +
#66560000000
0!
0'
#66570000000
1!
b10 %
1'
b10 +
#66580000000
0!
0'
#66590000000
1!
b11 %
1'
b11 +
#66600000000
0!
0'
#66610000000
1!
b100 %
1'
b100 +
#66620000000
0!
0'
#66630000000
1!
b101 %
1'
b101 +
#66640000000
0!
0'
#66650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#66660000000
0!
0'
#66670000000
1!
b111 %
1'
b111 +
#66680000000
0!
0'
#66690000000
1!
b1000 %
1'
b1000 +
#66700000000
0!
0'
#66710000000
1!
b1001 %
1'
b1001 +
#66720000000
0!
0'
#66730000000
1!
b0 %
1'
b0 +
#66740000000
0!
0'
#66750000000
1!
1$
b1 %
1'
1*
b1 +
#66760000000
0!
0'
#66770000000
1!
b10 %
1'
b10 +
#66780000000
0!
0'
#66790000000
1!
b11 %
1'
b11 +
#66800000000
0!
0'
#66810000000
1!
b100 %
1'
b100 +
#66820000000
0!
0'
#66830000000
1!
b101 %
1'
b101 +
#66840000000
0!
0'
#66850000000
1!
0$
b110 %
1'
0*
b110 +
#66860000000
1"
1(
#66870000000
0!
0"
b100 &
0'
0(
b100 ,
#66880000000
1!
1$
b111 %
1'
1*
b111 +
#66890000000
0!
0'
#66900000000
1!
0$
b1000 %
1'
0*
b1000 +
#66910000000
0!
0'
#66920000000
1!
b1001 %
1'
b1001 +
#66930000000
0!
0'
#66940000000
1!
b0 %
1'
b0 +
#66950000000
0!
0'
#66960000000
1!
1$
b1 %
1'
1*
b1 +
#66970000000
0!
0'
#66980000000
1!
b10 %
1'
b10 +
#66990000000
0!
0'
#67000000000
1!
b11 %
1'
b11 +
#67010000000
0!
0'
#67020000000
1!
b100 %
1'
b100 +
#67030000000
0!
0'
#67040000000
1!
b101 %
1'
b101 +
#67050000000
0!
0'
#67060000000
1!
b110 %
1'
b110 +
#67070000000
0!
0'
#67080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#67090000000
0!
0'
#67100000000
1!
b1000 %
1'
b1000 +
#67110000000
0!
0'
#67120000000
1!
b1001 %
1'
b1001 +
#67130000000
0!
0'
#67140000000
1!
b0 %
1'
b0 +
#67150000000
0!
0'
#67160000000
1!
1$
b1 %
1'
1*
b1 +
#67170000000
0!
0'
#67180000000
1!
b10 %
1'
b10 +
#67190000000
0!
0'
#67200000000
1!
b11 %
1'
b11 +
#67210000000
0!
0'
#67220000000
1!
b100 %
1'
b100 +
#67230000000
0!
0'
#67240000000
1!
b101 %
1'
b101 +
#67250000000
0!
0'
#67260000000
1!
0$
b110 %
1'
0*
b110 +
#67270000000
0!
0'
#67280000000
1!
b111 %
1'
b111 +
#67290000000
1"
1(
#67300000000
0!
0"
b100 &
0'
0(
b100 ,
#67310000000
1!
b1000 %
1'
b1000 +
#67320000000
0!
0'
#67330000000
1!
b1001 %
1'
b1001 +
#67340000000
0!
0'
#67350000000
1!
b0 %
1'
b0 +
#67360000000
0!
0'
#67370000000
1!
1$
b1 %
1'
1*
b1 +
#67380000000
0!
0'
#67390000000
1!
b10 %
1'
b10 +
#67400000000
0!
0'
#67410000000
1!
b11 %
1'
b11 +
#67420000000
0!
0'
#67430000000
1!
b100 %
1'
b100 +
#67440000000
0!
0'
#67450000000
1!
b101 %
1'
b101 +
#67460000000
0!
0'
#67470000000
1!
b110 %
1'
b110 +
#67480000000
0!
0'
#67490000000
1!
b111 %
1'
b111 +
#67500000000
0!
0'
#67510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#67520000000
0!
0'
#67530000000
1!
b1001 %
1'
b1001 +
#67540000000
0!
0'
#67550000000
1!
b0 %
1'
b0 +
#67560000000
0!
0'
#67570000000
1!
1$
b1 %
1'
1*
b1 +
#67580000000
0!
0'
#67590000000
1!
b10 %
1'
b10 +
#67600000000
0!
0'
#67610000000
1!
b11 %
1'
b11 +
#67620000000
0!
0'
#67630000000
1!
b100 %
1'
b100 +
#67640000000
0!
0'
#67650000000
1!
b101 %
1'
b101 +
#67660000000
0!
0'
#67670000000
1!
0$
b110 %
1'
0*
b110 +
#67680000000
0!
0'
#67690000000
1!
b111 %
1'
b111 +
#67700000000
0!
0'
#67710000000
1!
b1000 %
1'
b1000 +
#67720000000
1"
1(
#67730000000
0!
0"
b100 &
0'
0(
b100 ,
#67740000000
1!
b1001 %
1'
b1001 +
#67750000000
0!
0'
#67760000000
1!
b0 %
1'
b0 +
#67770000000
0!
0'
#67780000000
1!
1$
b1 %
1'
1*
b1 +
#67790000000
0!
0'
#67800000000
1!
b10 %
1'
b10 +
#67810000000
0!
0'
#67820000000
1!
b11 %
1'
b11 +
#67830000000
0!
0'
#67840000000
1!
b100 %
1'
b100 +
#67850000000
0!
0'
#67860000000
1!
b101 %
1'
b101 +
#67870000000
0!
0'
#67880000000
1!
b110 %
1'
b110 +
#67890000000
0!
0'
#67900000000
1!
b111 %
1'
b111 +
#67910000000
0!
0'
#67920000000
1!
0$
b1000 %
1'
0*
b1000 +
#67930000000
0!
0'
#67940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#67950000000
0!
0'
#67960000000
1!
b0 %
1'
b0 +
#67970000000
0!
0'
#67980000000
1!
1$
b1 %
1'
1*
b1 +
#67990000000
0!
0'
#68000000000
1!
b10 %
1'
b10 +
#68010000000
0!
0'
#68020000000
1!
b11 %
1'
b11 +
#68030000000
0!
0'
#68040000000
1!
b100 %
1'
b100 +
#68050000000
0!
0'
#68060000000
1!
b101 %
1'
b101 +
#68070000000
0!
0'
#68080000000
1!
0$
b110 %
1'
0*
b110 +
#68090000000
0!
0'
#68100000000
1!
b111 %
1'
b111 +
#68110000000
0!
0'
#68120000000
1!
b1000 %
1'
b1000 +
#68130000000
0!
0'
#68140000000
1!
b1001 %
1'
b1001 +
#68150000000
1"
1(
#68160000000
0!
0"
b100 &
0'
0(
b100 ,
#68170000000
1!
b0 %
1'
b0 +
#68180000000
0!
0'
#68190000000
1!
1$
b1 %
1'
1*
b1 +
#68200000000
0!
0'
#68210000000
1!
b10 %
1'
b10 +
#68220000000
0!
0'
#68230000000
1!
b11 %
1'
b11 +
#68240000000
0!
0'
#68250000000
1!
b100 %
1'
b100 +
#68260000000
0!
0'
#68270000000
1!
b101 %
1'
b101 +
#68280000000
0!
0'
#68290000000
1!
b110 %
1'
b110 +
#68300000000
0!
0'
#68310000000
1!
b111 %
1'
b111 +
#68320000000
0!
0'
#68330000000
1!
0$
b1000 %
1'
0*
b1000 +
#68340000000
0!
0'
#68350000000
1!
b1001 %
1'
b1001 +
#68360000000
0!
0'
#68370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#68380000000
0!
0'
#68390000000
1!
1$
b1 %
1'
1*
b1 +
#68400000000
0!
0'
#68410000000
1!
b10 %
1'
b10 +
#68420000000
0!
0'
#68430000000
1!
b11 %
1'
b11 +
#68440000000
0!
0'
#68450000000
1!
b100 %
1'
b100 +
#68460000000
0!
0'
#68470000000
1!
b101 %
1'
b101 +
#68480000000
0!
0'
#68490000000
1!
0$
b110 %
1'
0*
b110 +
#68500000000
0!
0'
#68510000000
1!
b111 %
1'
b111 +
#68520000000
0!
0'
#68530000000
1!
b1000 %
1'
b1000 +
#68540000000
0!
0'
#68550000000
1!
b1001 %
1'
b1001 +
#68560000000
0!
0'
#68570000000
1!
b0 %
1'
b0 +
#68580000000
1"
1(
#68590000000
0!
0"
b100 &
0'
0(
b100 ,
#68600000000
1!
1$
b1 %
1'
1*
b1 +
#68610000000
0!
0'
#68620000000
1!
b10 %
1'
b10 +
#68630000000
0!
0'
#68640000000
1!
b11 %
1'
b11 +
#68650000000
0!
0'
#68660000000
1!
b100 %
1'
b100 +
#68670000000
0!
0'
#68680000000
1!
b101 %
1'
b101 +
#68690000000
0!
0'
#68700000000
1!
b110 %
1'
b110 +
#68710000000
0!
0'
#68720000000
1!
b111 %
1'
b111 +
#68730000000
0!
0'
#68740000000
1!
0$
b1000 %
1'
0*
b1000 +
#68750000000
0!
0'
#68760000000
1!
b1001 %
1'
b1001 +
#68770000000
0!
0'
#68780000000
1!
b0 %
1'
b0 +
#68790000000
0!
0'
#68800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#68810000000
0!
0'
#68820000000
1!
b10 %
1'
b10 +
#68830000000
0!
0'
#68840000000
1!
b11 %
1'
b11 +
#68850000000
0!
0'
#68860000000
1!
b100 %
1'
b100 +
#68870000000
0!
0'
#68880000000
1!
b101 %
1'
b101 +
#68890000000
0!
0'
#68900000000
1!
0$
b110 %
1'
0*
b110 +
#68910000000
0!
0'
#68920000000
1!
b111 %
1'
b111 +
#68930000000
0!
0'
#68940000000
1!
b1000 %
1'
b1000 +
#68950000000
0!
0'
#68960000000
1!
b1001 %
1'
b1001 +
#68970000000
0!
0'
#68980000000
1!
b0 %
1'
b0 +
#68990000000
0!
0'
#69000000000
1!
1$
b1 %
1'
1*
b1 +
#69010000000
1"
1(
#69020000000
0!
0"
b100 &
0'
0(
b100 ,
#69030000000
1!
b10 %
1'
b10 +
#69040000000
0!
0'
#69050000000
1!
b11 %
1'
b11 +
#69060000000
0!
0'
#69070000000
1!
b100 %
1'
b100 +
#69080000000
0!
0'
#69090000000
1!
b101 %
1'
b101 +
#69100000000
0!
0'
#69110000000
1!
b110 %
1'
b110 +
#69120000000
0!
0'
#69130000000
1!
b111 %
1'
b111 +
#69140000000
0!
0'
#69150000000
1!
0$
b1000 %
1'
0*
b1000 +
#69160000000
0!
0'
#69170000000
1!
b1001 %
1'
b1001 +
#69180000000
0!
0'
#69190000000
1!
b0 %
1'
b0 +
#69200000000
0!
0'
#69210000000
1!
1$
b1 %
1'
1*
b1 +
#69220000000
0!
0'
#69230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#69240000000
0!
0'
#69250000000
1!
b11 %
1'
b11 +
#69260000000
0!
0'
#69270000000
1!
b100 %
1'
b100 +
#69280000000
0!
0'
#69290000000
1!
b101 %
1'
b101 +
#69300000000
0!
0'
#69310000000
1!
0$
b110 %
1'
0*
b110 +
#69320000000
0!
0'
#69330000000
1!
b111 %
1'
b111 +
#69340000000
0!
0'
#69350000000
1!
b1000 %
1'
b1000 +
#69360000000
0!
0'
#69370000000
1!
b1001 %
1'
b1001 +
#69380000000
0!
0'
#69390000000
1!
b0 %
1'
b0 +
#69400000000
0!
0'
#69410000000
1!
1$
b1 %
1'
1*
b1 +
#69420000000
0!
0'
#69430000000
1!
b10 %
1'
b10 +
#69440000000
1"
1(
#69450000000
0!
0"
b100 &
0'
0(
b100 ,
#69460000000
1!
b11 %
1'
b11 +
#69470000000
0!
0'
#69480000000
1!
b100 %
1'
b100 +
#69490000000
0!
0'
#69500000000
1!
b101 %
1'
b101 +
#69510000000
0!
0'
#69520000000
1!
b110 %
1'
b110 +
#69530000000
0!
0'
#69540000000
1!
b111 %
1'
b111 +
#69550000000
0!
0'
#69560000000
1!
0$
b1000 %
1'
0*
b1000 +
#69570000000
0!
0'
#69580000000
1!
b1001 %
1'
b1001 +
#69590000000
0!
0'
#69600000000
1!
b0 %
1'
b0 +
#69610000000
0!
0'
#69620000000
1!
1$
b1 %
1'
1*
b1 +
#69630000000
0!
0'
#69640000000
1!
b10 %
1'
b10 +
#69650000000
0!
0'
#69660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#69670000000
0!
0'
#69680000000
1!
b100 %
1'
b100 +
#69690000000
0!
0'
#69700000000
1!
b101 %
1'
b101 +
#69710000000
0!
0'
#69720000000
1!
0$
b110 %
1'
0*
b110 +
#69730000000
0!
0'
#69740000000
1!
b111 %
1'
b111 +
#69750000000
0!
0'
#69760000000
1!
b1000 %
1'
b1000 +
#69770000000
0!
0'
#69780000000
1!
b1001 %
1'
b1001 +
#69790000000
0!
0'
#69800000000
1!
b0 %
1'
b0 +
#69810000000
0!
0'
#69820000000
1!
1$
b1 %
1'
1*
b1 +
#69830000000
0!
0'
#69840000000
1!
b10 %
1'
b10 +
#69850000000
0!
0'
#69860000000
1!
b11 %
1'
b11 +
#69870000000
1"
1(
#69880000000
0!
0"
b100 &
0'
0(
b100 ,
#69890000000
1!
b100 %
1'
b100 +
#69900000000
0!
0'
#69910000000
1!
b101 %
1'
b101 +
#69920000000
0!
0'
#69930000000
1!
b110 %
1'
b110 +
#69940000000
0!
0'
#69950000000
1!
b111 %
1'
b111 +
#69960000000
0!
0'
#69970000000
1!
0$
b1000 %
1'
0*
b1000 +
#69980000000
0!
0'
#69990000000
1!
b1001 %
1'
b1001 +
#70000000000
0!
0'
#70010000000
1!
b0 %
1'
b0 +
#70020000000
0!
0'
#70030000000
1!
1$
b1 %
1'
1*
b1 +
#70040000000
0!
0'
#70050000000
1!
b10 %
1'
b10 +
#70060000000
0!
0'
#70070000000
1!
b11 %
1'
b11 +
#70080000000
0!
0'
#70090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#70100000000
0!
0'
#70110000000
1!
b101 %
1'
b101 +
#70120000000
0!
0'
#70130000000
1!
0$
b110 %
1'
0*
b110 +
#70140000000
0!
0'
#70150000000
1!
b111 %
1'
b111 +
#70160000000
0!
0'
#70170000000
1!
b1000 %
1'
b1000 +
#70180000000
0!
0'
#70190000000
1!
b1001 %
1'
b1001 +
#70200000000
0!
0'
#70210000000
1!
b0 %
1'
b0 +
#70220000000
0!
0'
#70230000000
1!
1$
b1 %
1'
1*
b1 +
#70240000000
0!
0'
#70250000000
1!
b10 %
1'
b10 +
#70260000000
0!
0'
#70270000000
1!
b11 %
1'
b11 +
#70280000000
0!
0'
#70290000000
1!
b100 %
1'
b100 +
#70300000000
1"
1(
#70310000000
0!
0"
b100 &
0'
0(
b100 ,
#70320000000
1!
b101 %
1'
b101 +
#70330000000
0!
0'
#70340000000
1!
b110 %
1'
b110 +
#70350000000
0!
0'
#70360000000
1!
b111 %
1'
b111 +
#70370000000
0!
0'
#70380000000
1!
0$
b1000 %
1'
0*
b1000 +
#70390000000
0!
0'
#70400000000
1!
b1001 %
1'
b1001 +
#70410000000
0!
0'
#70420000000
1!
b0 %
1'
b0 +
#70430000000
0!
0'
#70440000000
1!
1$
b1 %
1'
1*
b1 +
#70450000000
0!
0'
#70460000000
1!
b10 %
1'
b10 +
#70470000000
0!
0'
#70480000000
1!
b11 %
1'
b11 +
#70490000000
0!
0'
#70500000000
1!
b100 %
1'
b100 +
#70510000000
0!
0'
#70520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#70530000000
0!
0'
#70540000000
1!
0$
b110 %
1'
0*
b110 +
#70550000000
0!
0'
#70560000000
1!
b111 %
1'
b111 +
#70570000000
0!
0'
#70580000000
1!
b1000 %
1'
b1000 +
#70590000000
0!
0'
#70600000000
1!
b1001 %
1'
b1001 +
#70610000000
0!
0'
#70620000000
1!
b0 %
1'
b0 +
#70630000000
0!
0'
#70640000000
1!
1$
b1 %
1'
1*
b1 +
#70650000000
0!
0'
#70660000000
1!
b10 %
1'
b10 +
#70670000000
0!
0'
#70680000000
1!
b11 %
1'
b11 +
#70690000000
0!
0'
#70700000000
1!
b100 %
1'
b100 +
#70710000000
0!
0'
#70720000000
1!
b101 %
1'
b101 +
#70730000000
1"
1(
#70740000000
0!
0"
b100 &
0'
0(
b100 ,
#70750000000
1!
b110 %
1'
b110 +
#70760000000
0!
0'
#70770000000
1!
b111 %
1'
b111 +
#70780000000
0!
0'
#70790000000
1!
0$
b1000 %
1'
0*
b1000 +
#70800000000
0!
0'
#70810000000
1!
b1001 %
1'
b1001 +
#70820000000
0!
0'
#70830000000
1!
b0 %
1'
b0 +
#70840000000
0!
0'
#70850000000
1!
1$
b1 %
1'
1*
b1 +
#70860000000
0!
0'
#70870000000
1!
b10 %
1'
b10 +
#70880000000
0!
0'
#70890000000
1!
b11 %
1'
b11 +
#70900000000
0!
0'
#70910000000
1!
b100 %
1'
b100 +
#70920000000
0!
0'
#70930000000
1!
b101 %
1'
b101 +
#70940000000
0!
0'
#70950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#70960000000
0!
0'
#70970000000
1!
b111 %
1'
b111 +
#70980000000
0!
0'
#70990000000
1!
b1000 %
1'
b1000 +
#71000000000
0!
0'
#71010000000
1!
b1001 %
1'
b1001 +
#71020000000
0!
0'
#71030000000
1!
b0 %
1'
b0 +
#71040000000
0!
0'
#71050000000
1!
1$
b1 %
1'
1*
b1 +
#71060000000
0!
0'
#71070000000
1!
b10 %
1'
b10 +
#71080000000
0!
0'
#71090000000
1!
b11 %
1'
b11 +
#71100000000
0!
0'
#71110000000
1!
b100 %
1'
b100 +
#71120000000
0!
0'
#71130000000
1!
b101 %
1'
b101 +
#71140000000
0!
0'
#71150000000
1!
0$
b110 %
1'
0*
b110 +
#71160000000
1"
1(
#71170000000
0!
0"
b100 &
0'
0(
b100 ,
#71180000000
1!
1$
b111 %
1'
1*
b111 +
#71190000000
0!
0'
#71200000000
1!
0$
b1000 %
1'
0*
b1000 +
#71210000000
0!
0'
#71220000000
1!
b1001 %
1'
b1001 +
#71230000000
0!
0'
#71240000000
1!
b0 %
1'
b0 +
#71250000000
0!
0'
#71260000000
1!
1$
b1 %
1'
1*
b1 +
#71270000000
0!
0'
#71280000000
1!
b10 %
1'
b10 +
#71290000000
0!
0'
#71300000000
1!
b11 %
1'
b11 +
#71310000000
0!
0'
#71320000000
1!
b100 %
1'
b100 +
#71330000000
0!
0'
#71340000000
1!
b101 %
1'
b101 +
#71350000000
0!
0'
#71360000000
1!
b110 %
1'
b110 +
#71370000000
0!
0'
#71380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#71390000000
0!
0'
#71400000000
1!
b1000 %
1'
b1000 +
#71410000000
0!
0'
#71420000000
1!
b1001 %
1'
b1001 +
#71430000000
0!
0'
#71440000000
1!
b0 %
1'
b0 +
#71450000000
0!
0'
#71460000000
1!
1$
b1 %
1'
1*
b1 +
#71470000000
0!
0'
#71480000000
1!
b10 %
1'
b10 +
#71490000000
0!
0'
#71500000000
1!
b11 %
1'
b11 +
#71510000000
0!
0'
#71520000000
1!
b100 %
1'
b100 +
#71530000000
0!
0'
#71540000000
1!
b101 %
1'
b101 +
#71550000000
0!
0'
#71560000000
1!
0$
b110 %
1'
0*
b110 +
#71570000000
0!
0'
#71580000000
1!
b111 %
1'
b111 +
#71590000000
1"
1(
#71600000000
0!
0"
b100 &
0'
0(
b100 ,
#71610000000
1!
b1000 %
1'
b1000 +
#71620000000
0!
0'
#71630000000
1!
b1001 %
1'
b1001 +
#71640000000
0!
0'
#71650000000
1!
b0 %
1'
b0 +
#71660000000
0!
0'
#71670000000
1!
1$
b1 %
1'
1*
b1 +
#71680000000
0!
0'
#71690000000
1!
b10 %
1'
b10 +
#71700000000
0!
0'
#71710000000
1!
b11 %
1'
b11 +
#71720000000
0!
0'
#71730000000
1!
b100 %
1'
b100 +
#71740000000
0!
0'
#71750000000
1!
b101 %
1'
b101 +
#71760000000
0!
0'
#71770000000
1!
b110 %
1'
b110 +
#71780000000
0!
0'
#71790000000
1!
b111 %
1'
b111 +
#71800000000
0!
0'
#71810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#71820000000
0!
0'
#71830000000
1!
b1001 %
1'
b1001 +
#71840000000
0!
0'
#71850000000
1!
b0 %
1'
b0 +
#71860000000
0!
0'
#71870000000
1!
1$
b1 %
1'
1*
b1 +
#71880000000
0!
0'
#71890000000
1!
b10 %
1'
b10 +
#71900000000
0!
0'
#71910000000
1!
b11 %
1'
b11 +
#71920000000
0!
0'
#71930000000
1!
b100 %
1'
b100 +
#71940000000
0!
0'
#71950000000
1!
b101 %
1'
b101 +
#71960000000
0!
0'
#71970000000
1!
0$
b110 %
1'
0*
b110 +
#71980000000
0!
0'
#71990000000
1!
b111 %
1'
b111 +
#72000000000
0!
0'
#72010000000
1!
b1000 %
1'
b1000 +
#72020000000
1"
1(
#72030000000
0!
0"
b100 &
0'
0(
b100 ,
#72040000000
1!
b1001 %
1'
b1001 +
#72050000000
0!
0'
#72060000000
1!
b0 %
1'
b0 +
#72070000000
0!
0'
#72080000000
1!
1$
b1 %
1'
1*
b1 +
#72090000000
0!
0'
#72100000000
1!
b10 %
1'
b10 +
#72110000000
0!
0'
#72120000000
1!
b11 %
1'
b11 +
#72130000000
0!
0'
#72140000000
1!
b100 %
1'
b100 +
#72150000000
0!
0'
#72160000000
1!
b101 %
1'
b101 +
#72170000000
0!
0'
#72180000000
1!
b110 %
1'
b110 +
#72190000000
0!
0'
#72200000000
1!
b111 %
1'
b111 +
#72210000000
0!
0'
#72220000000
1!
0$
b1000 %
1'
0*
b1000 +
#72230000000
0!
0'
#72240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#72250000000
0!
0'
#72260000000
1!
b0 %
1'
b0 +
#72270000000
0!
0'
#72280000000
1!
1$
b1 %
1'
1*
b1 +
#72290000000
0!
0'
#72300000000
1!
b10 %
1'
b10 +
#72310000000
0!
0'
#72320000000
1!
b11 %
1'
b11 +
#72330000000
0!
0'
#72340000000
1!
b100 %
1'
b100 +
#72350000000
0!
0'
#72360000000
1!
b101 %
1'
b101 +
#72370000000
0!
0'
#72380000000
1!
0$
b110 %
1'
0*
b110 +
#72390000000
0!
0'
#72400000000
1!
b111 %
1'
b111 +
#72410000000
0!
0'
#72420000000
1!
b1000 %
1'
b1000 +
#72430000000
0!
0'
#72440000000
1!
b1001 %
1'
b1001 +
#72450000000
1"
1(
#72460000000
0!
0"
b100 &
0'
0(
b100 ,
#72470000000
1!
b0 %
1'
b0 +
#72480000000
0!
0'
#72490000000
1!
1$
b1 %
1'
1*
b1 +
#72500000000
0!
0'
#72510000000
1!
b10 %
1'
b10 +
#72520000000
0!
0'
#72530000000
1!
b11 %
1'
b11 +
#72540000000
0!
0'
#72550000000
1!
b100 %
1'
b100 +
#72560000000
0!
0'
#72570000000
1!
b101 %
1'
b101 +
#72580000000
0!
0'
#72590000000
1!
b110 %
1'
b110 +
#72600000000
0!
0'
#72610000000
1!
b111 %
1'
b111 +
#72620000000
0!
0'
#72630000000
1!
0$
b1000 %
1'
0*
b1000 +
#72640000000
0!
0'
#72650000000
1!
b1001 %
1'
b1001 +
#72660000000
0!
0'
#72670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#72680000000
0!
0'
#72690000000
1!
1$
b1 %
1'
1*
b1 +
#72700000000
0!
0'
#72710000000
1!
b10 %
1'
b10 +
#72720000000
0!
0'
#72730000000
1!
b11 %
1'
b11 +
#72740000000
0!
0'
#72750000000
1!
b100 %
1'
b100 +
#72760000000
0!
0'
#72770000000
1!
b101 %
1'
b101 +
#72780000000
0!
0'
#72790000000
1!
0$
b110 %
1'
0*
b110 +
#72800000000
0!
0'
#72810000000
1!
b111 %
1'
b111 +
#72820000000
0!
0'
#72830000000
1!
b1000 %
1'
b1000 +
#72840000000
0!
0'
#72850000000
1!
b1001 %
1'
b1001 +
#72860000000
0!
0'
#72870000000
1!
b0 %
1'
b0 +
#72880000000
1"
1(
#72890000000
0!
0"
b100 &
0'
0(
b100 ,
#72900000000
1!
1$
b1 %
1'
1*
b1 +
#72910000000
0!
0'
#72920000000
1!
b10 %
1'
b10 +
#72930000000
0!
0'
#72940000000
1!
b11 %
1'
b11 +
#72950000000
0!
0'
#72960000000
1!
b100 %
1'
b100 +
#72970000000
0!
0'
#72980000000
1!
b101 %
1'
b101 +
#72990000000
0!
0'
#73000000000
1!
b110 %
1'
b110 +
#73010000000
0!
0'
#73020000000
1!
b111 %
1'
b111 +
#73030000000
0!
0'
#73040000000
1!
0$
b1000 %
1'
0*
b1000 +
#73050000000
0!
0'
#73060000000
1!
b1001 %
1'
b1001 +
#73070000000
0!
0'
#73080000000
1!
b0 %
1'
b0 +
#73090000000
0!
0'
#73100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#73110000000
0!
0'
#73120000000
1!
b10 %
1'
b10 +
#73130000000
0!
0'
#73140000000
1!
b11 %
1'
b11 +
#73150000000
0!
0'
#73160000000
1!
b100 %
1'
b100 +
#73170000000
0!
0'
#73180000000
1!
b101 %
1'
b101 +
#73190000000
0!
0'
#73200000000
1!
0$
b110 %
1'
0*
b110 +
#73210000000
0!
0'
#73220000000
1!
b111 %
1'
b111 +
#73230000000
0!
0'
#73240000000
1!
b1000 %
1'
b1000 +
#73250000000
0!
0'
#73260000000
1!
b1001 %
1'
b1001 +
#73270000000
0!
0'
#73280000000
1!
b0 %
1'
b0 +
#73290000000
0!
0'
#73300000000
1!
1$
b1 %
1'
1*
b1 +
#73310000000
1"
1(
#73320000000
0!
0"
b100 &
0'
0(
b100 ,
#73330000000
1!
b10 %
1'
b10 +
#73340000000
0!
0'
#73350000000
1!
b11 %
1'
b11 +
#73360000000
0!
0'
#73370000000
1!
b100 %
1'
b100 +
#73380000000
0!
0'
#73390000000
1!
b101 %
1'
b101 +
#73400000000
0!
0'
#73410000000
1!
b110 %
1'
b110 +
#73420000000
0!
0'
#73430000000
1!
b111 %
1'
b111 +
#73440000000
0!
0'
#73450000000
1!
0$
b1000 %
1'
0*
b1000 +
#73460000000
0!
0'
#73470000000
1!
b1001 %
1'
b1001 +
#73480000000
0!
0'
#73490000000
1!
b0 %
1'
b0 +
#73500000000
0!
0'
#73510000000
1!
1$
b1 %
1'
1*
b1 +
#73520000000
0!
0'
#73530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#73540000000
0!
0'
#73550000000
1!
b11 %
1'
b11 +
#73560000000
0!
0'
#73570000000
1!
b100 %
1'
b100 +
#73580000000
0!
0'
#73590000000
1!
b101 %
1'
b101 +
#73600000000
0!
0'
#73610000000
1!
0$
b110 %
1'
0*
b110 +
#73620000000
0!
0'
#73630000000
1!
b111 %
1'
b111 +
#73640000000
0!
0'
#73650000000
1!
b1000 %
1'
b1000 +
#73660000000
0!
0'
#73670000000
1!
b1001 %
1'
b1001 +
#73680000000
0!
0'
#73690000000
1!
b0 %
1'
b0 +
#73700000000
0!
0'
#73710000000
1!
1$
b1 %
1'
1*
b1 +
#73720000000
0!
0'
#73730000000
1!
b10 %
1'
b10 +
#73740000000
1"
1(
#73750000000
0!
0"
b100 &
0'
0(
b100 ,
#73760000000
1!
b11 %
1'
b11 +
#73770000000
0!
0'
#73780000000
1!
b100 %
1'
b100 +
#73790000000
0!
0'
#73800000000
1!
b101 %
1'
b101 +
#73810000000
0!
0'
#73820000000
1!
b110 %
1'
b110 +
#73830000000
0!
0'
#73840000000
1!
b111 %
1'
b111 +
#73850000000
0!
0'
#73860000000
1!
0$
b1000 %
1'
0*
b1000 +
#73870000000
0!
0'
#73880000000
1!
b1001 %
1'
b1001 +
#73890000000
0!
0'
#73900000000
1!
b0 %
1'
b0 +
#73910000000
0!
0'
#73920000000
1!
1$
b1 %
1'
1*
b1 +
#73930000000
0!
0'
#73940000000
1!
b10 %
1'
b10 +
#73950000000
0!
0'
#73960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#73970000000
0!
0'
#73980000000
1!
b100 %
1'
b100 +
#73990000000
0!
0'
#74000000000
1!
b101 %
1'
b101 +
#74010000000
0!
0'
#74020000000
1!
0$
b110 %
1'
0*
b110 +
#74030000000
0!
0'
#74040000000
1!
b111 %
1'
b111 +
#74050000000
0!
0'
#74060000000
1!
b1000 %
1'
b1000 +
#74070000000
0!
0'
#74080000000
1!
b1001 %
1'
b1001 +
#74090000000
0!
0'
#74100000000
1!
b0 %
1'
b0 +
#74110000000
0!
0'
#74120000000
1!
1$
b1 %
1'
1*
b1 +
#74130000000
0!
0'
#74140000000
1!
b10 %
1'
b10 +
#74150000000
0!
0'
#74160000000
1!
b11 %
1'
b11 +
#74170000000
1"
1(
#74180000000
0!
0"
b100 &
0'
0(
b100 ,
#74190000000
1!
b100 %
1'
b100 +
#74200000000
0!
0'
#74210000000
1!
b101 %
1'
b101 +
#74220000000
0!
0'
#74230000000
1!
b110 %
1'
b110 +
#74240000000
0!
0'
#74250000000
1!
b111 %
1'
b111 +
#74260000000
0!
0'
#74270000000
1!
0$
b1000 %
1'
0*
b1000 +
#74280000000
0!
0'
#74290000000
1!
b1001 %
1'
b1001 +
#74300000000
0!
0'
#74310000000
1!
b0 %
1'
b0 +
#74320000000
0!
0'
#74330000000
1!
1$
b1 %
1'
1*
b1 +
#74340000000
0!
0'
#74350000000
1!
b10 %
1'
b10 +
#74360000000
0!
0'
#74370000000
1!
b11 %
1'
b11 +
#74380000000
0!
0'
#74390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#74400000000
0!
0'
#74410000000
1!
b101 %
1'
b101 +
#74420000000
0!
0'
#74430000000
1!
0$
b110 %
1'
0*
b110 +
#74440000000
0!
0'
#74450000000
1!
b111 %
1'
b111 +
#74460000000
0!
0'
#74470000000
1!
b1000 %
1'
b1000 +
#74480000000
0!
0'
#74490000000
1!
b1001 %
1'
b1001 +
#74500000000
0!
0'
#74510000000
1!
b0 %
1'
b0 +
#74520000000
0!
0'
#74530000000
1!
1$
b1 %
1'
1*
b1 +
#74540000000
0!
0'
#74550000000
1!
b10 %
1'
b10 +
#74560000000
0!
0'
#74570000000
1!
b11 %
1'
b11 +
#74580000000
0!
0'
#74590000000
1!
b100 %
1'
b100 +
#74600000000
1"
1(
#74610000000
0!
0"
b100 &
0'
0(
b100 ,
#74620000000
1!
b101 %
1'
b101 +
#74630000000
0!
0'
#74640000000
1!
b110 %
1'
b110 +
#74650000000
0!
0'
#74660000000
1!
b111 %
1'
b111 +
#74670000000
0!
0'
#74680000000
1!
0$
b1000 %
1'
0*
b1000 +
#74690000000
0!
0'
#74700000000
1!
b1001 %
1'
b1001 +
#74710000000
0!
0'
#74720000000
1!
b0 %
1'
b0 +
#74730000000
0!
0'
#74740000000
1!
1$
b1 %
1'
1*
b1 +
#74750000000
0!
0'
#74760000000
1!
b10 %
1'
b10 +
#74770000000
0!
0'
#74780000000
1!
b11 %
1'
b11 +
#74790000000
0!
0'
#74800000000
1!
b100 %
1'
b100 +
#74810000000
0!
0'
#74820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#74830000000
0!
0'
#74840000000
1!
0$
b110 %
1'
0*
b110 +
#74850000000
0!
0'
#74860000000
1!
b111 %
1'
b111 +
#74870000000
0!
0'
#74880000000
1!
b1000 %
1'
b1000 +
#74890000000
0!
0'
#74900000000
1!
b1001 %
1'
b1001 +
#74910000000
0!
0'
#74920000000
1!
b0 %
1'
b0 +
#74930000000
0!
0'
#74940000000
1!
1$
b1 %
1'
1*
b1 +
#74950000000
0!
0'
#74960000000
1!
b10 %
1'
b10 +
#74970000000
0!
0'
#74980000000
1!
b11 %
1'
b11 +
#74990000000
0!
0'
#75000000000
1!
b100 %
1'
b100 +
#75010000000
0!
0'
#75020000000
1!
b101 %
1'
b101 +
#75030000000
1"
1(
#75040000000
0!
0"
b100 &
0'
0(
b100 ,
#75050000000
1!
b110 %
1'
b110 +
#75060000000
0!
0'
#75070000000
1!
b111 %
1'
b111 +
#75080000000
0!
0'
#75090000000
1!
0$
b1000 %
1'
0*
b1000 +
#75100000000
0!
0'
#75110000000
1!
b1001 %
1'
b1001 +
#75120000000
0!
0'
#75130000000
1!
b0 %
1'
b0 +
#75140000000
0!
0'
#75150000000
1!
1$
b1 %
1'
1*
b1 +
#75160000000
0!
0'
#75170000000
1!
b10 %
1'
b10 +
#75180000000
0!
0'
#75190000000
1!
b11 %
1'
b11 +
#75200000000
0!
0'
#75210000000
1!
b100 %
1'
b100 +
#75220000000
0!
0'
#75230000000
1!
b101 %
1'
b101 +
#75240000000
0!
0'
#75250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#75260000000
0!
0'
#75270000000
1!
b111 %
1'
b111 +
#75280000000
0!
0'
#75290000000
1!
b1000 %
1'
b1000 +
#75300000000
0!
0'
#75310000000
1!
b1001 %
1'
b1001 +
#75320000000
0!
0'
#75330000000
1!
b0 %
1'
b0 +
#75340000000
0!
0'
#75350000000
1!
1$
b1 %
1'
1*
b1 +
#75360000000
0!
0'
#75370000000
1!
b10 %
1'
b10 +
#75380000000
0!
0'
#75390000000
1!
b11 %
1'
b11 +
#75400000000
0!
0'
#75410000000
1!
b100 %
1'
b100 +
#75420000000
0!
0'
#75430000000
1!
b101 %
1'
b101 +
#75440000000
0!
0'
#75450000000
1!
0$
b110 %
1'
0*
b110 +
#75460000000
1"
1(
#75470000000
0!
0"
b100 &
0'
0(
b100 ,
#75480000000
1!
1$
b111 %
1'
1*
b111 +
#75490000000
0!
0'
#75500000000
1!
0$
b1000 %
1'
0*
b1000 +
#75510000000
0!
0'
#75520000000
1!
b1001 %
1'
b1001 +
#75530000000
0!
0'
#75540000000
1!
b0 %
1'
b0 +
#75550000000
0!
0'
#75560000000
1!
1$
b1 %
1'
1*
b1 +
#75570000000
0!
0'
#75580000000
1!
b10 %
1'
b10 +
#75590000000
0!
0'
#75600000000
1!
b11 %
1'
b11 +
#75610000000
0!
0'
#75620000000
1!
b100 %
1'
b100 +
#75630000000
0!
0'
#75640000000
1!
b101 %
1'
b101 +
#75650000000
0!
0'
#75660000000
1!
b110 %
1'
b110 +
#75670000000
0!
0'
#75680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#75690000000
0!
0'
#75700000000
1!
b1000 %
1'
b1000 +
#75710000000
0!
0'
#75720000000
1!
b1001 %
1'
b1001 +
#75730000000
0!
0'
#75740000000
1!
b0 %
1'
b0 +
#75750000000
0!
0'
#75760000000
1!
1$
b1 %
1'
1*
b1 +
#75770000000
0!
0'
#75780000000
1!
b10 %
1'
b10 +
#75790000000
0!
0'
#75800000000
1!
b11 %
1'
b11 +
#75810000000
0!
0'
#75820000000
1!
b100 %
1'
b100 +
#75830000000
0!
0'
#75840000000
1!
b101 %
1'
b101 +
#75850000000
0!
0'
#75860000000
1!
0$
b110 %
1'
0*
b110 +
#75870000000
0!
0'
#75880000000
1!
b111 %
1'
b111 +
#75890000000
1"
1(
#75900000000
0!
0"
b100 &
0'
0(
b100 ,
#75910000000
1!
b1000 %
1'
b1000 +
#75920000000
0!
0'
#75930000000
1!
b1001 %
1'
b1001 +
#75940000000
0!
0'
#75950000000
1!
b0 %
1'
b0 +
#75960000000
0!
0'
#75970000000
1!
1$
b1 %
1'
1*
b1 +
#75980000000
0!
0'
#75990000000
1!
b10 %
1'
b10 +
#76000000000
0!
0'
#76010000000
1!
b11 %
1'
b11 +
#76020000000
0!
0'
#76030000000
1!
b100 %
1'
b100 +
#76040000000
0!
0'
#76050000000
1!
b101 %
1'
b101 +
#76060000000
0!
0'
#76070000000
1!
b110 %
1'
b110 +
#76080000000
0!
0'
#76090000000
1!
b111 %
1'
b111 +
#76100000000
0!
0'
#76110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#76120000000
0!
0'
#76130000000
1!
b1001 %
1'
b1001 +
#76140000000
0!
0'
#76150000000
1!
b0 %
1'
b0 +
#76160000000
0!
0'
#76170000000
1!
1$
b1 %
1'
1*
b1 +
#76180000000
0!
0'
#76190000000
1!
b10 %
1'
b10 +
#76200000000
0!
0'
#76210000000
1!
b11 %
1'
b11 +
#76220000000
0!
0'
#76230000000
1!
b100 %
1'
b100 +
#76240000000
0!
0'
#76250000000
1!
b101 %
1'
b101 +
#76260000000
0!
0'
#76270000000
1!
0$
b110 %
1'
0*
b110 +
#76280000000
0!
0'
#76290000000
1!
b111 %
1'
b111 +
#76300000000
0!
0'
#76310000000
1!
b1000 %
1'
b1000 +
#76320000000
1"
1(
#76330000000
0!
0"
b100 &
0'
0(
b100 ,
#76340000000
1!
b1001 %
1'
b1001 +
#76350000000
0!
0'
#76360000000
1!
b0 %
1'
b0 +
#76370000000
0!
0'
#76380000000
1!
1$
b1 %
1'
1*
b1 +
#76390000000
0!
0'
#76400000000
1!
b10 %
1'
b10 +
#76410000000
0!
0'
#76420000000
1!
b11 %
1'
b11 +
#76430000000
0!
0'
#76440000000
1!
b100 %
1'
b100 +
#76450000000
0!
0'
#76460000000
1!
b101 %
1'
b101 +
#76470000000
0!
0'
#76480000000
1!
b110 %
1'
b110 +
#76490000000
0!
0'
#76500000000
1!
b111 %
1'
b111 +
#76510000000
0!
0'
#76520000000
1!
0$
b1000 %
1'
0*
b1000 +
#76530000000
0!
0'
#76540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#76550000000
0!
0'
#76560000000
1!
b0 %
1'
b0 +
#76570000000
0!
0'
#76580000000
1!
1$
b1 %
1'
1*
b1 +
#76590000000
0!
0'
#76600000000
1!
b10 %
1'
b10 +
#76610000000
0!
0'
#76620000000
1!
b11 %
1'
b11 +
#76630000000
0!
0'
#76640000000
1!
b100 %
1'
b100 +
#76650000000
0!
0'
#76660000000
1!
b101 %
1'
b101 +
#76670000000
0!
0'
#76680000000
1!
0$
b110 %
1'
0*
b110 +
#76690000000
0!
0'
#76700000000
1!
b111 %
1'
b111 +
#76710000000
0!
0'
#76720000000
1!
b1000 %
1'
b1000 +
#76730000000
0!
0'
#76740000000
1!
b1001 %
1'
b1001 +
#76750000000
1"
1(
#76760000000
0!
0"
b100 &
0'
0(
b100 ,
#76770000000
1!
b0 %
1'
b0 +
#76780000000
0!
0'
#76790000000
1!
1$
b1 %
1'
1*
b1 +
#76800000000
0!
0'
#76810000000
1!
b10 %
1'
b10 +
#76820000000
0!
0'
#76830000000
1!
b11 %
1'
b11 +
#76840000000
0!
0'
#76850000000
1!
b100 %
1'
b100 +
#76860000000
0!
0'
#76870000000
1!
b101 %
1'
b101 +
#76880000000
0!
0'
#76890000000
1!
b110 %
1'
b110 +
#76900000000
0!
0'
#76910000000
1!
b111 %
1'
b111 +
#76920000000
0!
0'
#76930000000
1!
0$
b1000 %
1'
0*
b1000 +
#76940000000
0!
0'
#76950000000
1!
b1001 %
1'
b1001 +
#76960000000
0!
0'
#76970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#76980000000
0!
0'
#76990000000
1!
1$
b1 %
1'
1*
b1 +
#77000000000
0!
0'
#77010000000
1!
b10 %
1'
b10 +
#77020000000
0!
0'
#77030000000
1!
b11 %
1'
b11 +
#77040000000
0!
0'
#77050000000
1!
b100 %
1'
b100 +
#77060000000
0!
0'
#77070000000
1!
b101 %
1'
b101 +
#77080000000
0!
0'
#77090000000
1!
0$
b110 %
1'
0*
b110 +
#77100000000
0!
0'
#77110000000
1!
b111 %
1'
b111 +
#77120000000
0!
0'
#77130000000
1!
b1000 %
1'
b1000 +
#77140000000
0!
0'
#77150000000
1!
b1001 %
1'
b1001 +
#77160000000
0!
0'
#77170000000
1!
b0 %
1'
b0 +
#77180000000
1"
1(
#77190000000
0!
0"
b100 &
0'
0(
b100 ,
#77200000000
1!
1$
b1 %
1'
1*
b1 +
#77210000000
0!
0'
#77220000000
1!
b10 %
1'
b10 +
#77230000000
0!
0'
#77240000000
1!
b11 %
1'
b11 +
#77250000000
0!
0'
#77260000000
1!
b100 %
1'
b100 +
#77270000000
0!
0'
#77280000000
1!
b101 %
1'
b101 +
#77290000000
0!
0'
#77300000000
1!
b110 %
1'
b110 +
#77310000000
0!
0'
#77320000000
1!
b111 %
1'
b111 +
#77330000000
0!
0'
#77340000000
1!
0$
b1000 %
1'
0*
b1000 +
#77350000000
0!
0'
#77360000000
1!
b1001 %
1'
b1001 +
#77370000000
0!
0'
#77380000000
1!
b0 %
1'
b0 +
#77390000000
0!
0'
#77400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#77410000000
0!
0'
#77420000000
1!
b10 %
1'
b10 +
#77430000000
0!
0'
#77440000000
1!
b11 %
1'
b11 +
#77450000000
0!
0'
#77460000000
1!
b100 %
1'
b100 +
#77470000000
0!
0'
#77480000000
1!
b101 %
1'
b101 +
#77490000000
0!
0'
#77500000000
1!
0$
b110 %
1'
0*
b110 +
#77510000000
0!
0'
#77520000000
1!
b111 %
1'
b111 +
#77530000000
0!
0'
#77540000000
1!
b1000 %
1'
b1000 +
#77550000000
0!
0'
#77560000000
1!
b1001 %
1'
b1001 +
#77570000000
0!
0'
#77580000000
1!
b0 %
1'
b0 +
#77590000000
0!
0'
#77600000000
1!
1$
b1 %
1'
1*
b1 +
#77610000000
1"
1(
#77620000000
0!
0"
b100 &
0'
0(
b100 ,
#77630000000
1!
b10 %
1'
b10 +
#77640000000
0!
0'
#77650000000
1!
b11 %
1'
b11 +
#77660000000
0!
0'
#77670000000
1!
b100 %
1'
b100 +
#77680000000
0!
0'
#77690000000
1!
b101 %
1'
b101 +
#77700000000
0!
0'
#77710000000
1!
b110 %
1'
b110 +
#77720000000
0!
0'
#77730000000
1!
b111 %
1'
b111 +
#77740000000
0!
0'
#77750000000
1!
0$
b1000 %
1'
0*
b1000 +
#77760000000
0!
0'
#77770000000
1!
b1001 %
1'
b1001 +
#77780000000
0!
0'
#77790000000
1!
b0 %
1'
b0 +
#77800000000
0!
0'
#77810000000
1!
1$
b1 %
1'
1*
b1 +
#77820000000
0!
0'
#77830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#77840000000
0!
0'
#77850000000
1!
b11 %
1'
b11 +
#77860000000
0!
0'
#77870000000
1!
b100 %
1'
b100 +
#77880000000
0!
0'
#77890000000
1!
b101 %
1'
b101 +
#77900000000
0!
0'
#77910000000
1!
0$
b110 %
1'
0*
b110 +
#77920000000
0!
0'
#77930000000
1!
b111 %
1'
b111 +
#77940000000
0!
0'
#77950000000
1!
b1000 %
1'
b1000 +
#77960000000
0!
0'
#77970000000
1!
b1001 %
1'
b1001 +
#77980000000
0!
0'
#77990000000
1!
b0 %
1'
b0 +
#78000000000
0!
0'
#78010000000
1!
1$
b1 %
1'
1*
b1 +
#78020000000
0!
0'
#78030000000
1!
b10 %
1'
b10 +
#78040000000
1"
1(
#78050000000
0!
0"
b100 &
0'
0(
b100 ,
#78060000000
1!
b11 %
1'
b11 +
#78070000000
0!
0'
#78080000000
1!
b100 %
1'
b100 +
#78090000000
0!
0'
#78100000000
1!
b101 %
1'
b101 +
#78110000000
0!
0'
#78120000000
1!
b110 %
1'
b110 +
#78130000000
0!
0'
#78140000000
1!
b111 %
1'
b111 +
#78150000000
0!
0'
#78160000000
1!
0$
b1000 %
1'
0*
b1000 +
#78170000000
0!
0'
#78180000000
1!
b1001 %
1'
b1001 +
#78190000000
0!
0'
#78200000000
1!
b0 %
1'
b0 +
#78210000000
0!
0'
#78220000000
1!
1$
b1 %
1'
1*
b1 +
#78230000000
0!
0'
#78240000000
1!
b10 %
1'
b10 +
#78250000000
0!
0'
#78260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#78270000000
0!
0'
#78280000000
1!
b100 %
1'
b100 +
#78290000000
0!
0'
#78300000000
1!
b101 %
1'
b101 +
#78310000000
0!
0'
#78320000000
1!
0$
b110 %
1'
0*
b110 +
#78330000000
0!
0'
#78340000000
1!
b111 %
1'
b111 +
#78350000000
0!
0'
#78360000000
1!
b1000 %
1'
b1000 +
#78370000000
0!
0'
#78380000000
1!
b1001 %
1'
b1001 +
#78390000000
0!
0'
#78400000000
1!
b0 %
1'
b0 +
#78410000000
0!
0'
#78420000000
1!
1$
b1 %
1'
1*
b1 +
#78430000000
0!
0'
#78440000000
1!
b10 %
1'
b10 +
#78450000000
0!
0'
#78460000000
1!
b11 %
1'
b11 +
#78470000000
1"
1(
#78480000000
0!
0"
b100 &
0'
0(
b100 ,
#78490000000
1!
b100 %
1'
b100 +
#78500000000
0!
0'
#78510000000
1!
b101 %
1'
b101 +
#78520000000
0!
0'
#78530000000
1!
b110 %
1'
b110 +
#78540000000
0!
0'
#78550000000
1!
b111 %
1'
b111 +
#78560000000
0!
0'
#78570000000
1!
0$
b1000 %
1'
0*
b1000 +
#78580000000
0!
0'
#78590000000
1!
b1001 %
1'
b1001 +
#78600000000
0!
0'
#78610000000
1!
b0 %
1'
b0 +
#78620000000
0!
0'
#78630000000
1!
1$
b1 %
1'
1*
b1 +
#78640000000
0!
0'
#78650000000
1!
b10 %
1'
b10 +
#78660000000
0!
0'
#78670000000
1!
b11 %
1'
b11 +
#78680000000
0!
0'
#78690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#78700000000
0!
0'
#78710000000
1!
b101 %
1'
b101 +
#78720000000
0!
0'
#78730000000
1!
0$
b110 %
1'
0*
b110 +
#78740000000
0!
0'
#78750000000
1!
b111 %
1'
b111 +
#78760000000
0!
0'
#78770000000
1!
b1000 %
1'
b1000 +
#78780000000
0!
0'
#78790000000
1!
b1001 %
1'
b1001 +
#78800000000
0!
0'
#78810000000
1!
b0 %
1'
b0 +
#78820000000
0!
0'
#78830000000
1!
1$
b1 %
1'
1*
b1 +
#78840000000
0!
0'
#78850000000
1!
b10 %
1'
b10 +
#78860000000
0!
0'
#78870000000
1!
b11 %
1'
b11 +
#78880000000
0!
0'
#78890000000
1!
b100 %
1'
b100 +
#78900000000
1"
1(
#78910000000
0!
0"
b100 &
0'
0(
b100 ,
#78920000000
1!
b101 %
1'
b101 +
#78930000000
0!
0'
#78940000000
1!
b110 %
1'
b110 +
#78950000000
0!
0'
#78960000000
1!
b111 %
1'
b111 +
#78970000000
0!
0'
#78980000000
1!
0$
b1000 %
1'
0*
b1000 +
#78990000000
0!
0'
#79000000000
1!
b1001 %
1'
b1001 +
#79010000000
0!
0'
#79020000000
1!
b0 %
1'
b0 +
#79030000000
0!
0'
#79040000000
1!
1$
b1 %
1'
1*
b1 +
#79050000000
0!
0'
#79060000000
1!
b10 %
1'
b10 +
#79070000000
0!
0'
#79080000000
1!
b11 %
1'
b11 +
#79090000000
0!
0'
#79100000000
1!
b100 %
1'
b100 +
#79110000000
0!
0'
#79120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#79130000000
0!
0'
#79140000000
1!
0$
b110 %
1'
0*
b110 +
#79150000000
0!
0'
#79160000000
1!
b111 %
1'
b111 +
#79170000000
0!
0'
#79180000000
1!
b1000 %
1'
b1000 +
#79190000000
0!
0'
#79200000000
1!
b1001 %
1'
b1001 +
#79210000000
0!
0'
#79220000000
1!
b0 %
1'
b0 +
#79230000000
0!
0'
#79240000000
1!
1$
b1 %
1'
1*
b1 +
#79250000000
0!
0'
#79260000000
1!
b10 %
1'
b10 +
#79270000000
0!
0'
#79280000000
1!
b11 %
1'
b11 +
#79290000000
0!
0'
#79300000000
1!
b100 %
1'
b100 +
#79310000000
0!
0'
#79320000000
1!
b101 %
1'
b101 +
#79330000000
1"
1(
#79340000000
0!
0"
b100 &
0'
0(
b100 ,
#79350000000
1!
b110 %
1'
b110 +
#79360000000
0!
0'
#79370000000
1!
b111 %
1'
b111 +
#79380000000
0!
0'
#79390000000
1!
0$
b1000 %
1'
0*
b1000 +
#79400000000
0!
0'
#79410000000
1!
b1001 %
1'
b1001 +
#79420000000
0!
0'
#79430000000
1!
b0 %
1'
b0 +
#79440000000
0!
0'
#79450000000
1!
1$
b1 %
1'
1*
b1 +
#79460000000
0!
0'
#79470000000
1!
b10 %
1'
b10 +
#79480000000
0!
0'
#79490000000
1!
b11 %
1'
b11 +
#79500000000
0!
0'
#79510000000
1!
b100 %
1'
b100 +
#79520000000
0!
0'
#79530000000
1!
b101 %
1'
b101 +
#79540000000
0!
0'
#79550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#79560000000
0!
0'
#79570000000
1!
b111 %
1'
b111 +
#79580000000
0!
0'
#79590000000
1!
b1000 %
1'
b1000 +
#79600000000
0!
0'
#79610000000
1!
b1001 %
1'
b1001 +
#79620000000
0!
0'
#79630000000
1!
b0 %
1'
b0 +
#79640000000
0!
0'
#79650000000
1!
1$
b1 %
1'
1*
b1 +
#79660000000
0!
0'
#79670000000
1!
b10 %
1'
b10 +
#79680000000
0!
0'
#79690000000
1!
b11 %
1'
b11 +
#79700000000
0!
0'
#79710000000
1!
b100 %
1'
b100 +
#79720000000
0!
0'
#79730000000
1!
b101 %
1'
b101 +
#79740000000
0!
0'
#79750000000
1!
0$
b110 %
1'
0*
b110 +
#79760000000
1"
1(
#79770000000
0!
0"
b100 &
0'
0(
b100 ,
#79780000000
1!
1$
b111 %
1'
1*
b111 +
#79790000000
0!
0'
#79800000000
1!
0$
b1000 %
1'
0*
b1000 +
#79810000000
0!
0'
#79820000000
1!
b1001 %
1'
b1001 +
#79830000000
0!
0'
#79840000000
1!
b0 %
1'
b0 +
#79850000000
0!
0'
#79860000000
1!
1$
b1 %
1'
1*
b1 +
#79870000000
0!
0'
#79880000000
1!
b10 %
1'
b10 +
#79890000000
0!
0'
#79900000000
1!
b11 %
1'
b11 +
#79910000000
0!
0'
#79920000000
1!
b100 %
1'
b100 +
#79930000000
0!
0'
#79940000000
1!
b101 %
1'
b101 +
#79950000000
0!
0'
#79960000000
1!
b110 %
1'
b110 +
#79970000000
0!
0'
#79980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#79990000000
0!
0'
#80000000000
1!
b1000 %
1'
b1000 +
#80010000000
0!
0'
#80020000000
1!
b1001 %
1'
b1001 +
#80030000000
0!
0'
#80040000000
1!
b0 %
1'
b0 +
#80050000000
0!
0'
#80060000000
1!
1$
b1 %
1'
1*
b1 +
#80070000000
0!
0'
#80080000000
1!
b10 %
1'
b10 +
#80090000000
0!
0'
#80100000000
1!
b11 %
1'
b11 +
#80110000000
0!
0'
#80120000000
1!
b100 %
1'
b100 +
#80130000000
0!
0'
#80140000000
1!
b101 %
1'
b101 +
#80150000000
0!
0'
#80160000000
1!
0$
b110 %
1'
0*
b110 +
#80170000000
0!
0'
#80180000000
1!
b111 %
1'
b111 +
#80190000000
1"
1(
#80200000000
0!
0"
b100 &
0'
0(
b100 ,
#80210000000
1!
b1000 %
1'
b1000 +
#80220000000
0!
0'
#80230000000
1!
b1001 %
1'
b1001 +
#80240000000
0!
0'
#80250000000
1!
b0 %
1'
b0 +
#80260000000
0!
0'
#80270000000
1!
1$
b1 %
1'
1*
b1 +
#80280000000
0!
0'
#80290000000
1!
b10 %
1'
b10 +
#80300000000
0!
0'
#80310000000
1!
b11 %
1'
b11 +
#80320000000
0!
0'
#80330000000
1!
b100 %
1'
b100 +
#80340000000
0!
0'
#80350000000
1!
b101 %
1'
b101 +
#80360000000
0!
0'
#80370000000
1!
b110 %
1'
b110 +
#80380000000
0!
0'
#80390000000
1!
b111 %
1'
b111 +
#80400000000
0!
0'
#80410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#80420000000
0!
0'
#80430000000
1!
b1001 %
1'
b1001 +
#80440000000
0!
0'
#80450000000
1!
b0 %
1'
b0 +
#80460000000
0!
0'
#80470000000
1!
1$
b1 %
1'
1*
b1 +
#80480000000
0!
0'
#80490000000
1!
b10 %
1'
b10 +
#80500000000
0!
0'
#80510000000
1!
b11 %
1'
b11 +
#80520000000
0!
0'
#80530000000
1!
b100 %
1'
b100 +
#80540000000
0!
0'
#80550000000
1!
b101 %
1'
b101 +
#80560000000
0!
0'
#80570000000
1!
0$
b110 %
1'
0*
b110 +
#80580000000
0!
0'
#80590000000
1!
b111 %
1'
b111 +
#80600000000
0!
0'
#80610000000
1!
b1000 %
1'
b1000 +
#80620000000
1"
1(
#80630000000
0!
0"
b100 &
0'
0(
b100 ,
#80640000000
1!
b1001 %
1'
b1001 +
#80650000000
0!
0'
#80660000000
1!
b0 %
1'
b0 +
#80670000000
0!
0'
#80680000000
1!
1$
b1 %
1'
1*
b1 +
#80690000000
0!
0'
#80700000000
1!
b10 %
1'
b10 +
#80710000000
0!
0'
#80720000000
1!
b11 %
1'
b11 +
#80730000000
0!
0'
#80740000000
1!
b100 %
1'
b100 +
#80750000000
0!
0'
#80760000000
1!
b101 %
1'
b101 +
#80770000000
0!
0'
#80780000000
1!
b110 %
1'
b110 +
#80790000000
0!
0'
#80800000000
1!
b111 %
1'
b111 +
#80810000000
0!
0'
#80820000000
1!
0$
b1000 %
1'
0*
b1000 +
#80830000000
0!
0'
#80840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#80850000000
0!
0'
#80860000000
1!
b0 %
1'
b0 +
#80870000000
0!
0'
#80880000000
1!
1$
b1 %
1'
1*
b1 +
#80890000000
0!
0'
#80900000000
1!
b10 %
1'
b10 +
#80910000000
0!
0'
#80920000000
1!
b11 %
1'
b11 +
#80930000000
0!
0'
#80940000000
1!
b100 %
1'
b100 +
#80950000000
0!
0'
#80960000000
1!
b101 %
1'
b101 +
#80970000000
0!
0'
#80980000000
1!
0$
b110 %
1'
0*
b110 +
#80990000000
0!
0'
#81000000000
1!
b111 %
1'
b111 +
#81010000000
0!
0'
#81020000000
1!
b1000 %
1'
b1000 +
#81030000000
0!
0'
#81040000000
1!
b1001 %
1'
b1001 +
#81050000000
1"
1(
#81060000000
0!
0"
b100 &
0'
0(
b100 ,
#81070000000
1!
b0 %
1'
b0 +
#81080000000
0!
0'
#81090000000
1!
1$
b1 %
1'
1*
b1 +
#81100000000
0!
0'
#81110000000
1!
b10 %
1'
b10 +
#81120000000
0!
0'
#81130000000
1!
b11 %
1'
b11 +
#81140000000
0!
0'
#81150000000
1!
b100 %
1'
b100 +
#81160000000
0!
0'
#81170000000
1!
b101 %
1'
b101 +
#81180000000
0!
0'
#81190000000
1!
b110 %
1'
b110 +
#81200000000
0!
0'
#81210000000
1!
b111 %
1'
b111 +
#81220000000
0!
0'
#81230000000
1!
0$
b1000 %
1'
0*
b1000 +
#81240000000
0!
0'
#81250000000
1!
b1001 %
1'
b1001 +
#81260000000
0!
0'
#81270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#81280000000
0!
0'
#81290000000
1!
1$
b1 %
1'
1*
b1 +
#81300000000
0!
0'
#81310000000
1!
b10 %
1'
b10 +
#81320000000
0!
0'
#81330000000
1!
b11 %
1'
b11 +
#81340000000
0!
0'
#81350000000
1!
b100 %
1'
b100 +
#81360000000
0!
0'
#81370000000
1!
b101 %
1'
b101 +
#81380000000
0!
0'
#81390000000
1!
0$
b110 %
1'
0*
b110 +
#81400000000
0!
0'
#81410000000
1!
b111 %
1'
b111 +
#81420000000
0!
0'
#81430000000
1!
b1000 %
1'
b1000 +
#81440000000
0!
0'
#81450000000
1!
b1001 %
1'
b1001 +
#81460000000
0!
0'
#81470000000
1!
b0 %
1'
b0 +
#81480000000
1"
1(
#81490000000
0!
0"
b100 &
0'
0(
b100 ,
#81500000000
1!
1$
b1 %
1'
1*
b1 +
#81510000000
0!
0'
#81520000000
1!
b10 %
1'
b10 +
#81530000000
0!
0'
#81540000000
1!
b11 %
1'
b11 +
#81550000000
0!
0'
#81560000000
1!
b100 %
1'
b100 +
#81570000000
0!
0'
#81580000000
1!
b101 %
1'
b101 +
#81590000000
0!
0'
#81600000000
1!
b110 %
1'
b110 +
#81610000000
0!
0'
#81620000000
1!
b111 %
1'
b111 +
#81630000000
0!
0'
#81640000000
1!
0$
b1000 %
1'
0*
b1000 +
#81650000000
0!
0'
#81660000000
1!
b1001 %
1'
b1001 +
#81670000000
0!
0'
#81680000000
1!
b0 %
1'
b0 +
#81690000000
0!
0'
#81700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#81710000000
0!
0'
#81720000000
1!
b10 %
1'
b10 +
#81730000000
0!
0'
#81740000000
1!
b11 %
1'
b11 +
#81750000000
0!
0'
#81760000000
1!
b100 %
1'
b100 +
#81770000000
0!
0'
#81780000000
1!
b101 %
1'
b101 +
#81790000000
0!
0'
#81800000000
1!
0$
b110 %
1'
0*
b110 +
#81810000000
0!
0'
#81820000000
1!
b111 %
1'
b111 +
#81830000000
0!
0'
#81840000000
1!
b1000 %
1'
b1000 +
#81850000000
0!
0'
#81860000000
1!
b1001 %
1'
b1001 +
#81870000000
0!
0'
#81880000000
1!
b0 %
1'
b0 +
#81890000000
0!
0'
#81900000000
1!
1$
b1 %
1'
1*
b1 +
#81910000000
1"
1(
#81920000000
0!
0"
b100 &
0'
0(
b100 ,
#81930000000
1!
b10 %
1'
b10 +
#81940000000
0!
0'
#81950000000
1!
b11 %
1'
b11 +
#81960000000
0!
0'
#81970000000
1!
b100 %
1'
b100 +
#81980000000
0!
0'
#81990000000
1!
b101 %
1'
b101 +
#82000000000
0!
0'
#82010000000
1!
b110 %
1'
b110 +
#82020000000
0!
0'
#82030000000
1!
b111 %
1'
b111 +
#82040000000
0!
0'
#82050000000
1!
0$
b1000 %
1'
0*
b1000 +
#82060000000
0!
0'
#82070000000
1!
b1001 %
1'
b1001 +
#82080000000
0!
0'
#82090000000
1!
b0 %
1'
b0 +
#82100000000
0!
0'
#82110000000
1!
1$
b1 %
1'
1*
b1 +
#82120000000
0!
0'
#82130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#82140000000
0!
0'
#82150000000
1!
b11 %
1'
b11 +
#82160000000
0!
0'
#82170000000
1!
b100 %
1'
b100 +
#82180000000
0!
0'
#82190000000
1!
b101 %
1'
b101 +
#82200000000
0!
0'
#82210000000
1!
0$
b110 %
1'
0*
b110 +
#82220000000
0!
0'
#82230000000
1!
b111 %
1'
b111 +
#82240000000
0!
0'
#82250000000
1!
b1000 %
1'
b1000 +
#82260000000
0!
0'
#82270000000
1!
b1001 %
1'
b1001 +
#82280000000
0!
0'
#82290000000
1!
b0 %
1'
b0 +
#82300000000
0!
0'
#82310000000
1!
1$
b1 %
1'
1*
b1 +
#82320000000
0!
0'
#82330000000
1!
b10 %
1'
b10 +
#82340000000
1"
1(
#82350000000
0!
0"
b100 &
0'
0(
b100 ,
#82360000000
1!
b11 %
1'
b11 +
#82370000000
0!
0'
#82380000000
1!
b100 %
1'
b100 +
#82390000000
0!
0'
#82400000000
1!
b101 %
1'
b101 +
#82410000000
0!
0'
#82420000000
1!
b110 %
1'
b110 +
#82430000000
0!
0'
#82440000000
1!
b111 %
1'
b111 +
#82450000000
0!
0'
#82460000000
1!
0$
b1000 %
1'
0*
b1000 +
#82470000000
0!
0'
#82480000000
1!
b1001 %
1'
b1001 +
#82490000000
0!
0'
#82500000000
1!
b0 %
1'
b0 +
#82510000000
0!
0'
#82520000000
1!
1$
b1 %
1'
1*
b1 +
#82530000000
0!
0'
#82540000000
1!
b10 %
1'
b10 +
#82550000000
0!
0'
#82560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#82570000000
0!
0'
#82580000000
1!
b100 %
1'
b100 +
#82590000000
0!
0'
#82600000000
1!
b101 %
1'
b101 +
#82610000000
0!
0'
#82620000000
1!
0$
b110 %
1'
0*
b110 +
#82630000000
0!
0'
#82640000000
1!
b111 %
1'
b111 +
#82650000000
0!
0'
#82660000000
1!
b1000 %
1'
b1000 +
#82670000000
0!
0'
#82680000000
1!
b1001 %
1'
b1001 +
#82690000000
0!
0'
#82700000000
1!
b0 %
1'
b0 +
#82710000000
0!
0'
#82720000000
1!
1$
b1 %
1'
1*
b1 +
#82730000000
0!
0'
#82740000000
1!
b10 %
1'
b10 +
#82750000000
0!
0'
#82760000000
1!
b11 %
1'
b11 +
#82770000000
1"
1(
#82780000000
0!
0"
b100 &
0'
0(
b100 ,
#82790000000
1!
b100 %
1'
b100 +
#82800000000
0!
0'
#82810000000
1!
b101 %
1'
b101 +
#82820000000
0!
0'
#82830000000
1!
b110 %
1'
b110 +
#82840000000
0!
0'
#82850000000
1!
b111 %
1'
b111 +
#82860000000
0!
0'
#82870000000
1!
0$
b1000 %
1'
0*
b1000 +
#82880000000
0!
0'
#82890000000
1!
b1001 %
1'
b1001 +
#82900000000
0!
0'
#82910000000
1!
b0 %
1'
b0 +
#82920000000
0!
0'
#82930000000
1!
1$
b1 %
1'
1*
b1 +
#82940000000
0!
0'
#82950000000
1!
b10 %
1'
b10 +
#82960000000
0!
0'
#82970000000
1!
b11 %
1'
b11 +
#82980000000
0!
0'
#82990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#83000000000
0!
0'
#83010000000
1!
b101 %
1'
b101 +
#83020000000
0!
0'
#83030000000
1!
0$
b110 %
1'
0*
b110 +
#83040000000
0!
0'
#83050000000
1!
b111 %
1'
b111 +
#83060000000
0!
0'
#83070000000
1!
b1000 %
1'
b1000 +
#83080000000
0!
0'
#83090000000
1!
b1001 %
1'
b1001 +
#83100000000
0!
0'
#83110000000
1!
b0 %
1'
b0 +
#83120000000
0!
0'
#83130000000
1!
1$
b1 %
1'
1*
b1 +
#83140000000
0!
0'
#83150000000
1!
b10 %
1'
b10 +
#83160000000
0!
0'
#83170000000
1!
b11 %
1'
b11 +
#83180000000
0!
0'
#83190000000
1!
b100 %
1'
b100 +
#83200000000
1"
1(
#83210000000
0!
0"
b100 &
0'
0(
b100 ,
#83220000000
1!
b101 %
1'
b101 +
#83230000000
0!
0'
#83240000000
1!
b110 %
1'
b110 +
#83250000000
0!
0'
#83260000000
1!
b111 %
1'
b111 +
#83270000000
0!
0'
#83280000000
1!
0$
b1000 %
1'
0*
b1000 +
#83290000000
0!
0'
#83300000000
1!
b1001 %
1'
b1001 +
#83310000000
0!
0'
#83320000000
1!
b0 %
1'
b0 +
#83330000000
0!
0'
#83340000000
1!
1$
b1 %
1'
1*
b1 +
#83350000000
0!
0'
#83360000000
1!
b10 %
1'
b10 +
#83370000000
0!
0'
#83380000000
1!
b11 %
1'
b11 +
#83390000000
0!
0'
#83400000000
1!
b100 %
1'
b100 +
#83410000000
0!
0'
#83420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#83430000000
0!
0'
#83440000000
1!
0$
b110 %
1'
0*
b110 +
#83450000000
0!
0'
#83460000000
1!
b111 %
1'
b111 +
#83470000000
0!
0'
#83480000000
1!
b1000 %
1'
b1000 +
#83490000000
0!
0'
#83500000000
1!
b1001 %
1'
b1001 +
#83510000000
0!
0'
#83520000000
1!
b0 %
1'
b0 +
#83530000000
0!
0'
#83540000000
1!
1$
b1 %
1'
1*
b1 +
#83550000000
0!
0'
#83560000000
1!
b10 %
1'
b10 +
#83570000000
0!
0'
#83580000000
1!
b11 %
1'
b11 +
#83590000000
0!
0'
#83600000000
1!
b100 %
1'
b100 +
#83610000000
0!
0'
#83620000000
1!
b101 %
1'
b101 +
#83630000000
1"
1(
#83640000000
0!
0"
b100 &
0'
0(
b100 ,
#83650000000
1!
b110 %
1'
b110 +
#83660000000
0!
0'
#83670000000
1!
b111 %
1'
b111 +
#83680000000
0!
0'
#83690000000
1!
0$
b1000 %
1'
0*
b1000 +
#83700000000
0!
0'
#83710000000
1!
b1001 %
1'
b1001 +
#83720000000
0!
0'
#83730000000
1!
b0 %
1'
b0 +
#83740000000
0!
0'
#83750000000
1!
1$
b1 %
1'
1*
b1 +
#83760000000
0!
0'
#83770000000
1!
b10 %
1'
b10 +
#83780000000
0!
0'
#83790000000
1!
b11 %
1'
b11 +
#83800000000
0!
0'
#83810000000
1!
b100 %
1'
b100 +
#83820000000
0!
0'
#83830000000
1!
b101 %
1'
b101 +
#83840000000
0!
0'
#83850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#83860000000
0!
0'
#83870000000
1!
b111 %
1'
b111 +
#83880000000
0!
0'
#83890000000
1!
b1000 %
1'
b1000 +
#83900000000
0!
0'
#83910000000
1!
b1001 %
1'
b1001 +
#83920000000
0!
0'
#83930000000
1!
b0 %
1'
b0 +
#83940000000
0!
0'
#83950000000
1!
1$
b1 %
1'
1*
b1 +
#83960000000
0!
0'
#83970000000
1!
b10 %
1'
b10 +
#83980000000
0!
0'
#83990000000
1!
b11 %
1'
b11 +
#84000000000
0!
0'
#84010000000
1!
b100 %
1'
b100 +
#84020000000
0!
0'
#84030000000
1!
b101 %
1'
b101 +
#84040000000
0!
0'
#84050000000
1!
0$
b110 %
1'
0*
b110 +
#84060000000
1"
1(
#84070000000
0!
0"
b100 &
0'
0(
b100 ,
#84080000000
1!
1$
b111 %
1'
1*
b111 +
#84090000000
0!
0'
#84100000000
1!
0$
b1000 %
1'
0*
b1000 +
#84110000000
0!
0'
#84120000000
1!
b1001 %
1'
b1001 +
#84130000000
0!
0'
#84140000000
1!
b0 %
1'
b0 +
#84150000000
0!
0'
#84160000000
1!
1$
b1 %
1'
1*
b1 +
#84170000000
0!
0'
#84180000000
1!
b10 %
1'
b10 +
#84190000000
0!
0'
#84200000000
1!
b11 %
1'
b11 +
#84210000000
0!
0'
#84220000000
1!
b100 %
1'
b100 +
#84230000000
0!
0'
#84240000000
1!
b101 %
1'
b101 +
#84250000000
0!
0'
#84260000000
1!
b110 %
1'
b110 +
#84270000000
0!
0'
#84280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#84290000000
0!
0'
#84300000000
1!
b1000 %
1'
b1000 +
#84310000000
0!
0'
#84320000000
1!
b1001 %
1'
b1001 +
#84330000000
0!
0'
#84340000000
1!
b0 %
1'
b0 +
#84350000000
0!
0'
#84360000000
1!
1$
b1 %
1'
1*
b1 +
#84370000000
0!
0'
#84380000000
1!
b10 %
1'
b10 +
#84390000000
0!
0'
#84400000000
1!
b11 %
1'
b11 +
#84410000000
0!
0'
#84420000000
1!
b100 %
1'
b100 +
#84430000000
0!
0'
#84440000000
1!
b101 %
1'
b101 +
#84450000000
0!
0'
#84460000000
1!
0$
b110 %
1'
0*
b110 +
#84470000000
0!
0'
#84480000000
1!
b111 %
1'
b111 +
#84490000000
1"
1(
#84500000000
0!
0"
b100 &
0'
0(
b100 ,
#84510000000
1!
b1000 %
1'
b1000 +
#84520000000
0!
0'
#84530000000
1!
b1001 %
1'
b1001 +
#84540000000
0!
0'
#84550000000
1!
b0 %
1'
b0 +
#84560000000
0!
0'
#84570000000
1!
1$
b1 %
1'
1*
b1 +
#84580000000
0!
0'
#84590000000
1!
b10 %
1'
b10 +
#84600000000
0!
0'
#84610000000
1!
b11 %
1'
b11 +
#84620000000
0!
0'
#84630000000
1!
b100 %
1'
b100 +
#84640000000
0!
0'
#84650000000
1!
b101 %
1'
b101 +
#84660000000
0!
0'
#84670000000
1!
b110 %
1'
b110 +
#84680000000
0!
0'
#84690000000
1!
b111 %
1'
b111 +
#84700000000
0!
0'
#84710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#84720000000
0!
0'
#84730000000
1!
b1001 %
1'
b1001 +
#84740000000
0!
0'
#84750000000
1!
b0 %
1'
b0 +
#84760000000
0!
0'
#84770000000
1!
1$
b1 %
1'
1*
b1 +
#84780000000
0!
0'
#84790000000
1!
b10 %
1'
b10 +
#84800000000
0!
0'
#84810000000
1!
b11 %
1'
b11 +
#84820000000
0!
0'
#84830000000
1!
b100 %
1'
b100 +
#84840000000
0!
0'
#84850000000
1!
b101 %
1'
b101 +
#84860000000
0!
0'
#84870000000
1!
0$
b110 %
1'
0*
b110 +
#84880000000
0!
0'
#84890000000
1!
b111 %
1'
b111 +
#84900000000
0!
0'
#84910000000
1!
b1000 %
1'
b1000 +
#84920000000
1"
1(
#84930000000
0!
0"
b100 &
0'
0(
b100 ,
#84940000000
1!
b1001 %
1'
b1001 +
#84950000000
0!
0'
#84960000000
1!
b0 %
1'
b0 +
#84970000000
0!
0'
#84980000000
1!
1$
b1 %
1'
1*
b1 +
#84990000000
0!
0'
#85000000000
1!
b10 %
1'
b10 +
#85010000000
0!
0'
#85020000000
1!
b11 %
1'
b11 +
#85030000000
0!
0'
#85040000000
1!
b100 %
1'
b100 +
#85050000000
0!
0'
#85060000000
1!
b101 %
1'
b101 +
#85070000000
0!
0'
#85080000000
1!
b110 %
1'
b110 +
#85090000000
0!
0'
#85100000000
1!
b111 %
1'
b111 +
#85110000000
0!
0'
#85120000000
1!
0$
b1000 %
1'
0*
b1000 +
#85130000000
0!
0'
#85140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#85150000000
0!
0'
#85160000000
1!
b0 %
1'
b0 +
#85170000000
0!
0'
#85180000000
1!
1$
b1 %
1'
1*
b1 +
#85190000000
0!
0'
#85200000000
1!
b10 %
1'
b10 +
#85210000000
0!
0'
#85220000000
1!
b11 %
1'
b11 +
#85230000000
0!
0'
#85240000000
1!
b100 %
1'
b100 +
#85250000000
0!
0'
#85260000000
1!
b101 %
1'
b101 +
#85270000000
0!
0'
#85280000000
1!
0$
b110 %
1'
0*
b110 +
#85290000000
0!
0'
#85300000000
1!
b111 %
1'
b111 +
#85310000000
0!
0'
#85320000000
1!
b1000 %
1'
b1000 +
#85330000000
0!
0'
#85340000000
1!
b1001 %
1'
b1001 +
#85350000000
1"
1(
#85360000000
0!
0"
b100 &
0'
0(
b100 ,
#85370000000
1!
b0 %
1'
b0 +
#85380000000
0!
0'
#85390000000
1!
1$
b1 %
1'
1*
b1 +
#85400000000
0!
0'
#85410000000
1!
b10 %
1'
b10 +
#85420000000
0!
0'
#85430000000
1!
b11 %
1'
b11 +
#85440000000
0!
0'
#85450000000
1!
b100 %
1'
b100 +
#85460000000
0!
0'
#85470000000
1!
b101 %
1'
b101 +
#85480000000
0!
0'
#85490000000
1!
b110 %
1'
b110 +
#85500000000
0!
0'
#85510000000
1!
b111 %
1'
b111 +
#85520000000
0!
0'
#85530000000
1!
0$
b1000 %
1'
0*
b1000 +
#85540000000
0!
0'
#85550000000
1!
b1001 %
1'
b1001 +
#85560000000
0!
0'
#85570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#85580000000
0!
0'
#85590000000
1!
1$
b1 %
1'
1*
b1 +
#85600000000
0!
0'
#85610000000
1!
b10 %
1'
b10 +
#85620000000
0!
0'
#85630000000
1!
b11 %
1'
b11 +
#85640000000
0!
0'
#85650000000
1!
b100 %
1'
b100 +
#85660000000
0!
0'
#85670000000
1!
b101 %
1'
b101 +
#85680000000
0!
0'
#85690000000
1!
0$
b110 %
1'
0*
b110 +
#85700000000
0!
0'
#85710000000
1!
b111 %
1'
b111 +
#85720000000
0!
0'
#85730000000
1!
b1000 %
1'
b1000 +
#85740000000
0!
0'
#85750000000
1!
b1001 %
1'
b1001 +
#85760000000
0!
0'
#85770000000
1!
b0 %
1'
b0 +
#85780000000
1"
1(
#85790000000
0!
0"
b100 &
0'
0(
b100 ,
#85800000000
1!
1$
b1 %
1'
1*
b1 +
#85810000000
0!
0'
#85820000000
1!
b10 %
1'
b10 +
#85830000000
0!
0'
#85840000000
1!
b11 %
1'
b11 +
#85850000000
0!
0'
#85860000000
1!
b100 %
1'
b100 +
#85870000000
0!
0'
#85880000000
1!
b101 %
1'
b101 +
#85890000000
0!
0'
#85900000000
1!
b110 %
1'
b110 +
#85910000000
0!
0'
#85920000000
1!
b111 %
1'
b111 +
#85930000000
0!
0'
#85940000000
1!
0$
b1000 %
1'
0*
b1000 +
#85950000000
0!
0'
#85960000000
1!
b1001 %
1'
b1001 +
#85970000000
0!
0'
#85980000000
1!
b0 %
1'
b0 +
#85990000000
0!
0'
#86000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#86010000000
0!
0'
#86020000000
1!
b10 %
1'
b10 +
#86030000000
0!
0'
#86040000000
1!
b11 %
1'
b11 +
#86050000000
0!
0'
#86060000000
1!
b100 %
1'
b100 +
#86070000000
0!
0'
#86080000000
1!
b101 %
1'
b101 +
#86090000000
0!
0'
#86100000000
1!
0$
b110 %
1'
0*
b110 +
#86110000000
0!
0'
#86120000000
1!
b111 %
1'
b111 +
#86130000000
0!
0'
#86140000000
1!
b1000 %
1'
b1000 +
#86150000000
0!
0'
#86160000000
1!
b1001 %
1'
b1001 +
#86170000000
0!
0'
#86180000000
1!
b0 %
1'
b0 +
#86190000000
0!
0'
#86200000000
1!
1$
b1 %
1'
1*
b1 +
#86210000000
1"
1(
#86220000000
0!
0"
b100 &
0'
0(
b100 ,
#86230000000
1!
b10 %
1'
b10 +
#86240000000
0!
0'
#86250000000
1!
b11 %
1'
b11 +
#86260000000
0!
0'
#86270000000
1!
b100 %
1'
b100 +
#86280000000
0!
0'
#86290000000
1!
b101 %
1'
b101 +
#86300000000
0!
0'
#86310000000
1!
b110 %
1'
b110 +
#86320000000
0!
0'
#86330000000
1!
b111 %
1'
b111 +
#86340000000
0!
0'
#86350000000
1!
0$
b1000 %
1'
0*
b1000 +
#86360000000
0!
0'
#86370000000
1!
b1001 %
1'
b1001 +
#86380000000
0!
0'
#86390000000
1!
b0 %
1'
b0 +
#86400000000
0!
0'
#86410000000
1!
1$
b1 %
1'
1*
b1 +
#86420000000
0!
0'
#86430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#86440000000
0!
0'
#86450000000
1!
b11 %
1'
b11 +
#86460000000
0!
0'
#86470000000
1!
b100 %
1'
b100 +
#86480000000
0!
0'
#86490000000
1!
b101 %
1'
b101 +
#86500000000
0!
0'
#86510000000
1!
0$
b110 %
1'
0*
b110 +
#86520000000
0!
0'
#86530000000
1!
b111 %
1'
b111 +
#86540000000
0!
0'
#86550000000
1!
b1000 %
1'
b1000 +
#86560000000
0!
0'
#86570000000
1!
b1001 %
1'
b1001 +
#86580000000
0!
0'
#86590000000
1!
b0 %
1'
b0 +
#86600000000
0!
0'
#86610000000
1!
1$
b1 %
1'
1*
b1 +
#86620000000
0!
0'
#86630000000
1!
b10 %
1'
b10 +
#86640000000
1"
1(
#86650000000
0!
0"
b100 &
0'
0(
b100 ,
#86660000000
1!
b11 %
1'
b11 +
#86670000000
0!
0'
#86680000000
1!
b100 %
1'
b100 +
#86690000000
0!
0'
#86700000000
1!
b101 %
1'
b101 +
#86710000000
0!
0'
#86720000000
1!
b110 %
1'
b110 +
#86730000000
0!
0'
#86740000000
1!
b111 %
1'
b111 +
#86750000000
0!
0'
#86760000000
1!
0$
b1000 %
1'
0*
b1000 +
#86770000000
0!
0'
#86780000000
1!
b1001 %
1'
b1001 +
#86790000000
0!
0'
#86800000000
1!
b0 %
1'
b0 +
#86810000000
0!
0'
#86820000000
1!
1$
b1 %
1'
1*
b1 +
#86830000000
0!
0'
#86840000000
1!
b10 %
1'
b10 +
#86850000000
0!
0'
#86860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#86870000000
0!
0'
#86880000000
1!
b100 %
1'
b100 +
#86890000000
0!
0'
#86900000000
1!
b101 %
1'
b101 +
#86910000000
0!
0'
#86920000000
1!
0$
b110 %
1'
0*
b110 +
#86930000000
0!
0'
#86940000000
1!
b111 %
1'
b111 +
#86950000000
0!
0'
#86960000000
1!
b1000 %
1'
b1000 +
#86970000000
0!
0'
#86980000000
1!
b1001 %
1'
b1001 +
#86990000000
0!
0'
#87000000000
1!
b0 %
1'
b0 +
#87010000000
0!
0'
#87020000000
1!
1$
b1 %
1'
1*
b1 +
#87030000000
0!
0'
#87040000000
1!
b10 %
1'
b10 +
#87050000000
0!
0'
#87060000000
1!
b11 %
1'
b11 +
#87070000000
1"
1(
#87080000000
0!
0"
b100 &
0'
0(
b100 ,
#87090000000
1!
b100 %
1'
b100 +
#87100000000
0!
0'
#87110000000
1!
b101 %
1'
b101 +
#87120000000
0!
0'
#87130000000
1!
b110 %
1'
b110 +
#87140000000
0!
0'
#87150000000
1!
b111 %
1'
b111 +
#87160000000
0!
0'
#87170000000
1!
0$
b1000 %
1'
0*
b1000 +
#87180000000
0!
0'
#87190000000
1!
b1001 %
1'
b1001 +
#87200000000
0!
0'
#87210000000
1!
b0 %
1'
b0 +
#87220000000
0!
0'
#87230000000
1!
1$
b1 %
1'
1*
b1 +
#87240000000
0!
0'
#87250000000
1!
b10 %
1'
b10 +
#87260000000
0!
0'
#87270000000
1!
b11 %
1'
b11 +
#87280000000
0!
0'
#87290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#87300000000
0!
0'
#87310000000
1!
b101 %
1'
b101 +
#87320000000
0!
0'
#87330000000
1!
0$
b110 %
1'
0*
b110 +
#87340000000
0!
0'
#87350000000
1!
b111 %
1'
b111 +
#87360000000
0!
0'
#87370000000
1!
b1000 %
1'
b1000 +
#87380000000
0!
0'
#87390000000
1!
b1001 %
1'
b1001 +
#87400000000
0!
0'
#87410000000
1!
b0 %
1'
b0 +
#87420000000
0!
0'
#87430000000
1!
1$
b1 %
1'
1*
b1 +
#87440000000
0!
0'
#87450000000
1!
b10 %
1'
b10 +
#87460000000
0!
0'
#87470000000
1!
b11 %
1'
b11 +
#87480000000
0!
0'
#87490000000
1!
b100 %
1'
b100 +
#87500000000
1"
1(
#87510000000
0!
0"
b100 &
0'
0(
b100 ,
#87520000000
1!
b101 %
1'
b101 +
#87530000000
0!
0'
#87540000000
1!
b110 %
1'
b110 +
#87550000000
0!
0'
#87560000000
1!
b111 %
1'
b111 +
#87570000000
0!
0'
#87580000000
1!
0$
b1000 %
1'
0*
b1000 +
#87590000000
0!
0'
#87600000000
1!
b1001 %
1'
b1001 +
#87610000000
0!
0'
#87620000000
1!
b0 %
1'
b0 +
#87630000000
0!
0'
#87640000000
1!
1$
b1 %
1'
1*
b1 +
#87650000000
0!
0'
#87660000000
1!
b10 %
1'
b10 +
#87670000000
0!
0'
#87680000000
1!
b11 %
1'
b11 +
#87690000000
0!
0'
#87700000000
1!
b100 %
1'
b100 +
#87710000000
0!
0'
#87720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#87730000000
0!
0'
#87740000000
1!
0$
b110 %
1'
0*
b110 +
#87750000000
0!
0'
#87760000000
1!
b111 %
1'
b111 +
#87770000000
0!
0'
#87780000000
1!
b1000 %
1'
b1000 +
#87790000000
0!
0'
#87800000000
1!
b1001 %
1'
b1001 +
#87810000000
0!
0'
#87820000000
1!
b0 %
1'
b0 +
#87830000000
0!
0'
#87840000000
1!
1$
b1 %
1'
1*
b1 +
#87850000000
0!
0'
#87860000000
1!
b10 %
1'
b10 +
#87870000000
0!
0'
#87880000000
1!
b11 %
1'
b11 +
#87890000000
0!
0'
#87900000000
1!
b100 %
1'
b100 +
#87910000000
0!
0'
#87920000000
1!
b101 %
1'
b101 +
#87930000000
1"
1(
#87940000000
0!
0"
b100 &
0'
0(
b100 ,
#87950000000
1!
b110 %
1'
b110 +
#87960000000
0!
0'
#87970000000
1!
b111 %
1'
b111 +
#87980000000
0!
0'
#87990000000
1!
0$
b1000 %
1'
0*
b1000 +
#88000000000
0!
0'
#88010000000
1!
b1001 %
1'
b1001 +
#88020000000
0!
0'
#88030000000
1!
b0 %
1'
b0 +
#88040000000
0!
0'
#88050000000
1!
1$
b1 %
1'
1*
b1 +
#88060000000
0!
0'
#88070000000
1!
b10 %
1'
b10 +
#88080000000
0!
0'
#88090000000
1!
b11 %
1'
b11 +
#88100000000
0!
0'
#88110000000
1!
b100 %
1'
b100 +
#88120000000
0!
0'
#88130000000
1!
b101 %
1'
b101 +
#88140000000
0!
0'
#88150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#88160000000
0!
0'
#88170000000
1!
b111 %
1'
b111 +
#88180000000
0!
0'
#88190000000
1!
b1000 %
1'
b1000 +
#88200000000
0!
0'
#88210000000
1!
b1001 %
1'
b1001 +
#88220000000
0!
0'
#88230000000
1!
b0 %
1'
b0 +
#88240000000
0!
0'
#88250000000
1!
1$
b1 %
1'
1*
b1 +
#88260000000
0!
0'
#88270000000
1!
b10 %
1'
b10 +
#88280000000
0!
0'
#88290000000
1!
b11 %
1'
b11 +
#88300000000
0!
0'
#88310000000
1!
b100 %
1'
b100 +
#88320000000
0!
0'
#88330000000
1!
b101 %
1'
b101 +
#88340000000
0!
0'
#88350000000
1!
0$
b110 %
1'
0*
b110 +
#88360000000
1"
1(
#88370000000
0!
0"
b100 &
0'
0(
b100 ,
#88380000000
1!
1$
b111 %
1'
1*
b111 +
#88390000000
0!
0'
#88400000000
1!
0$
b1000 %
1'
0*
b1000 +
#88410000000
0!
0'
#88420000000
1!
b1001 %
1'
b1001 +
#88430000000
0!
0'
#88440000000
1!
b0 %
1'
b0 +
#88450000000
0!
0'
#88460000000
1!
1$
b1 %
1'
1*
b1 +
#88470000000
0!
0'
#88480000000
1!
b10 %
1'
b10 +
#88490000000
0!
0'
#88500000000
1!
b11 %
1'
b11 +
#88510000000
0!
0'
#88520000000
1!
b100 %
1'
b100 +
#88530000000
0!
0'
#88540000000
1!
b101 %
1'
b101 +
#88550000000
0!
0'
#88560000000
1!
b110 %
1'
b110 +
#88570000000
0!
0'
#88580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#88590000000
0!
0'
#88600000000
1!
b1000 %
1'
b1000 +
#88610000000
0!
0'
#88620000000
1!
b1001 %
1'
b1001 +
#88630000000
0!
0'
#88640000000
1!
b0 %
1'
b0 +
#88650000000
0!
0'
#88660000000
1!
1$
b1 %
1'
1*
b1 +
#88670000000
0!
0'
#88680000000
1!
b10 %
1'
b10 +
#88690000000
0!
0'
#88700000000
1!
b11 %
1'
b11 +
#88710000000
0!
0'
#88720000000
1!
b100 %
1'
b100 +
#88730000000
0!
0'
#88740000000
1!
b101 %
1'
b101 +
#88750000000
0!
0'
#88760000000
1!
0$
b110 %
1'
0*
b110 +
#88770000000
0!
0'
#88780000000
1!
b111 %
1'
b111 +
#88790000000
1"
1(
#88800000000
0!
0"
b100 &
0'
0(
b100 ,
#88810000000
1!
b1000 %
1'
b1000 +
#88820000000
0!
0'
#88830000000
1!
b1001 %
1'
b1001 +
#88840000000
0!
0'
#88850000000
1!
b0 %
1'
b0 +
#88860000000
0!
0'
#88870000000
1!
1$
b1 %
1'
1*
b1 +
#88880000000
0!
0'
#88890000000
1!
b10 %
1'
b10 +
#88900000000
0!
0'
#88910000000
1!
b11 %
1'
b11 +
#88920000000
0!
0'
#88930000000
1!
b100 %
1'
b100 +
#88940000000
0!
0'
#88950000000
1!
b101 %
1'
b101 +
#88960000000
0!
0'
#88970000000
1!
b110 %
1'
b110 +
#88980000000
0!
0'
#88990000000
1!
b111 %
1'
b111 +
#89000000000
0!
0'
#89010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#89020000000
0!
0'
#89030000000
1!
b1001 %
1'
b1001 +
#89040000000
0!
0'
#89050000000
1!
b0 %
1'
b0 +
#89060000000
0!
0'
#89070000000
1!
1$
b1 %
1'
1*
b1 +
#89080000000
0!
0'
#89090000000
1!
b10 %
1'
b10 +
#89100000000
0!
0'
#89110000000
1!
b11 %
1'
b11 +
#89120000000
0!
0'
#89130000000
1!
b100 %
1'
b100 +
#89140000000
0!
0'
#89150000000
1!
b101 %
1'
b101 +
#89160000000
0!
0'
#89170000000
1!
0$
b110 %
1'
0*
b110 +
#89180000000
0!
0'
#89190000000
1!
b111 %
1'
b111 +
#89200000000
0!
0'
#89210000000
1!
b1000 %
1'
b1000 +
#89220000000
1"
1(
#89230000000
0!
0"
b100 &
0'
0(
b100 ,
#89240000000
1!
b1001 %
1'
b1001 +
#89250000000
0!
0'
#89260000000
1!
b0 %
1'
b0 +
#89270000000
0!
0'
#89280000000
1!
1$
b1 %
1'
1*
b1 +
#89290000000
0!
0'
#89300000000
1!
b10 %
1'
b10 +
#89310000000
0!
0'
#89320000000
1!
b11 %
1'
b11 +
#89330000000
0!
0'
#89340000000
1!
b100 %
1'
b100 +
#89350000000
0!
0'
#89360000000
1!
b101 %
1'
b101 +
#89370000000
0!
0'
#89380000000
1!
b110 %
1'
b110 +
#89390000000
0!
0'
#89400000000
1!
b111 %
1'
b111 +
#89410000000
0!
0'
#89420000000
1!
0$
b1000 %
1'
0*
b1000 +
#89430000000
0!
0'
#89440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#89450000000
0!
0'
#89460000000
1!
b0 %
1'
b0 +
#89470000000
0!
0'
#89480000000
1!
1$
b1 %
1'
1*
b1 +
#89490000000
0!
0'
#89500000000
1!
b10 %
1'
b10 +
#89510000000
0!
0'
#89520000000
1!
b11 %
1'
b11 +
#89530000000
0!
0'
#89540000000
1!
b100 %
1'
b100 +
#89550000000
0!
0'
#89560000000
1!
b101 %
1'
b101 +
#89570000000
0!
0'
#89580000000
1!
0$
b110 %
1'
0*
b110 +
#89590000000
0!
0'
#89600000000
1!
b111 %
1'
b111 +
#89610000000
0!
0'
#89620000000
1!
b1000 %
1'
b1000 +
#89630000000
0!
0'
#89640000000
1!
b1001 %
1'
b1001 +
#89650000000
1"
1(
#89660000000
0!
0"
b100 &
0'
0(
b100 ,
#89670000000
1!
b0 %
1'
b0 +
#89680000000
0!
0'
#89690000000
1!
1$
b1 %
1'
1*
b1 +
#89700000000
0!
0'
#89710000000
1!
b10 %
1'
b10 +
#89720000000
0!
0'
#89730000000
1!
b11 %
1'
b11 +
#89740000000
0!
0'
#89750000000
1!
b100 %
1'
b100 +
#89760000000
0!
0'
#89770000000
1!
b101 %
1'
b101 +
#89780000000
0!
0'
#89790000000
1!
b110 %
1'
b110 +
#89800000000
0!
0'
#89810000000
1!
b111 %
1'
b111 +
#89820000000
0!
0'
#89830000000
1!
0$
b1000 %
1'
0*
b1000 +
#89840000000
0!
0'
#89850000000
1!
b1001 %
1'
b1001 +
#89860000000
0!
0'
#89870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#89880000000
0!
0'
#89890000000
1!
1$
b1 %
1'
1*
b1 +
#89900000000
0!
0'
#89910000000
1!
b10 %
1'
b10 +
#89920000000
0!
0'
#89930000000
1!
b11 %
1'
b11 +
#89940000000
0!
0'
#89950000000
1!
b100 %
1'
b100 +
#89960000000
0!
0'
#89970000000
1!
b101 %
1'
b101 +
#89980000000
0!
0'
#89990000000
1!
0$
b110 %
1'
0*
b110 +
#90000000000
0!
0'
#90010000000
1!
b111 %
1'
b111 +
#90020000000
0!
0'
#90030000000
1!
b1000 %
1'
b1000 +
#90040000000
0!
0'
#90050000000
1!
b1001 %
1'
b1001 +
#90060000000
0!
0'
#90070000000
1!
b0 %
1'
b0 +
#90080000000
1"
1(
#90090000000
0!
0"
b100 &
0'
0(
b100 ,
#90100000000
1!
1$
b1 %
1'
1*
b1 +
#90110000000
0!
0'
#90120000000
1!
b10 %
1'
b10 +
#90130000000
0!
0'
#90140000000
1!
b11 %
1'
b11 +
#90150000000
0!
0'
#90160000000
1!
b100 %
1'
b100 +
#90170000000
0!
0'
#90180000000
1!
b101 %
1'
b101 +
#90190000000
0!
0'
#90200000000
1!
b110 %
1'
b110 +
#90210000000
0!
0'
#90220000000
1!
b111 %
1'
b111 +
#90230000000
0!
0'
#90240000000
1!
0$
b1000 %
1'
0*
b1000 +
#90250000000
0!
0'
#90260000000
1!
b1001 %
1'
b1001 +
#90270000000
0!
0'
#90280000000
1!
b0 %
1'
b0 +
#90290000000
0!
0'
#90300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#90310000000
0!
0'
#90320000000
1!
b10 %
1'
b10 +
#90330000000
0!
0'
#90340000000
1!
b11 %
1'
b11 +
#90350000000
0!
0'
#90360000000
1!
b100 %
1'
b100 +
#90370000000
0!
0'
#90380000000
1!
b101 %
1'
b101 +
#90390000000
0!
0'
#90400000000
1!
0$
b110 %
1'
0*
b110 +
#90410000000
0!
0'
#90420000000
1!
b111 %
1'
b111 +
#90430000000
0!
0'
#90440000000
1!
b1000 %
1'
b1000 +
#90450000000
0!
0'
#90460000000
1!
b1001 %
1'
b1001 +
#90470000000
0!
0'
#90480000000
1!
b0 %
1'
b0 +
#90490000000
0!
0'
#90500000000
1!
1$
b1 %
1'
1*
b1 +
#90510000000
1"
1(
#90520000000
0!
0"
b100 &
0'
0(
b100 ,
#90530000000
1!
b10 %
1'
b10 +
#90540000000
0!
0'
#90550000000
1!
b11 %
1'
b11 +
#90560000000
0!
0'
#90570000000
1!
b100 %
1'
b100 +
#90580000000
0!
0'
#90590000000
1!
b101 %
1'
b101 +
#90600000000
0!
0'
#90610000000
1!
b110 %
1'
b110 +
#90620000000
0!
0'
#90630000000
1!
b111 %
1'
b111 +
#90640000000
0!
0'
#90650000000
1!
0$
b1000 %
1'
0*
b1000 +
#90660000000
0!
0'
#90670000000
1!
b1001 %
1'
b1001 +
#90680000000
0!
0'
#90690000000
1!
b0 %
1'
b0 +
#90700000000
0!
0'
#90710000000
1!
1$
b1 %
1'
1*
b1 +
#90720000000
0!
0'
#90730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#90740000000
0!
0'
#90750000000
1!
b11 %
1'
b11 +
#90760000000
0!
0'
#90770000000
1!
b100 %
1'
b100 +
#90780000000
0!
0'
#90790000000
1!
b101 %
1'
b101 +
#90800000000
0!
0'
#90810000000
1!
0$
b110 %
1'
0*
b110 +
#90820000000
0!
0'
#90830000000
1!
b111 %
1'
b111 +
#90840000000
0!
0'
#90850000000
1!
b1000 %
1'
b1000 +
#90860000000
0!
0'
#90870000000
1!
b1001 %
1'
b1001 +
#90880000000
0!
0'
#90890000000
1!
b0 %
1'
b0 +
#90900000000
0!
0'
#90910000000
1!
1$
b1 %
1'
1*
b1 +
#90920000000
0!
0'
#90930000000
1!
b10 %
1'
b10 +
#90940000000
1"
1(
#90950000000
0!
0"
b100 &
0'
0(
b100 ,
#90960000000
1!
b11 %
1'
b11 +
#90970000000
0!
0'
#90980000000
1!
b100 %
1'
b100 +
#90990000000
0!
0'
#91000000000
1!
b101 %
1'
b101 +
#91010000000
0!
0'
#91020000000
1!
b110 %
1'
b110 +
#91030000000
0!
0'
#91040000000
1!
b111 %
1'
b111 +
#91050000000
0!
0'
#91060000000
1!
0$
b1000 %
1'
0*
b1000 +
#91070000000
0!
0'
#91080000000
1!
b1001 %
1'
b1001 +
#91090000000
0!
0'
#91100000000
1!
b0 %
1'
b0 +
#91110000000
0!
0'
#91120000000
1!
1$
b1 %
1'
1*
b1 +
#91130000000
0!
0'
#91140000000
1!
b10 %
1'
b10 +
#91150000000
0!
0'
#91160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#91170000000
0!
0'
#91180000000
1!
b100 %
1'
b100 +
#91190000000
0!
0'
#91200000000
1!
b101 %
1'
b101 +
#91210000000
0!
0'
#91220000000
1!
0$
b110 %
1'
0*
b110 +
#91230000000
0!
0'
#91240000000
1!
b111 %
1'
b111 +
#91250000000
0!
0'
#91260000000
1!
b1000 %
1'
b1000 +
#91270000000
0!
0'
#91280000000
1!
b1001 %
1'
b1001 +
#91290000000
0!
0'
#91300000000
1!
b0 %
1'
b0 +
#91310000000
0!
0'
#91320000000
1!
1$
b1 %
1'
1*
b1 +
#91330000000
0!
0'
#91340000000
1!
b10 %
1'
b10 +
#91350000000
0!
0'
#91360000000
1!
b11 %
1'
b11 +
#91370000000
1"
1(
#91380000000
0!
0"
b100 &
0'
0(
b100 ,
#91390000000
1!
b100 %
1'
b100 +
#91400000000
0!
0'
#91410000000
1!
b101 %
1'
b101 +
#91420000000
0!
0'
#91430000000
1!
b110 %
1'
b110 +
#91440000000
0!
0'
#91450000000
1!
b111 %
1'
b111 +
#91460000000
0!
0'
#91470000000
1!
0$
b1000 %
1'
0*
b1000 +
#91480000000
0!
0'
#91490000000
1!
b1001 %
1'
b1001 +
#91500000000
0!
0'
#91510000000
1!
b0 %
1'
b0 +
#91520000000
0!
0'
#91530000000
1!
1$
b1 %
1'
1*
b1 +
#91540000000
0!
0'
#91550000000
1!
b10 %
1'
b10 +
#91560000000
0!
0'
#91570000000
1!
b11 %
1'
b11 +
#91580000000
0!
0'
#91590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#91600000000
0!
0'
#91610000000
1!
b101 %
1'
b101 +
#91620000000
0!
0'
#91630000000
1!
0$
b110 %
1'
0*
b110 +
#91640000000
0!
0'
#91650000000
1!
b111 %
1'
b111 +
#91660000000
0!
0'
#91670000000
1!
b1000 %
1'
b1000 +
#91680000000
0!
0'
#91690000000
1!
b1001 %
1'
b1001 +
#91700000000
0!
0'
#91710000000
1!
b0 %
1'
b0 +
#91720000000
0!
0'
#91730000000
1!
1$
b1 %
1'
1*
b1 +
#91740000000
0!
0'
#91750000000
1!
b10 %
1'
b10 +
#91760000000
0!
0'
#91770000000
1!
b11 %
1'
b11 +
#91780000000
0!
0'
#91790000000
1!
b100 %
1'
b100 +
#91800000000
1"
1(
#91810000000
0!
0"
b100 &
0'
0(
b100 ,
#91820000000
1!
b101 %
1'
b101 +
#91830000000
0!
0'
#91840000000
1!
b110 %
1'
b110 +
#91850000000
0!
0'
#91860000000
1!
b111 %
1'
b111 +
#91870000000
0!
0'
#91880000000
1!
0$
b1000 %
1'
0*
b1000 +
#91890000000
0!
0'
#91900000000
1!
b1001 %
1'
b1001 +
#91910000000
0!
0'
#91920000000
1!
b0 %
1'
b0 +
#91930000000
0!
0'
#91940000000
1!
1$
b1 %
1'
1*
b1 +
#91950000000
0!
0'
#91960000000
1!
b10 %
1'
b10 +
#91970000000
0!
0'
#91980000000
1!
b11 %
1'
b11 +
#91990000000
0!
0'
#92000000000
1!
b100 %
1'
b100 +
#92010000000
0!
0'
#92020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#92030000000
0!
0'
#92040000000
1!
0$
b110 %
1'
0*
b110 +
#92050000000
0!
0'
#92060000000
1!
b111 %
1'
b111 +
#92070000000
0!
0'
#92080000000
1!
b1000 %
1'
b1000 +
#92090000000
0!
0'
#92100000000
1!
b1001 %
1'
b1001 +
#92110000000
0!
0'
#92120000000
1!
b0 %
1'
b0 +
#92130000000
0!
0'
#92140000000
1!
1$
b1 %
1'
1*
b1 +
#92150000000
0!
0'
#92160000000
1!
b10 %
1'
b10 +
#92170000000
0!
0'
#92180000000
1!
b11 %
1'
b11 +
#92190000000
0!
0'
#92200000000
1!
b100 %
1'
b100 +
#92210000000
0!
0'
#92220000000
1!
b101 %
1'
b101 +
#92230000000
1"
1(
#92240000000
0!
0"
b100 &
0'
0(
b100 ,
#92250000000
1!
b110 %
1'
b110 +
#92260000000
0!
0'
#92270000000
1!
b111 %
1'
b111 +
#92280000000
0!
0'
#92290000000
1!
0$
b1000 %
1'
0*
b1000 +
#92300000000
0!
0'
#92310000000
1!
b1001 %
1'
b1001 +
#92320000000
0!
0'
#92330000000
1!
b0 %
1'
b0 +
#92340000000
0!
0'
#92350000000
1!
1$
b1 %
1'
1*
b1 +
#92360000000
0!
0'
#92370000000
1!
b10 %
1'
b10 +
#92380000000
0!
0'
#92390000000
1!
b11 %
1'
b11 +
#92400000000
0!
0'
#92410000000
1!
b100 %
1'
b100 +
#92420000000
0!
0'
#92430000000
1!
b101 %
1'
b101 +
#92440000000
0!
0'
#92450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#92460000000
0!
0'
#92470000000
1!
b111 %
1'
b111 +
#92480000000
0!
0'
#92490000000
1!
b1000 %
1'
b1000 +
#92500000000
0!
0'
#92510000000
1!
b1001 %
1'
b1001 +
#92520000000
0!
0'
#92530000000
1!
b0 %
1'
b0 +
#92540000000
0!
0'
#92550000000
1!
1$
b1 %
1'
1*
b1 +
#92560000000
0!
0'
#92570000000
1!
b10 %
1'
b10 +
#92580000000
0!
0'
#92590000000
1!
b11 %
1'
b11 +
#92600000000
0!
0'
#92610000000
1!
b100 %
1'
b100 +
#92620000000
0!
0'
#92630000000
1!
b101 %
1'
b101 +
#92640000000
0!
0'
#92650000000
1!
0$
b110 %
1'
0*
b110 +
#92660000000
1"
1(
#92670000000
0!
0"
b100 &
0'
0(
b100 ,
#92680000000
1!
1$
b111 %
1'
1*
b111 +
#92690000000
0!
0'
#92700000000
1!
0$
b1000 %
1'
0*
b1000 +
#92710000000
0!
0'
#92720000000
1!
b1001 %
1'
b1001 +
#92730000000
0!
0'
#92740000000
1!
b0 %
1'
b0 +
#92750000000
0!
0'
#92760000000
1!
1$
b1 %
1'
1*
b1 +
#92770000000
0!
0'
#92780000000
1!
b10 %
1'
b10 +
#92790000000
0!
0'
#92800000000
1!
b11 %
1'
b11 +
#92810000000
0!
0'
#92820000000
1!
b100 %
1'
b100 +
#92830000000
0!
0'
#92840000000
1!
b101 %
1'
b101 +
#92850000000
0!
0'
#92860000000
1!
b110 %
1'
b110 +
#92870000000
0!
0'
#92880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#92890000000
0!
0'
#92900000000
1!
b1000 %
1'
b1000 +
#92910000000
0!
0'
#92920000000
1!
b1001 %
1'
b1001 +
#92930000000
0!
0'
#92940000000
1!
b0 %
1'
b0 +
#92950000000
0!
0'
#92960000000
1!
1$
b1 %
1'
1*
b1 +
#92970000000
0!
0'
#92980000000
1!
b10 %
1'
b10 +
#92990000000
0!
0'
#93000000000
1!
b11 %
1'
b11 +
#93010000000
0!
0'
#93020000000
1!
b100 %
1'
b100 +
#93030000000
0!
0'
#93040000000
1!
b101 %
1'
b101 +
#93050000000
0!
0'
#93060000000
1!
0$
b110 %
1'
0*
b110 +
#93070000000
0!
0'
#93080000000
1!
b111 %
1'
b111 +
#93090000000
1"
1(
#93100000000
0!
0"
b100 &
0'
0(
b100 ,
#93110000000
1!
b1000 %
1'
b1000 +
#93120000000
0!
0'
#93130000000
1!
b1001 %
1'
b1001 +
#93140000000
0!
0'
#93150000000
1!
b0 %
1'
b0 +
#93160000000
0!
0'
#93170000000
1!
1$
b1 %
1'
1*
b1 +
#93180000000
0!
0'
#93190000000
1!
b10 %
1'
b10 +
#93200000000
0!
0'
#93210000000
1!
b11 %
1'
b11 +
#93220000000
0!
0'
#93230000000
1!
b100 %
1'
b100 +
#93240000000
0!
0'
#93250000000
1!
b101 %
1'
b101 +
#93260000000
0!
0'
#93270000000
1!
b110 %
1'
b110 +
#93280000000
0!
0'
#93290000000
1!
b111 %
1'
b111 +
#93300000000
0!
0'
#93310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#93320000000
0!
0'
#93330000000
1!
b1001 %
1'
b1001 +
#93340000000
0!
0'
#93350000000
1!
b0 %
1'
b0 +
#93360000000
0!
0'
#93370000000
1!
1$
b1 %
1'
1*
b1 +
#93380000000
0!
0'
#93390000000
1!
b10 %
1'
b10 +
#93400000000
0!
0'
#93410000000
1!
b11 %
1'
b11 +
#93420000000
0!
0'
#93430000000
1!
b100 %
1'
b100 +
#93440000000
0!
0'
#93450000000
1!
b101 %
1'
b101 +
#93460000000
0!
0'
#93470000000
1!
0$
b110 %
1'
0*
b110 +
#93480000000
0!
0'
#93490000000
1!
b111 %
1'
b111 +
#93500000000
0!
0'
#93510000000
1!
b1000 %
1'
b1000 +
#93520000000
1"
1(
#93530000000
0!
0"
b100 &
0'
0(
b100 ,
#93540000000
1!
b1001 %
1'
b1001 +
#93550000000
0!
0'
#93560000000
1!
b0 %
1'
b0 +
#93570000000
0!
0'
#93580000000
1!
1$
b1 %
1'
1*
b1 +
#93590000000
0!
0'
#93600000000
1!
b10 %
1'
b10 +
#93610000000
0!
0'
#93620000000
1!
b11 %
1'
b11 +
#93630000000
0!
0'
#93640000000
1!
b100 %
1'
b100 +
#93650000000
0!
0'
#93660000000
1!
b101 %
1'
b101 +
#93670000000
0!
0'
#93680000000
1!
b110 %
1'
b110 +
#93690000000
0!
0'
#93700000000
1!
b111 %
1'
b111 +
#93710000000
0!
0'
#93720000000
1!
0$
b1000 %
1'
0*
b1000 +
#93730000000
0!
0'
#93740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#93750000000
0!
0'
#93760000000
1!
b0 %
1'
b0 +
#93770000000
0!
0'
#93780000000
1!
1$
b1 %
1'
1*
b1 +
#93790000000
0!
0'
#93800000000
1!
b10 %
1'
b10 +
#93810000000
0!
0'
#93820000000
1!
b11 %
1'
b11 +
#93830000000
0!
0'
#93840000000
1!
b100 %
1'
b100 +
#93850000000
0!
0'
#93860000000
1!
b101 %
1'
b101 +
#93870000000
0!
0'
#93880000000
1!
0$
b110 %
1'
0*
b110 +
#93890000000
0!
0'
#93900000000
1!
b111 %
1'
b111 +
#93910000000
0!
0'
#93920000000
1!
b1000 %
1'
b1000 +
#93930000000
0!
0'
#93940000000
1!
b1001 %
1'
b1001 +
#93950000000
1"
1(
#93960000000
0!
0"
b100 &
0'
0(
b100 ,
#93970000000
1!
b0 %
1'
b0 +
#93980000000
0!
0'
#93990000000
1!
1$
b1 %
1'
1*
b1 +
#94000000000
0!
0'
#94010000000
1!
b10 %
1'
b10 +
#94020000000
0!
0'
#94030000000
1!
b11 %
1'
b11 +
#94040000000
0!
0'
#94050000000
1!
b100 %
1'
b100 +
#94060000000
0!
0'
#94070000000
1!
b101 %
1'
b101 +
#94080000000
0!
0'
#94090000000
1!
b110 %
1'
b110 +
#94100000000
0!
0'
#94110000000
1!
b111 %
1'
b111 +
#94120000000
0!
0'
#94130000000
1!
0$
b1000 %
1'
0*
b1000 +
#94140000000
0!
0'
#94150000000
1!
b1001 %
1'
b1001 +
#94160000000
0!
0'
#94170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#94180000000
0!
0'
#94190000000
1!
1$
b1 %
1'
1*
b1 +
#94200000000
0!
0'
#94210000000
1!
b10 %
1'
b10 +
#94220000000
0!
0'
#94230000000
1!
b11 %
1'
b11 +
#94240000000
0!
0'
#94250000000
1!
b100 %
1'
b100 +
#94260000000
0!
0'
#94270000000
1!
b101 %
1'
b101 +
#94280000000
0!
0'
#94290000000
1!
0$
b110 %
1'
0*
b110 +
#94300000000
0!
0'
#94310000000
1!
b111 %
1'
b111 +
#94320000000
0!
0'
#94330000000
1!
b1000 %
1'
b1000 +
#94340000000
0!
0'
#94350000000
1!
b1001 %
1'
b1001 +
#94360000000
0!
0'
#94370000000
1!
b0 %
1'
b0 +
#94380000000
1"
1(
#94390000000
0!
0"
b100 &
0'
0(
b100 ,
#94400000000
1!
1$
b1 %
1'
1*
b1 +
#94410000000
0!
0'
#94420000000
1!
b10 %
1'
b10 +
#94430000000
0!
0'
#94440000000
1!
b11 %
1'
b11 +
#94450000000
0!
0'
#94460000000
1!
b100 %
1'
b100 +
#94470000000
0!
0'
#94480000000
1!
b101 %
1'
b101 +
#94490000000
0!
0'
#94500000000
1!
b110 %
1'
b110 +
#94510000000
0!
0'
#94520000000
1!
b111 %
1'
b111 +
#94530000000
0!
0'
#94540000000
1!
0$
b1000 %
1'
0*
b1000 +
#94550000000
0!
0'
#94560000000
1!
b1001 %
1'
b1001 +
#94570000000
0!
0'
#94580000000
1!
b0 %
1'
b0 +
#94590000000
0!
0'
#94600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#94610000000
0!
0'
#94620000000
1!
b10 %
1'
b10 +
#94630000000
0!
0'
#94640000000
1!
b11 %
1'
b11 +
#94650000000
0!
0'
#94660000000
1!
b100 %
1'
b100 +
#94670000000
0!
0'
#94680000000
1!
b101 %
1'
b101 +
#94690000000
0!
0'
#94700000000
1!
0$
b110 %
1'
0*
b110 +
#94710000000
0!
0'
#94720000000
1!
b111 %
1'
b111 +
#94730000000
0!
0'
#94740000000
1!
b1000 %
1'
b1000 +
#94750000000
0!
0'
#94760000000
1!
b1001 %
1'
b1001 +
#94770000000
0!
0'
#94780000000
1!
b0 %
1'
b0 +
#94790000000
0!
0'
#94800000000
1!
1$
b1 %
1'
1*
b1 +
#94810000000
1"
1(
#94820000000
0!
0"
b100 &
0'
0(
b100 ,
#94830000000
1!
b10 %
1'
b10 +
#94840000000
0!
0'
#94850000000
1!
b11 %
1'
b11 +
#94860000000
0!
0'
#94870000000
1!
b100 %
1'
b100 +
#94880000000
0!
0'
#94890000000
1!
b101 %
1'
b101 +
#94900000000
0!
0'
#94910000000
1!
b110 %
1'
b110 +
#94920000000
0!
0'
#94930000000
1!
b111 %
1'
b111 +
#94940000000
0!
0'
#94950000000
1!
0$
b1000 %
1'
0*
b1000 +
#94960000000
0!
0'
#94970000000
1!
b1001 %
1'
b1001 +
#94980000000
0!
0'
#94990000000
1!
b0 %
1'
b0 +
#95000000000
0!
0'
#95010000000
1!
1$
b1 %
1'
1*
b1 +
#95020000000
0!
0'
#95030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#95040000000
0!
0'
#95050000000
1!
b11 %
1'
b11 +
#95060000000
0!
0'
#95070000000
1!
b100 %
1'
b100 +
#95080000000
0!
0'
#95090000000
1!
b101 %
1'
b101 +
#95100000000
0!
0'
#95110000000
1!
0$
b110 %
1'
0*
b110 +
#95120000000
0!
0'
#95130000000
1!
b111 %
1'
b111 +
#95140000000
0!
0'
#95150000000
1!
b1000 %
1'
b1000 +
#95160000000
0!
0'
#95170000000
1!
b1001 %
1'
b1001 +
#95180000000
0!
0'
#95190000000
1!
b0 %
1'
b0 +
#95200000000
0!
0'
#95210000000
1!
1$
b1 %
1'
1*
b1 +
#95220000000
0!
0'
#95230000000
1!
b10 %
1'
b10 +
#95240000000
1"
1(
#95250000000
0!
0"
b100 &
0'
0(
b100 ,
#95260000000
1!
b11 %
1'
b11 +
#95270000000
0!
0'
#95280000000
1!
b100 %
1'
b100 +
#95290000000
0!
0'
#95300000000
1!
b101 %
1'
b101 +
#95310000000
0!
0'
#95320000000
1!
b110 %
1'
b110 +
#95330000000
0!
0'
#95340000000
1!
b111 %
1'
b111 +
#95350000000
0!
0'
#95360000000
1!
0$
b1000 %
1'
0*
b1000 +
#95370000000
0!
0'
#95380000000
1!
b1001 %
1'
b1001 +
#95390000000
0!
0'
#95400000000
1!
b0 %
1'
b0 +
#95410000000
0!
0'
#95420000000
1!
1$
b1 %
1'
1*
b1 +
#95430000000
0!
0'
#95440000000
1!
b10 %
1'
b10 +
#95450000000
0!
0'
#95460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#95470000000
0!
0'
#95480000000
1!
b100 %
1'
b100 +
#95490000000
0!
0'
#95500000000
1!
b101 %
1'
b101 +
#95510000000
0!
0'
#95520000000
1!
0$
b110 %
1'
0*
b110 +
#95530000000
0!
0'
#95540000000
1!
b111 %
1'
b111 +
#95550000000
0!
0'
#95560000000
1!
b1000 %
1'
b1000 +
#95570000000
0!
0'
#95580000000
1!
b1001 %
1'
b1001 +
#95590000000
0!
0'
#95600000000
1!
b0 %
1'
b0 +
#95610000000
0!
0'
#95620000000
1!
1$
b1 %
1'
1*
b1 +
#95630000000
0!
0'
#95640000000
1!
b10 %
1'
b10 +
#95650000000
0!
0'
#95660000000
1!
b11 %
1'
b11 +
#95670000000
1"
1(
#95680000000
0!
0"
b100 &
0'
0(
b100 ,
#95690000000
1!
b100 %
1'
b100 +
#95700000000
0!
0'
#95710000000
1!
b101 %
1'
b101 +
#95720000000
0!
0'
#95730000000
1!
b110 %
1'
b110 +
#95740000000
0!
0'
#95750000000
1!
b111 %
1'
b111 +
#95760000000
0!
0'
#95770000000
1!
0$
b1000 %
1'
0*
b1000 +
#95780000000
0!
0'
#95790000000
1!
b1001 %
1'
b1001 +
#95800000000
0!
0'
#95810000000
1!
b0 %
1'
b0 +
#95820000000
0!
0'
#95830000000
1!
1$
b1 %
1'
1*
b1 +
#95840000000
0!
0'
#95850000000
1!
b10 %
1'
b10 +
#95860000000
0!
0'
#95870000000
1!
b11 %
1'
b11 +
#95880000000
0!
0'
#95890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#95900000000
0!
0'
#95910000000
1!
b101 %
1'
b101 +
#95920000000
0!
0'
#95930000000
1!
0$
b110 %
1'
0*
b110 +
#95940000000
0!
0'
#95950000000
1!
b111 %
1'
b111 +
#95960000000
0!
0'
#95970000000
1!
b1000 %
1'
b1000 +
#95980000000
0!
0'
#95990000000
1!
b1001 %
1'
b1001 +
#96000000000
0!
0'
#96010000000
1!
b0 %
1'
b0 +
#96020000000
0!
0'
#96030000000
1!
1$
b1 %
1'
1*
b1 +
#96040000000
0!
0'
#96050000000
1!
b10 %
1'
b10 +
#96060000000
0!
0'
#96070000000
1!
b11 %
1'
b11 +
#96080000000
0!
0'
#96090000000
1!
b100 %
1'
b100 +
#96100000000
1"
1(
#96110000000
0!
0"
b100 &
0'
0(
b100 ,
#96120000000
1!
b101 %
1'
b101 +
#96130000000
0!
0'
#96140000000
1!
b110 %
1'
b110 +
#96150000000
0!
0'
#96160000000
1!
b111 %
1'
b111 +
#96170000000
0!
0'
#96180000000
1!
0$
b1000 %
1'
0*
b1000 +
#96190000000
0!
0'
#96200000000
1!
b1001 %
1'
b1001 +
#96210000000
0!
0'
#96220000000
1!
b0 %
1'
b0 +
#96230000000
0!
0'
#96240000000
1!
1$
b1 %
1'
1*
b1 +
#96250000000
0!
0'
#96260000000
1!
b10 %
1'
b10 +
#96270000000
0!
0'
#96280000000
1!
b11 %
1'
b11 +
#96290000000
0!
0'
#96300000000
1!
b100 %
1'
b100 +
#96310000000
0!
0'
#96320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#96330000000
0!
0'
#96340000000
1!
0$
b110 %
1'
0*
b110 +
#96350000000
0!
0'
#96360000000
1!
b111 %
1'
b111 +
#96370000000
0!
0'
#96380000000
1!
b1000 %
1'
b1000 +
#96390000000
0!
0'
#96400000000
1!
b1001 %
1'
b1001 +
#96410000000
0!
0'
#96420000000
1!
b0 %
1'
b0 +
#96430000000
0!
0'
#96440000000
1!
1$
b1 %
1'
1*
b1 +
#96450000000
0!
0'
#96460000000
1!
b10 %
1'
b10 +
#96470000000
0!
0'
#96480000000
1!
b11 %
1'
b11 +
#96490000000
0!
0'
#96500000000
1!
b100 %
1'
b100 +
#96510000000
0!
0'
#96520000000
1!
b101 %
1'
b101 +
#96530000000
1"
1(
#96540000000
0!
0"
b100 &
0'
0(
b100 ,
#96550000000
1!
b110 %
1'
b110 +
#96560000000
0!
0'
#96570000000
1!
b111 %
1'
b111 +
#96580000000
0!
0'
#96590000000
1!
0$
b1000 %
1'
0*
b1000 +
#96600000000
0!
0'
#96610000000
1!
b1001 %
1'
b1001 +
#96620000000
0!
0'
#96630000000
1!
b0 %
1'
b0 +
#96640000000
0!
0'
#96650000000
1!
1$
b1 %
1'
1*
b1 +
#96660000000
0!
0'
#96670000000
1!
b10 %
1'
b10 +
#96680000000
0!
0'
#96690000000
1!
b11 %
1'
b11 +
#96700000000
0!
0'
#96710000000
1!
b100 %
1'
b100 +
#96720000000
0!
0'
#96730000000
1!
b101 %
1'
b101 +
#96740000000
0!
0'
#96750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#96760000000
0!
0'
#96770000000
1!
b111 %
1'
b111 +
#96780000000
0!
0'
#96790000000
1!
b1000 %
1'
b1000 +
#96800000000
0!
0'
#96810000000
1!
b1001 %
1'
b1001 +
#96820000000
0!
0'
#96830000000
1!
b0 %
1'
b0 +
#96840000000
0!
0'
#96850000000
1!
1$
b1 %
1'
1*
b1 +
#96860000000
0!
0'
#96870000000
1!
b10 %
1'
b10 +
#96880000000
0!
0'
#96890000000
1!
b11 %
1'
b11 +
#96900000000
0!
0'
#96910000000
1!
b100 %
1'
b100 +
#96920000000
0!
0'
#96930000000
1!
b101 %
1'
b101 +
#96940000000
0!
0'
#96950000000
1!
0$
b110 %
1'
0*
b110 +
#96960000000
1"
1(
#96970000000
0!
0"
b100 &
0'
0(
b100 ,
#96980000000
1!
1$
b111 %
1'
1*
b111 +
#96990000000
0!
0'
#97000000000
1!
0$
b1000 %
1'
0*
b1000 +
#97010000000
0!
0'
#97020000000
1!
b1001 %
1'
b1001 +
#97030000000
0!
0'
#97040000000
1!
b0 %
1'
b0 +
#97050000000
0!
0'
#97060000000
1!
1$
b1 %
1'
1*
b1 +
#97070000000
0!
0'
#97080000000
1!
b10 %
1'
b10 +
#97090000000
0!
0'
#97100000000
1!
b11 %
1'
b11 +
#97110000000
0!
0'
#97120000000
1!
b100 %
1'
b100 +
#97130000000
0!
0'
#97140000000
1!
b101 %
1'
b101 +
#97150000000
0!
0'
#97160000000
1!
b110 %
1'
b110 +
#97170000000
0!
0'
#97180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#97190000000
0!
0'
#97200000000
1!
b1000 %
1'
b1000 +
#97210000000
0!
0'
#97220000000
1!
b1001 %
1'
b1001 +
#97230000000
0!
0'
#97240000000
1!
b0 %
1'
b0 +
#97250000000
0!
0'
#97260000000
1!
1$
b1 %
1'
1*
b1 +
#97270000000
0!
0'
#97280000000
1!
b10 %
1'
b10 +
#97290000000
0!
0'
#97300000000
1!
b11 %
1'
b11 +
#97310000000
0!
0'
#97320000000
1!
b100 %
1'
b100 +
#97330000000
0!
0'
#97340000000
1!
b101 %
1'
b101 +
#97350000000
0!
0'
#97360000000
1!
0$
b110 %
1'
0*
b110 +
#97370000000
0!
0'
#97380000000
1!
b111 %
1'
b111 +
#97390000000
1"
1(
#97400000000
0!
0"
b100 &
0'
0(
b100 ,
#97410000000
1!
b1000 %
1'
b1000 +
#97420000000
0!
0'
#97430000000
1!
b1001 %
1'
b1001 +
#97440000000
0!
0'
#97450000000
1!
b0 %
1'
b0 +
#97460000000
0!
0'
#97470000000
1!
1$
b1 %
1'
1*
b1 +
#97480000000
0!
0'
#97490000000
1!
b10 %
1'
b10 +
#97500000000
0!
0'
#97510000000
1!
b11 %
1'
b11 +
#97520000000
0!
0'
#97530000000
1!
b100 %
1'
b100 +
#97540000000
0!
0'
#97550000000
1!
b101 %
1'
b101 +
#97560000000
0!
0'
#97570000000
1!
b110 %
1'
b110 +
#97580000000
0!
0'
#97590000000
1!
b111 %
1'
b111 +
#97600000000
0!
0'
#97610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#97620000000
0!
0'
#97630000000
1!
b1001 %
1'
b1001 +
#97640000000
0!
0'
#97650000000
1!
b0 %
1'
b0 +
#97660000000
0!
0'
#97670000000
1!
1$
b1 %
1'
1*
b1 +
#97680000000
0!
0'
#97690000000
1!
b10 %
1'
b10 +
#97700000000
0!
0'
#97710000000
1!
b11 %
1'
b11 +
#97720000000
0!
0'
#97730000000
1!
b100 %
1'
b100 +
#97740000000
0!
0'
#97750000000
1!
b101 %
1'
b101 +
#97760000000
0!
0'
#97770000000
1!
0$
b110 %
1'
0*
b110 +
#97780000000
0!
0'
#97790000000
1!
b111 %
1'
b111 +
#97800000000
0!
0'
#97810000000
1!
b1000 %
1'
b1000 +
#97820000000
1"
1(
#97830000000
0!
0"
b100 &
0'
0(
b100 ,
#97840000000
1!
b1001 %
1'
b1001 +
#97850000000
0!
0'
#97860000000
1!
b0 %
1'
b0 +
#97870000000
0!
0'
#97880000000
1!
1$
b1 %
1'
1*
b1 +
#97890000000
0!
0'
#97900000000
1!
b10 %
1'
b10 +
#97910000000
0!
0'
#97920000000
1!
b11 %
1'
b11 +
#97930000000
0!
0'
#97940000000
1!
b100 %
1'
b100 +
#97950000000
0!
0'
#97960000000
1!
b101 %
1'
b101 +
#97970000000
0!
0'
#97980000000
1!
b110 %
1'
b110 +
#97990000000
0!
0'
#98000000000
1!
b111 %
1'
b111 +
#98010000000
0!
0'
#98020000000
1!
0$
b1000 %
1'
0*
b1000 +
#98030000000
0!
0'
#98040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#98050000000
0!
0'
#98060000000
1!
b0 %
1'
b0 +
#98070000000
0!
0'
#98080000000
1!
1$
b1 %
1'
1*
b1 +
#98090000000
0!
0'
#98100000000
1!
b10 %
1'
b10 +
#98110000000
0!
0'
#98120000000
1!
b11 %
1'
b11 +
#98130000000
0!
0'
#98140000000
1!
b100 %
1'
b100 +
#98150000000
0!
0'
#98160000000
1!
b101 %
1'
b101 +
#98170000000
0!
0'
#98180000000
1!
0$
b110 %
1'
0*
b110 +
#98190000000
0!
0'
#98200000000
1!
b111 %
1'
b111 +
#98210000000
0!
0'
#98220000000
1!
b1000 %
1'
b1000 +
#98230000000
0!
0'
#98240000000
1!
b1001 %
1'
b1001 +
#98250000000
1"
1(
#98260000000
0!
0"
b100 &
0'
0(
b100 ,
#98270000000
1!
b0 %
1'
b0 +
#98280000000
0!
0'
#98290000000
1!
1$
b1 %
1'
1*
b1 +
#98300000000
0!
0'
#98310000000
1!
b10 %
1'
b10 +
#98320000000
0!
0'
#98330000000
1!
b11 %
1'
b11 +
#98340000000
0!
0'
#98350000000
1!
b100 %
1'
b100 +
#98360000000
0!
0'
#98370000000
1!
b101 %
1'
b101 +
#98380000000
0!
0'
#98390000000
1!
b110 %
1'
b110 +
#98400000000
0!
0'
#98410000000
1!
b111 %
1'
b111 +
#98420000000
0!
0'
#98430000000
1!
0$
b1000 %
1'
0*
b1000 +
#98440000000
0!
0'
#98450000000
1!
b1001 %
1'
b1001 +
#98460000000
0!
0'
#98470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#98480000000
0!
0'
#98490000000
1!
1$
b1 %
1'
1*
b1 +
#98500000000
0!
0'
#98510000000
1!
b10 %
1'
b10 +
#98520000000
0!
0'
#98530000000
1!
b11 %
1'
b11 +
#98540000000
0!
0'
#98550000000
1!
b100 %
1'
b100 +
#98560000000
0!
0'
#98570000000
1!
b101 %
1'
b101 +
#98580000000
0!
0'
#98590000000
1!
0$
b110 %
1'
0*
b110 +
#98600000000
0!
0'
#98610000000
1!
b111 %
1'
b111 +
#98620000000
0!
0'
#98630000000
1!
b1000 %
1'
b1000 +
#98640000000
0!
0'
#98650000000
1!
b1001 %
1'
b1001 +
#98660000000
0!
0'
#98670000000
1!
b0 %
1'
b0 +
#98680000000
1"
1(
#98690000000
0!
0"
b100 &
0'
0(
b100 ,
#98700000000
1!
1$
b1 %
1'
1*
b1 +
#98710000000
0!
0'
#98720000000
1!
b10 %
1'
b10 +
#98730000000
0!
0'
#98740000000
1!
b11 %
1'
b11 +
#98750000000
0!
0'
#98760000000
1!
b100 %
1'
b100 +
#98770000000
0!
0'
#98780000000
1!
b101 %
1'
b101 +
#98790000000
0!
0'
#98800000000
1!
b110 %
1'
b110 +
#98810000000
0!
0'
#98820000000
1!
b111 %
1'
b111 +
#98830000000
0!
0'
#98840000000
1!
0$
b1000 %
1'
0*
b1000 +
#98850000000
0!
0'
#98860000000
1!
b1001 %
1'
b1001 +
#98870000000
0!
0'
#98880000000
1!
b0 %
1'
b0 +
#98890000000
0!
0'
#98900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#98910000000
0!
0'
#98920000000
1!
b10 %
1'
b10 +
#98930000000
0!
0'
#98940000000
1!
b11 %
1'
b11 +
#98950000000
0!
0'
#98960000000
1!
b100 %
1'
b100 +
#98970000000
0!
0'
#98980000000
1!
b101 %
1'
b101 +
#98990000000
0!
0'
#99000000000
1!
0$
b110 %
1'
0*
b110 +
#99010000000
0!
0'
#99020000000
1!
b111 %
1'
b111 +
#99030000000
0!
0'
#99040000000
1!
b1000 %
1'
b1000 +
#99050000000
0!
0'
#99060000000
1!
b1001 %
1'
b1001 +
#99070000000
0!
0'
#99080000000
1!
b0 %
1'
b0 +
#99090000000
0!
0'
#99100000000
1!
1$
b1 %
1'
1*
b1 +
#99110000000
1"
1(
#99120000000
0!
0"
b100 &
0'
0(
b100 ,
#99130000000
1!
b10 %
1'
b10 +
#99140000000
0!
0'
#99150000000
1!
b11 %
1'
b11 +
#99160000000
0!
0'
#99170000000
1!
b100 %
1'
b100 +
#99180000000
0!
0'
#99190000000
1!
b101 %
1'
b101 +
#99200000000
0!
0'
#99210000000
1!
b110 %
1'
b110 +
#99220000000
0!
0'
#99230000000
1!
b111 %
1'
b111 +
#99240000000
0!
0'
#99250000000
1!
0$
b1000 %
1'
0*
b1000 +
#99260000000
0!
0'
#99270000000
1!
b1001 %
1'
b1001 +
#99280000000
0!
0'
#99290000000
1!
b0 %
1'
b0 +
#99300000000
0!
0'
#99310000000
1!
1$
b1 %
1'
1*
b1 +
#99320000000
0!
0'
#99330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#99340000000
0!
0'
#99350000000
1!
b11 %
1'
b11 +
#99360000000
0!
0'
#99370000000
1!
b100 %
1'
b100 +
#99380000000
0!
0'
#99390000000
1!
b101 %
1'
b101 +
#99400000000
0!
0'
#99410000000
1!
0$
b110 %
1'
0*
b110 +
#99420000000
0!
0'
#99430000000
1!
b111 %
1'
b111 +
#99440000000
0!
0'
#99450000000
1!
b1000 %
1'
b1000 +
#99460000000
0!
0'
#99470000000
1!
b1001 %
1'
b1001 +
#99480000000
0!
0'
#99490000000
1!
b0 %
1'
b0 +
#99500000000
0!
0'
#99510000000
1!
1$
b1 %
1'
1*
b1 +
#99520000000
0!
0'
#99530000000
1!
b10 %
1'
b10 +
#99540000000
1"
1(
#99550000000
0!
0"
b100 &
0'
0(
b100 ,
#99560000000
1!
b11 %
1'
b11 +
#99570000000
0!
0'
#99580000000
1!
b100 %
1'
b100 +
#99590000000
0!
0'
#99600000000
1!
b101 %
1'
b101 +
#99610000000
0!
0'
#99620000000
1!
b110 %
1'
b110 +
#99630000000
0!
0'
#99640000000
1!
b111 %
1'
b111 +
#99650000000
0!
0'
#99660000000
1!
0$
b1000 %
1'
0*
b1000 +
#99670000000
0!
0'
#99680000000
1!
b1001 %
1'
b1001 +
#99690000000
0!
0'
#99700000000
1!
b0 %
1'
b0 +
#99710000000
0!
0'
#99720000000
1!
1$
b1 %
1'
1*
b1 +
#99730000000
0!
0'
#99740000000
1!
b10 %
1'
b10 +
#99750000000
0!
0'
#99760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#99770000000
0!
0'
#99780000000
1!
b100 %
1'
b100 +
#99790000000
0!
0'
#99800000000
1!
b101 %
1'
b101 +
#99810000000
0!
0'
#99820000000
1!
0$
b110 %
1'
0*
b110 +
#99830000000
0!
0'
#99840000000
1!
b111 %
1'
b111 +
#99850000000
0!
0'
#99860000000
1!
b1000 %
1'
b1000 +
#99870000000
0!
0'
#99880000000
1!
b1001 %
1'
b1001 +
#99890000000
0!
0'
#99900000000
1!
b0 %
1'
b0 +
#99910000000
0!
0'
#99920000000
1!
1$
b1 %
1'
1*
b1 +
#99930000000
0!
0'
#99940000000
1!
b10 %
1'
b10 +
#99950000000
0!
0'
#99960000000
1!
b11 %
1'
b11 +
#99970000000
1"
1(
#99980000000
0!
0"
b100 &
0'
0(
b100 ,
#99990000000
1!
b100 %
1'
b100 +
#100000000000
0!
0'
#100010000000
1!
b101 %
1'
b101 +
#100020000000
0!
0'
#100030000000
1!
b110 %
1'
b110 +
#100040000000
0!
0'
#100050000000
1!
b111 %
1'
b111 +
#100060000000
0!
0'
#100070000000
1!
0$
b1000 %
1'
0*
b1000 +
#100080000000
0!
0'
#100090000000
1!
b1001 %
1'
b1001 +
#100100000000
0!
0'
#100110000000
1!
b0 %
1'
b0 +
#100120000000
0!
0'
#100130000000
1!
1$
b1 %
1'
1*
b1 +
#100140000000
0!
0'
#100150000000
1!
b10 %
1'
b10 +
#100160000000
0!
0'
#100170000000
1!
b11 %
1'
b11 +
#100180000000
0!
0'
#100190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#100200000000
0!
0'
#100210000000
1!
b101 %
1'
b101 +
#100220000000
0!
0'
#100230000000
1!
0$
b110 %
1'
0*
b110 +
#100240000000
0!
0'
#100250000000
1!
b111 %
1'
b111 +
#100260000000
0!
0'
#100270000000
1!
b1000 %
1'
b1000 +
#100280000000
0!
0'
#100290000000
1!
b1001 %
1'
b1001 +
#100300000000
0!
0'
#100310000000
1!
b0 %
1'
b0 +
#100320000000
0!
0'
#100330000000
1!
1$
b1 %
1'
1*
b1 +
#100340000000
0!
0'
#100350000000
1!
b10 %
1'
b10 +
#100360000000
0!
0'
#100370000000
1!
b11 %
1'
b11 +
#100380000000
0!
0'
#100390000000
1!
b100 %
1'
b100 +
#100400000000
1"
1(
#100410000000
0!
0"
b100 &
0'
0(
b100 ,
#100420000000
1!
b101 %
1'
b101 +
#100430000000
0!
0'
#100440000000
1!
b110 %
1'
b110 +
#100450000000
0!
0'
#100460000000
1!
b111 %
1'
b111 +
#100470000000
0!
0'
#100480000000
1!
0$
b1000 %
1'
0*
b1000 +
#100490000000
0!
0'
#100500000000
1!
b1001 %
1'
b1001 +
#100510000000
0!
0'
#100520000000
1!
b0 %
1'
b0 +
#100530000000
0!
0'
#100540000000
1!
1$
b1 %
1'
1*
b1 +
#100550000000
0!
0'
#100560000000
1!
b10 %
1'
b10 +
#100570000000
0!
0'
#100580000000
1!
b11 %
1'
b11 +
#100590000000
0!
0'
#100600000000
1!
b100 %
1'
b100 +
#100610000000
0!
0'
#100620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#100630000000
0!
0'
#100640000000
1!
0$
b110 %
1'
0*
b110 +
#100650000000
0!
0'
#100660000000
1!
b111 %
1'
b111 +
#100670000000
0!
0'
#100680000000
1!
b1000 %
1'
b1000 +
#100690000000
0!
0'
#100700000000
1!
b1001 %
1'
b1001 +
#100710000000
0!
0'
#100720000000
1!
b0 %
1'
b0 +
#100730000000
0!
0'
#100740000000
1!
1$
b1 %
1'
1*
b1 +
#100750000000
0!
0'
#100760000000
1!
b10 %
1'
b10 +
#100770000000
0!
0'
#100780000000
1!
b11 %
1'
b11 +
#100790000000
0!
0'
#100800000000
1!
b100 %
1'
b100 +
#100810000000
0!
0'
#100820000000
1!
b101 %
1'
b101 +
#100830000000
1"
1(
#100840000000
0!
0"
b100 &
0'
0(
b100 ,
#100850000000
1!
b110 %
1'
b110 +
#100860000000
0!
0'
#100870000000
1!
b111 %
1'
b111 +
#100880000000
0!
0'
#100890000000
1!
0$
b1000 %
1'
0*
b1000 +
#100900000000
0!
0'
#100910000000
1!
b1001 %
1'
b1001 +
#100920000000
0!
0'
#100930000000
1!
b0 %
1'
b0 +
#100940000000
0!
0'
#100950000000
1!
1$
b1 %
1'
1*
b1 +
#100960000000
0!
0'
#100970000000
1!
b10 %
1'
b10 +
#100980000000
0!
0'
#100990000000
1!
b11 %
1'
b11 +
#101000000000
0!
0'
#101010000000
1!
b100 %
1'
b100 +
#101020000000
0!
0'
#101030000000
1!
b101 %
1'
b101 +
#101040000000
0!
0'
#101050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#101060000000
0!
0'
#101070000000
1!
b111 %
1'
b111 +
#101080000000
0!
0'
#101090000000
1!
b1000 %
1'
b1000 +
#101100000000
0!
0'
#101110000000
1!
b1001 %
1'
b1001 +
#101120000000
0!
0'
#101130000000
1!
b0 %
1'
b0 +
#101140000000
0!
0'
#101150000000
1!
1$
b1 %
1'
1*
b1 +
#101160000000
0!
0'
#101170000000
1!
b10 %
1'
b10 +
#101180000000
0!
0'
#101190000000
1!
b11 %
1'
b11 +
#101200000000
0!
0'
#101210000000
1!
b100 %
1'
b100 +
#101220000000
0!
0'
#101230000000
1!
b101 %
1'
b101 +
#101240000000
0!
0'
#101250000000
1!
0$
b110 %
1'
0*
b110 +
#101260000000
1"
1(
#101270000000
0!
0"
b100 &
0'
0(
b100 ,
#101280000000
1!
1$
b111 %
1'
1*
b111 +
#101290000000
0!
0'
#101300000000
1!
0$
b1000 %
1'
0*
b1000 +
#101310000000
0!
0'
#101320000000
1!
b1001 %
1'
b1001 +
#101330000000
0!
0'
#101340000000
1!
b0 %
1'
b0 +
#101350000000
0!
0'
#101360000000
1!
1$
b1 %
1'
1*
b1 +
#101370000000
0!
0'
#101380000000
1!
b10 %
1'
b10 +
#101390000000
0!
0'
#101400000000
1!
b11 %
1'
b11 +
#101410000000
0!
0'
#101420000000
1!
b100 %
1'
b100 +
#101430000000
0!
0'
#101440000000
1!
b101 %
1'
b101 +
#101450000000
0!
0'
#101460000000
1!
b110 %
1'
b110 +
#101470000000
0!
0'
#101480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#101490000000
0!
0'
#101500000000
1!
b1000 %
1'
b1000 +
#101510000000
0!
0'
#101520000000
1!
b1001 %
1'
b1001 +
#101530000000
0!
0'
#101540000000
1!
b0 %
1'
b0 +
#101550000000
0!
0'
#101560000000
1!
1$
b1 %
1'
1*
b1 +
#101570000000
0!
0'
#101580000000
1!
b10 %
1'
b10 +
#101590000000
0!
0'
#101600000000
1!
b11 %
1'
b11 +
#101610000000
0!
0'
#101620000000
1!
b100 %
1'
b100 +
#101630000000
0!
0'
#101640000000
1!
b101 %
1'
b101 +
#101650000000
0!
0'
#101660000000
1!
0$
b110 %
1'
0*
b110 +
#101670000000
0!
0'
#101680000000
1!
b111 %
1'
b111 +
#101690000000
1"
1(
#101700000000
0!
0"
b100 &
0'
0(
b100 ,
#101710000000
1!
b1000 %
1'
b1000 +
#101720000000
0!
0'
#101730000000
1!
b1001 %
1'
b1001 +
#101740000000
0!
0'
#101750000000
1!
b0 %
1'
b0 +
#101760000000
0!
0'
#101770000000
1!
1$
b1 %
1'
1*
b1 +
#101780000000
0!
0'
#101790000000
1!
b10 %
1'
b10 +
#101800000000
0!
0'
#101810000000
1!
b11 %
1'
b11 +
#101820000000
0!
0'
#101830000000
1!
b100 %
1'
b100 +
#101840000000
0!
0'
#101850000000
1!
b101 %
1'
b101 +
#101860000000
0!
0'
#101870000000
1!
b110 %
1'
b110 +
#101880000000
0!
0'
#101890000000
1!
b111 %
1'
b111 +
#101900000000
0!
0'
#101910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#101920000000
0!
0'
#101930000000
1!
b1001 %
1'
b1001 +
#101940000000
0!
0'
#101950000000
1!
b0 %
1'
b0 +
#101960000000
0!
0'
#101970000000
1!
1$
b1 %
1'
1*
b1 +
#101980000000
0!
0'
#101990000000
1!
b10 %
1'
b10 +
#102000000000
0!
0'
#102010000000
1!
b11 %
1'
b11 +
#102020000000
0!
0'
#102030000000
1!
b100 %
1'
b100 +
#102040000000
0!
0'
#102050000000
1!
b101 %
1'
b101 +
#102060000000
0!
0'
#102070000000
1!
0$
b110 %
1'
0*
b110 +
#102080000000
0!
0'
#102090000000
1!
b111 %
1'
b111 +
#102100000000
0!
0'
#102110000000
1!
b1000 %
1'
b1000 +
#102120000000
1"
1(
#102130000000
0!
0"
b100 &
0'
0(
b100 ,
#102140000000
1!
b1001 %
1'
b1001 +
#102150000000
0!
0'
#102160000000
1!
b0 %
1'
b0 +
#102170000000
0!
0'
#102180000000
1!
1$
b1 %
1'
1*
b1 +
#102190000000
0!
0'
#102200000000
1!
b10 %
1'
b10 +
#102210000000
0!
0'
#102220000000
1!
b11 %
1'
b11 +
#102230000000
0!
0'
#102240000000
1!
b100 %
1'
b100 +
#102250000000
0!
0'
#102260000000
1!
b101 %
1'
b101 +
#102270000000
0!
0'
#102280000000
1!
b110 %
1'
b110 +
#102290000000
0!
0'
#102300000000
1!
b111 %
1'
b111 +
#102310000000
0!
0'
#102320000000
1!
0$
b1000 %
1'
0*
b1000 +
#102330000000
0!
0'
#102340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#102350000000
0!
0'
#102360000000
1!
b0 %
1'
b0 +
#102370000000
0!
0'
#102380000000
1!
1$
b1 %
1'
1*
b1 +
#102390000000
0!
0'
#102400000000
1!
b10 %
1'
b10 +
#102410000000
0!
0'
#102420000000
1!
b11 %
1'
b11 +
#102430000000
0!
0'
#102440000000
1!
b100 %
1'
b100 +
#102450000000
0!
0'
#102460000000
1!
b101 %
1'
b101 +
#102470000000
0!
0'
#102480000000
1!
0$
b110 %
1'
0*
b110 +
#102490000000
0!
0'
#102500000000
1!
b111 %
1'
b111 +
#102510000000
0!
0'
#102520000000
1!
b1000 %
1'
b1000 +
#102530000000
0!
0'
#102540000000
1!
b1001 %
1'
b1001 +
#102550000000
1"
1(
#102560000000
0!
0"
b100 &
0'
0(
b100 ,
#102570000000
1!
b0 %
1'
b0 +
#102580000000
0!
0'
#102590000000
1!
1$
b1 %
1'
1*
b1 +
#102600000000
0!
0'
#102610000000
1!
b10 %
1'
b10 +
#102620000000
0!
0'
#102630000000
1!
b11 %
1'
b11 +
#102640000000
0!
0'
#102650000000
1!
b100 %
1'
b100 +
#102660000000
0!
0'
#102670000000
1!
b101 %
1'
b101 +
#102680000000
0!
0'
#102690000000
1!
b110 %
1'
b110 +
#102700000000
0!
0'
#102710000000
1!
b111 %
1'
b111 +
#102720000000
0!
0'
#102730000000
1!
0$
b1000 %
1'
0*
b1000 +
#102740000000
0!
0'
#102750000000
1!
b1001 %
1'
b1001 +
#102760000000
0!
0'
#102770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#102780000000
0!
0'
#102790000000
1!
1$
b1 %
1'
1*
b1 +
#102800000000
0!
0'
#102810000000
1!
b10 %
1'
b10 +
#102820000000
0!
0'
#102830000000
1!
b11 %
1'
b11 +
#102840000000
0!
0'
#102850000000
1!
b100 %
1'
b100 +
#102860000000
0!
0'
#102870000000
1!
b101 %
1'
b101 +
#102880000000
0!
0'
#102890000000
1!
0$
b110 %
1'
0*
b110 +
#102900000000
0!
0'
#102910000000
1!
b111 %
1'
b111 +
#102920000000
0!
0'
#102930000000
1!
b1000 %
1'
b1000 +
#102940000000
0!
0'
#102950000000
1!
b1001 %
1'
b1001 +
#102960000000
0!
0'
#102970000000
1!
b0 %
1'
b0 +
#102980000000
1"
1(
#102990000000
0!
0"
b100 &
0'
0(
b100 ,
#103000000000
1!
1$
b1 %
1'
1*
b1 +
#103010000000
0!
0'
#103020000000
1!
b10 %
1'
b10 +
#103030000000
0!
0'
#103040000000
1!
b11 %
1'
b11 +
#103050000000
0!
0'
#103060000000
1!
b100 %
1'
b100 +
#103070000000
0!
0'
#103080000000
1!
b101 %
1'
b101 +
#103090000000
0!
0'
#103100000000
1!
b110 %
1'
b110 +
#103110000000
0!
0'
#103120000000
1!
b111 %
1'
b111 +
#103130000000
0!
0'
#103140000000
1!
0$
b1000 %
1'
0*
b1000 +
#103150000000
0!
0'
#103160000000
1!
b1001 %
1'
b1001 +
#103170000000
0!
0'
#103180000000
1!
b0 %
1'
b0 +
#103190000000
0!
0'
#103200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#103210000000
0!
0'
#103220000000
1!
b10 %
1'
b10 +
#103230000000
0!
0'
#103240000000
1!
b11 %
1'
b11 +
#103250000000
0!
0'
#103260000000
1!
b100 %
1'
b100 +
#103270000000
0!
0'
#103280000000
1!
b101 %
1'
b101 +
#103290000000
0!
0'
#103300000000
1!
0$
b110 %
1'
0*
b110 +
#103310000000
0!
0'
#103320000000
1!
b111 %
1'
b111 +
#103330000000
0!
0'
#103340000000
1!
b1000 %
1'
b1000 +
#103350000000
0!
0'
#103360000000
1!
b1001 %
1'
b1001 +
#103370000000
0!
0'
#103380000000
1!
b0 %
1'
b0 +
#103390000000
0!
0'
#103400000000
1!
1$
b1 %
1'
1*
b1 +
#103410000000
1"
1(
#103420000000
0!
0"
b100 &
0'
0(
b100 ,
#103430000000
1!
b10 %
1'
b10 +
#103440000000
0!
0'
#103450000000
1!
b11 %
1'
b11 +
#103460000000
0!
0'
#103470000000
1!
b100 %
1'
b100 +
#103480000000
0!
0'
#103490000000
1!
b101 %
1'
b101 +
#103500000000
0!
0'
#103510000000
1!
b110 %
1'
b110 +
#103520000000
0!
0'
#103530000000
1!
b111 %
1'
b111 +
#103540000000
0!
0'
#103550000000
1!
0$
b1000 %
1'
0*
b1000 +
#103560000000
0!
0'
#103570000000
1!
b1001 %
1'
b1001 +
#103580000000
0!
0'
#103590000000
1!
b0 %
1'
b0 +
#103600000000
0!
0'
#103610000000
1!
1$
b1 %
1'
1*
b1 +
#103620000000
0!
0'
#103630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#103640000000
0!
0'
#103650000000
1!
b11 %
1'
b11 +
#103660000000
0!
0'
#103670000000
1!
b100 %
1'
b100 +
#103680000000
0!
0'
#103690000000
1!
b101 %
1'
b101 +
#103700000000
0!
0'
#103710000000
1!
0$
b110 %
1'
0*
b110 +
#103720000000
0!
0'
#103730000000
1!
b111 %
1'
b111 +
#103740000000
0!
0'
#103750000000
1!
b1000 %
1'
b1000 +
#103760000000
0!
0'
#103770000000
1!
b1001 %
1'
b1001 +
#103780000000
0!
0'
#103790000000
1!
b0 %
1'
b0 +
#103800000000
0!
0'
#103810000000
1!
1$
b1 %
1'
1*
b1 +
#103820000000
0!
0'
#103830000000
1!
b10 %
1'
b10 +
#103840000000
1"
1(
#103850000000
0!
0"
b100 &
0'
0(
b100 ,
#103860000000
1!
b11 %
1'
b11 +
#103870000000
0!
0'
#103880000000
1!
b100 %
1'
b100 +
#103890000000
0!
0'
#103900000000
1!
b101 %
1'
b101 +
#103910000000
0!
0'
#103920000000
1!
b110 %
1'
b110 +
#103930000000
0!
0'
#103940000000
1!
b111 %
1'
b111 +
#103950000000
0!
0'
#103960000000
1!
0$
b1000 %
1'
0*
b1000 +
#103970000000
0!
0'
#103980000000
1!
b1001 %
1'
b1001 +
#103990000000
0!
0'
#104000000000
1!
b0 %
1'
b0 +
#104010000000
0!
0'
#104020000000
1!
1$
b1 %
1'
1*
b1 +
#104030000000
0!
0'
#104040000000
1!
b10 %
1'
b10 +
#104050000000
0!
0'
#104060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#104070000000
0!
0'
#104080000000
1!
b100 %
1'
b100 +
#104090000000
0!
0'
#104100000000
1!
b101 %
1'
b101 +
#104110000000
0!
0'
#104120000000
1!
0$
b110 %
1'
0*
b110 +
#104130000000
0!
0'
#104140000000
1!
b111 %
1'
b111 +
#104150000000
0!
0'
#104160000000
1!
b1000 %
1'
b1000 +
#104170000000
0!
0'
#104180000000
1!
b1001 %
1'
b1001 +
#104190000000
0!
0'
#104200000000
1!
b0 %
1'
b0 +
#104210000000
0!
0'
#104220000000
1!
1$
b1 %
1'
1*
b1 +
#104230000000
0!
0'
#104240000000
1!
b10 %
1'
b10 +
#104250000000
0!
0'
#104260000000
1!
b11 %
1'
b11 +
#104270000000
1"
1(
#104280000000
0!
0"
b100 &
0'
0(
b100 ,
#104290000000
1!
b100 %
1'
b100 +
#104300000000
0!
0'
#104310000000
1!
b101 %
1'
b101 +
#104320000000
0!
0'
#104330000000
1!
b110 %
1'
b110 +
#104340000000
0!
0'
#104350000000
1!
b111 %
1'
b111 +
#104360000000
0!
0'
#104370000000
1!
0$
b1000 %
1'
0*
b1000 +
#104380000000
0!
0'
#104390000000
1!
b1001 %
1'
b1001 +
#104400000000
0!
0'
#104410000000
1!
b0 %
1'
b0 +
#104420000000
0!
0'
#104430000000
1!
1$
b1 %
1'
1*
b1 +
#104440000000
0!
0'
#104450000000
1!
b10 %
1'
b10 +
#104460000000
0!
0'
#104470000000
1!
b11 %
1'
b11 +
#104480000000
0!
0'
#104490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#104500000000
0!
0'
#104510000000
1!
b101 %
1'
b101 +
#104520000000
0!
0'
#104530000000
1!
0$
b110 %
1'
0*
b110 +
#104540000000
0!
0'
#104550000000
1!
b111 %
1'
b111 +
#104560000000
0!
0'
#104570000000
1!
b1000 %
1'
b1000 +
#104580000000
0!
0'
#104590000000
1!
b1001 %
1'
b1001 +
#104600000000
0!
0'
#104610000000
1!
b0 %
1'
b0 +
#104620000000
0!
0'
#104630000000
1!
1$
b1 %
1'
1*
b1 +
#104640000000
0!
0'
#104650000000
1!
b10 %
1'
b10 +
#104660000000
0!
0'
#104670000000
1!
b11 %
1'
b11 +
#104680000000
0!
0'
#104690000000
1!
b100 %
1'
b100 +
#104700000000
1"
1(
#104710000000
0!
0"
b100 &
0'
0(
b100 ,
#104720000000
1!
b101 %
1'
b101 +
#104730000000
0!
0'
#104740000000
1!
b110 %
1'
b110 +
#104750000000
0!
0'
#104760000000
1!
b111 %
1'
b111 +
#104770000000
0!
0'
#104780000000
1!
0$
b1000 %
1'
0*
b1000 +
#104790000000
0!
0'
#104800000000
1!
b1001 %
1'
b1001 +
#104810000000
0!
0'
#104820000000
1!
b0 %
1'
b0 +
#104830000000
0!
0'
#104840000000
1!
1$
b1 %
1'
1*
b1 +
#104850000000
0!
0'
#104860000000
1!
b10 %
1'
b10 +
#104870000000
0!
0'
#104880000000
1!
b11 %
1'
b11 +
#104890000000
0!
0'
#104900000000
1!
b100 %
1'
b100 +
#104910000000
0!
0'
#104920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#104930000000
0!
0'
#104940000000
1!
0$
b110 %
1'
0*
b110 +
#104950000000
0!
0'
#104960000000
1!
b111 %
1'
b111 +
#104970000000
0!
0'
#104980000000
1!
b1000 %
1'
b1000 +
#104990000000
0!
0'
#105000000000
1!
b1001 %
1'
b1001 +
#105010000000
0!
0'
#105020000000
1!
b0 %
1'
b0 +
#105030000000
0!
0'
#105040000000
1!
1$
b1 %
1'
1*
b1 +
#105050000000
0!
0'
#105060000000
1!
b10 %
1'
b10 +
#105070000000
0!
0'
#105080000000
1!
b11 %
1'
b11 +
#105090000000
0!
0'
#105100000000
1!
b100 %
1'
b100 +
#105110000000
0!
0'
#105120000000
1!
b101 %
1'
b101 +
#105130000000
1"
1(
#105140000000
0!
0"
b100 &
0'
0(
b100 ,
#105150000000
1!
b110 %
1'
b110 +
#105160000000
0!
0'
#105170000000
1!
b111 %
1'
b111 +
#105180000000
0!
0'
#105190000000
1!
0$
b1000 %
1'
0*
b1000 +
#105200000000
0!
0'
#105210000000
1!
b1001 %
1'
b1001 +
#105220000000
0!
0'
#105230000000
1!
b0 %
1'
b0 +
#105240000000
0!
0'
#105250000000
1!
1$
b1 %
1'
1*
b1 +
#105260000000
0!
0'
#105270000000
1!
b10 %
1'
b10 +
#105280000000
0!
0'
#105290000000
1!
b11 %
1'
b11 +
#105300000000
0!
0'
#105310000000
1!
b100 %
1'
b100 +
#105320000000
0!
0'
#105330000000
1!
b101 %
1'
b101 +
#105340000000
0!
0'
#105350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#105360000000
0!
0'
#105370000000
1!
b111 %
1'
b111 +
#105380000000
0!
0'
#105390000000
1!
b1000 %
1'
b1000 +
#105400000000
0!
0'
#105410000000
1!
b1001 %
1'
b1001 +
#105420000000
0!
0'
#105430000000
1!
b0 %
1'
b0 +
#105440000000
0!
0'
#105450000000
1!
1$
b1 %
1'
1*
b1 +
#105460000000
0!
0'
#105470000000
1!
b10 %
1'
b10 +
#105480000000
0!
0'
#105490000000
1!
b11 %
1'
b11 +
#105500000000
0!
0'
#105510000000
1!
b100 %
1'
b100 +
#105520000000
0!
0'
#105530000000
1!
b101 %
1'
b101 +
#105540000000
0!
0'
#105550000000
1!
0$
b110 %
1'
0*
b110 +
#105560000000
1"
1(
#105570000000
0!
0"
b100 &
0'
0(
b100 ,
#105580000000
1!
1$
b111 %
1'
1*
b111 +
#105590000000
0!
0'
#105600000000
1!
0$
b1000 %
1'
0*
b1000 +
#105610000000
0!
0'
#105620000000
1!
b1001 %
1'
b1001 +
#105630000000
0!
0'
#105640000000
1!
b0 %
1'
b0 +
#105650000000
0!
0'
#105660000000
1!
1$
b1 %
1'
1*
b1 +
#105670000000
0!
0'
#105680000000
1!
b10 %
1'
b10 +
#105690000000
0!
0'
#105700000000
1!
b11 %
1'
b11 +
#105710000000
0!
0'
#105720000000
1!
b100 %
1'
b100 +
#105730000000
0!
0'
#105740000000
1!
b101 %
1'
b101 +
#105750000000
0!
0'
#105760000000
1!
b110 %
1'
b110 +
#105770000000
0!
0'
#105780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#105790000000
0!
0'
#105800000000
1!
b1000 %
1'
b1000 +
#105810000000
0!
0'
#105820000000
1!
b1001 %
1'
b1001 +
#105830000000
0!
0'
#105840000000
1!
b0 %
1'
b0 +
#105850000000
0!
0'
#105860000000
1!
1$
b1 %
1'
1*
b1 +
#105870000000
0!
0'
#105880000000
1!
b10 %
1'
b10 +
#105890000000
0!
0'
#105900000000
1!
b11 %
1'
b11 +
#105910000000
0!
0'
#105920000000
1!
b100 %
1'
b100 +
#105930000000
0!
0'
#105940000000
1!
b101 %
1'
b101 +
#105950000000
0!
0'
#105960000000
1!
0$
b110 %
1'
0*
b110 +
#105970000000
0!
0'
#105980000000
1!
b111 %
1'
b111 +
#105990000000
1"
1(
#106000000000
0!
0"
b100 &
0'
0(
b100 ,
#106010000000
1!
b1000 %
1'
b1000 +
#106020000000
0!
0'
#106030000000
1!
b1001 %
1'
b1001 +
#106040000000
0!
0'
#106050000000
1!
b0 %
1'
b0 +
#106060000000
0!
0'
#106070000000
1!
1$
b1 %
1'
1*
b1 +
#106080000000
0!
0'
#106090000000
1!
b10 %
1'
b10 +
#106100000000
0!
0'
#106110000000
1!
b11 %
1'
b11 +
#106120000000
0!
0'
#106130000000
1!
b100 %
1'
b100 +
#106140000000
0!
0'
#106150000000
1!
b101 %
1'
b101 +
#106160000000
0!
0'
#106170000000
1!
b110 %
1'
b110 +
#106180000000
0!
0'
#106190000000
1!
b111 %
1'
b111 +
#106200000000
0!
0'
#106210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#106220000000
0!
0'
#106230000000
1!
b1001 %
1'
b1001 +
#106240000000
0!
0'
#106250000000
1!
b0 %
1'
b0 +
#106260000000
0!
0'
#106270000000
1!
1$
b1 %
1'
1*
b1 +
#106280000000
0!
0'
#106290000000
1!
b10 %
1'
b10 +
#106300000000
0!
0'
#106310000000
1!
b11 %
1'
b11 +
#106320000000
0!
0'
#106330000000
1!
b100 %
1'
b100 +
#106340000000
0!
0'
#106350000000
1!
b101 %
1'
b101 +
#106360000000
0!
0'
#106370000000
1!
0$
b110 %
1'
0*
b110 +
#106380000000
0!
0'
#106390000000
1!
b111 %
1'
b111 +
#106400000000
0!
0'
#106410000000
1!
b1000 %
1'
b1000 +
#106420000000
1"
1(
#106430000000
0!
0"
b100 &
0'
0(
b100 ,
#106440000000
1!
b1001 %
1'
b1001 +
#106450000000
0!
0'
#106460000000
1!
b0 %
1'
b0 +
#106470000000
0!
0'
#106480000000
1!
1$
b1 %
1'
1*
b1 +
#106490000000
0!
0'
#106500000000
1!
b10 %
1'
b10 +
#106510000000
0!
0'
#106520000000
1!
b11 %
1'
b11 +
#106530000000
0!
0'
#106540000000
1!
b100 %
1'
b100 +
#106550000000
0!
0'
#106560000000
1!
b101 %
1'
b101 +
#106570000000
0!
0'
#106580000000
1!
b110 %
1'
b110 +
#106590000000
0!
0'
#106600000000
1!
b111 %
1'
b111 +
#106610000000
0!
0'
#106620000000
1!
0$
b1000 %
1'
0*
b1000 +
#106630000000
0!
0'
#106640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#106650000000
0!
0'
#106660000000
1!
b0 %
1'
b0 +
#106670000000
0!
0'
#106680000000
1!
1$
b1 %
1'
1*
b1 +
#106690000000
0!
0'
#106700000000
1!
b10 %
1'
b10 +
#106710000000
0!
0'
#106720000000
1!
b11 %
1'
b11 +
#106730000000
0!
0'
#106740000000
1!
b100 %
1'
b100 +
#106750000000
0!
0'
#106760000000
1!
b101 %
1'
b101 +
#106770000000
0!
0'
#106780000000
1!
0$
b110 %
1'
0*
b110 +
#106790000000
0!
0'
#106800000000
1!
b111 %
1'
b111 +
#106810000000
0!
0'
#106820000000
1!
b1000 %
1'
b1000 +
#106830000000
0!
0'
#106840000000
1!
b1001 %
1'
b1001 +
#106850000000
1"
1(
#106860000000
0!
0"
b100 &
0'
0(
b100 ,
#106870000000
1!
b0 %
1'
b0 +
#106880000000
0!
0'
#106890000000
1!
1$
b1 %
1'
1*
b1 +
#106900000000
0!
0'
#106910000000
1!
b10 %
1'
b10 +
#106920000000
0!
0'
#106930000000
1!
b11 %
1'
b11 +
#106940000000
0!
0'
#106950000000
1!
b100 %
1'
b100 +
#106960000000
0!
0'
#106970000000
1!
b101 %
1'
b101 +
#106980000000
0!
0'
#106990000000
1!
b110 %
1'
b110 +
#107000000000
0!
0'
#107010000000
1!
b111 %
1'
b111 +
#107020000000
0!
0'
#107030000000
1!
0$
b1000 %
1'
0*
b1000 +
#107040000000
0!
0'
#107050000000
1!
b1001 %
1'
b1001 +
#107060000000
0!
0'
#107070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#107080000000
0!
0'
#107090000000
1!
1$
b1 %
1'
1*
b1 +
#107100000000
0!
0'
#107110000000
1!
b10 %
1'
b10 +
#107120000000
0!
0'
#107130000000
1!
b11 %
1'
b11 +
#107140000000
0!
0'
#107150000000
1!
b100 %
1'
b100 +
#107160000000
0!
0'
#107170000000
1!
b101 %
1'
b101 +
#107180000000
0!
0'
#107190000000
1!
0$
b110 %
1'
0*
b110 +
#107200000000
0!
0'
#107210000000
1!
b111 %
1'
b111 +
#107220000000
0!
0'
#107230000000
1!
b1000 %
1'
b1000 +
#107240000000
0!
0'
#107250000000
1!
b1001 %
1'
b1001 +
#107260000000
0!
0'
#107270000000
1!
b0 %
1'
b0 +
#107280000000
1"
1(
#107290000000
0!
0"
b100 &
0'
0(
b100 ,
#107300000000
1!
1$
b1 %
1'
1*
b1 +
#107310000000
0!
0'
#107320000000
1!
b10 %
1'
b10 +
#107330000000
0!
0'
#107340000000
1!
b11 %
1'
b11 +
#107350000000
0!
0'
#107360000000
1!
b100 %
1'
b100 +
#107370000000
0!
0'
#107380000000
1!
b101 %
1'
b101 +
#107390000000
0!
0'
#107400000000
1!
b110 %
1'
b110 +
#107410000000
0!
0'
#107420000000
1!
b111 %
1'
b111 +
#107430000000
0!
0'
#107440000000
1!
0$
b1000 %
1'
0*
b1000 +
#107450000000
0!
0'
#107460000000
1!
b1001 %
1'
b1001 +
#107470000000
0!
0'
#107480000000
1!
b0 %
1'
b0 +
#107490000000
0!
0'
#107500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#107510000000
0!
0'
#107520000000
1!
b10 %
1'
b10 +
#107530000000
0!
0'
#107540000000
1!
b11 %
1'
b11 +
#107550000000
0!
0'
#107560000000
1!
b100 %
1'
b100 +
#107570000000
0!
0'
#107580000000
1!
b101 %
1'
b101 +
#107590000000
0!
0'
#107600000000
1!
0$
b110 %
1'
0*
b110 +
#107610000000
0!
0'
#107620000000
1!
b111 %
1'
b111 +
#107630000000
0!
0'
#107640000000
1!
b1000 %
1'
b1000 +
#107650000000
0!
0'
#107660000000
1!
b1001 %
1'
b1001 +
#107670000000
0!
0'
#107680000000
1!
b0 %
1'
b0 +
#107690000000
0!
0'
#107700000000
1!
1$
b1 %
1'
1*
b1 +
#107710000000
1"
1(
#107720000000
0!
0"
b100 &
0'
0(
b100 ,
#107730000000
1!
b10 %
1'
b10 +
#107740000000
0!
0'
#107750000000
1!
b11 %
1'
b11 +
#107760000000
0!
0'
#107770000000
1!
b100 %
1'
b100 +
#107780000000
0!
0'
#107790000000
1!
b101 %
1'
b101 +
#107800000000
0!
0'
#107810000000
1!
b110 %
1'
b110 +
#107820000000
0!
0'
#107830000000
1!
b111 %
1'
b111 +
#107840000000
0!
0'
#107850000000
1!
0$
b1000 %
1'
0*
b1000 +
#107860000000
0!
0'
#107870000000
1!
b1001 %
1'
b1001 +
#107880000000
0!
0'
#107890000000
1!
b0 %
1'
b0 +
#107900000000
0!
0'
#107910000000
1!
1$
b1 %
1'
1*
b1 +
#107920000000
0!
0'
#107930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#107940000000
0!
0'
#107950000000
1!
b11 %
1'
b11 +
#107960000000
0!
0'
#107970000000
1!
b100 %
1'
b100 +
#107980000000
0!
0'
#107990000000
1!
b101 %
1'
b101 +
#108000000000
0!
0'
#108010000000
1!
0$
b110 %
1'
0*
b110 +
#108020000000
0!
0'
#108030000000
1!
b111 %
1'
b111 +
#108040000000
0!
0'
#108050000000
1!
b1000 %
1'
b1000 +
#108060000000
0!
0'
#108070000000
1!
b1001 %
1'
b1001 +
#108080000000
0!
0'
#108090000000
1!
b0 %
1'
b0 +
#108100000000
0!
0'
#108110000000
1!
1$
b1 %
1'
1*
b1 +
#108120000000
0!
0'
#108130000000
1!
b10 %
1'
b10 +
#108140000000
1"
1(
#108150000000
0!
0"
b100 &
0'
0(
b100 ,
#108160000000
1!
b11 %
1'
b11 +
#108170000000
0!
0'
#108180000000
1!
b100 %
1'
b100 +
#108190000000
0!
0'
#108200000000
1!
b101 %
1'
b101 +
#108210000000
0!
0'
#108220000000
1!
b110 %
1'
b110 +
#108230000000
0!
0'
#108240000000
1!
b111 %
1'
b111 +
#108250000000
0!
0'
#108260000000
1!
0$
b1000 %
1'
0*
b1000 +
#108270000000
0!
0'
#108280000000
1!
b1001 %
1'
b1001 +
#108290000000
0!
0'
#108300000000
1!
b0 %
1'
b0 +
#108310000000
0!
0'
#108320000000
1!
1$
b1 %
1'
1*
b1 +
#108330000000
0!
0'
#108340000000
1!
b10 %
1'
b10 +
#108350000000
0!
0'
#108360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#108370000000
0!
0'
#108380000000
1!
b100 %
1'
b100 +
#108390000000
0!
0'
#108400000000
1!
b101 %
1'
b101 +
#108410000000
0!
0'
#108420000000
1!
0$
b110 %
1'
0*
b110 +
#108430000000
0!
0'
#108440000000
1!
b111 %
1'
b111 +
#108450000000
0!
0'
#108460000000
1!
b1000 %
1'
b1000 +
#108470000000
0!
0'
#108480000000
1!
b1001 %
1'
b1001 +
#108490000000
0!
0'
#108500000000
1!
b0 %
1'
b0 +
#108510000000
0!
0'
#108520000000
1!
1$
b1 %
1'
1*
b1 +
#108530000000
0!
0'
#108540000000
1!
b10 %
1'
b10 +
#108550000000
0!
0'
#108560000000
1!
b11 %
1'
b11 +
#108570000000
1"
1(
#108580000000
0!
0"
b100 &
0'
0(
b100 ,
#108590000000
1!
b100 %
1'
b100 +
#108600000000
0!
0'
#108610000000
1!
b101 %
1'
b101 +
#108620000000
0!
0'
#108630000000
1!
b110 %
1'
b110 +
#108640000000
0!
0'
#108650000000
1!
b111 %
1'
b111 +
#108660000000
0!
0'
#108670000000
1!
0$
b1000 %
1'
0*
b1000 +
#108680000000
0!
0'
#108690000000
1!
b1001 %
1'
b1001 +
#108700000000
0!
0'
#108710000000
1!
b0 %
1'
b0 +
#108720000000
0!
0'
#108730000000
1!
1$
b1 %
1'
1*
b1 +
#108740000000
0!
0'
#108750000000
1!
b10 %
1'
b10 +
#108760000000
0!
0'
#108770000000
1!
b11 %
1'
b11 +
#108780000000
0!
0'
#108790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#108800000000
0!
0'
#108810000000
1!
b101 %
1'
b101 +
#108820000000
0!
0'
#108830000000
1!
0$
b110 %
1'
0*
b110 +
#108840000000
0!
0'
#108850000000
1!
b111 %
1'
b111 +
#108860000000
0!
0'
#108870000000
1!
b1000 %
1'
b1000 +
#108880000000
0!
0'
#108890000000
1!
b1001 %
1'
b1001 +
#108900000000
0!
0'
#108910000000
1!
b0 %
1'
b0 +
#108920000000
0!
0'
#108930000000
1!
1$
b1 %
1'
1*
b1 +
#108940000000
0!
0'
#108950000000
1!
b10 %
1'
b10 +
#108960000000
0!
0'
#108970000000
1!
b11 %
1'
b11 +
#108980000000
0!
0'
#108990000000
1!
b100 %
1'
b100 +
#109000000000
1"
1(
#109010000000
0!
0"
b100 &
0'
0(
b100 ,
#109020000000
1!
b101 %
1'
b101 +
#109030000000
0!
0'
#109040000000
1!
b110 %
1'
b110 +
#109050000000
0!
0'
#109060000000
1!
b111 %
1'
b111 +
#109070000000
0!
0'
#109080000000
1!
0$
b1000 %
1'
0*
b1000 +
#109090000000
0!
0'
#109100000000
1!
b1001 %
1'
b1001 +
#109110000000
0!
0'
#109120000000
1!
b0 %
1'
b0 +
#109130000000
0!
0'
#109140000000
1!
1$
b1 %
1'
1*
b1 +
#109150000000
0!
0'
#109160000000
1!
b10 %
1'
b10 +
#109170000000
0!
0'
#109180000000
1!
b11 %
1'
b11 +
#109190000000
0!
0'
#109200000000
1!
b100 %
1'
b100 +
#109210000000
0!
0'
#109220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#109230000000
0!
0'
#109240000000
1!
0$
b110 %
1'
0*
b110 +
#109250000000
0!
0'
#109260000000
1!
b111 %
1'
b111 +
#109270000000
0!
0'
#109280000000
1!
b1000 %
1'
b1000 +
#109290000000
0!
0'
#109300000000
1!
b1001 %
1'
b1001 +
#109310000000
0!
0'
#109320000000
1!
b0 %
1'
b0 +
#109330000000
0!
0'
#109340000000
1!
1$
b1 %
1'
1*
b1 +
#109350000000
0!
0'
#109360000000
1!
b10 %
1'
b10 +
#109370000000
0!
0'
#109380000000
1!
b11 %
1'
b11 +
#109390000000
0!
0'
#109400000000
1!
b100 %
1'
b100 +
#109410000000
0!
0'
#109420000000
1!
b101 %
1'
b101 +
#109430000000
1"
1(
#109440000000
0!
0"
b100 &
0'
0(
b100 ,
#109450000000
1!
b110 %
1'
b110 +
#109460000000
0!
0'
#109470000000
1!
b111 %
1'
b111 +
#109480000000
0!
0'
#109490000000
1!
0$
b1000 %
1'
0*
b1000 +
#109500000000
0!
0'
#109510000000
1!
b1001 %
1'
b1001 +
#109520000000
0!
0'
#109530000000
1!
b0 %
1'
b0 +
#109540000000
0!
0'
#109550000000
1!
1$
b1 %
1'
1*
b1 +
#109560000000
0!
0'
#109570000000
1!
b10 %
1'
b10 +
#109580000000
0!
0'
#109590000000
1!
b11 %
1'
b11 +
#109600000000
0!
0'
#109610000000
1!
b100 %
1'
b100 +
#109620000000
0!
0'
#109630000000
1!
b101 %
1'
b101 +
#109640000000
0!
0'
#109650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#109660000000
0!
0'
#109670000000
1!
b111 %
1'
b111 +
#109680000000
0!
0'
#109690000000
1!
b1000 %
1'
b1000 +
#109700000000
0!
0'
#109710000000
1!
b1001 %
1'
b1001 +
#109720000000
0!
0'
#109730000000
1!
b0 %
1'
b0 +
#109740000000
0!
0'
#109750000000
1!
1$
b1 %
1'
1*
b1 +
#109760000000
0!
0'
#109770000000
1!
b10 %
1'
b10 +
#109780000000
0!
0'
#109790000000
1!
b11 %
1'
b11 +
#109800000000
0!
0'
#109810000000
1!
b100 %
1'
b100 +
#109820000000
0!
0'
#109830000000
1!
b101 %
1'
b101 +
#109840000000
0!
0'
#109850000000
1!
0$
b110 %
1'
0*
b110 +
#109860000000
1"
1(
#109870000000
0!
0"
b100 &
0'
0(
b100 ,
#109880000000
1!
1$
b111 %
1'
1*
b111 +
#109890000000
0!
0'
#109900000000
1!
0$
b1000 %
1'
0*
b1000 +
#109910000000
0!
0'
#109920000000
1!
b1001 %
1'
b1001 +
#109930000000
0!
0'
#109940000000
1!
b0 %
1'
b0 +
#109950000000
0!
0'
#109960000000
1!
1$
b1 %
1'
1*
b1 +
#109970000000
0!
0'
#109980000000
1!
b10 %
1'
b10 +
#109990000000
0!
0'
#110000000000
1!
b11 %
1'
b11 +
#110010000000
0!
0'
#110020000000
1!
b100 %
1'
b100 +
#110030000000
0!
0'
#110040000000
1!
b101 %
1'
b101 +
#110050000000
0!
0'
#110060000000
1!
b110 %
1'
b110 +
#110070000000
0!
0'
#110080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#110090000000
0!
0'
#110100000000
1!
b1000 %
1'
b1000 +
#110110000000
0!
0'
#110120000000
1!
b1001 %
1'
b1001 +
#110130000000
0!
0'
#110140000000
1!
b0 %
1'
b0 +
#110150000000
0!
0'
#110160000000
1!
1$
b1 %
1'
1*
b1 +
#110170000000
0!
0'
#110180000000
1!
b10 %
1'
b10 +
#110190000000
0!
0'
#110200000000
1!
b11 %
1'
b11 +
#110210000000
0!
0'
#110220000000
1!
b100 %
1'
b100 +
#110230000000
0!
0'
#110240000000
1!
b101 %
1'
b101 +
#110250000000
0!
0'
#110260000000
1!
0$
b110 %
1'
0*
b110 +
#110270000000
0!
0'
#110280000000
1!
b111 %
1'
b111 +
#110290000000
1"
1(
#110300000000
0!
0"
b100 &
0'
0(
b100 ,
#110310000000
1!
b1000 %
1'
b1000 +
#110320000000
0!
0'
#110330000000
1!
b1001 %
1'
b1001 +
#110340000000
0!
0'
#110350000000
1!
b0 %
1'
b0 +
#110360000000
0!
0'
#110370000000
1!
1$
b1 %
1'
1*
b1 +
#110380000000
0!
0'
#110390000000
1!
b10 %
1'
b10 +
#110400000000
0!
0'
#110410000000
1!
b11 %
1'
b11 +
#110420000000
0!
0'
#110430000000
1!
b100 %
1'
b100 +
#110440000000
0!
0'
#110450000000
1!
b101 %
1'
b101 +
#110460000000
0!
0'
#110470000000
1!
b110 %
1'
b110 +
#110480000000
0!
0'
#110490000000
1!
b111 %
1'
b111 +
#110500000000
0!
0'
#110510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#110520000000
0!
0'
#110530000000
1!
b1001 %
1'
b1001 +
#110540000000
0!
0'
#110550000000
1!
b0 %
1'
b0 +
#110560000000
0!
0'
#110570000000
1!
1$
b1 %
1'
1*
b1 +
#110580000000
0!
0'
#110590000000
1!
b10 %
1'
b10 +
#110600000000
0!
0'
#110610000000
1!
b11 %
1'
b11 +
#110620000000
0!
0'
#110630000000
1!
b100 %
1'
b100 +
#110640000000
0!
0'
#110650000000
1!
b101 %
1'
b101 +
#110660000000
0!
0'
#110670000000
1!
0$
b110 %
1'
0*
b110 +
#110680000000
0!
0'
#110690000000
1!
b111 %
1'
b111 +
#110700000000
0!
0'
#110710000000
1!
b1000 %
1'
b1000 +
#110720000000
1"
1(
#110730000000
0!
0"
b100 &
0'
0(
b100 ,
#110740000000
1!
b1001 %
1'
b1001 +
#110750000000
0!
0'
#110760000000
1!
b0 %
1'
b0 +
#110770000000
0!
0'
#110780000000
1!
1$
b1 %
1'
1*
b1 +
#110790000000
0!
0'
#110800000000
1!
b10 %
1'
b10 +
#110810000000
0!
0'
#110820000000
1!
b11 %
1'
b11 +
#110830000000
0!
0'
#110840000000
1!
b100 %
1'
b100 +
#110850000000
0!
0'
#110860000000
1!
b101 %
1'
b101 +
#110870000000
0!
0'
#110880000000
1!
b110 %
1'
b110 +
#110890000000
0!
0'
#110900000000
1!
b111 %
1'
b111 +
#110910000000
0!
0'
#110920000000
1!
0$
b1000 %
1'
0*
b1000 +
#110930000000
0!
0'
#110940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#110950000000
0!
0'
#110960000000
1!
b0 %
1'
b0 +
#110970000000
0!
0'
#110980000000
1!
1$
b1 %
1'
1*
b1 +
#110990000000
0!
0'
#111000000000
1!
b10 %
1'
b10 +
#111010000000
0!
0'
#111020000000
1!
b11 %
1'
b11 +
#111030000000
0!
0'
#111040000000
1!
b100 %
1'
b100 +
#111050000000
0!
0'
#111060000000
1!
b101 %
1'
b101 +
#111070000000
0!
0'
#111080000000
1!
0$
b110 %
1'
0*
b110 +
#111090000000
0!
0'
#111100000000
1!
b111 %
1'
b111 +
#111110000000
0!
0'
#111120000000
1!
b1000 %
1'
b1000 +
#111130000000
0!
0'
#111140000000
1!
b1001 %
1'
b1001 +
#111150000000
1"
1(
#111160000000
0!
0"
b100 &
0'
0(
b100 ,
#111170000000
1!
b0 %
1'
b0 +
#111180000000
0!
0'
#111190000000
1!
1$
b1 %
1'
1*
b1 +
#111200000000
0!
0'
#111210000000
1!
b10 %
1'
b10 +
#111220000000
0!
0'
#111230000000
1!
b11 %
1'
b11 +
#111240000000
0!
0'
#111250000000
1!
b100 %
1'
b100 +
#111260000000
0!
0'
#111270000000
1!
b101 %
1'
b101 +
#111280000000
0!
0'
#111290000000
1!
b110 %
1'
b110 +
#111300000000
0!
0'
#111310000000
1!
b111 %
1'
b111 +
#111320000000
0!
0'
#111330000000
1!
0$
b1000 %
1'
0*
b1000 +
#111340000000
0!
0'
#111350000000
1!
b1001 %
1'
b1001 +
#111360000000
0!
0'
#111370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#111380000000
0!
0'
#111390000000
1!
1$
b1 %
1'
1*
b1 +
#111400000000
0!
0'
#111410000000
1!
b10 %
1'
b10 +
#111420000000
0!
0'
#111430000000
1!
b11 %
1'
b11 +
#111440000000
0!
0'
#111450000000
1!
b100 %
1'
b100 +
#111460000000
0!
0'
#111470000000
1!
b101 %
1'
b101 +
#111480000000
0!
0'
#111490000000
1!
0$
b110 %
1'
0*
b110 +
#111500000000
0!
0'
#111510000000
1!
b111 %
1'
b111 +
#111520000000
0!
0'
#111530000000
1!
b1000 %
1'
b1000 +
#111540000000
0!
0'
#111550000000
1!
b1001 %
1'
b1001 +
#111560000000
0!
0'
#111570000000
1!
b0 %
1'
b0 +
#111580000000
1"
1(
#111590000000
0!
0"
b100 &
0'
0(
b100 ,
#111600000000
1!
1$
b1 %
1'
1*
b1 +
#111610000000
0!
0'
#111620000000
1!
b10 %
1'
b10 +
#111630000000
0!
0'
#111640000000
1!
b11 %
1'
b11 +
#111650000000
0!
0'
#111660000000
1!
b100 %
1'
b100 +
#111670000000
0!
0'
#111680000000
1!
b101 %
1'
b101 +
#111690000000
0!
0'
#111700000000
1!
b110 %
1'
b110 +
#111710000000
0!
0'
#111720000000
1!
b111 %
1'
b111 +
#111730000000
0!
0'
#111740000000
1!
0$
b1000 %
1'
0*
b1000 +
#111750000000
0!
0'
#111760000000
1!
b1001 %
1'
b1001 +
#111770000000
0!
0'
#111780000000
1!
b0 %
1'
b0 +
#111790000000
0!
0'
#111800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#111810000000
0!
0'
#111820000000
1!
b10 %
1'
b10 +
#111830000000
0!
0'
#111840000000
1!
b11 %
1'
b11 +
#111850000000
0!
0'
#111860000000
1!
b100 %
1'
b100 +
#111870000000
0!
0'
#111880000000
1!
b101 %
1'
b101 +
#111890000000
0!
0'
#111900000000
1!
0$
b110 %
1'
0*
b110 +
#111910000000
0!
0'
#111920000000
1!
b111 %
1'
b111 +
#111930000000
0!
0'
#111940000000
1!
b1000 %
1'
b1000 +
#111950000000
0!
0'
#111960000000
1!
b1001 %
1'
b1001 +
#111970000000
0!
0'
#111980000000
1!
b0 %
1'
b0 +
#111990000000
0!
0'
#112000000000
1!
1$
b1 %
1'
1*
b1 +
#112010000000
1"
1(
#112020000000
0!
0"
b100 &
0'
0(
b100 ,
#112030000000
1!
b10 %
1'
b10 +
#112040000000
0!
0'
#112050000000
1!
b11 %
1'
b11 +
#112060000000
0!
0'
#112070000000
1!
b100 %
1'
b100 +
#112080000000
0!
0'
#112090000000
1!
b101 %
1'
b101 +
#112100000000
0!
0'
#112110000000
1!
b110 %
1'
b110 +
#112120000000
0!
0'
#112130000000
1!
b111 %
1'
b111 +
#112140000000
0!
0'
#112150000000
1!
0$
b1000 %
1'
0*
b1000 +
#112160000000
0!
0'
#112170000000
1!
b1001 %
1'
b1001 +
#112180000000
0!
0'
#112190000000
1!
b0 %
1'
b0 +
#112200000000
0!
0'
#112210000000
1!
1$
b1 %
1'
1*
b1 +
#112220000000
0!
0'
#112230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#112240000000
0!
0'
#112250000000
1!
b11 %
1'
b11 +
#112260000000
0!
0'
#112270000000
1!
b100 %
1'
b100 +
#112280000000
0!
0'
#112290000000
1!
b101 %
1'
b101 +
#112300000000
0!
0'
#112310000000
1!
0$
b110 %
1'
0*
b110 +
#112320000000
0!
0'
#112330000000
1!
b111 %
1'
b111 +
#112340000000
0!
0'
#112350000000
1!
b1000 %
1'
b1000 +
#112360000000
0!
0'
#112370000000
1!
b1001 %
1'
b1001 +
#112380000000
0!
0'
#112390000000
1!
b0 %
1'
b0 +
#112400000000
0!
0'
#112410000000
1!
1$
b1 %
1'
1*
b1 +
#112420000000
0!
0'
#112430000000
1!
b10 %
1'
b10 +
#112440000000
1"
1(
#112450000000
0!
0"
b100 &
0'
0(
b100 ,
#112460000000
1!
b11 %
1'
b11 +
#112470000000
0!
0'
#112480000000
1!
b100 %
1'
b100 +
#112490000000
0!
0'
#112500000000
1!
b101 %
1'
b101 +
#112510000000
0!
0'
#112520000000
1!
b110 %
1'
b110 +
#112530000000
0!
0'
#112540000000
1!
b111 %
1'
b111 +
#112550000000
0!
0'
#112560000000
1!
0$
b1000 %
1'
0*
b1000 +
#112570000000
0!
0'
#112580000000
1!
b1001 %
1'
b1001 +
#112590000000
0!
0'
#112600000000
1!
b0 %
1'
b0 +
#112610000000
0!
0'
#112620000000
1!
1$
b1 %
1'
1*
b1 +
#112630000000
0!
0'
#112640000000
1!
b10 %
1'
b10 +
#112650000000
0!
0'
#112660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#112670000000
0!
0'
#112680000000
1!
b100 %
1'
b100 +
#112690000000
0!
0'
#112700000000
1!
b101 %
1'
b101 +
#112710000000
0!
0'
#112720000000
1!
0$
b110 %
1'
0*
b110 +
#112730000000
0!
0'
#112740000000
1!
b111 %
1'
b111 +
#112750000000
0!
0'
#112760000000
1!
b1000 %
1'
b1000 +
#112770000000
0!
0'
#112780000000
1!
b1001 %
1'
b1001 +
#112790000000
0!
0'
#112800000000
1!
b0 %
1'
b0 +
#112810000000
0!
0'
#112820000000
1!
1$
b1 %
1'
1*
b1 +
#112830000000
0!
0'
#112840000000
1!
b10 %
1'
b10 +
#112850000000
0!
0'
#112860000000
1!
b11 %
1'
b11 +
#112870000000
1"
1(
#112880000000
0!
0"
b100 &
0'
0(
b100 ,
#112890000000
1!
b100 %
1'
b100 +
#112900000000
0!
0'
#112910000000
1!
b101 %
1'
b101 +
#112920000000
0!
0'
#112930000000
1!
b110 %
1'
b110 +
#112940000000
0!
0'
#112950000000
1!
b111 %
1'
b111 +
#112960000000
0!
0'
#112970000000
1!
0$
b1000 %
1'
0*
b1000 +
#112980000000
0!
0'
#112990000000
1!
b1001 %
1'
b1001 +
#113000000000
0!
0'
#113010000000
1!
b0 %
1'
b0 +
#113020000000
0!
0'
#113030000000
1!
1$
b1 %
1'
1*
b1 +
#113040000000
0!
0'
#113050000000
1!
b10 %
1'
b10 +
#113060000000
0!
0'
#113070000000
1!
b11 %
1'
b11 +
#113080000000
0!
0'
#113090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#113100000000
0!
0'
#113110000000
1!
b101 %
1'
b101 +
#113120000000
0!
0'
#113130000000
1!
0$
b110 %
1'
0*
b110 +
#113140000000
0!
0'
#113150000000
1!
b111 %
1'
b111 +
#113160000000
0!
0'
#113170000000
1!
b1000 %
1'
b1000 +
#113180000000
0!
0'
#113190000000
1!
b1001 %
1'
b1001 +
#113200000000
0!
0'
#113210000000
1!
b0 %
1'
b0 +
#113220000000
0!
0'
#113230000000
1!
1$
b1 %
1'
1*
b1 +
#113240000000
0!
0'
#113250000000
1!
b10 %
1'
b10 +
#113260000000
0!
0'
#113270000000
1!
b11 %
1'
b11 +
#113280000000
0!
0'
#113290000000
1!
b100 %
1'
b100 +
#113300000000
1"
1(
#113310000000
0!
0"
b100 &
0'
0(
b100 ,
#113320000000
1!
b101 %
1'
b101 +
#113330000000
0!
0'
#113340000000
1!
b110 %
1'
b110 +
#113350000000
0!
0'
#113360000000
1!
b111 %
1'
b111 +
#113370000000
0!
0'
#113380000000
1!
0$
b1000 %
1'
0*
b1000 +
#113390000000
0!
0'
#113400000000
1!
b1001 %
1'
b1001 +
#113410000000
0!
0'
#113420000000
1!
b0 %
1'
b0 +
#113430000000
0!
0'
#113440000000
1!
1$
b1 %
1'
1*
b1 +
#113450000000
0!
0'
#113460000000
1!
b10 %
1'
b10 +
#113470000000
0!
0'
#113480000000
1!
b11 %
1'
b11 +
#113490000000
0!
0'
#113500000000
1!
b100 %
1'
b100 +
#113510000000
0!
0'
#113520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#113530000000
0!
0'
#113540000000
1!
0$
b110 %
1'
0*
b110 +
#113550000000
0!
0'
#113560000000
1!
b111 %
1'
b111 +
#113570000000
0!
0'
#113580000000
1!
b1000 %
1'
b1000 +
#113590000000
0!
0'
#113600000000
1!
b1001 %
1'
b1001 +
#113610000000
0!
0'
#113620000000
1!
b0 %
1'
b0 +
#113630000000
0!
0'
#113640000000
1!
1$
b1 %
1'
1*
b1 +
#113650000000
0!
0'
#113660000000
1!
b10 %
1'
b10 +
#113670000000
0!
0'
#113680000000
1!
b11 %
1'
b11 +
#113690000000
0!
0'
#113700000000
1!
b100 %
1'
b100 +
#113710000000
0!
0'
#113720000000
1!
b101 %
1'
b101 +
#113730000000
1"
1(
#113740000000
0!
0"
b100 &
0'
0(
b100 ,
#113750000000
1!
b110 %
1'
b110 +
#113760000000
0!
0'
#113770000000
1!
b111 %
1'
b111 +
#113780000000
0!
0'
#113790000000
1!
0$
b1000 %
1'
0*
b1000 +
#113800000000
0!
0'
#113810000000
1!
b1001 %
1'
b1001 +
#113820000000
0!
0'
#113830000000
1!
b0 %
1'
b0 +
#113840000000
0!
0'
#113850000000
1!
1$
b1 %
1'
1*
b1 +
#113860000000
0!
0'
#113870000000
1!
b10 %
1'
b10 +
#113880000000
0!
0'
#113890000000
1!
b11 %
1'
b11 +
#113900000000
0!
0'
#113910000000
1!
b100 %
1'
b100 +
#113920000000
0!
0'
#113930000000
1!
b101 %
1'
b101 +
#113940000000
0!
0'
#113950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#113960000000
0!
0'
#113970000000
1!
b111 %
1'
b111 +
#113980000000
0!
0'
#113990000000
1!
b1000 %
1'
b1000 +
#114000000000
0!
0'
#114010000000
1!
b1001 %
1'
b1001 +
#114020000000
0!
0'
#114030000000
1!
b0 %
1'
b0 +
#114040000000
0!
0'
#114050000000
1!
1$
b1 %
1'
1*
b1 +
#114060000000
0!
0'
#114070000000
1!
b10 %
1'
b10 +
#114080000000
0!
0'
#114090000000
1!
b11 %
1'
b11 +
#114100000000
0!
0'
#114110000000
1!
b100 %
1'
b100 +
#114120000000
0!
0'
#114130000000
1!
b101 %
1'
b101 +
#114140000000
0!
0'
#114150000000
1!
0$
b110 %
1'
0*
b110 +
#114160000000
1"
1(
#114170000000
0!
0"
b100 &
0'
0(
b100 ,
#114180000000
1!
1$
b111 %
1'
1*
b111 +
#114190000000
0!
0'
#114200000000
1!
0$
b1000 %
1'
0*
b1000 +
#114210000000
0!
0'
#114220000000
1!
b1001 %
1'
b1001 +
#114230000000
0!
0'
#114240000000
1!
b0 %
1'
b0 +
#114250000000
0!
0'
#114260000000
1!
1$
b1 %
1'
1*
b1 +
#114270000000
0!
0'
#114280000000
1!
b10 %
1'
b10 +
#114290000000
0!
0'
#114300000000
1!
b11 %
1'
b11 +
#114310000000
0!
0'
#114320000000
1!
b100 %
1'
b100 +
#114330000000
0!
0'
#114340000000
1!
b101 %
1'
b101 +
#114350000000
0!
0'
#114360000000
1!
b110 %
1'
b110 +
#114370000000
0!
0'
#114380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#114390000000
0!
0'
#114400000000
1!
b1000 %
1'
b1000 +
#114410000000
0!
0'
#114420000000
1!
b1001 %
1'
b1001 +
#114430000000
0!
0'
#114440000000
1!
b0 %
1'
b0 +
#114450000000
0!
0'
#114460000000
1!
1$
b1 %
1'
1*
b1 +
#114470000000
0!
0'
#114480000000
1!
b10 %
1'
b10 +
#114490000000
0!
0'
#114500000000
1!
b11 %
1'
b11 +
#114510000000
0!
0'
#114520000000
1!
b100 %
1'
b100 +
#114530000000
0!
0'
#114540000000
1!
b101 %
1'
b101 +
#114550000000
0!
0'
#114560000000
1!
0$
b110 %
1'
0*
b110 +
#114570000000
0!
0'
#114580000000
1!
b111 %
1'
b111 +
#114590000000
1"
1(
#114600000000
0!
0"
b100 &
0'
0(
b100 ,
#114610000000
1!
b1000 %
1'
b1000 +
#114620000000
0!
0'
#114630000000
1!
b1001 %
1'
b1001 +
#114640000000
0!
0'
#114650000000
1!
b0 %
1'
b0 +
#114660000000
0!
0'
#114670000000
1!
1$
b1 %
1'
1*
b1 +
#114680000000
0!
0'
#114690000000
1!
b10 %
1'
b10 +
#114700000000
0!
0'
#114710000000
1!
b11 %
1'
b11 +
#114720000000
0!
0'
#114730000000
1!
b100 %
1'
b100 +
#114740000000
0!
0'
#114750000000
1!
b101 %
1'
b101 +
#114760000000
0!
0'
#114770000000
1!
b110 %
1'
b110 +
#114780000000
0!
0'
#114790000000
1!
b111 %
1'
b111 +
#114800000000
0!
0'
#114810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#114820000000
0!
0'
#114830000000
1!
b1001 %
1'
b1001 +
#114840000000
0!
0'
#114850000000
1!
b0 %
1'
b0 +
#114860000000
0!
0'
#114870000000
1!
1$
b1 %
1'
1*
b1 +
#114880000000
0!
0'
#114890000000
1!
b10 %
1'
b10 +
#114900000000
0!
0'
#114910000000
1!
b11 %
1'
b11 +
#114920000000
0!
0'
#114930000000
1!
b100 %
1'
b100 +
#114940000000
0!
0'
#114950000000
1!
b101 %
1'
b101 +
#114960000000
0!
0'
#114970000000
1!
0$
b110 %
1'
0*
b110 +
#114980000000
0!
0'
#114990000000
1!
b111 %
1'
b111 +
#115000000000
0!
0'
#115010000000
1!
b1000 %
1'
b1000 +
#115020000000
1"
1(
#115030000000
0!
0"
b100 &
0'
0(
b100 ,
#115040000000
1!
b1001 %
1'
b1001 +
#115050000000
0!
0'
#115060000000
1!
b0 %
1'
b0 +
#115070000000
0!
0'
#115080000000
1!
1$
b1 %
1'
1*
b1 +
#115090000000
0!
0'
#115100000000
1!
b10 %
1'
b10 +
#115110000000
0!
0'
#115120000000
1!
b11 %
1'
b11 +
#115130000000
0!
0'
#115140000000
1!
b100 %
1'
b100 +
#115150000000
0!
0'
#115160000000
1!
b101 %
1'
b101 +
#115170000000
0!
0'
#115180000000
1!
b110 %
1'
b110 +
#115190000000
0!
0'
#115200000000
1!
b111 %
1'
b111 +
#115210000000
0!
0'
#115220000000
1!
0$
b1000 %
1'
0*
b1000 +
#115230000000
0!
0'
#115240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#115250000000
0!
0'
#115260000000
1!
b0 %
1'
b0 +
#115270000000
0!
0'
#115280000000
1!
1$
b1 %
1'
1*
b1 +
#115290000000
0!
0'
#115300000000
1!
b10 %
1'
b10 +
#115310000000
0!
0'
#115320000000
1!
b11 %
1'
b11 +
#115330000000
0!
0'
#115340000000
1!
b100 %
1'
b100 +
#115350000000
0!
0'
#115360000000
1!
b101 %
1'
b101 +
#115370000000
0!
0'
#115380000000
1!
0$
b110 %
1'
0*
b110 +
#115390000000
0!
0'
#115400000000
1!
b111 %
1'
b111 +
#115410000000
0!
0'
#115420000000
1!
b1000 %
1'
b1000 +
#115430000000
0!
0'
#115440000000
1!
b1001 %
1'
b1001 +
#115450000000
1"
1(
#115460000000
0!
0"
b100 &
0'
0(
b100 ,
#115470000000
1!
b0 %
1'
b0 +
#115480000000
0!
0'
#115490000000
1!
1$
b1 %
1'
1*
b1 +
#115500000000
0!
0'
#115510000000
1!
b10 %
1'
b10 +
#115520000000
0!
0'
#115530000000
1!
b11 %
1'
b11 +
#115540000000
0!
0'
#115550000000
1!
b100 %
1'
b100 +
#115560000000
0!
0'
#115570000000
1!
b101 %
1'
b101 +
#115580000000
0!
0'
#115590000000
1!
b110 %
1'
b110 +
#115600000000
0!
0'
#115610000000
1!
b111 %
1'
b111 +
#115620000000
0!
0'
#115630000000
1!
0$
b1000 %
1'
0*
b1000 +
#115640000000
0!
0'
#115650000000
1!
b1001 %
1'
b1001 +
#115660000000
0!
0'
#115670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#115680000000
0!
0'
#115690000000
1!
1$
b1 %
1'
1*
b1 +
#115700000000
0!
0'
#115710000000
1!
b10 %
1'
b10 +
#115720000000
0!
0'
#115730000000
1!
b11 %
1'
b11 +
#115740000000
0!
0'
#115750000000
1!
b100 %
1'
b100 +
#115760000000
0!
0'
#115770000000
1!
b101 %
1'
b101 +
#115780000000
0!
0'
#115790000000
1!
0$
b110 %
1'
0*
b110 +
#115800000000
0!
0'
#115810000000
1!
b111 %
1'
b111 +
#115820000000
0!
0'
#115830000000
1!
b1000 %
1'
b1000 +
#115840000000
0!
0'
#115850000000
1!
b1001 %
1'
b1001 +
#115860000000
0!
0'
#115870000000
1!
b0 %
1'
b0 +
#115880000000
1"
1(
#115890000000
0!
0"
b100 &
0'
0(
b100 ,
#115900000000
1!
1$
b1 %
1'
1*
b1 +
#115910000000
0!
0'
#115920000000
1!
b10 %
1'
b10 +
#115930000000
0!
0'
#115940000000
1!
b11 %
1'
b11 +
#115950000000
0!
0'
#115960000000
1!
b100 %
1'
b100 +
#115970000000
0!
0'
#115980000000
1!
b101 %
1'
b101 +
#115990000000
0!
0'
#116000000000
1!
b110 %
1'
b110 +
#116010000000
0!
0'
#116020000000
1!
b111 %
1'
b111 +
#116030000000
0!
0'
#116040000000
1!
0$
b1000 %
1'
0*
b1000 +
#116050000000
0!
0'
#116060000000
1!
b1001 %
1'
b1001 +
#116070000000
0!
0'
#116080000000
1!
b0 %
1'
b0 +
#116090000000
0!
0'
#116100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#116110000000
0!
0'
#116120000000
1!
b10 %
1'
b10 +
#116130000000
0!
0'
#116140000000
1!
b11 %
1'
b11 +
#116150000000
0!
0'
#116160000000
1!
b100 %
1'
b100 +
#116170000000
0!
0'
#116180000000
1!
b101 %
1'
b101 +
#116190000000
0!
0'
#116200000000
1!
0$
b110 %
1'
0*
b110 +
#116210000000
0!
0'
#116220000000
1!
b111 %
1'
b111 +
#116230000000
0!
0'
#116240000000
1!
b1000 %
1'
b1000 +
#116250000000
0!
0'
#116260000000
1!
b1001 %
1'
b1001 +
#116270000000
0!
0'
#116280000000
1!
b0 %
1'
b0 +
#116290000000
0!
0'
#116300000000
1!
1$
b1 %
1'
1*
b1 +
#116310000000
1"
1(
#116320000000
0!
0"
b100 &
0'
0(
b100 ,
#116330000000
1!
b10 %
1'
b10 +
#116340000000
0!
0'
#116350000000
1!
b11 %
1'
b11 +
#116360000000
0!
0'
#116370000000
1!
b100 %
1'
b100 +
#116380000000
0!
0'
#116390000000
1!
b101 %
1'
b101 +
#116400000000
0!
0'
#116410000000
1!
b110 %
1'
b110 +
#116420000000
0!
0'
#116430000000
1!
b111 %
1'
b111 +
#116440000000
0!
0'
#116450000000
1!
0$
b1000 %
1'
0*
b1000 +
#116460000000
0!
0'
#116470000000
1!
b1001 %
1'
b1001 +
#116480000000
0!
0'
#116490000000
1!
b0 %
1'
b0 +
#116500000000
0!
0'
#116510000000
1!
1$
b1 %
1'
1*
b1 +
#116520000000
0!
0'
#116530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#116540000000
0!
0'
#116550000000
1!
b11 %
1'
b11 +
#116560000000
0!
0'
#116570000000
1!
b100 %
1'
b100 +
#116580000000
0!
0'
#116590000000
1!
b101 %
1'
b101 +
#116600000000
0!
0'
#116610000000
1!
0$
b110 %
1'
0*
b110 +
#116620000000
0!
0'
#116630000000
1!
b111 %
1'
b111 +
#116640000000
0!
0'
#116650000000
1!
b1000 %
1'
b1000 +
#116660000000
0!
0'
#116670000000
1!
b1001 %
1'
b1001 +
#116680000000
0!
0'
#116690000000
1!
b0 %
1'
b0 +
#116700000000
0!
0'
#116710000000
1!
1$
b1 %
1'
1*
b1 +
#116720000000
0!
0'
#116730000000
1!
b10 %
1'
b10 +
#116740000000
1"
1(
#116750000000
0!
0"
b100 &
0'
0(
b100 ,
#116760000000
1!
b11 %
1'
b11 +
#116770000000
0!
0'
#116780000000
1!
b100 %
1'
b100 +
#116790000000
0!
0'
#116800000000
1!
b101 %
1'
b101 +
#116810000000
0!
0'
#116820000000
1!
b110 %
1'
b110 +
#116830000000
0!
0'
#116840000000
1!
b111 %
1'
b111 +
#116850000000
0!
0'
#116860000000
1!
0$
b1000 %
1'
0*
b1000 +
#116870000000
0!
0'
#116880000000
1!
b1001 %
1'
b1001 +
#116890000000
0!
0'
#116900000000
1!
b0 %
1'
b0 +
#116910000000
0!
0'
#116920000000
1!
1$
b1 %
1'
1*
b1 +
#116930000000
0!
0'
#116940000000
1!
b10 %
1'
b10 +
#116950000000
0!
0'
#116960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#116970000000
0!
0'
#116980000000
1!
b100 %
1'
b100 +
#116990000000
0!
0'
#117000000000
1!
b101 %
1'
b101 +
#117010000000
0!
0'
#117020000000
1!
0$
b110 %
1'
0*
b110 +
#117030000000
0!
0'
#117040000000
1!
b111 %
1'
b111 +
#117050000000
0!
0'
#117060000000
1!
b1000 %
1'
b1000 +
#117070000000
0!
0'
#117080000000
1!
b1001 %
1'
b1001 +
#117090000000
0!
0'
#117100000000
1!
b0 %
1'
b0 +
#117110000000
0!
0'
#117120000000
1!
1$
b1 %
1'
1*
b1 +
#117130000000
0!
0'
#117140000000
1!
b10 %
1'
b10 +
#117150000000
0!
0'
#117160000000
1!
b11 %
1'
b11 +
#117170000000
1"
1(
#117180000000
0!
0"
b100 &
0'
0(
b100 ,
#117190000000
1!
b100 %
1'
b100 +
#117200000000
0!
0'
#117210000000
1!
b101 %
1'
b101 +
#117220000000
0!
0'
#117230000000
1!
b110 %
1'
b110 +
#117240000000
0!
0'
#117250000000
1!
b111 %
1'
b111 +
#117260000000
0!
0'
#117270000000
1!
0$
b1000 %
1'
0*
b1000 +
#117280000000
0!
0'
#117290000000
1!
b1001 %
1'
b1001 +
#117300000000
0!
0'
#117310000000
1!
b0 %
1'
b0 +
#117320000000
0!
0'
#117330000000
1!
1$
b1 %
1'
1*
b1 +
#117340000000
0!
0'
#117350000000
1!
b10 %
1'
b10 +
#117360000000
0!
0'
#117370000000
1!
b11 %
1'
b11 +
#117380000000
0!
0'
#117390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#117400000000
0!
0'
#117410000000
1!
b101 %
1'
b101 +
#117420000000
0!
0'
#117430000000
1!
0$
b110 %
1'
0*
b110 +
#117440000000
0!
0'
#117450000000
1!
b111 %
1'
b111 +
#117460000000
0!
0'
#117470000000
1!
b1000 %
1'
b1000 +
#117480000000
0!
0'
#117490000000
1!
b1001 %
1'
b1001 +
#117500000000
0!
0'
#117510000000
1!
b0 %
1'
b0 +
#117520000000
0!
0'
#117530000000
1!
1$
b1 %
1'
1*
b1 +
#117540000000
0!
0'
#117550000000
1!
b10 %
1'
b10 +
#117560000000
0!
0'
#117570000000
1!
b11 %
1'
b11 +
#117580000000
0!
0'
#117590000000
1!
b100 %
1'
b100 +
#117600000000
1"
1(
#117610000000
0!
0"
b100 &
0'
0(
b100 ,
#117620000000
1!
b101 %
1'
b101 +
#117630000000
0!
0'
#117640000000
1!
b110 %
1'
b110 +
#117650000000
0!
0'
#117660000000
1!
b111 %
1'
b111 +
#117670000000
0!
0'
#117680000000
1!
0$
b1000 %
1'
0*
b1000 +
#117690000000
0!
0'
#117700000000
1!
b1001 %
1'
b1001 +
#117710000000
0!
0'
#117720000000
1!
b0 %
1'
b0 +
#117730000000
0!
0'
#117740000000
1!
1$
b1 %
1'
1*
b1 +
#117750000000
0!
0'
#117760000000
1!
b10 %
1'
b10 +
#117770000000
0!
0'
#117780000000
1!
b11 %
1'
b11 +
#117790000000
0!
0'
#117800000000
1!
b100 %
1'
b100 +
#117810000000
0!
0'
#117820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#117830000000
0!
0'
#117840000000
1!
0$
b110 %
1'
0*
b110 +
#117850000000
0!
0'
#117860000000
1!
b111 %
1'
b111 +
#117870000000
0!
0'
#117880000000
1!
b1000 %
1'
b1000 +
#117890000000
0!
0'
#117900000000
1!
b1001 %
1'
b1001 +
#117910000000
0!
0'
#117920000000
1!
b0 %
1'
b0 +
#117930000000
0!
0'
#117940000000
1!
1$
b1 %
1'
1*
b1 +
#117950000000
0!
0'
#117960000000
1!
b10 %
1'
b10 +
#117970000000
0!
0'
#117980000000
1!
b11 %
1'
b11 +
#117990000000
0!
0'
#118000000000
1!
b100 %
1'
b100 +
#118010000000
0!
0'
#118020000000
1!
b101 %
1'
b101 +
#118030000000
1"
1(
#118040000000
0!
0"
b100 &
0'
0(
b100 ,
#118050000000
1!
b110 %
1'
b110 +
#118060000000
0!
0'
#118070000000
1!
b111 %
1'
b111 +
#118080000000
0!
0'
#118090000000
1!
0$
b1000 %
1'
0*
b1000 +
#118100000000
0!
0'
#118110000000
1!
b1001 %
1'
b1001 +
#118120000000
0!
0'
#118130000000
1!
b0 %
1'
b0 +
#118140000000
0!
0'
#118150000000
1!
1$
b1 %
1'
1*
b1 +
#118160000000
0!
0'
#118170000000
1!
b10 %
1'
b10 +
#118180000000
0!
0'
#118190000000
1!
b11 %
1'
b11 +
#118200000000
0!
0'
#118210000000
1!
b100 %
1'
b100 +
#118220000000
0!
0'
#118230000000
1!
b101 %
1'
b101 +
#118240000000
0!
0'
#118250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#118260000000
0!
0'
#118270000000
1!
b111 %
1'
b111 +
#118280000000
0!
0'
#118290000000
1!
b1000 %
1'
b1000 +
#118300000000
0!
0'
#118310000000
1!
b1001 %
1'
b1001 +
#118320000000
0!
0'
#118330000000
1!
b0 %
1'
b0 +
#118340000000
0!
0'
#118350000000
1!
1$
b1 %
1'
1*
b1 +
#118360000000
0!
0'
#118370000000
1!
b10 %
1'
b10 +
#118380000000
0!
0'
#118390000000
1!
b11 %
1'
b11 +
#118400000000
0!
0'
#118410000000
1!
b100 %
1'
b100 +
#118420000000
0!
0'
#118430000000
1!
b101 %
1'
b101 +
#118440000000
0!
0'
#118450000000
1!
0$
b110 %
1'
0*
b110 +
#118460000000
1"
1(
#118470000000
0!
0"
b100 &
0'
0(
b100 ,
#118480000000
1!
1$
b111 %
1'
1*
b111 +
#118490000000
0!
0'
#118500000000
1!
0$
b1000 %
1'
0*
b1000 +
#118510000000
0!
0'
#118520000000
1!
b1001 %
1'
b1001 +
#118530000000
0!
0'
#118540000000
1!
b0 %
1'
b0 +
#118550000000
0!
0'
#118560000000
1!
1$
b1 %
1'
1*
b1 +
#118570000000
0!
0'
#118580000000
1!
b10 %
1'
b10 +
#118590000000
0!
0'
#118600000000
1!
b11 %
1'
b11 +
#118610000000
0!
0'
#118620000000
1!
b100 %
1'
b100 +
#118630000000
0!
0'
#118640000000
1!
b101 %
1'
b101 +
#118650000000
0!
0'
#118660000000
1!
b110 %
1'
b110 +
#118670000000
0!
0'
#118680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#118690000000
0!
0'
#118700000000
1!
b1000 %
1'
b1000 +
#118710000000
0!
0'
#118720000000
1!
b1001 %
1'
b1001 +
#118730000000
0!
0'
#118740000000
1!
b0 %
1'
b0 +
#118750000000
0!
0'
#118760000000
1!
1$
b1 %
1'
1*
b1 +
#118770000000
0!
0'
#118780000000
1!
b10 %
1'
b10 +
#118790000000
0!
0'
#118800000000
1!
b11 %
1'
b11 +
#118810000000
0!
0'
#118820000000
1!
b100 %
1'
b100 +
#118830000000
0!
0'
#118840000000
1!
b101 %
1'
b101 +
#118850000000
0!
0'
#118860000000
1!
0$
b110 %
1'
0*
b110 +
#118870000000
0!
0'
#118880000000
1!
b111 %
1'
b111 +
#118890000000
1"
1(
#118900000000
0!
0"
b100 &
0'
0(
b100 ,
#118910000000
1!
b1000 %
1'
b1000 +
#118920000000
0!
0'
#118930000000
1!
b1001 %
1'
b1001 +
#118940000000
0!
0'
#118950000000
1!
b0 %
1'
b0 +
#118960000000
0!
0'
#118970000000
1!
1$
b1 %
1'
1*
b1 +
#118980000000
0!
0'
#118990000000
1!
b10 %
1'
b10 +
#119000000000
0!
0'
#119010000000
1!
b11 %
1'
b11 +
#119020000000
0!
0'
#119030000000
1!
b100 %
1'
b100 +
#119040000000
0!
0'
#119050000000
1!
b101 %
1'
b101 +
#119060000000
0!
0'
#119070000000
1!
b110 %
1'
b110 +
#119080000000
0!
0'
#119090000000
1!
b111 %
1'
b111 +
#119100000000
0!
0'
#119110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#119120000000
0!
0'
#119130000000
1!
b1001 %
1'
b1001 +
#119140000000
0!
0'
#119150000000
1!
b0 %
1'
b0 +
#119160000000
0!
0'
#119170000000
1!
1$
b1 %
1'
1*
b1 +
#119180000000
0!
0'
#119190000000
1!
b10 %
1'
b10 +
#119200000000
0!
0'
#119210000000
1!
b11 %
1'
b11 +
#119220000000
0!
0'
#119230000000
1!
b100 %
1'
b100 +
#119240000000
0!
0'
#119250000000
1!
b101 %
1'
b101 +
#119260000000
0!
0'
#119270000000
1!
0$
b110 %
1'
0*
b110 +
#119280000000
0!
0'
#119290000000
1!
b111 %
1'
b111 +
#119300000000
0!
0'
#119310000000
1!
b1000 %
1'
b1000 +
#119320000000
1"
1(
#119330000000
0!
0"
b100 &
0'
0(
b100 ,
#119340000000
1!
b1001 %
1'
b1001 +
#119350000000
0!
0'
#119360000000
1!
b0 %
1'
b0 +
#119370000000
0!
0'
#119380000000
1!
1$
b1 %
1'
1*
b1 +
#119390000000
0!
0'
#119400000000
1!
b10 %
1'
b10 +
#119410000000
0!
0'
#119420000000
1!
b11 %
1'
b11 +
#119430000000
0!
0'
#119440000000
1!
b100 %
1'
b100 +
#119450000000
0!
0'
#119460000000
1!
b101 %
1'
b101 +
#119470000000
0!
0'
#119480000000
1!
b110 %
1'
b110 +
#119490000000
0!
0'
#119500000000
1!
b111 %
1'
b111 +
#119510000000
0!
0'
#119520000000
1!
0$
b1000 %
1'
0*
b1000 +
#119530000000
0!
0'
#119540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#119550000000
0!
0'
#119560000000
1!
b0 %
1'
b0 +
#119570000000
0!
0'
#119580000000
1!
1$
b1 %
1'
1*
b1 +
#119590000000
0!
0'
#119600000000
1!
b10 %
1'
b10 +
#119610000000
0!
0'
#119620000000
1!
b11 %
1'
b11 +
#119630000000
0!
0'
#119640000000
1!
b100 %
1'
b100 +
#119650000000
0!
0'
#119660000000
1!
b101 %
1'
b101 +
#119670000000
0!
0'
#119680000000
1!
0$
b110 %
1'
0*
b110 +
#119690000000
0!
0'
#119700000000
1!
b111 %
1'
b111 +
#119710000000
0!
0'
#119720000000
1!
b1000 %
1'
b1000 +
#119730000000
0!
0'
#119740000000
1!
b1001 %
1'
b1001 +
#119750000000
1"
1(
#119760000000
0!
0"
b100 &
0'
0(
b100 ,
#119770000000
1!
b0 %
1'
b0 +
#119780000000
0!
0'
#119790000000
1!
1$
b1 %
1'
1*
b1 +
#119800000000
0!
0'
#119810000000
1!
b10 %
1'
b10 +
#119820000000
0!
0'
#119830000000
1!
b11 %
1'
b11 +
#119840000000
0!
0'
#119850000000
1!
b100 %
1'
b100 +
#119860000000
0!
0'
#119870000000
1!
b101 %
1'
b101 +
#119880000000
0!
0'
#119890000000
1!
b110 %
1'
b110 +
#119900000000
0!
0'
#119910000000
1!
b111 %
1'
b111 +
#119920000000
0!
0'
#119930000000
1!
0$
b1000 %
1'
0*
b1000 +
#119940000000
0!
0'
#119950000000
1!
b1001 %
1'
b1001 +
#119960000000
0!
0'
#119970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#119980000000
0!
0'
#119990000000
1!
1$
b1 %
1'
1*
b1 +
#120000000000
0!
0'
#120010000000
1!
b10 %
1'
b10 +
#120020000000
0!
0'
#120030000000
1!
b11 %
1'
b11 +
#120040000000
0!
0'
#120050000000
1!
b100 %
1'
b100 +
#120060000000
0!
0'
#120070000000
1!
b101 %
1'
b101 +
#120080000000
0!
0'
#120090000000
1!
0$
b110 %
1'
0*
b110 +
#120100000000
0!
0'
#120110000000
1!
b111 %
1'
b111 +
#120120000000
0!
0'
#120130000000
1!
b1000 %
1'
b1000 +
#120140000000
0!
0'
#120150000000
1!
b1001 %
1'
b1001 +
#120160000000
0!
0'
#120170000000
1!
b0 %
1'
b0 +
#120180000000
1"
1(
#120190000000
0!
0"
b100 &
0'
0(
b100 ,
#120200000000
1!
1$
b1 %
1'
1*
b1 +
#120210000000
0!
0'
#120220000000
1!
b10 %
1'
b10 +
#120230000000
0!
0'
#120240000000
1!
b11 %
1'
b11 +
#120250000000
0!
0'
#120260000000
1!
b100 %
1'
b100 +
#120270000000
0!
0'
#120280000000
1!
b101 %
1'
b101 +
#120290000000
0!
0'
#120300000000
1!
b110 %
1'
b110 +
#120310000000
0!
0'
#120320000000
1!
b111 %
1'
b111 +
#120330000000
0!
0'
#120340000000
1!
0$
b1000 %
1'
0*
b1000 +
#120350000000
0!
0'
#120360000000
1!
b1001 %
1'
b1001 +
#120370000000
0!
0'
#120380000000
1!
b0 %
1'
b0 +
#120390000000
0!
0'
#120400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#120410000000
0!
0'
#120420000000
1!
b10 %
1'
b10 +
#120430000000
0!
0'
#120440000000
1!
b11 %
1'
b11 +
#120450000000
0!
0'
#120460000000
1!
b100 %
1'
b100 +
#120470000000
0!
0'
#120480000000
1!
b101 %
1'
b101 +
#120490000000
0!
0'
#120500000000
1!
0$
b110 %
1'
0*
b110 +
#120510000000
0!
0'
#120520000000
1!
b111 %
1'
b111 +
#120530000000
0!
0'
#120540000000
1!
b1000 %
1'
b1000 +
#120550000000
0!
0'
#120560000000
1!
b1001 %
1'
b1001 +
#120570000000
0!
0'
#120580000000
1!
b0 %
1'
b0 +
#120590000000
0!
0'
#120600000000
1!
1$
b1 %
1'
1*
b1 +
#120610000000
1"
1(
#120620000000
0!
0"
b100 &
0'
0(
b100 ,
#120630000000
1!
b10 %
1'
b10 +
#120640000000
0!
0'
#120650000000
1!
b11 %
1'
b11 +
#120660000000
0!
0'
#120670000000
1!
b100 %
1'
b100 +
#120680000000
0!
0'
#120690000000
1!
b101 %
1'
b101 +
#120700000000
0!
0'
#120710000000
1!
b110 %
1'
b110 +
#120720000000
0!
0'
#120730000000
1!
b111 %
1'
b111 +
#120740000000
0!
0'
#120750000000
1!
0$
b1000 %
1'
0*
b1000 +
#120760000000
0!
0'
#120770000000
1!
b1001 %
1'
b1001 +
#120780000000
0!
0'
#120790000000
1!
b0 %
1'
b0 +
#120800000000
0!
0'
#120810000000
1!
1$
b1 %
1'
1*
b1 +
#120820000000
0!
0'
#120830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#120840000000
0!
0'
#120850000000
1!
b11 %
1'
b11 +
#120860000000
0!
0'
#120870000000
1!
b100 %
1'
b100 +
#120880000000
0!
0'
#120890000000
1!
b101 %
1'
b101 +
#120900000000
0!
0'
#120910000000
1!
0$
b110 %
1'
0*
b110 +
#120920000000
0!
0'
#120930000000
1!
b111 %
1'
b111 +
#120940000000
0!
0'
#120950000000
1!
b1000 %
1'
b1000 +
#120960000000
0!
0'
#120970000000
1!
b1001 %
1'
b1001 +
#120980000000
0!
0'
#120990000000
1!
b0 %
1'
b0 +
#121000000000
0!
0'
#121010000000
1!
1$
b1 %
1'
1*
b1 +
#121020000000
0!
0'
#121030000000
1!
b10 %
1'
b10 +
#121040000000
1"
1(
#121050000000
0!
0"
b100 &
0'
0(
b100 ,
#121060000000
1!
b11 %
1'
b11 +
#121070000000
0!
0'
#121080000000
1!
b100 %
1'
b100 +
#121090000000
0!
0'
#121100000000
1!
b101 %
1'
b101 +
#121110000000
0!
0'
#121120000000
1!
b110 %
1'
b110 +
#121130000000
0!
0'
#121140000000
1!
b111 %
1'
b111 +
#121150000000
0!
0'
#121160000000
1!
0$
b1000 %
1'
0*
b1000 +
#121170000000
0!
0'
#121180000000
1!
b1001 %
1'
b1001 +
#121190000000
0!
0'
#121200000000
1!
b0 %
1'
b0 +
#121210000000
0!
0'
#121220000000
1!
1$
b1 %
1'
1*
b1 +
#121230000000
0!
0'
#121240000000
1!
b10 %
1'
b10 +
#121250000000
0!
0'
#121260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#121270000000
0!
0'
#121280000000
1!
b100 %
1'
b100 +
#121290000000
0!
0'
#121300000000
1!
b101 %
1'
b101 +
#121310000000
0!
0'
#121320000000
1!
0$
b110 %
1'
0*
b110 +
#121330000000
0!
0'
#121340000000
1!
b111 %
1'
b111 +
#121350000000
0!
0'
#121360000000
1!
b1000 %
1'
b1000 +
#121370000000
0!
0'
#121380000000
1!
b1001 %
1'
b1001 +
#121390000000
0!
0'
#121400000000
1!
b0 %
1'
b0 +
#121410000000
0!
0'
#121420000000
1!
1$
b1 %
1'
1*
b1 +
#121430000000
0!
0'
#121440000000
1!
b10 %
1'
b10 +
#121450000000
0!
0'
#121460000000
1!
b11 %
1'
b11 +
#121470000000
1"
1(
#121480000000
0!
0"
b100 &
0'
0(
b100 ,
#121490000000
1!
b100 %
1'
b100 +
#121500000000
0!
0'
#121510000000
1!
b101 %
1'
b101 +
#121520000000
0!
0'
#121530000000
1!
b110 %
1'
b110 +
#121540000000
0!
0'
#121550000000
1!
b111 %
1'
b111 +
#121560000000
0!
0'
#121570000000
1!
0$
b1000 %
1'
0*
b1000 +
#121580000000
0!
0'
#121590000000
1!
b1001 %
1'
b1001 +
#121600000000
0!
0'
#121610000000
1!
b0 %
1'
b0 +
#121620000000
0!
0'
#121630000000
1!
1$
b1 %
1'
1*
b1 +
#121640000000
0!
0'
#121650000000
1!
b10 %
1'
b10 +
#121660000000
0!
0'
#121670000000
1!
b11 %
1'
b11 +
#121680000000
0!
0'
#121690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#121700000000
0!
0'
#121710000000
1!
b101 %
1'
b101 +
#121720000000
0!
0'
#121730000000
1!
0$
b110 %
1'
0*
b110 +
#121740000000
0!
0'
#121750000000
1!
b111 %
1'
b111 +
#121760000000
0!
0'
#121770000000
1!
b1000 %
1'
b1000 +
#121780000000
0!
0'
#121790000000
1!
b1001 %
1'
b1001 +
#121800000000
0!
0'
#121810000000
1!
b0 %
1'
b0 +
#121820000000
0!
0'
#121830000000
1!
1$
b1 %
1'
1*
b1 +
#121840000000
0!
0'
#121850000000
1!
b10 %
1'
b10 +
#121860000000
0!
0'
#121870000000
1!
b11 %
1'
b11 +
#121880000000
0!
0'
#121890000000
1!
b100 %
1'
b100 +
#121900000000
1"
1(
#121910000000
0!
0"
b100 &
0'
0(
b100 ,
#121920000000
1!
b101 %
1'
b101 +
#121930000000
0!
0'
#121940000000
1!
b110 %
1'
b110 +
#121950000000
0!
0'
#121960000000
1!
b111 %
1'
b111 +
#121970000000
0!
0'
#121980000000
1!
0$
b1000 %
1'
0*
b1000 +
#121990000000
0!
0'
#122000000000
1!
b1001 %
1'
b1001 +
#122010000000
0!
0'
#122020000000
1!
b0 %
1'
b0 +
#122030000000
0!
0'
#122040000000
1!
1$
b1 %
1'
1*
b1 +
#122050000000
0!
0'
#122060000000
1!
b10 %
1'
b10 +
#122070000000
0!
0'
#122080000000
1!
b11 %
1'
b11 +
#122090000000
0!
0'
#122100000000
1!
b100 %
1'
b100 +
#122110000000
0!
0'
#122120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#122130000000
0!
0'
#122140000000
1!
0$
b110 %
1'
0*
b110 +
#122150000000
0!
0'
#122160000000
1!
b111 %
1'
b111 +
#122170000000
0!
0'
#122180000000
1!
b1000 %
1'
b1000 +
#122190000000
0!
0'
#122200000000
1!
b1001 %
1'
b1001 +
#122210000000
0!
0'
#122220000000
1!
b0 %
1'
b0 +
#122230000000
0!
0'
#122240000000
1!
1$
b1 %
1'
1*
b1 +
#122250000000
0!
0'
#122260000000
1!
b10 %
1'
b10 +
#122270000000
0!
0'
#122280000000
1!
b11 %
1'
b11 +
#122290000000
0!
0'
#122300000000
1!
b100 %
1'
b100 +
#122310000000
0!
0'
#122320000000
1!
b101 %
1'
b101 +
#122330000000
1"
1(
#122340000000
0!
0"
b100 &
0'
0(
b100 ,
#122350000000
1!
b110 %
1'
b110 +
#122360000000
0!
0'
#122370000000
1!
b111 %
1'
b111 +
#122380000000
0!
0'
#122390000000
1!
0$
b1000 %
1'
0*
b1000 +
#122400000000
0!
0'
#122410000000
1!
b1001 %
1'
b1001 +
#122420000000
0!
0'
#122430000000
1!
b0 %
1'
b0 +
#122440000000
0!
0'
#122450000000
1!
1$
b1 %
1'
1*
b1 +
#122460000000
0!
0'
#122470000000
1!
b10 %
1'
b10 +
#122480000000
0!
0'
#122490000000
1!
b11 %
1'
b11 +
#122500000000
0!
0'
#122510000000
1!
b100 %
1'
b100 +
#122520000000
0!
0'
#122530000000
1!
b101 %
1'
b101 +
#122540000000
0!
0'
#122550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#122560000000
0!
0'
#122570000000
1!
b111 %
1'
b111 +
#122580000000
0!
0'
#122590000000
1!
b1000 %
1'
b1000 +
#122600000000
0!
0'
#122610000000
1!
b1001 %
1'
b1001 +
#122620000000
0!
0'
#122630000000
1!
b0 %
1'
b0 +
#122640000000
0!
0'
#122650000000
1!
1$
b1 %
1'
1*
b1 +
#122660000000
0!
0'
#122670000000
1!
b10 %
1'
b10 +
#122680000000
0!
0'
#122690000000
1!
b11 %
1'
b11 +
#122700000000
0!
0'
#122710000000
1!
b100 %
1'
b100 +
#122720000000
0!
0'
#122730000000
1!
b101 %
1'
b101 +
#122740000000
0!
0'
#122750000000
1!
0$
b110 %
1'
0*
b110 +
#122760000000
1"
1(
#122770000000
0!
0"
b100 &
0'
0(
b100 ,
#122780000000
1!
1$
b111 %
1'
1*
b111 +
#122790000000
0!
0'
#122800000000
1!
0$
b1000 %
1'
0*
b1000 +
#122810000000
0!
0'
#122820000000
1!
b1001 %
1'
b1001 +
#122830000000
0!
0'
#122840000000
1!
b0 %
1'
b0 +
#122850000000
0!
0'
#122860000000
1!
1$
b1 %
1'
1*
b1 +
#122870000000
0!
0'
#122880000000
1!
b10 %
1'
b10 +
#122890000000
0!
0'
#122900000000
1!
b11 %
1'
b11 +
#122910000000
0!
0'
#122920000000
1!
b100 %
1'
b100 +
#122930000000
0!
0'
#122940000000
1!
b101 %
1'
b101 +
#122950000000
0!
0'
#122960000000
1!
b110 %
1'
b110 +
#122970000000
0!
0'
#122980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#122990000000
0!
0'
#123000000000
1!
b1000 %
1'
b1000 +
#123010000000
0!
0'
#123020000000
1!
b1001 %
1'
b1001 +
#123030000000
0!
0'
#123040000000
1!
b0 %
1'
b0 +
#123050000000
0!
0'
#123060000000
1!
1$
b1 %
1'
1*
b1 +
#123070000000
0!
0'
#123080000000
1!
b10 %
1'
b10 +
#123090000000
0!
0'
#123100000000
1!
b11 %
1'
b11 +
#123110000000
0!
0'
#123120000000
1!
b100 %
1'
b100 +
#123130000000
0!
0'
#123140000000
1!
b101 %
1'
b101 +
#123150000000
0!
0'
#123160000000
1!
0$
b110 %
1'
0*
b110 +
#123170000000
0!
0'
#123180000000
1!
b111 %
1'
b111 +
#123190000000
1"
1(
#123200000000
0!
0"
b100 &
0'
0(
b100 ,
#123210000000
1!
b1000 %
1'
b1000 +
#123220000000
0!
0'
#123230000000
1!
b1001 %
1'
b1001 +
#123240000000
0!
0'
#123250000000
1!
b0 %
1'
b0 +
#123260000000
0!
0'
#123270000000
1!
1$
b1 %
1'
1*
b1 +
#123280000000
0!
0'
#123290000000
1!
b10 %
1'
b10 +
#123300000000
0!
0'
#123310000000
1!
b11 %
1'
b11 +
#123320000000
0!
0'
#123330000000
1!
b100 %
1'
b100 +
#123340000000
0!
0'
#123350000000
1!
b101 %
1'
b101 +
#123360000000
0!
0'
#123370000000
1!
b110 %
1'
b110 +
#123380000000
0!
0'
#123390000000
1!
b111 %
1'
b111 +
#123400000000
0!
0'
#123410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#123420000000
0!
0'
#123430000000
1!
b1001 %
1'
b1001 +
#123440000000
0!
0'
#123450000000
1!
b0 %
1'
b0 +
#123460000000
0!
0'
#123470000000
1!
1$
b1 %
1'
1*
b1 +
#123480000000
0!
0'
#123490000000
1!
b10 %
1'
b10 +
#123500000000
0!
0'
#123510000000
1!
b11 %
1'
b11 +
#123520000000
0!
0'
#123530000000
1!
b100 %
1'
b100 +
#123540000000
0!
0'
#123550000000
1!
b101 %
1'
b101 +
#123560000000
0!
0'
#123570000000
1!
0$
b110 %
1'
0*
b110 +
#123580000000
0!
0'
#123590000000
1!
b111 %
1'
b111 +
#123600000000
0!
0'
#123610000000
1!
b1000 %
1'
b1000 +
#123620000000
1"
1(
#123630000000
0!
0"
b100 &
0'
0(
b100 ,
#123640000000
1!
b1001 %
1'
b1001 +
#123650000000
0!
0'
#123660000000
1!
b0 %
1'
b0 +
#123670000000
0!
0'
#123680000000
1!
1$
b1 %
1'
1*
b1 +
#123690000000
0!
0'
#123700000000
1!
b10 %
1'
b10 +
#123710000000
0!
0'
#123720000000
1!
b11 %
1'
b11 +
#123730000000
0!
0'
#123740000000
1!
b100 %
1'
b100 +
#123750000000
0!
0'
#123760000000
1!
b101 %
1'
b101 +
#123770000000
0!
0'
#123780000000
1!
b110 %
1'
b110 +
#123790000000
0!
0'
#123800000000
1!
b111 %
1'
b111 +
#123810000000
0!
0'
#123820000000
1!
0$
b1000 %
1'
0*
b1000 +
#123830000000
0!
0'
#123840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#123850000000
0!
0'
#123860000000
1!
b0 %
1'
b0 +
#123870000000
0!
0'
#123880000000
1!
1$
b1 %
1'
1*
b1 +
#123890000000
0!
0'
#123900000000
1!
b10 %
1'
b10 +
#123910000000
0!
0'
#123920000000
1!
b11 %
1'
b11 +
#123930000000
0!
0'
#123940000000
1!
b100 %
1'
b100 +
#123950000000
0!
0'
#123960000000
1!
b101 %
1'
b101 +
#123970000000
0!
0'
#123980000000
1!
0$
b110 %
1'
0*
b110 +
#123990000000
0!
0'
#124000000000
1!
b111 %
1'
b111 +
#124010000000
0!
0'
#124020000000
1!
b1000 %
1'
b1000 +
#124030000000
0!
0'
#124040000000
1!
b1001 %
1'
b1001 +
#124050000000
1"
1(
#124060000000
0!
0"
b100 &
0'
0(
b100 ,
#124070000000
1!
b0 %
1'
b0 +
#124080000000
0!
0'
#124090000000
1!
1$
b1 %
1'
1*
b1 +
#124100000000
0!
0'
#124110000000
1!
b10 %
1'
b10 +
#124120000000
0!
0'
#124130000000
1!
b11 %
1'
b11 +
#124140000000
0!
0'
#124150000000
1!
b100 %
1'
b100 +
#124160000000
0!
0'
#124170000000
1!
b101 %
1'
b101 +
#124180000000
0!
0'
#124190000000
1!
b110 %
1'
b110 +
#124200000000
0!
0'
#124210000000
1!
b111 %
1'
b111 +
#124220000000
0!
0'
#124230000000
1!
0$
b1000 %
1'
0*
b1000 +
#124240000000
0!
0'
#124250000000
1!
b1001 %
1'
b1001 +
#124260000000
0!
0'
#124270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#124280000000
0!
0'
#124290000000
1!
1$
b1 %
1'
1*
b1 +
#124300000000
0!
0'
#124310000000
1!
b10 %
1'
b10 +
#124320000000
0!
0'
#124330000000
1!
b11 %
1'
b11 +
#124340000000
0!
0'
#124350000000
1!
b100 %
1'
b100 +
#124360000000
0!
0'
#124370000000
1!
b101 %
1'
b101 +
#124380000000
0!
0'
#124390000000
1!
0$
b110 %
1'
0*
b110 +
#124400000000
0!
0'
#124410000000
1!
b111 %
1'
b111 +
#124420000000
0!
0'
#124430000000
1!
b1000 %
1'
b1000 +
#124440000000
0!
0'
#124450000000
1!
b1001 %
1'
b1001 +
#124460000000
0!
0'
#124470000000
1!
b0 %
1'
b0 +
#124480000000
1"
1(
#124490000000
0!
0"
b100 &
0'
0(
b100 ,
#124500000000
1!
1$
b1 %
1'
1*
b1 +
#124510000000
0!
0'
#124520000000
1!
b10 %
1'
b10 +
#124530000000
0!
0'
#124540000000
1!
b11 %
1'
b11 +
#124550000000
0!
0'
#124560000000
1!
b100 %
1'
b100 +
#124570000000
0!
0'
#124580000000
1!
b101 %
1'
b101 +
#124590000000
0!
0'
#124600000000
1!
b110 %
1'
b110 +
#124610000000
0!
0'
#124620000000
1!
b111 %
1'
b111 +
#124630000000
0!
0'
#124640000000
1!
0$
b1000 %
1'
0*
b1000 +
#124650000000
0!
0'
#124660000000
1!
b1001 %
1'
b1001 +
#124670000000
0!
0'
#124680000000
1!
b0 %
1'
b0 +
#124690000000
0!
0'
#124700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#124710000000
0!
0'
#124720000000
1!
b10 %
1'
b10 +
#124730000000
0!
0'
#124740000000
1!
b11 %
1'
b11 +
#124750000000
0!
0'
#124760000000
1!
b100 %
1'
b100 +
#124770000000
0!
0'
#124780000000
1!
b101 %
1'
b101 +
#124790000000
0!
0'
#124800000000
1!
0$
b110 %
1'
0*
b110 +
#124810000000
0!
0'
#124820000000
1!
b111 %
1'
b111 +
#124830000000
0!
0'
#124840000000
1!
b1000 %
1'
b1000 +
#124850000000
0!
0'
#124860000000
1!
b1001 %
1'
b1001 +
#124870000000
0!
0'
#124880000000
1!
b0 %
1'
b0 +
#124890000000
0!
0'
#124900000000
1!
1$
b1 %
1'
1*
b1 +
#124910000000
1"
1(
#124920000000
0!
0"
b100 &
0'
0(
b100 ,
#124930000000
1!
b10 %
1'
b10 +
#124940000000
0!
0'
#124950000000
1!
b11 %
1'
b11 +
#124960000000
0!
0'
#124970000000
1!
b100 %
1'
b100 +
#124980000000
0!
0'
#124990000000
1!
b101 %
1'
b101 +
#125000000000
0!
0'
#125010000000
1!
b110 %
1'
b110 +
#125020000000
0!
0'
#125030000000
1!
b111 %
1'
b111 +
#125040000000
0!
0'
#125050000000
1!
0$
b1000 %
1'
0*
b1000 +
#125060000000
0!
0'
#125070000000
1!
b1001 %
1'
b1001 +
#125080000000
0!
0'
#125090000000
1!
b0 %
1'
b0 +
#125100000000
0!
0'
#125110000000
1!
1$
b1 %
1'
1*
b1 +
#125120000000
0!
0'
#125130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#125140000000
0!
0'
#125150000000
1!
b11 %
1'
b11 +
#125160000000
0!
0'
#125170000000
1!
b100 %
1'
b100 +
#125180000000
0!
0'
#125190000000
1!
b101 %
1'
b101 +
#125200000000
0!
0'
#125210000000
1!
0$
b110 %
1'
0*
b110 +
#125220000000
0!
0'
#125230000000
1!
b111 %
1'
b111 +
#125240000000
0!
0'
#125250000000
1!
b1000 %
1'
b1000 +
#125260000000
0!
0'
#125270000000
1!
b1001 %
1'
b1001 +
#125280000000
0!
0'
#125290000000
1!
b0 %
1'
b0 +
#125300000000
0!
0'
#125310000000
1!
1$
b1 %
1'
1*
b1 +
#125320000000
0!
0'
#125330000000
1!
b10 %
1'
b10 +
#125340000000
1"
1(
#125350000000
0!
0"
b100 &
0'
0(
b100 ,
#125360000000
1!
b11 %
1'
b11 +
#125370000000
0!
0'
#125380000000
1!
b100 %
1'
b100 +
#125390000000
0!
0'
#125400000000
1!
b101 %
1'
b101 +
#125410000000
0!
0'
#125420000000
1!
b110 %
1'
b110 +
#125430000000
0!
0'
#125440000000
1!
b111 %
1'
b111 +
#125450000000
0!
0'
#125460000000
1!
0$
b1000 %
1'
0*
b1000 +
#125470000000
0!
0'
#125480000000
1!
b1001 %
1'
b1001 +
#125490000000
0!
0'
#125500000000
1!
b0 %
1'
b0 +
#125510000000
0!
0'
#125520000000
1!
1$
b1 %
1'
1*
b1 +
#125530000000
0!
0'
#125540000000
1!
b10 %
1'
b10 +
#125550000000
0!
0'
#125560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#125570000000
0!
0'
#125580000000
1!
b100 %
1'
b100 +
#125590000000
0!
0'
#125600000000
1!
b101 %
1'
b101 +
#125610000000
0!
0'
#125620000000
1!
0$
b110 %
1'
0*
b110 +
#125630000000
0!
0'
#125640000000
1!
b111 %
1'
b111 +
#125650000000
0!
0'
#125660000000
1!
b1000 %
1'
b1000 +
#125670000000
0!
0'
#125680000000
1!
b1001 %
1'
b1001 +
#125690000000
0!
0'
#125700000000
1!
b0 %
1'
b0 +
#125710000000
0!
0'
#125720000000
1!
1$
b1 %
1'
1*
b1 +
#125730000000
0!
0'
#125740000000
1!
b10 %
1'
b10 +
#125750000000
0!
0'
#125760000000
1!
b11 %
1'
b11 +
#125770000000
1"
1(
#125780000000
0!
0"
b100 &
0'
0(
b100 ,
#125790000000
1!
b100 %
1'
b100 +
#125800000000
0!
0'
#125810000000
1!
b101 %
1'
b101 +
#125820000000
0!
0'
#125830000000
1!
b110 %
1'
b110 +
#125840000000
0!
0'
#125850000000
1!
b111 %
1'
b111 +
#125860000000
0!
0'
#125870000000
1!
0$
b1000 %
1'
0*
b1000 +
#125880000000
0!
0'
#125890000000
1!
b1001 %
1'
b1001 +
#125900000000
0!
0'
#125910000000
1!
b0 %
1'
b0 +
#125920000000
0!
0'
#125930000000
1!
1$
b1 %
1'
1*
b1 +
#125940000000
0!
0'
#125950000000
1!
b10 %
1'
b10 +
#125960000000
0!
0'
#125970000000
1!
b11 %
1'
b11 +
#125980000000
0!
0'
#125990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#126000000000
0!
0'
#126010000000
1!
b101 %
1'
b101 +
#126020000000
0!
0'
#126030000000
1!
0$
b110 %
1'
0*
b110 +
#126040000000
0!
0'
#126050000000
1!
b111 %
1'
b111 +
#126060000000
0!
0'
#126070000000
1!
b1000 %
1'
b1000 +
#126080000000
0!
0'
#126090000000
1!
b1001 %
1'
b1001 +
#126100000000
0!
0'
#126110000000
1!
b0 %
1'
b0 +
#126120000000
0!
0'
#126130000000
1!
1$
b1 %
1'
1*
b1 +
#126140000000
0!
0'
#126150000000
1!
b10 %
1'
b10 +
#126160000000
0!
0'
#126170000000
1!
b11 %
1'
b11 +
#126180000000
0!
0'
#126190000000
1!
b100 %
1'
b100 +
#126200000000
1"
1(
#126210000000
0!
0"
b100 &
0'
0(
b100 ,
#126220000000
1!
b101 %
1'
b101 +
#126230000000
0!
0'
#126240000000
1!
b110 %
1'
b110 +
#126250000000
0!
0'
#126260000000
1!
b111 %
1'
b111 +
#126270000000
0!
0'
#126280000000
1!
0$
b1000 %
1'
0*
b1000 +
#126290000000
0!
0'
#126300000000
1!
b1001 %
1'
b1001 +
#126310000000
0!
0'
#126320000000
1!
b0 %
1'
b0 +
#126330000000
0!
0'
#126340000000
1!
1$
b1 %
1'
1*
b1 +
#126350000000
0!
0'
#126360000000
1!
b10 %
1'
b10 +
#126370000000
0!
0'
#126380000000
1!
b11 %
1'
b11 +
#126390000000
0!
0'
#126400000000
1!
b100 %
1'
b100 +
#126410000000
0!
0'
#126420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#126430000000
0!
0'
#126440000000
1!
0$
b110 %
1'
0*
b110 +
#126450000000
0!
0'
#126460000000
1!
b111 %
1'
b111 +
#126470000000
0!
0'
#126480000000
1!
b1000 %
1'
b1000 +
#126490000000
0!
0'
#126500000000
1!
b1001 %
1'
b1001 +
#126510000000
0!
0'
#126520000000
1!
b0 %
1'
b0 +
#126530000000
0!
0'
#126540000000
1!
1$
b1 %
1'
1*
b1 +
#126550000000
0!
0'
#126560000000
1!
b10 %
1'
b10 +
#126570000000
0!
0'
#126580000000
1!
b11 %
1'
b11 +
#126590000000
0!
0'
#126600000000
1!
b100 %
1'
b100 +
#126610000000
0!
0'
#126620000000
1!
b101 %
1'
b101 +
#126630000000
1"
1(
#126640000000
0!
0"
b100 &
0'
0(
b100 ,
#126650000000
1!
b110 %
1'
b110 +
#126660000000
0!
0'
#126670000000
1!
b111 %
1'
b111 +
#126680000000
0!
0'
#126690000000
1!
0$
b1000 %
1'
0*
b1000 +
#126700000000
0!
0'
#126710000000
1!
b1001 %
1'
b1001 +
#126720000000
0!
0'
#126730000000
1!
b0 %
1'
b0 +
#126740000000
0!
0'
#126750000000
1!
1$
b1 %
1'
1*
b1 +
#126760000000
0!
0'
#126770000000
1!
b10 %
1'
b10 +
#126780000000
0!
0'
#126790000000
1!
b11 %
1'
b11 +
#126800000000
0!
0'
#126810000000
1!
b100 %
1'
b100 +
#126820000000
0!
0'
#126830000000
1!
b101 %
1'
b101 +
#126840000000
0!
0'
#126850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#126860000000
0!
0'
#126870000000
1!
b111 %
1'
b111 +
#126880000000
0!
0'
#126890000000
1!
b1000 %
1'
b1000 +
#126900000000
0!
0'
#126910000000
1!
b1001 %
1'
b1001 +
#126920000000
0!
0'
#126930000000
1!
b0 %
1'
b0 +
#126940000000
0!
0'
#126950000000
1!
1$
b1 %
1'
1*
b1 +
#126960000000
0!
0'
#126970000000
1!
b10 %
1'
b10 +
#126980000000
0!
0'
#126990000000
1!
b11 %
1'
b11 +
#127000000000
0!
0'
#127010000000
1!
b100 %
1'
b100 +
#127020000000
0!
0'
#127030000000
1!
b101 %
1'
b101 +
#127040000000
0!
0'
#127050000000
1!
0$
b110 %
1'
0*
b110 +
#127060000000
1"
1(
#127070000000
0!
0"
b100 &
0'
0(
b100 ,
#127080000000
1!
1$
b111 %
1'
1*
b111 +
#127090000000
0!
0'
#127100000000
1!
0$
b1000 %
1'
0*
b1000 +
#127110000000
0!
0'
#127120000000
1!
b1001 %
1'
b1001 +
#127130000000
0!
0'
#127140000000
1!
b0 %
1'
b0 +
#127150000000
0!
0'
#127160000000
1!
1$
b1 %
1'
1*
b1 +
#127170000000
0!
0'
#127180000000
1!
b10 %
1'
b10 +
#127190000000
0!
0'
#127200000000
1!
b11 %
1'
b11 +
#127210000000
0!
0'
#127220000000
1!
b100 %
1'
b100 +
#127230000000
0!
0'
#127240000000
1!
b101 %
1'
b101 +
#127250000000
0!
0'
#127260000000
1!
b110 %
1'
b110 +
#127270000000
0!
0'
#127280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#127290000000
0!
0'
#127300000000
1!
b1000 %
1'
b1000 +
#127310000000
0!
0'
#127320000000
1!
b1001 %
1'
b1001 +
#127330000000
0!
0'
#127340000000
1!
b0 %
1'
b0 +
#127350000000
0!
0'
#127360000000
1!
1$
b1 %
1'
1*
b1 +
#127370000000
0!
0'
#127380000000
1!
b10 %
1'
b10 +
#127390000000
0!
0'
#127400000000
1!
b11 %
1'
b11 +
#127410000000
0!
0'
#127420000000
1!
b100 %
1'
b100 +
#127430000000
0!
0'
#127440000000
1!
b101 %
1'
b101 +
#127450000000
0!
0'
#127460000000
1!
0$
b110 %
1'
0*
b110 +
#127470000000
0!
0'
#127480000000
1!
b111 %
1'
b111 +
#127490000000
1"
1(
#127500000000
0!
0"
b100 &
0'
0(
b100 ,
#127510000000
1!
b1000 %
1'
b1000 +
#127520000000
0!
0'
#127530000000
1!
b1001 %
1'
b1001 +
#127540000000
0!
0'
#127550000000
1!
b0 %
1'
b0 +
#127560000000
0!
0'
#127570000000
1!
1$
b1 %
1'
1*
b1 +
#127580000000
0!
0'
#127590000000
1!
b10 %
1'
b10 +
#127600000000
0!
0'
#127610000000
1!
b11 %
1'
b11 +
#127620000000
0!
0'
#127630000000
1!
b100 %
1'
b100 +
#127640000000
0!
0'
#127650000000
1!
b101 %
1'
b101 +
#127660000000
0!
0'
#127670000000
1!
b110 %
1'
b110 +
#127680000000
0!
0'
#127690000000
1!
b111 %
1'
b111 +
#127700000000
0!
0'
#127710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#127720000000
0!
0'
#127730000000
1!
b1001 %
1'
b1001 +
#127740000000
0!
0'
#127750000000
1!
b0 %
1'
b0 +
#127760000000
0!
0'
#127770000000
1!
1$
b1 %
1'
1*
b1 +
#127780000000
0!
0'
#127790000000
1!
b10 %
1'
b10 +
#127800000000
0!
0'
#127810000000
1!
b11 %
1'
b11 +
#127820000000
0!
0'
#127830000000
1!
b100 %
1'
b100 +
#127840000000
0!
0'
#127850000000
1!
b101 %
1'
b101 +
#127860000000
0!
0'
#127870000000
1!
0$
b110 %
1'
0*
b110 +
#127880000000
0!
0'
#127890000000
1!
b111 %
1'
b111 +
#127900000000
0!
0'
#127910000000
1!
b1000 %
1'
b1000 +
#127920000000
1"
1(
#127930000000
0!
0"
b100 &
0'
0(
b100 ,
#127940000000
1!
b1001 %
1'
b1001 +
#127950000000
0!
0'
#127960000000
1!
b0 %
1'
b0 +
#127970000000
0!
0'
#127980000000
1!
1$
b1 %
1'
1*
b1 +
#127990000000
0!
0'
#128000000000
1!
b10 %
1'
b10 +
#128010000000
0!
0'
#128020000000
1!
b11 %
1'
b11 +
#128030000000
0!
0'
#128040000000
1!
b100 %
1'
b100 +
#128050000000
0!
0'
#128060000000
1!
b101 %
1'
b101 +
#128070000000
0!
0'
#128080000000
1!
b110 %
1'
b110 +
#128090000000
0!
0'
#128100000000
1!
b111 %
1'
b111 +
#128110000000
0!
0'
#128120000000
1!
0$
b1000 %
1'
0*
b1000 +
#128130000000
0!
0'
#128140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#128150000000
0!
0'
#128160000000
1!
b0 %
1'
b0 +
#128170000000
0!
0'
#128180000000
1!
1$
b1 %
1'
1*
b1 +
#128190000000
0!
0'
#128200000000
1!
b10 %
1'
b10 +
#128210000000
0!
0'
#128220000000
1!
b11 %
1'
b11 +
#128230000000
0!
0'
#128240000000
1!
b100 %
1'
b100 +
#128250000000
0!
0'
#128260000000
1!
b101 %
1'
b101 +
#128270000000
0!
0'
#128280000000
1!
0$
b110 %
1'
0*
b110 +
#128290000000
0!
0'
#128300000000
1!
b111 %
1'
b111 +
#128310000000
0!
0'
#128320000000
1!
b1000 %
1'
b1000 +
#128330000000
0!
0'
#128340000000
1!
b1001 %
1'
b1001 +
#128350000000
1"
1(
#128360000000
0!
0"
b100 &
0'
0(
b100 ,
#128370000000
1!
b0 %
1'
b0 +
#128380000000
0!
0'
#128390000000
1!
1$
b1 %
1'
1*
b1 +
#128400000000
0!
0'
#128410000000
1!
b10 %
1'
b10 +
#128420000000
0!
0'
#128430000000
1!
b11 %
1'
b11 +
#128440000000
0!
0'
#128450000000
1!
b100 %
1'
b100 +
#128460000000
0!
0'
#128470000000
1!
b101 %
1'
b101 +
#128480000000
0!
0'
#128490000000
1!
b110 %
1'
b110 +
#128500000000
0!
0'
#128510000000
1!
b111 %
1'
b111 +
#128520000000
0!
0'
#128530000000
1!
0$
b1000 %
1'
0*
b1000 +
#128540000000
0!
0'
#128550000000
1!
b1001 %
1'
b1001 +
#128560000000
0!
0'
#128570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#128580000000
0!
0'
#128590000000
1!
1$
b1 %
1'
1*
b1 +
#128600000000
0!
0'
#128610000000
1!
b10 %
1'
b10 +
#128620000000
0!
0'
#128630000000
1!
b11 %
1'
b11 +
#128640000000
0!
0'
#128650000000
1!
b100 %
1'
b100 +
#128660000000
0!
0'
#128670000000
1!
b101 %
1'
b101 +
#128680000000
0!
0'
#128690000000
1!
0$
b110 %
1'
0*
b110 +
#128700000000
0!
0'
#128710000000
1!
b111 %
1'
b111 +
#128720000000
0!
0'
#128730000000
1!
b1000 %
1'
b1000 +
#128740000000
0!
0'
#128750000000
1!
b1001 %
1'
b1001 +
#128760000000
0!
0'
#128770000000
1!
b0 %
1'
b0 +
#128780000000
1"
1(
#128790000000
0!
0"
b100 &
0'
0(
b100 ,
#128800000000
1!
1$
b1 %
1'
1*
b1 +
#128810000000
0!
0'
#128820000000
1!
b10 %
1'
b10 +
#128830000000
0!
0'
#128840000000
1!
b11 %
1'
b11 +
#128850000000
0!
0'
#128860000000
1!
b100 %
1'
b100 +
#128870000000
0!
0'
#128880000000
1!
b101 %
1'
b101 +
#128890000000
0!
0'
#128900000000
1!
b110 %
1'
b110 +
#128910000000
0!
0'
#128920000000
1!
b111 %
1'
b111 +
#128930000000
0!
0'
#128940000000
1!
0$
b1000 %
1'
0*
b1000 +
#128950000000
0!
0'
#128960000000
1!
b1001 %
1'
b1001 +
#128970000000
0!
0'
#128980000000
1!
b0 %
1'
b0 +
#128990000000
0!
0'
#129000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#129010000000
0!
0'
#129020000000
1!
b10 %
1'
b10 +
#129030000000
0!
0'
#129040000000
1!
b11 %
1'
b11 +
#129050000000
0!
0'
#129060000000
1!
b100 %
1'
b100 +
#129070000000
0!
0'
#129080000000
1!
b101 %
1'
b101 +
#129090000000
0!
0'
#129100000000
1!
0$
b110 %
1'
0*
b110 +
#129110000000
0!
0'
#129120000000
1!
b111 %
1'
b111 +
#129130000000
0!
0'
#129140000000
1!
b1000 %
1'
b1000 +
#129150000000
0!
0'
#129160000000
1!
b1001 %
1'
b1001 +
#129170000000
0!
0'
#129180000000
1!
b0 %
1'
b0 +
#129190000000
0!
0'
#129200000000
1!
1$
b1 %
1'
1*
b1 +
#129210000000
1"
1(
#129220000000
0!
0"
b100 &
0'
0(
b100 ,
#129230000000
1!
b10 %
1'
b10 +
#129240000000
0!
0'
#129250000000
1!
b11 %
1'
b11 +
#129260000000
0!
0'
#129270000000
1!
b100 %
1'
b100 +
#129280000000
0!
0'
#129290000000
1!
b101 %
1'
b101 +
#129300000000
0!
0'
#129310000000
1!
b110 %
1'
b110 +
#129320000000
0!
0'
#129330000000
1!
b111 %
1'
b111 +
#129340000000
0!
0'
#129350000000
1!
0$
b1000 %
1'
0*
b1000 +
#129360000000
0!
0'
#129370000000
1!
b1001 %
1'
b1001 +
#129380000000
0!
0'
#129390000000
1!
b0 %
1'
b0 +
#129400000000
0!
0'
#129410000000
1!
1$
b1 %
1'
1*
b1 +
#129420000000
0!
0'
#129430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#129440000000
0!
0'
#129450000000
1!
b11 %
1'
b11 +
#129460000000
0!
0'
#129470000000
1!
b100 %
1'
b100 +
#129480000000
0!
0'
#129490000000
1!
b101 %
1'
b101 +
#129500000000
0!
0'
#129510000000
1!
0$
b110 %
1'
0*
b110 +
#129520000000
0!
0'
#129530000000
1!
b111 %
1'
b111 +
#129540000000
0!
0'
#129550000000
1!
b1000 %
1'
b1000 +
#129560000000
0!
0'
#129570000000
1!
b1001 %
1'
b1001 +
#129580000000
0!
0'
#129590000000
1!
b0 %
1'
b0 +
#129600000000
0!
0'
#129610000000
1!
1$
b1 %
1'
1*
b1 +
#129620000000
0!
0'
#129630000000
1!
b10 %
1'
b10 +
#129640000000
1"
1(
#129650000000
0!
0"
b100 &
0'
0(
b100 ,
#129660000000
1!
b11 %
1'
b11 +
#129670000000
0!
0'
#129680000000
1!
b100 %
1'
b100 +
#129690000000
0!
0'
#129700000000
1!
b101 %
1'
b101 +
#129710000000
0!
0'
#129720000000
1!
b110 %
1'
b110 +
#129730000000
0!
0'
#129740000000
1!
b111 %
1'
b111 +
#129750000000
0!
0'
#129760000000
1!
0$
b1000 %
1'
0*
b1000 +
#129770000000
0!
0'
#129780000000
1!
b1001 %
1'
b1001 +
#129790000000
0!
0'
#129800000000
1!
b0 %
1'
b0 +
#129810000000
0!
0'
#129820000000
1!
1$
b1 %
1'
1*
b1 +
#129830000000
0!
0'
#129840000000
1!
b10 %
1'
b10 +
#129850000000
0!
0'
#129860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#129870000000
0!
0'
#129880000000
1!
b100 %
1'
b100 +
#129890000000
0!
0'
#129900000000
1!
b101 %
1'
b101 +
#129910000000
0!
0'
#129920000000
1!
0$
b110 %
1'
0*
b110 +
#129930000000
0!
0'
#129940000000
1!
b111 %
1'
b111 +
#129950000000
0!
0'
#129960000000
1!
b1000 %
1'
b1000 +
#129970000000
0!
0'
#129980000000
1!
b1001 %
1'
b1001 +
#129990000000
0!
0'
#130000000000
1!
b0 %
1'
b0 +
#130010000000
0!
0'
#130020000000
1!
1$
b1 %
1'
1*
b1 +
#130030000000
0!
0'
#130040000000
1!
b10 %
1'
b10 +
#130050000000
0!
0'
#130060000000
1!
b11 %
1'
b11 +
#130070000000
1"
1(
#130080000000
0!
0"
b100 &
0'
0(
b100 ,
#130090000000
1!
b100 %
1'
b100 +
#130100000000
0!
0'
#130110000000
1!
b101 %
1'
b101 +
#130120000000
0!
0'
#130130000000
1!
b110 %
1'
b110 +
#130140000000
0!
0'
#130150000000
1!
b111 %
1'
b111 +
#130160000000
0!
0'
#130170000000
1!
0$
b1000 %
1'
0*
b1000 +
#130180000000
0!
0'
#130190000000
1!
b1001 %
1'
b1001 +
#130200000000
0!
0'
#130210000000
1!
b0 %
1'
b0 +
#130220000000
0!
0'
#130230000000
1!
1$
b1 %
1'
1*
b1 +
#130240000000
0!
0'
#130250000000
1!
b10 %
1'
b10 +
#130260000000
0!
0'
#130270000000
1!
b11 %
1'
b11 +
#130280000000
0!
0'
#130290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#130300000000
0!
0'
#130310000000
1!
b101 %
1'
b101 +
#130320000000
0!
0'
#130330000000
1!
0$
b110 %
1'
0*
b110 +
#130340000000
0!
0'
#130350000000
1!
b111 %
1'
b111 +
#130360000000
0!
0'
#130370000000
1!
b1000 %
1'
b1000 +
#130380000000
0!
0'
#130390000000
1!
b1001 %
1'
b1001 +
#130400000000
0!
0'
#130410000000
1!
b0 %
1'
b0 +
#130420000000
0!
0'
#130430000000
1!
1$
b1 %
1'
1*
b1 +
#130440000000
0!
0'
#130450000000
1!
b10 %
1'
b10 +
#130460000000
0!
0'
#130470000000
1!
b11 %
1'
b11 +
#130480000000
0!
0'
#130490000000
1!
b100 %
1'
b100 +
#130500000000
1"
1(
#130510000000
0!
0"
b100 &
0'
0(
b100 ,
#130520000000
1!
b101 %
1'
b101 +
#130530000000
0!
0'
#130540000000
1!
b110 %
1'
b110 +
#130550000000
0!
0'
#130560000000
1!
b111 %
1'
b111 +
#130570000000
0!
0'
#130580000000
1!
0$
b1000 %
1'
0*
b1000 +
#130590000000
0!
0'
#130600000000
1!
b1001 %
1'
b1001 +
#130610000000
0!
0'
#130620000000
1!
b0 %
1'
b0 +
#130630000000
0!
0'
#130640000000
1!
1$
b1 %
1'
1*
b1 +
#130650000000
0!
0'
#130660000000
1!
b10 %
1'
b10 +
#130670000000
0!
0'
#130680000000
1!
b11 %
1'
b11 +
#130690000000
0!
0'
#130700000000
1!
b100 %
1'
b100 +
#130710000000
0!
0'
#130720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#130730000000
0!
0'
#130740000000
1!
0$
b110 %
1'
0*
b110 +
#130750000000
0!
0'
#130760000000
1!
b111 %
1'
b111 +
#130770000000
0!
0'
#130780000000
1!
b1000 %
1'
b1000 +
#130790000000
0!
0'
#130800000000
1!
b1001 %
1'
b1001 +
#130810000000
0!
0'
#130820000000
1!
b0 %
1'
b0 +
#130830000000
0!
0'
#130840000000
1!
1$
b1 %
1'
1*
b1 +
#130850000000
0!
0'
#130860000000
1!
b10 %
1'
b10 +
#130870000000
0!
0'
#130880000000
1!
b11 %
1'
b11 +
#130890000000
0!
0'
#130900000000
1!
b100 %
1'
b100 +
#130910000000
0!
0'
#130920000000
1!
b101 %
1'
b101 +
#130930000000
1"
1(
#130940000000
0!
0"
b100 &
0'
0(
b100 ,
#130950000000
1!
b110 %
1'
b110 +
#130960000000
0!
0'
#130970000000
1!
b111 %
1'
b111 +
#130980000000
0!
0'
#130990000000
1!
0$
b1000 %
1'
0*
b1000 +
#131000000000
0!
0'
#131010000000
1!
b1001 %
1'
b1001 +
#131020000000
0!
0'
#131030000000
1!
b0 %
1'
b0 +
#131040000000
0!
0'
#131050000000
1!
1$
b1 %
1'
1*
b1 +
#131060000000
0!
0'
#131070000000
1!
b10 %
1'
b10 +
#131080000000
0!
0'
#131090000000
1!
b11 %
1'
b11 +
#131100000000
0!
0'
#131110000000
1!
b100 %
1'
b100 +
#131120000000
0!
0'
#131130000000
1!
b101 %
1'
b101 +
#131140000000
0!
0'
#131150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#131160000000
0!
0'
#131170000000
1!
b111 %
1'
b111 +
#131180000000
0!
0'
#131190000000
1!
b1000 %
1'
b1000 +
#131200000000
0!
0'
#131210000000
1!
b1001 %
1'
b1001 +
#131220000000
0!
0'
#131230000000
1!
b0 %
1'
b0 +
#131240000000
0!
0'
#131250000000
1!
1$
b1 %
1'
1*
b1 +
#131260000000
0!
0'
#131270000000
1!
b10 %
1'
b10 +
#131280000000
0!
0'
#131290000000
1!
b11 %
1'
b11 +
#131300000000
0!
0'
#131310000000
1!
b100 %
1'
b100 +
#131320000000
0!
0'
#131330000000
1!
b101 %
1'
b101 +
#131340000000
0!
0'
#131350000000
1!
0$
b110 %
1'
0*
b110 +
#131360000000
1"
1(
#131370000000
0!
0"
b100 &
0'
0(
b100 ,
#131380000000
1!
1$
b111 %
1'
1*
b111 +
#131390000000
0!
0'
#131400000000
1!
0$
b1000 %
1'
0*
b1000 +
#131410000000
0!
0'
#131420000000
1!
b1001 %
1'
b1001 +
#131430000000
0!
0'
#131440000000
1!
b0 %
1'
b0 +
#131450000000
0!
0'
#131460000000
1!
1$
b1 %
1'
1*
b1 +
#131470000000
0!
0'
#131480000000
1!
b10 %
1'
b10 +
#131490000000
0!
0'
#131500000000
1!
b11 %
1'
b11 +
#131510000000
0!
0'
#131520000000
1!
b100 %
1'
b100 +
#131530000000
0!
0'
#131540000000
1!
b101 %
1'
b101 +
#131550000000
0!
0'
#131560000000
1!
b110 %
1'
b110 +
#131570000000
0!
0'
#131580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#131590000000
0!
0'
#131600000000
1!
b1000 %
1'
b1000 +
#131610000000
0!
0'
#131620000000
1!
b1001 %
1'
b1001 +
#131630000000
0!
0'
#131640000000
1!
b0 %
1'
b0 +
#131650000000
0!
0'
#131660000000
1!
1$
b1 %
1'
1*
b1 +
#131670000000
0!
0'
#131680000000
1!
b10 %
1'
b10 +
#131690000000
0!
0'
#131700000000
1!
b11 %
1'
b11 +
#131710000000
0!
0'
#131720000000
1!
b100 %
1'
b100 +
#131730000000
0!
0'
#131740000000
1!
b101 %
1'
b101 +
#131750000000
0!
0'
#131760000000
1!
0$
b110 %
1'
0*
b110 +
#131770000000
0!
0'
#131780000000
1!
b111 %
1'
b111 +
#131790000000
1"
1(
#131800000000
0!
0"
b100 &
0'
0(
b100 ,
#131810000000
1!
b1000 %
1'
b1000 +
#131820000000
0!
0'
#131830000000
1!
b1001 %
1'
b1001 +
#131840000000
0!
0'
#131850000000
1!
b0 %
1'
b0 +
#131860000000
0!
0'
#131870000000
1!
1$
b1 %
1'
1*
b1 +
#131880000000
0!
0'
#131890000000
1!
b10 %
1'
b10 +
#131900000000
0!
0'
#131910000000
1!
b11 %
1'
b11 +
#131920000000
0!
0'
#131930000000
1!
b100 %
1'
b100 +
#131940000000
0!
0'
#131950000000
1!
b101 %
1'
b101 +
#131960000000
0!
0'
#131970000000
1!
b110 %
1'
b110 +
#131980000000
0!
0'
#131990000000
1!
b111 %
1'
b111 +
#132000000000
0!
0'
#132010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#132020000000
0!
0'
#132030000000
1!
b1001 %
1'
b1001 +
#132040000000
0!
0'
#132050000000
1!
b0 %
1'
b0 +
#132060000000
0!
0'
#132070000000
1!
1$
b1 %
1'
1*
b1 +
#132080000000
0!
0'
#132090000000
1!
b10 %
1'
b10 +
#132100000000
0!
0'
#132110000000
1!
b11 %
1'
b11 +
#132120000000
0!
0'
#132130000000
1!
b100 %
1'
b100 +
#132140000000
0!
0'
#132150000000
1!
b101 %
1'
b101 +
#132160000000
0!
0'
#132170000000
1!
0$
b110 %
1'
0*
b110 +
#132180000000
0!
0'
#132190000000
1!
b111 %
1'
b111 +
#132200000000
0!
0'
#132210000000
1!
b1000 %
1'
b1000 +
#132220000000
1"
1(
#132230000000
0!
0"
b100 &
0'
0(
b100 ,
#132240000000
1!
b1001 %
1'
b1001 +
#132250000000
0!
0'
#132260000000
1!
b0 %
1'
b0 +
#132270000000
0!
0'
#132280000000
1!
1$
b1 %
1'
1*
b1 +
#132290000000
0!
0'
#132300000000
1!
b10 %
1'
b10 +
#132310000000
0!
0'
#132320000000
1!
b11 %
1'
b11 +
#132330000000
0!
0'
#132340000000
1!
b100 %
1'
b100 +
#132350000000
0!
0'
#132360000000
1!
b101 %
1'
b101 +
#132370000000
0!
0'
#132380000000
1!
b110 %
1'
b110 +
#132390000000
0!
0'
#132400000000
1!
b111 %
1'
b111 +
#132410000000
0!
0'
#132420000000
1!
0$
b1000 %
1'
0*
b1000 +
#132430000000
0!
0'
#132440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#132450000000
0!
0'
#132460000000
1!
b0 %
1'
b0 +
#132470000000
0!
0'
#132480000000
1!
1$
b1 %
1'
1*
b1 +
#132490000000
0!
0'
#132500000000
1!
b10 %
1'
b10 +
#132510000000
0!
0'
#132520000000
1!
b11 %
1'
b11 +
#132530000000
0!
0'
#132540000000
1!
b100 %
1'
b100 +
#132550000000
0!
0'
#132560000000
1!
b101 %
1'
b101 +
#132570000000
0!
0'
#132580000000
1!
0$
b110 %
1'
0*
b110 +
#132590000000
0!
0'
#132600000000
1!
b111 %
1'
b111 +
#132610000000
0!
0'
#132620000000
1!
b1000 %
1'
b1000 +
#132630000000
0!
0'
#132640000000
1!
b1001 %
1'
b1001 +
#132650000000
1"
1(
#132660000000
0!
0"
b100 &
0'
0(
b100 ,
#132670000000
1!
b0 %
1'
b0 +
#132680000000
0!
0'
#132690000000
1!
1$
b1 %
1'
1*
b1 +
#132700000000
0!
0'
#132710000000
1!
b10 %
1'
b10 +
#132720000000
0!
0'
#132730000000
1!
b11 %
1'
b11 +
#132740000000
0!
0'
#132750000000
1!
b100 %
1'
b100 +
#132760000000
0!
0'
#132770000000
1!
b101 %
1'
b101 +
#132780000000
0!
0'
#132790000000
1!
b110 %
1'
b110 +
#132800000000
0!
0'
#132810000000
1!
b111 %
1'
b111 +
#132820000000
0!
0'
#132830000000
1!
0$
b1000 %
1'
0*
b1000 +
#132840000000
0!
0'
#132850000000
1!
b1001 %
1'
b1001 +
#132860000000
0!
0'
#132870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#132880000000
0!
0'
#132890000000
1!
1$
b1 %
1'
1*
b1 +
#132900000000
0!
0'
#132910000000
1!
b10 %
1'
b10 +
#132920000000
0!
0'
#132930000000
1!
b11 %
1'
b11 +
#132940000000
0!
0'
#132950000000
1!
b100 %
1'
b100 +
#132960000000
0!
0'
#132970000000
1!
b101 %
1'
b101 +
#132980000000
0!
0'
#132990000000
1!
0$
b110 %
1'
0*
b110 +
#133000000000
0!
0'
#133010000000
1!
b111 %
1'
b111 +
#133020000000
0!
0'
#133030000000
1!
b1000 %
1'
b1000 +
#133040000000
0!
0'
#133050000000
1!
b1001 %
1'
b1001 +
#133060000000
0!
0'
#133070000000
1!
b0 %
1'
b0 +
#133080000000
1"
1(
#133090000000
0!
0"
b100 &
0'
0(
b100 ,
#133100000000
1!
1$
b1 %
1'
1*
b1 +
#133110000000
0!
0'
#133120000000
1!
b10 %
1'
b10 +
#133130000000
0!
0'
#133140000000
1!
b11 %
1'
b11 +
#133150000000
0!
0'
#133160000000
1!
b100 %
1'
b100 +
#133170000000
0!
0'
#133180000000
1!
b101 %
1'
b101 +
#133190000000
0!
0'
#133200000000
1!
b110 %
1'
b110 +
#133210000000
0!
0'
#133220000000
1!
b111 %
1'
b111 +
#133230000000
0!
0'
#133240000000
1!
0$
b1000 %
1'
0*
b1000 +
#133250000000
0!
0'
#133260000000
1!
b1001 %
1'
b1001 +
#133270000000
0!
0'
#133280000000
1!
b0 %
1'
b0 +
#133290000000
0!
0'
#133300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#133310000000
0!
0'
#133320000000
1!
b10 %
1'
b10 +
#133330000000
0!
0'
#133340000000
1!
b11 %
1'
b11 +
#133350000000
0!
0'
#133360000000
1!
b100 %
1'
b100 +
#133370000000
0!
0'
#133380000000
1!
b101 %
1'
b101 +
#133390000000
0!
0'
#133400000000
1!
0$
b110 %
1'
0*
b110 +
#133410000000
0!
0'
#133420000000
1!
b111 %
1'
b111 +
#133430000000
0!
0'
#133440000000
1!
b1000 %
1'
b1000 +
#133450000000
0!
0'
#133460000000
1!
b1001 %
1'
b1001 +
#133470000000
0!
0'
#133480000000
1!
b0 %
1'
b0 +
#133490000000
0!
0'
#133500000000
1!
1$
b1 %
1'
1*
b1 +
#133510000000
1"
1(
#133520000000
0!
0"
b100 &
0'
0(
b100 ,
#133530000000
1!
b10 %
1'
b10 +
#133540000000
0!
0'
#133550000000
1!
b11 %
1'
b11 +
#133560000000
0!
0'
#133570000000
1!
b100 %
1'
b100 +
#133580000000
0!
0'
#133590000000
1!
b101 %
1'
b101 +
#133600000000
0!
0'
#133610000000
1!
b110 %
1'
b110 +
#133620000000
0!
0'
#133630000000
1!
b111 %
1'
b111 +
#133640000000
0!
0'
#133650000000
1!
0$
b1000 %
1'
0*
b1000 +
#133660000000
0!
0'
#133670000000
1!
b1001 %
1'
b1001 +
#133680000000
0!
0'
#133690000000
1!
b0 %
1'
b0 +
#133700000000
0!
0'
#133710000000
1!
1$
b1 %
1'
1*
b1 +
#133720000000
0!
0'
#133730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#133740000000
0!
0'
#133750000000
1!
b11 %
1'
b11 +
#133760000000
0!
0'
#133770000000
1!
b100 %
1'
b100 +
#133780000000
0!
0'
#133790000000
1!
b101 %
1'
b101 +
#133800000000
0!
0'
#133810000000
1!
0$
b110 %
1'
0*
b110 +
#133820000000
0!
0'
#133830000000
1!
b111 %
1'
b111 +
#133840000000
0!
0'
#133850000000
1!
b1000 %
1'
b1000 +
#133860000000
0!
0'
#133870000000
1!
b1001 %
1'
b1001 +
#133880000000
0!
0'
#133890000000
1!
b0 %
1'
b0 +
#133900000000
0!
0'
#133910000000
1!
1$
b1 %
1'
1*
b1 +
#133920000000
0!
0'
#133930000000
1!
b10 %
1'
b10 +
#133940000000
1"
1(
#133950000000
0!
0"
b100 &
0'
0(
b100 ,
#133960000000
1!
b11 %
1'
b11 +
#133970000000
0!
0'
#133980000000
1!
b100 %
1'
b100 +
#133990000000
0!
0'
#134000000000
1!
b101 %
1'
b101 +
#134010000000
0!
0'
#134020000000
1!
b110 %
1'
b110 +
#134030000000
0!
0'
#134040000000
1!
b111 %
1'
b111 +
#134050000000
0!
0'
#134060000000
1!
0$
b1000 %
1'
0*
b1000 +
#134070000000
0!
0'
#134080000000
1!
b1001 %
1'
b1001 +
#134090000000
0!
0'
#134100000000
1!
b0 %
1'
b0 +
#134110000000
0!
0'
#134120000000
1!
1$
b1 %
1'
1*
b1 +
#134130000000
0!
0'
#134140000000
1!
b10 %
1'
b10 +
#134150000000
0!
0'
#134160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#134170000000
0!
0'
#134180000000
1!
b100 %
1'
b100 +
#134190000000
0!
0'
#134200000000
1!
b101 %
1'
b101 +
#134210000000
0!
0'
#134220000000
1!
0$
b110 %
1'
0*
b110 +
#134230000000
0!
0'
#134240000000
1!
b111 %
1'
b111 +
#134250000000
0!
0'
#134260000000
1!
b1000 %
1'
b1000 +
#134270000000
0!
0'
#134280000000
1!
b1001 %
1'
b1001 +
#134290000000
0!
0'
#134300000000
1!
b0 %
1'
b0 +
#134310000000
0!
0'
#134320000000
1!
1$
b1 %
1'
1*
b1 +
#134330000000
0!
0'
#134340000000
1!
b10 %
1'
b10 +
#134350000000
0!
0'
#134360000000
1!
b11 %
1'
b11 +
#134370000000
1"
1(
#134380000000
0!
0"
b100 &
0'
0(
b100 ,
#134390000000
1!
b100 %
1'
b100 +
#134400000000
0!
0'
#134410000000
1!
b101 %
1'
b101 +
#134420000000
0!
0'
#134430000000
1!
b110 %
1'
b110 +
#134440000000
0!
0'
#134450000000
1!
b111 %
1'
b111 +
#134460000000
0!
0'
#134470000000
1!
0$
b1000 %
1'
0*
b1000 +
#134480000000
0!
0'
#134490000000
1!
b1001 %
1'
b1001 +
#134500000000
0!
0'
#134510000000
1!
b0 %
1'
b0 +
#134520000000
0!
0'
#134530000000
1!
1$
b1 %
1'
1*
b1 +
#134540000000
0!
0'
#134550000000
1!
b10 %
1'
b10 +
#134560000000
0!
0'
#134570000000
1!
b11 %
1'
b11 +
#134580000000
0!
0'
#134590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#134600000000
0!
0'
#134610000000
1!
b101 %
1'
b101 +
#134620000000
0!
0'
#134630000000
1!
0$
b110 %
1'
0*
b110 +
#134640000000
0!
0'
#134650000000
1!
b111 %
1'
b111 +
#134660000000
0!
0'
#134670000000
1!
b1000 %
1'
b1000 +
#134680000000
0!
0'
#134690000000
1!
b1001 %
1'
b1001 +
#134700000000
0!
0'
#134710000000
1!
b0 %
1'
b0 +
#134720000000
0!
0'
#134730000000
1!
1$
b1 %
1'
1*
b1 +
#134740000000
0!
0'
#134750000000
1!
b10 %
1'
b10 +
#134760000000
0!
0'
#134770000000
1!
b11 %
1'
b11 +
#134780000000
0!
0'
#134790000000
1!
b100 %
1'
b100 +
#134800000000
1"
1(
#134810000000
0!
0"
b100 &
0'
0(
b100 ,
#134820000000
1!
b101 %
1'
b101 +
#134830000000
0!
0'
#134840000000
1!
b110 %
1'
b110 +
#134850000000
0!
0'
#134860000000
1!
b111 %
1'
b111 +
#134870000000
0!
0'
#134880000000
1!
0$
b1000 %
1'
0*
b1000 +
#134890000000
0!
0'
#134900000000
1!
b1001 %
1'
b1001 +
#134910000000
0!
0'
#134920000000
1!
b0 %
1'
b0 +
#134930000000
0!
0'
#134940000000
1!
1$
b1 %
1'
1*
b1 +
#134950000000
0!
0'
#134960000000
1!
b10 %
1'
b10 +
#134970000000
0!
0'
#134980000000
1!
b11 %
1'
b11 +
#134990000000
0!
0'
#135000000000
1!
b100 %
1'
b100 +
#135010000000
0!
0'
#135020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#135030000000
0!
0'
#135040000000
1!
0$
b110 %
1'
0*
b110 +
#135050000000
0!
0'
#135060000000
1!
b111 %
1'
b111 +
#135070000000
0!
0'
#135080000000
1!
b1000 %
1'
b1000 +
#135090000000
0!
0'
#135100000000
1!
b1001 %
1'
b1001 +
#135110000000
0!
0'
#135120000000
1!
b0 %
1'
b0 +
#135130000000
0!
0'
#135140000000
1!
1$
b1 %
1'
1*
b1 +
#135150000000
0!
0'
#135160000000
1!
b10 %
1'
b10 +
#135170000000
0!
0'
#135180000000
1!
b11 %
1'
b11 +
#135190000000
0!
0'
#135200000000
1!
b100 %
1'
b100 +
#135210000000
0!
0'
#135220000000
1!
b101 %
1'
b101 +
#135230000000
1"
1(
#135240000000
0!
0"
b100 &
0'
0(
b100 ,
#135250000000
1!
b110 %
1'
b110 +
#135260000000
0!
0'
#135270000000
1!
b111 %
1'
b111 +
#135280000000
0!
0'
#135290000000
1!
0$
b1000 %
1'
0*
b1000 +
#135300000000
0!
0'
#135310000000
1!
b1001 %
1'
b1001 +
#135320000000
0!
0'
#135330000000
1!
b0 %
1'
b0 +
#135340000000
0!
0'
#135350000000
1!
1$
b1 %
1'
1*
b1 +
#135360000000
0!
0'
#135370000000
1!
b10 %
1'
b10 +
#135380000000
0!
0'
#135390000000
1!
b11 %
1'
b11 +
#135400000000
0!
0'
#135410000000
1!
b100 %
1'
b100 +
#135420000000
0!
0'
#135430000000
1!
b101 %
1'
b101 +
#135440000000
0!
0'
#135450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#135460000000
0!
0'
#135470000000
1!
b111 %
1'
b111 +
#135480000000
0!
0'
#135490000000
1!
b1000 %
1'
b1000 +
#135500000000
0!
0'
#135510000000
1!
b1001 %
1'
b1001 +
#135520000000
0!
0'
#135530000000
1!
b0 %
1'
b0 +
#135540000000
0!
0'
#135550000000
1!
1$
b1 %
1'
1*
b1 +
#135560000000
0!
0'
#135570000000
1!
b10 %
1'
b10 +
#135580000000
0!
0'
#135590000000
1!
b11 %
1'
b11 +
#135600000000
0!
0'
#135610000000
1!
b100 %
1'
b100 +
#135620000000
0!
0'
#135630000000
1!
b101 %
1'
b101 +
#135640000000
0!
0'
#135650000000
1!
0$
b110 %
1'
0*
b110 +
#135660000000
1"
1(
#135670000000
0!
0"
b100 &
0'
0(
b100 ,
#135680000000
1!
1$
b111 %
1'
1*
b111 +
#135690000000
0!
0'
#135700000000
1!
0$
b1000 %
1'
0*
b1000 +
#135710000000
0!
0'
#135720000000
1!
b1001 %
1'
b1001 +
#135730000000
0!
0'
#135740000000
1!
b0 %
1'
b0 +
#135750000000
0!
0'
#135760000000
1!
1$
b1 %
1'
1*
b1 +
#135770000000
0!
0'
#135780000000
1!
b10 %
1'
b10 +
#135790000000
0!
0'
#135800000000
1!
b11 %
1'
b11 +
#135810000000
0!
0'
#135820000000
1!
b100 %
1'
b100 +
#135830000000
0!
0'
#135840000000
1!
b101 %
1'
b101 +
#135850000000
0!
0'
#135860000000
1!
b110 %
1'
b110 +
#135870000000
0!
0'
#135880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#135890000000
0!
0'
#135900000000
1!
b1000 %
1'
b1000 +
#135910000000
0!
0'
#135920000000
1!
b1001 %
1'
b1001 +
#135930000000
0!
0'
#135940000000
1!
b0 %
1'
b0 +
#135950000000
0!
0'
#135960000000
1!
1$
b1 %
1'
1*
b1 +
#135970000000
0!
0'
#135980000000
1!
b10 %
1'
b10 +
#135990000000
0!
0'
#136000000000
1!
b11 %
1'
b11 +
#136010000000
0!
0'
#136020000000
1!
b100 %
1'
b100 +
#136030000000
0!
0'
#136040000000
1!
b101 %
1'
b101 +
#136050000000
0!
0'
#136060000000
1!
0$
b110 %
1'
0*
b110 +
#136070000000
0!
0'
#136080000000
1!
b111 %
1'
b111 +
#136090000000
1"
1(
#136100000000
0!
0"
b100 &
0'
0(
b100 ,
#136110000000
1!
b1000 %
1'
b1000 +
#136120000000
0!
0'
#136130000000
1!
b1001 %
1'
b1001 +
#136140000000
0!
0'
#136150000000
1!
b0 %
1'
b0 +
#136160000000
0!
0'
#136170000000
1!
1$
b1 %
1'
1*
b1 +
#136180000000
0!
0'
#136190000000
1!
b10 %
1'
b10 +
#136200000000
0!
0'
#136210000000
1!
b11 %
1'
b11 +
#136220000000
0!
0'
#136230000000
1!
b100 %
1'
b100 +
#136240000000
0!
0'
#136250000000
1!
b101 %
1'
b101 +
#136260000000
0!
0'
#136270000000
1!
b110 %
1'
b110 +
#136280000000
0!
0'
#136290000000
1!
b111 %
1'
b111 +
#136300000000
0!
0'
#136310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#136320000000
0!
0'
#136330000000
1!
b1001 %
1'
b1001 +
#136340000000
0!
0'
#136350000000
1!
b0 %
1'
b0 +
#136360000000
0!
0'
#136370000000
1!
1$
b1 %
1'
1*
b1 +
#136380000000
0!
0'
#136390000000
1!
b10 %
1'
b10 +
#136400000000
0!
0'
#136410000000
1!
b11 %
1'
b11 +
#136420000000
0!
0'
#136430000000
1!
b100 %
1'
b100 +
#136440000000
0!
0'
#136450000000
1!
b101 %
1'
b101 +
#136460000000
0!
0'
#136470000000
1!
0$
b110 %
1'
0*
b110 +
#136480000000
0!
0'
#136490000000
1!
b111 %
1'
b111 +
#136500000000
0!
0'
#136510000000
1!
b1000 %
1'
b1000 +
#136520000000
1"
1(
#136530000000
0!
0"
b100 &
0'
0(
b100 ,
#136540000000
1!
b1001 %
1'
b1001 +
#136550000000
0!
0'
#136560000000
1!
b0 %
1'
b0 +
#136570000000
0!
0'
#136580000000
1!
1$
b1 %
1'
1*
b1 +
#136590000000
0!
0'
#136600000000
1!
b10 %
1'
b10 +
#136610000000
0!
0'
#136620000000
1!
b11 %
1'
b11 +
#136630000000
0!
0'
#136640000000
1!
b100 %
1'
b100 +
#136650000000
0!
0'
#136660000000
1!
b101 %
1'
b101 +
#136670000000
0!
0'
#136680000000
1!
b110 %
1'
b110 +
#136690000000
0!
0'
#136700000000
1!
b111 %
1'
b111 +
#136710000000
0!
0'
#136720000000
1!
0$
b1000 %
1'
0*
b1000 +
#136730000000
0!
0'
#136740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#136750000000
0!
0'
#136760000000
1!
b0 %
1'
b0 +
#136770000000
0!
0'
#136780000000
1!
1$
b1 %
1'
1*
b1 +
#136790000000
0!
0'
#136800000000
1!
b10 %
1'
b10 +
#136810000000
0!
0'
#136820000000
1!
b11 %
1'
b11 +
#136830000000
0!
0'
#136840000000
1!
b100 %
1'
b100 +
#136850000000
0!
0'
#136860000000
1!
b101 %
1'
b101 +
#136870000000
0!
0'
#136880000000
1!
0$
b110 %
1'
0*
b110 +
#136890000000
0!
0'
#136900000000
1!
b111 %
1'
b111 +
#136910000000
0!
0'
#136920000000
1!
b1000 %
1'
b1000 +
#136930000000
0!
0'
#136940000000
1!
b1001 %
1'
b1001 +
#136950000000
1"
1(
#136960000000
0!
0"
b100 &
0'
0(
b100 ,
#136970000000
1!
b0 %
1'
b0 +
#136980000000
0!
0'
#136990000000
1!
1$
b1 %
1'
1*
b1 +
#137000000000
0!
0'
#137010000000
1!
b10 %
1'
b10 +
#137020000000
0!
0'
#137030000000
1!
b11 %
1'
b11 +
#137040000000
0!
0'
#137050000000
1!
b100 %
1'
b100 +
#137060000000
0!
0'
#137070000000
1!
b101 %
1'
b101 +
#137080000000
0!
0'
#137090000000
1!
b110 %
1'
b110 +
#137100000000
0!
0'
#137110000000
1!
b111 %
1'
b111 +
#137120000000
0!
0'
#137130000000
1!
0$
b1000 %
1'
0*
b1000 +
#137140000000
0!
0'
#137150000000
1!
b1001 %
1'
b1001 +
#137160000000
0!
0'
#137170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#137180000000
0!
0'
#137190000000
1!
1$
b1 %
1'
1*
b1 +
#137200000000
0!
0'
#137210000000
1!
b10 %
1'
b10 +
#137220000000
0!
0'
#137230000000
1!
b11 %
1'
b11 +
#137240000000
0!
0'
#137250000000
1!
b100 %
1'
b100 +
#137260000000
0!
0'
#137270000000
1!
b101 %
1'
b101 +
#137280000000
0!
0'
#137290000000
1!
0$
b110 %
1'
0*
b110 +
#137300000000
0!
0'
#137310000000
1!
b111 %
1'
b111 +
#137320000000
0!
0'
#137330000000
1!
b1000 %
1'
b1000 +
#137340000000
0!
0'
#137350000000
1!
b1001 %
1'
b1001 +
#137360000000
0!
0'
#137370000000
1!
b0 %
1'
b0 +
#137380000000
1"
1(
#137390000000
0!
0"
b100 &
0'
0(
b100 ,
#137400000000
1!
1$
b1 %
1'
1*
b1 +
#137410000000
0!
0'
#137420000000
1!
b10 %
1'
b10 +
#137430000000
0!
0'
#137440000000
1!
b11 %
1'
b11 +
#137450000000
0!
0'
#137460000000
1!
b100 %
1'
b100 +
#137470000000
0!
0'
#137480000000
1!
b101 %
1'
b101 +
#137490000000
0!
0'
#137500000000
1!
b110 %
1'
b110 +
#137510000000
0!
0'
#137520000000
1!
b111 %
1'
b111 +
#137530000000
0!
0'
#137540000000
1!
0$
b1000 %
1'
0*
b1000 +
#137550000000
0!
0'
#137560000000
1!
b1001 %
1'
b1001 +
#137570000000
0!
0'
#137580000000
1!
b0 %
1'
b0 +
#137590000000
0!
0'
#137600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#137610000000
0!
0'
#137620000000
1!
b10 %
1'
b10 +
#137630000000
0!
0'
#137640000000
1!
b11 %
1'
b11 +
#137650000000
0!
0'
#137660000000
1!
b100 %
1'
b100 +
#137670000000
0!
0'
#137680000000
1!
b101 %
1'
b101 +
#137690000000
0!
0'
#137700000000
1!
0$
b110 %
1'
0*
b110 +
#137710000000
0!
0'
#137720000000
1!
b111 %
1'
b111 +
#137730000000
0!
0'
#137740000000
1!
b1000 %
1'
b1000 +
#137750000000
0!
0'
#137760000000
1!
b1001 %
1'
b1001 +
#137770000000
0!
0'
#137780000000
1!
b0 %
1'
b0 +
#137790000000
0!
0'
#137800000000
1!
1$
b1 %
1'
1*
b1 +
#137810000000
1"
1(
#137820000000
0!
0"
b100 &
0'
0(
b100 ,
#137830000000
1!
b10 %
1'
b10 +
#137840000000
0!
0'
#137850000000
1!
b11 %
1'
b11 +
#137860000000
0!
0'
#137870000000
1!
b100 %
1'
b100 +
#137880000000
0!
0'
#137890000000
1!
b101 %
1'
b101 +
#137900000000
0!
0'
#137910000000
1!
b110 %
1'
b110 +
#137920000000
0!
0'
#137930000000
1!
b111 %
1'
b111 +
#137940000000
0!
0'
#137950000000
1!
0$
b1000 %
1'
0*
b1000 +
#137960000000
0!
0'
#137970000000
1!
b1001 %
1'
b1001 +
#137980000000
0!
0'
#137990000000
1!
b0 %
1'
b0 +
#138000000000
0!
0'
#138010000000
1!
1$
b1 %
1'
1*
b1 +
#138020000000
0!
0'
#138030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#138040000000
0!
0'
#138050000000
1!
b11 %
1'
b11 +
#138060000000
0!
0'
#138070000000
1!
b100 %
1'
b100 +
#138080000000
0!
0'
#138090000000
1!
b101 %
1'
b101 +
#138100000000
0!
0'
#138110000000
1!
0$
b110 %
1'
0*
b110 +
#138120000000
0!
0'
#138130000000
1!
b111 %
1'
b111 +
#138140000000
0!
0'
#138150000000
1!
b1000 %
1'
b1000 +
#138160000000
0!
0'
#138170000000
1!
b1001 %
1'
b1001 +
#138180000000
0!
0'
#138190000000
1!
b0 %
1'
b0 +
#138200000000
0!
0'
#138210000000
1!
1$
b1 %
1'
1*
b1 +
#138220000000
0!
0'
#138230000000
1!
b10 %
1'
b10 +
#138240000000
1"
1(
#138250000000
0!
0"
b100 &
0'
0(
b100 ,
#138260000000
1!
b11 %
1'
b11 +
#138270000000
0!
0'
#138280000000
1!
b100 %
1'
b100 +
#138290000000
0!
0'
#138300000000
1!
b101 %
1'
b101 +
#138310000000
0!
0'
#138320000000
1!
b110 %
1'
b110 +
#138330000000
0!
0'
#138340000000
1!
b111 %
1'
b111 +
#138350000000
0!
0'
#138360000000
1!
0$
b1000 %
1'
0*
b1000 +
#138370000000
0!
0'
#138380000000
1!
b1001 %
1'
b1001 +
#138390000000
0!
0'
#138400000000
1!
b0 %
1'
b0 +
#138410000000
0!
0'
#138420000000
1!
1$
b1 %
1'
1*
b1 +
#138430000000
0!
0'
#138440000000
1!
b10 %
1'
b10 +
#138450000000
0!
0'
#138460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#138470000000
0!
0'
#138480000000
1!
b100 %
1'
b100 +
#138490000000
0!
0'
#138500000000
1!
b101 %
1'
b101 +
#138510000000
0!
0'
#138520000000
1!
0$
b110 %
1'
0*
b110 +
#138530000000
0!
0'
#138540000000
1!
b111 %
1'
b111 +
#138550000000
0!
0'
#138560000000
1!
b1000 %
1'
b1000 +
#138570000000
0!
0'
#138580000000
1!
b1001 %
1'
b1001 +
#138590000000
0!
0'
#138600000000
1!
b0 %
1'
b0 +
#138610000000
0!
0'
#138620000000
1!
1$
b1 %
1'
1*
b1 +
#138630000000
0!
0'
#138640000000
1!
b10 %
1'
b10 +
#138650000000
0!
0'
#138660000000
1!
b11 %
1'
b11 +
#138670000000
1"
1(
#138680000000
0!
0"
b100 &
0'
0(
b100 ,
#138690000000
1!
b100 %
1'
b100 +
#138700000000
0!
0'
#138710000000
1!
b101 %
1'
b101 +
#138720000000
0!
0'
#138730000000
1!
b110 %
1'
b110 +
#138740000000
0!
0'
#138750000000
1!
b111 %
1'
b111 +
#138760000000
0!
0'
#138770000000
1!
0$
b1000 %
1'
0*
b1000 +
#138780000000
0!
0'
#138790000000
1!
b1001 %
1'
b1001 +
#138800000000
0!
0'
#138810000000
1!
b0 %
1'
b0 +
#138820000000
0!
0'
#138830000000
1!
1$
b1 %
1'
1*
b1 +
#138840000000
0!
0'
#138850000000
1!
b10 %
1'
b10 +
#138860000000
0!
0'
#138870000000
1!
b11 %
1'
b11 +
#138880000000
0!
0'
#138890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#138900000000
0!
0'
#138910000000
1!
b101 %
1'
b101 +
#138920000000
0!
0'
#138930000000
1!
0$
b110 %
1'
0*
b110 +
#138940000000
0!
0'
#138950000000
1!
b111 %
1'
b111 +
#138960000000
0!
0'
#138970000000
1!
b1000 %
1'
b1000 +
#138980000000
0!
0'
#138990000000
1!
b1001 %
1'
b1001 +
#139000000000
0!
0'
#139010000000
1!
b0 %
1'
b0 +
#139020000000
0!
0'
#139030000000
1!
1$
b1 %
1'
1*
b1 +
#139040000000
0!
0'
#139050000000
1!
b10 %
1'
b10 +
#139060000000
0!
0'
#139070000000
1!
b11 %
1'
b11 +
#139080000000
0!
0'
#139090000000
1!
b100 %
1'
b100 +
#139100000000
1"
1(
#139110000000
0!
0"
b100 &
0'
0(
b100 ,
#139120000000
1!
b101 %
1'
b101 +
#139130000000
0!
0'
#139140000000
1!
b110 %
1'
b110 +
#139150000000
0!
0'
#139160000000
1!
b111 %
1'
b111 +
#139170000000
0!
0'
#139180000000
1!
0$
b1000 %
1'
0*
b1000 +
#139190000000
0!
0'
#139200000000
1!
b1001 %
1'
b1001 +
#139210000000
0!
0'
#139220000000
1!
b0 %
1'
b0 +
#139230000000
0!
0'
#139240000000
1!
1$
b1 %
1'
1*
b1 +
#139250000000
0!
0'
#139260000000
1!
b10 %
1'
b10 +
#139270000000
0!
0'
#139280000000
1!
b11 %
1'
b11 +
#139290000000
0!
0'
#139300000000
1!
b100 %
1'
b100 +
#139310000000
0!
0'
#139320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#139330000000
0!
0'
#139340000000
1!
0$
b110 %
1'
0*
b110 +
#139350000000
0!
0'
#139360000000
1!
b111 %
1'
b111 +
#139370000000
0!
0'
#139380000000
1!
b1000 %
1'
b1000 +
#139390000000
0!
0'
#139400000000
1!
b1001 %
1'
b1001 +
#139410000000
0!
0'
#139420000000
1!
b0 %
1'
b0 +
#139430000000
0!
0'
#139440000000
1!
1$
b1 %
1'
1*
b1 +
#139450000000
0!
0'
#139460000000
1!
b10 %
1'
b10 +
#139470000000
0!
0'
#139480000000
1!
b11 %
1'
b11 +
#139490000000
0!
0'
#139500000000
1!
b100 %
1'
b100 +
#139510000000
0!
0'
#139520000000
1!
b101 %
1'
b101 +
#139530000000
1"
1(
#139540000000
0!
0"
b100 &
0'
0(
b100 ,
#139550000000
1!
b110 %
1'
b110 +
#139560000000
0!
0'
#139570000000
1!
b111 %
1'
b111 +
#139580000000
0!
0'
#139590000000
1!
0$
b1000 %
1'
0*
b1000 +
#139600000000
0!
0'
#139610000000
1!
b1001 %
1'
b1001 +
#139620000000
0!
0'
#139630000000
1!
b0 %
1'
b0 +
#139640000000
0!
0'
#139650000000
1!
1$
b1 %
1'
1*
b1 +
#139660000000
0!
0'
#139670000000
1!
b10 %
1'
b10 +
#139680000000
0!
0'
#139690000000
1!
b11 %
1'
b11 +
#139700000000
0!
0'
#139710000000
1!
b100 %
1'
b100 +
#139720000000
0!
0'
#139730000000
1!
b101 %
1'
b101 +
#139740000000
0!
0'
#139750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#139760000000
0!
0'
#139770000000
1!
b111 %
1'
b111 +
#139780000000
0!
0'
#139790000000
1!
b1000 %
1'
b1000 +
#139800000000
0!
0'
#139810000000
1!
b1001 %
1'
b1001 +
#139820000000
0!
0'
#139830000000
1!
b0 %
1'
b0 +
#139840000000
0!
0'
#139850000000
1!
1$
b1 %
1'
1*
b1 +
#139860000000
0!
0'
#139870000000
1!
b10 %
1'
b10 +
#139880000000
0!
0'
#139890000000
1!
b11 %
1'
b11 +
#139900000000
0!
0'
#139910000000
1!
b100 %
1'
b100 +
#139920000000
0!
0'
#139930000000
1!
b101 %
1'
b101 +
#139940000000
0!
0'
#139950000000
1!
0$
b110 %
1'
0*
b110 +
#139960000000
1"
1(
#139970000000
0!
0"
b100 &
0'
0(
b100 ,
#139980000000
1!
1$
b111 %
1'
1*
b111 +
#139990000000
0!
0'
#140000000000
1!
0$
b1000 %
1'
0*
b1000 +
#140010000000
0!
0'
#140020000000
1!
b1001 %
1'
b1001 +
#140030000000
0!
0'
#140040000000
1!
b0 %
1'
b0 +
#140050000000
0!
0'
#140060000000
1!
1$
b1 %
1'
1*
b1 +
#140070000000
0!
0'
#140080000000
1!
b10 %
1'
b10 +
#140090000000
0!
0'
#140100000000
1!
b11 %
1'
b11 +
#140110000000
0!
0'
#140120000000
1!
b100 %
1'
b100 +
#140130000000
0!
0'
#140140000000
1!
b101 %
1'
b101 +
#140150000000
0!
0'
#140160000000
1!
b110 %
1'
b110 +
#140170000000
0!
0'
#140180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#140190000000
0!
0'
#140200000000
1!
b1000 %
1'
b1000 +
#140210000000
0!
0'
#140220000000
1!
b1001 %
1'
b1001 +
#140230000000
0!
0'
#140240000000
1!
b0 %
1'
b0 +
#140250000000
0!
0'
#140260000000
1!
1$
b1 %
1'
1*
b1 +
#140270000000
0!
0'
#140280000000
1!
b10 %
1'
b10 +
#140290000000
0!
0'
#140300000000
1!
b11 %
1'
b11 +
#140310000000
0!
0'
#140320000000
1!
b100 %
1'
b100 +
#140330000000
0!
0'
#140340000000
1!
b101 %
1'
b101 +
#140350000000
0!
0'
#140360000000
1!
0$
b110 %
1'
0*
b110 +
#140370000000
0!
0'
#140380000000
1!
b111 %
1'
b111 +
#140390000000
1"
1(
#140400000000
0!
0"
b100 &
0'
0(
b100 ,
#140410000000
1!
b1000 %
1'
b1000 +
#140420000000
0!
0'
#140430000000
1!
b1001 %
1'
b1001 +
#140440000000
0!
0'
#140450000000
1!
b0 %
1'
b0 +
#140460000000
0!
0'
#140470000000
1!
1$
b1 %
1'
1*
b1 +
#140480000000
0!
0'
#140490000000
1!
b10 %
1'
b10 +
#140500000000
0!
0'
#140510000000
1!
b11 %
1'
b11 +
#140520000000
0!
0'
#140530000000
1!
b100 %
1'
b100 +
#140540000000
0!
0'
#140550000000
1!
b101 %
1'
b101 +
#140560000000
0!
0'
#140570000000
1!
b110 %
1'
b110 +
#140580000000
0!
0'
#140590000000
1!
b111 %
1'
b111 +
#140600000000
0!
0'
#140610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#140620000000
0!
0'
#140630000000
1!
b1001 %
1'
b1001 +
#140640000000
0!
0'
#140650000000
1!
b0 %
1'
b0 +
#140660000000
0!
0'
#140670000000
1!
1$
b1 %
1'
1*
b1 +
#140680000000
0!
0'
#140690000000
1!
b10 %
1'
b10 +
#140700000000
0!
0'
#140710000000
1!
b11 %
1'
b11 +
#140720000000
0!
0'
#140730000000
1!
b100 %
1'
b100 +
#140740000000
0!
0'
#140750000000
1!
b101 %
1'
b101 +
#140760000000
0!
0'
#140770000000
1!
0$
b110 %
1'
0*
b110 +
#140780000000
0!
0'
#140790000000
1!
b111 %
1'
b111 +
#140800000000
0!
0'
#140810000000
1!
b1000 %
1'
b1000 +
#140820000000
1"
1(
#140830000000
0!
0"
b100 &
0'
0(
b100 ,
#140840000000
1!
b1001 %
1'
b1001 +
#140850000000
0!
0'
#140860000000
1!
b0 %
1'
b0 +
#140870000000
0!
0'
#140880000000
1!
1$
b1 %
1'
1*
b1 +
#140890000000
0!
0'
#140900000000
1!
b10 %
1'
b10 +
#140910000000
0!
0'
#140920000000
1!
b11 %
1'
b11 +
#140930000000
0!
0'
#140940000000
1!
b100 %
1'
b100 +
#140950000000
0!
0'
#140960000000
1!
b101 %
1'
b101 +
#140970000000
0!
0'
#140980000000
1!
b110 %
1'
b110 +
#140990000000
0!
0'
#141000000000
1!
b111 %
1'
b111 +
#141010000000
0!
0'
#141020000000
1!
0$
b1000 %
1'
0*
b1000 +
#141030000000
0!
0'
#141040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#141050000000
0!
0'
#141060000000
1!
b0 %
1'
b0 +
#141070000000
0!
0'
#141080000000
1!
1$
b1 %
1'
1*
b1 +
#141090000000
0!
0'
#141100000000
1!
b10 %
1'
b10 +
#141110000000
0!
0'
#141120000000
1!
b11 %
1'
b11 +
#141130000000
0!
0'
#141140000000
1!
b100 %
1'
b100 +
#141150000000
0!
0'
#141160000000
1!
b101 %
1'
b101 +
#141170000000
0!
0'
#141180000000
1!
0$
b110 %
1'
0*
b110 +
#141190000000
0!
0'
#141200000000
1!
b111 %
1'
b111 +
#141210000000
0!
0'
#141220000000
1!
b1000 %
1'
b1000 +
#141230000000
0!
0'
#141240000000
1!
b1001 %
1'
b1001 +
#141250000000
1"
1(
#141260000000
0!
0"
b100 &
0'
0(
b100 ,
#141270000000
1!
b0 %
1'
b0 +
#141280000000
0!
0'
#141290000000
1!
1$
b1 %
1'
1*
b1 +
#141300000000
0!
0'
#141310000000
1!
b10 %
1'
b10 +
#141320000000
0!
0'
#141330000000
1!
b11 %
1'
b11 +
#141340000000
0!
0'
#141350000000
1!
b100 %
1'
b100 +
#141360000000
0!
0'
#141370000000
1!
b101 %
1'
b101 +
#141380000000
0!
0'
#141390000000
1!
b110 %
1'
b110 +
#141400000000
0!
0'
#141410000000
1!
b111 %
1'
b111 +
#141420000000
0!
0'
#141430000000
1!
0$
b1000 %
1'
0*
b1000 +
#141440000000
0!
0'
#141450000000
1!
b1001 %
1'
b1001 +
#141460000000
0!
0'
#141470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#141480000000
0!
0'
#141490000000
1!
1$
b1 %
1'
1*
b1 +
#141500000000
0!
0'
#141510000000
1!
b10 %
1'
b10 +
#141520000000
0!
0'
#141530000000
1!
b11 %
1'
b11 +
#141540000000
0!
0'
#141550000000
1!
b100 %
1'
b100 +
#141560000000
0!
0'
#141570000000
1!
b101 %
1'
b101 +
#141580000000
0!
0'
#141590000000
1!
0$
b110 %
1'
0*
b110 +
#141600000000
0!
0'
#141610000000
1!
b111 %
1'
b111 +
#141620000000
0!
0'
#141630000000
1!
b1000 %
1'
b1000 +
#141640000000
0!
0'
#141650000000
1!
b1001 %
1'
b1001 +
#141660000000
0!
0'
#141670000000
1!
b0 %
1'
b0 +
#141680000000
1"
1(
#141690000000
0!
0"
b100 &
0'
0(
b100 ,
#141700000000
1!
1$
b1 %
1'
1*
b1 +
#141710000000
0!
0'
#141720000000
1!
b10 %
1'
b10 +
#141730000000
0!
0'
#141740000000
1!
b11 %
1'
b11 +
#141750000000
0!
0'
#141760000000
1!
b100 %
1'
b100 +
#141770000000
0!
0'
#141780000000
1!
b101 %
1'
b101 +
#141790000000
0!
0'
#141800000000
1!
b110 %
1'
b110 +
#141810000000
0!
0'
#141820000000
1!
b111 %
1'
b111 +
#141830000000
0!
0'
#141840000000
1!
0$
b1000 %
1'
0*
b1000 +
#141850000000
0!
0'
#141860000000
1!
b1001 %
1'
b1001 +
#141870000000
0!
0'
#141880000000
1!
b0 %
1'
b0 +
#141890000000
0!
0'
#141900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#141910000000
0!
0'
#141920000000
1!
b10 %
1'
b10 +
#141930000000
0!
0'
#141940000000
1!
b11 %
1'
b11 +
#141950000000
0!
0'
#141960000000
1!
b100 %
1'
b100 +
#141970000000
0!
0'
#141980000000
1!
b101 %
1'
b101 +
#141990000000
0!
0'
#142000000000
1!
0$
b110 %
1'
0*
b110 +
#142010000000
0!
0'
#142020000000
1!
b111 %
1'
b111 +
#142030000000
0!
0'
#142040000000
1!
b1000 %
1'
b1000 +
#142050000000
0!
0'
#142060000000
1!
b1001 %
1'
b1001 +
#142070000000
0!
0'
#142080000000
1!
b0 %
1'
b0 +
#142090000000
0!
0'
#142100000000
1!
1$
b1 %
1'
1*
b1 +
#142110000000
1"
1(
#142120000000
0!
0"
b100 &
0'
0(
b100 ,
#142130000000
1!
b10 %
1'
b10 +
#142140000000
0!
0'
#142150000000
1!
b11 %
1'
b11 +
#142160000000
0!
0'
#142170000000
1!
b100 %
1'
b100 +
#142180000000
0!
0'
#142190000000
1!
b101 %
1'
b101 +
#142200000000
0!
0'
#142210000000
1!
b110 %
1'
b110 +
#142220000000
0!
0'
#142230000000
1!
b111 %
1'
b111 +
#142240000000
0!
0'
#142250000000
1!
0$
b1000 %
1'
0*
b1000 +
#142260000000
0!
0'
#142270000000
1!
b1001 %
1'
b1001 +
#142280000000
0!
0'
#142290000000
1!
b0 %
1'
b0 +
#142300000000
0!
0'
#142310000000
1!
1$
b1 %
1'
1*
b1 +
#142320000000
0!
0'
#142330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#142340000000
0!
0'
#142350000000
1!
b11 %
1'
b11 +
#142360000000
0!
0'
#142370000000
1!
b100 %
1'
b100 +
#142380000000
0!
0'
#142390000000
1!
b101 %
1'
b101 +
#142400000000
0!
0'
#142410000000
1!
0$
b110 %
1'
0*
b110 +
#142420000000
0!
0'
#142430000000
1!
b111 %
1'
b111 +
#142440000000
0!
0'
#142450000000
1!
b1000 %
1'
b1000 +
#142460000000
0!
0'
#142470000000
1!
b1001 %
1'
b1001 +
#142480000000
0!
0'
#142490000000
1!
b0 %
1'
b0 +
#142500000000
0!
0'
#142510000000
1!
1$
b1 %
1'
1*
b1 +
#142520000000
0!
0'
#142530000000
1!
b10 %
1'
b10 +
#142540000000
1"
1(
#142550000000
0!
0"
b100 &
0'
0(
b100 ,
#142560000000
1!
b11 %
1'
b11 +
#142570000000
0!
0'
#142580000000
1!
b100 %
1'
b100 +
#142590000000
0!
0'
#142600000000
1!
b101 %
1'
b101 +
#142610000000
0!
0'
#142620000000
1!
b110 %
1'
b110 +
#142630000000
0!
0'
#142640000000
1!
b111 %
1'
b111 +
#142650000000
0!
0'
#142660000000
1!
0$
b1000 %
1'
0*
b1000 +
#142670000000
0!
0'
#142680000000
1!
b1001 %
1'
b1001 +
#142690000000
0!
0'
#142700000000
1!
b0 %
1'
b0 +
#142710000000
0!
0'
#142720000000
1!
1$
b1 %
1'
1*
b1 +
#142730000000
0!
0'
#142740000000
1!
b10 %
1'
b10 +
#142750000000
0!
0'
#142760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#142770000000
0!
0'
#142780000000
1!
b100 %
1'
b100 +
#142790000000
0!
0'
#142800000000
1!
b101 %
1'
b101 +
#142810000000
0!
0'
#142820000000
1!
0$
b110 %
1'
0*
b110 +
#142830000000
0!
0'
#142840000000
1!
b111 %
1'
b111 +
#142850000000
0!
0'
#142860000000
1!
b1000 %
1'
b1000 +
#142870000000
0!
0'
#142880000000
1!
b1001 %
1'
b1001 +
#142890000000
0!
0'
#142900000000
1!
b0 %
1'
b0 +
#142910000000
0!
0'
#142920000000
1!
1$
b1 %
1'
1*
b1 +
#142930000000
0!
0'
#142940000000
1!
b10 %
1'
b10 +
#142950000000
0!
0'
#142960000000
1!
b11 %
1'
b11 +
#142970000000
1"
1(
#142980000000
0!
0"
b100 &
0'
0(
b100 ,
#142990000000
1!
b100 %
1'
b100 +
#143000000000
0!
0'
#143010000000
1!
b101 %
1'
b101 +
#143020000000
0!
0'
#143030000000
1!
b110 %
1'
b110 +
#143040000000
0!
0'
#143050000000
1!
b111 %
1'
b111 +
#143060000000
0!
0'
#143070000000
1!
0$
b1000 %
1'
0*
b1000 +
#143080000000
0!
0'
#143090000000
1!
b1001 %
1'
b1001 +
#143100000000
0!
0'
#143110000000
1!
b0 %
1'
b0 +
#143120000000
0!
0'
#143130000000
1!
1$
b1 %
1'
1*
b1 +
#143140000000
0!
0'
#143150000000
1!
b10 %
1'
b10 +
#143160000000
0!
0'
#143170000000
1!
b11 %
1'
b11 +
#143180000000
0!
0'
#143190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#143200000000
0!
0'
#143210000000
1!
b101 %
1'
b101 +
#143220000000
0!
0'
#143230000000
1!
0$
b110 %
1'
0*
b110 +
#143240000000
0!
0'
#143250000000
1!
b111 %
1'
b111 +
#143260000000
0!
0'
#143270000000
1!
b1000 %
1'
b1000 +
#143280000000
0!
0'
#143290000000
1!
b1001 %
1'
b1001 +
#143300000000
0!
0'
#143310000000
1!
b0 %
1'
b0 +
#143320000000
0!
0'
#143330000000
1!
1$
b1 %
1'
1*
b1 +
#143340000000
0!
0'
#143350000000
1!
b10 %
1'
b10 +
#143360000000
0!
0'
#143370000000
1!
b11 %
1'
b11 +
#143380000000
0!
0'
#143390000000
1!
b100 %
1'
b100 +
#143400000000
1"
1(
#143410000000
0!
0"
b100 &
0'
0(
b100 ,
#143420000000
1!
b101 %
1'
b101 +
#143430000000
0!
0'
#143440000000
1!
b110 %
1'
b110 +
#143450000000
0!
0'
#143460000000
1!
b111 %
1'
b111 +
#143470000000
0!
0'
#143480000000
1!
0$
b1000 %
1'
0*
b1000 +
#143490000000
0!
0'
#143500000000
1!
b1001 %
1'
b1001 +
#143510000000
0!
0'
#143520000000
1!
b0 %
1'
b0 +
#143530000000
0!
0'
#143540000000
1!
1$
b1 %
1'
1*
b1 +
#143550000000
0!
0'
#143560000000
1!
b10 %
1'
b10 +
#143570000000
0!
0'
#143580000000
1!
b11 %
1'
b11 +
#143590000000
0!
0'
#143600000000
1!
b100 %
1'
b100 +
#143610000000
0!
0'
#143620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#143630000000
0!
0'
#143640000000
1!
0$
b110 %
1'
0*
b110 +
#143650000000
0!
0'
#143660000000
1!
b111 %
1'
b111 +
#143670000000
0!
0'
#143680000000
1!
b1000 %
1'
b1000 +
#143690000000
0!
0'
#143700000000
1!
b1001 %
1'
b1001 +
#143710000000
0!
0'
#143720000000
1!
b0 %
1'
b0 +
#143730000000
0!
0'
#143740000000
1!
1$
b1 %
1'
1*
b1 +
#143750000000
0!
0'
#143760000000
1!
b10 %
1'
b10 +
#143770000000
0!
0'
#143780000000
1!
b11 %
1'
b11 +
#143790000000
0!
0'
#143800000000
1!
b100 %
1'
b100 +
#143810000000
0!
0'
#143820000000
1!
b101 %
1'
b101 +
#143830000000
1"
1(
#143840000000
0!
0"
b100 &
0'
0(
b100 ,
#143850000000
1!
b110 %
1'
b110 +
#143860000000
0!
0'
#143870000000
1!
b111 %
1'
b111 +
#143880000000
0!
0'
#143890000000
1!
0$
b1000 %
1'
0*
b1000 +
#143900000000
0!
0'
#143910000000
1!
b1001 %
1'
b1001 +
#143920000000
0!
0'
#143930000000
1!
b0 %
1'
b0 +
#143940000000
0!
0'
#143950000000
1!
1$
b1 %
1'
1*
b1 +
#143960000000
0!
0'
#143970000000
1!
b10 %
1'
b10 +
#143980000000
0!
0'
#143990000000
1!
b11 %
1'
b11 +
#144000000000
0!
0'
#144010000000
1!
b100 %
1'
b100 +
#144020000000
0!
0'
#144030000000
1!
b101 %
1'
b101 +
#144040000000
0!
0'
#144050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#144060000000
0!
0'
#144070000000
1!
b111 %
1'
b111 +
#144080000000
0!
0'
#144090000000
1!
b1000 %
1'
b1000 +
#144100000000
0!
0'
#144110000000
1!
b1001 %
1'
b1001 +
#144120000000
0!
0'
#144130000000
1!
b0 %
1'
b0 +
#144140000000
0!
0'
#144150000000
1!
1$
b1 %
1'
1*
b1 +
#144160000000
0!
0'
#144170000000
1!
b10 %
1'
b10 +
#144180000000
0!
0'
#144190000000
1!
b11 %
1'
b11 +
#144200000000
0!
0'
#144210000000
1!
b100 %
1'
b100 +
#144220000000
0!
0'
#144230000000
1!
b101 %
1'
b101 +
#144240000000
0!
0'
#144250000000
1!
0$
b110 %
1'
0*
b110 +
#144260000000
1"
1(
#144270000000
0!
0"
b100 &
0'
0(
b100 ,
#144280000000
1!
1$
b111 %
1'
1*
b111 +
#144290000000
0!
0'
#144300000000
1!
0$
b1000 %
1'
0*
b1000 +
#144310000000
0!
0'
#144320000000
1!
b1001 %
1'
b1001 +
#144330000000
0!
0'
#144340000000
1!
b0 %
1'
b0 +
#144350000000
0!
0'
#144360000000
1!
1$
b1 %
1'
1*
b1 +
#144370000000
0!
0'
#144380000000
1!
b10 %
1'
b10 +
#144390000000
0!
0'
#144400000000
1!
b11 %
1'
b11 +
#144410000000
0!
0'
#144420000000
1!
b100 %
1'
b100 +
#144430000000
0!
0'
#144440000000
1!
b101 %
1'
b101 +
#144450000000
0!
0'
#144460000000
1!
b110 %
1'
b110 +
#144470000000
0!
0'
#144480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#144490000000
0!
0'
#144500000000
1!
b1000 %
1'
b1000 +
#144510000000
0!
0'
#144520000000
1!
b1001 %
1'
b1001 +
#144530000000
0!
0'
#144540000000
1!
b0 %
1'
b0 +
#144550000000
0!
0'
#144560000000
1!
1$
b1 %
1'
1*
b1 +
#144570000000
0!
0'
#144580000000
1!
b10 %
1'
b10 +
#144590000000
0!
0'
#144600000000
1!
b11 %
1'
b11 +
#144610000000
0!
0'
#144620000000
1!
b100 %
1'
b100 +
#144630000000
0!
0'
#144640000000
1!
b101 %
1'
b101 +
#144650000000
0!
0'
#144660000000
1!
0$
b110 %
1'
0*
b110 +
#144670000000
0!
0'
#144680000000
1!
b111 %
1'
b111 +
#144690000000
1"
1(
#144700000000
0!
0"
b100 &
0'
0(
b100 ,
#144710000000
1!
b1000 %
1'
b1000 +
#144720000000
0!
0'
#144730000000
1!
b1001 %
1'
b1001 +
#144740000000
0!
0'
#144750000000
1!
b0 %
1'
b0 +
#144760000000
0!
0'
#144770000000
1!
1$
b1 %
1'
1*
b1 +
#144780000000
0!
0'
#144790000000
1!
b10 %
1'
b10 +
#144800000000
0!
0'
#144810000000
1!
b11 %
1'
b11 +
#144820000000
0!
0'
#144830000000
1!
b100 %
1'
b100 +
#144840000000
0!
0'
#144850000000
1!
b101 %
1'
b101 +
#144860000000
0!
0'
#144870000000
1!
b110 %
1'
b110 +
#144880000000
0!
0'
#144890000000
1!
b111 %
1'
b111 +
#144900000000
0!
0'
#144910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#144920000000
0!
0'
#144930000000
1!
b1001 %
1'
b1001 +
#144940000000
0!
0'
#144950000000
1!
b0 %
1'
b0 +
#144960000000
0!
0'
#144970000000
1!
1$
b1 %
1'
1*
b1 +
#144980000000
0!
0'
#144990000000
1!
b10 %
1'
b10 +
#145000000000
0!
0'
#145010000000
1!
b11 %
1'
b11 +
#145020000000
0!
0'
#145030000000
1!
b100 %
1'
b100 +
#145040000000
0!
0'
#145050000000
1!
b101 %
1'
b101 +
#145060000000
0!
0'
#145070000000
1!
0$
b110 %
1'
0*
b110 +
#145080000000
0!
0'
#145090000000
1!
b111 %
1'
b111 +
#145100000000
0!
0'
#145110000000
1!
b1000 %
1'
b1000 +
#145120000000
1"
1(
#145130000000
0!
0"
b100 &
0'
0(
b100 ,
#145140000000
1!
b1001 %
1'
b1001 +
#145150000000
0!
0'
#145160000000
1!
b0 %
1'
b0 +
#145170000000
0!
0'
#145180000000
1!
1$
b1 %
1'
1*
b1 +
#145190000000
0!
0'
#145200000000
1!
b10 %
1'
b10 +
#145210000000
0!
0'
#145220000000
1!
b11 %
1'
b11 +
#145230000000
0!
0'
#145240000000
1!
b100 %
1'
b100 +
#145250000000
0!
0'
#145260000000
1!
b101 %
1'
b101 +
#145270000000
0!
0'
#145280000000
1!
b110 %
1'
b110 +
#145290000000
0!
0'
#145300000000
1!
b111 %
1'
b111 +
#145310000000
0!
0'
#145320000000
1!
0$
b1000 %
1'
0*
b1000 +
#145330000000
0!
0'
#145340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#145350000000
0!
0'
#145360000000
1!
b0 %
1'
b0 +
#145370000000
0!
0'
#145380000000
1!
1$
b1 %
1'
1*
b1 +
#145390000000
0!
0'
#145400000000
1!
b10 %
1'
b10 +
#145410000000
0!
0'
#145420000000
1!
b11 %
1'
b11 +
#145430000000
0!
0'
#145440000000
1!
b100 %
1'
b100 +
#145450000000
0!
0'
#145460000000
1!
b101 %
1'
b101 +
#145470000000
0!
0'
#145480000000
1!
0$
b110 %
1'
0*
b110 +
#145490000000
0!
0'
#145500000000
1!
b111 %
1'
b111 +
#145510000000
0!
0'
#145520000000
1!
b1000 %
1'
b1000 +
#145530000000
0!
0'
#145540000000
1!
b1001 %
1'
b1001 +
#145550000000
1"
1(
#145560000000
0!
0"
b100 &
0'
0(
b100 ,
#145570000000
1!
b0 %
1'
b0 +
#145580000000
0!
0'
#145590000000
1!
1$
b1 %
1'
1*
b1 +
#145600000000
0!
0'
#145610000000
1!
b10 %
1'
b10 +
#145620000000
0!
0'
#145630000000
1!
b11 %
1'
b11 +
#145640000000
0!
0'
#145650000000
1!
b100 %
1'
b100 +
#145660000000
0!
0'
#145670000000
1!
b101 %
1'
b101 +
#145680000000
0!
0'
#145690000000
1!
b110 %
1'
b110 +
#145700000000
0!
0'
#145710000000
1!
b111 %
1'
b111 +
#145720000000
0!
0'
#145730000000
1!
0$
b1000 %
1'
0*
b1000 +
#145740000000
0!
0'
#145750000000
1!
b1001 %
1'
b1001 +
#145760000000
0!
0'
#145770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#145780000000
0!
0'
#145790000000
1!
1$
b1 %
1'
1*
b1 +
#145800000000
0!
0'
#145810000000
1!
b10 %
1'
b10 +
#145820000000
0!
0'
#145830000000
1!
b11 %
1'
b11 +
#145840000000
0!
0'
#145850000000
1!
b100 %
1'
b100 +
#145860000000
0!
0'
#145870000000
1!
b101 %
1'
b101 +
#145880000000
0!
0'
#145890000000
1!
0$
b110 %
1'
0*
b110 +
#145900000000
0!
0'
#145910000000
1!
b111 %
1'
b111 +
#145920000000
0!
0'
#145930000000
1!
b1000 %
1'
b1000 +
#145940000000
0!
0'
#145950000000
1!
b1001 %
1'
b1001 +
#145960000000
0!
0'
#145970000000
1!
b0 %
1'
b0 +
#145980000000
1"
1(
#145990000000
0!
0"
b100 &
0'
0(
b100 ,
#146000000000
1!
1$
b1 %
1'
1*
b1 +
#146010000000
0!
0'
#146020000000
1!
b10 %
1'
b10 +
#146030000000
0!
0'
#146040000000
1!
b11 %
1'
b11 +
#146050000000
0!
0'
#146060000000
1!
b100 %
1'
b100 +
#146070000000
0!
0'
#146080000000
1!
b101 %
1'
b101 +
#146090000000
0!
0'
#146100000000
1!
b110 %
1'
b110 +
#146110000000
0!
0'
#146120000000
1!
b111 %
1'
b111 +
#146130000000
0!
0'
#146140000000
1!
0$
b1000 %
1'
0*
b1000 +
#146150000000
0!
0'
#146160000000
1!
b1001 %
1'
b1001 +
#146170000000
0!
0'
#146180000000
1!
b0 %
1'
b0 +
#146190000000
0!
0'
#146200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#146210000000
0!
0'
#146220000000
1!
b10 %
1'
b10 +
#146230000000
0!
0'
#146240000000
1!
b11 %
1'
b11 +
#146250000000
0!
0'
#146260000000
1!
b100 %
1'
b100 +
#146270000000
0!
0'
#146280000000
1!
b101 %
1'
b101 +
#146290000000
0!
0'
#146300000000
1!
0$
b110 %
1'
0*
b110 +
#146310000000
0!
0'
#146320000000
1!
b111 %
1'
b111 +
#146330000000
0!
0'
#146340000000
1!
b1000 %
1'
b1000 +
#146350000000
0!
0'
#146360000000
1!
b1001 %
1'
b1001 +
#146370000000
0!
0'
#146380000000
1!
b0 %
1'
b0 +
#146390000000
0!
0'
#146400000000
1!
1$
b1 %
1'
1*
b1 +
#146410000000
1"
1(
#146420000000
0!
0"
b100 &
0'
0(
b100 ,
#146430000000
1!
b10 %
1'
b10 +
#146440000000
0!
0'
#146450000000
1!
b11 %
1'
b11 +
#146460000000
0!
0'
#146470000000
1!
b100 %
1'
b100 +
#146480000000
0!
0'
#146490000000
1!
b101 %
1'
b101 +
#146500000000
0!
0'
#146510000000
1!
b110 %
1'
b110 +
#146520000000
0!
0'
#146530000000
1!
b111 %
1'
b111 +
#146540000000
0!
0'
#146550000000
1!
0$
b1000 %
1'
0*
b1000 +
#146560000000
0!
0'
#146570000000
1!
b1001 %
1'
b1001 +
#146580000000
0!
0'
#146590000000
1!
b0 %
1'
b0 +
#146600000000
0!
0'
#146610000000
1!
1$
b1 %
1'
1*
b1 +
#146620000000
0!
0'
#146630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#146640000000
0!
0'
#146650000000
1!
b11 %
1'
b11 +
#146660000000
0!
0'
#146670000000
1!
b100 %
1'
b100 +
#146680000000
0!
0'
#146690000000
1!
b101 %
1'
b101 +
#146700000000
0!
0'
#146710000000
1!
0$
b110 %
1'
0*
b110 +
#146720000000
0!
0'
#146730000000
1!
b111 %
1'
b111 +
#146740000000
0!
0'
#146750000000
1!
b1000 %
1'
b1000 +
#146760000000
0!
0'
#146770000000
1!
b1001 %
1'
b1001 +
#146780000000
0!
0'
#146790000000
1!
b0 %
1'
b0 +
#146800000000
0!
0'
#146810000000
1!
1$
b1 %
1'
1*
b1 +
#146820000000
0!
0'
#146830000000
1!
b10 %
1'
b10 +
#146840000000
1"
1(
#146850000000
0!
0"
b100 &
0'
0(
b100 ,
#146860000000
1!
b11 %
1'
b11 +
#146870000000
0!
0'
#146880000000
1!
b100 %
1'
b100 +
#146890000000
0!
0'
#146900000000
1!
b101 %
1'
b101 +
#146910000000
0!
0'
#146920000000
1!
b110 %
1'
b110 +
#146930000000
0!
0'
#146940000000
1!
b111 %
1'
b111 +
#146950000000
0!
0'
#146960000000
1!
0$
b1000 %
1'
0*
b1000 +
#146970000000
0!
0'
#146980000000
1!
b1001 %
1'
b1001 +
#146990000000
0!
0'
#147000000000
1!
b0 %
1'
b0 +
#147010000000
0!
0'
#147020000000
1!
1$
b1 %
1'
1*
b1 +
#147030000000
0!
0'
#147040000000
1!
b10 %
1'
b10 +
#147050000000
0!
0'
#147060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#147070000000
0!
0'
#147080000000
1!
b100 %
1'
b100 +
#147090000000
0!
0'
#147100000000
1!
b101 %
1'
b101 +
#147110000000
0!
0'
#147120000000
1!
0$
b110 %
1'
0*
b110 +
#147130000000
0!
0'
#147140000000
1!
b111 %
1'
b111 +
#147150000000
0!
0'
#147160000000
1!
b1000 %
1'
b1000 +
#147170000000
0!
0'
#147180000000
1!
b1001 %
1'
b1001 +
#147190000000
0!
0'
#147200000000
1!
b0 %
1'
b0 +
#147210000000
0!
0'
#147220000000
1!
1$
b1 %
1'
1*
b1 +
#147230000000
0!
0'
#147240000000
1!
b10 %
1'
b10 +
#147250000000
0!
0'
#147260000000
1!
b11 %
1'
b11 +
#147270000000
1"
1(
#147280000000
0!
0"
b100 &
0'
0(
b100 ,
#147290000000
1!
b100 %
1'
b100 +
#147300000000
0!
0'
#147310000000
1!
b101 %
1'
b101 +
#147320000000
0!
0'
#147330000000
1!
b110 %
1'
b110 +
#147340000000
0!
0'
#147350000000
1!
b111 %
1'
b111 +
#147360000000
0!
0'
#147370000000
1!
0$
b1000 %
1'
0*
b1000 +
#147380000000
0!
0'
#147390000000
1!
b1001 %
1'
b1001 +
#147400000000
0!
0'
#147410000000
1!
b0 %
1'
b0 +
#147420000000
0!
0'
#147430000000
1!
1$
b1 %
1'
1*
b1 +
#147440000000
0!
0'
#147450000000
1!
b10 %
1'
b10 +
#147460000000
0!
0'
#147470000000
1!
b11 %
1'
b11 +
#147480000000
0!
0'
#147490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#147500000000
0!
0'
#147510000000
1!
b101 %
1'
b101 +
#147520000000
0!
0'
#147530000000
1!
0$
b110 %
1'
0*
b110 +
#147540000000
0!
0'
#147550000000
1!
b111 %
1'
b111 +
#147560000000
0!
0'
#147570000000
1!
b1000 %
1'
b1000 +
#147580000000
0!
0'
#147590000000
1!
b1001 %
1'
b1001 +
#147600000000
0!
0'
#147610000000
1!
b0 %
1'
b0 +
#147620000000
0!
0'
#147630000000
1!
1$
b1 %
1'
1*
b1 +
#147640000000
0!
0'
#147650000000
1!
b10 %
1'
b10 +
#147660000000
0!
0'
#147670000000
1!
b11 %
1'
b11 +
#147680000000
0!
0'
#147690000000
1!
b100 %
1'
b100 +
#147700000000
1"
1(
#147710000000
0!
0"
b100 &
0'
0(
b100 ,
#147720000000
1!
b101 %
1'
b101 +
#147730000000
0!
0'
#147740000000
1!
b110 %
1'
b110 +
#147750000000
0!
0'
#147760000000
1!
b111 %
1'
b111 +
#147770000000
0!
0'
#147780000000
1!
0$
b1000 %
1'
0*
b1000 +
#147790000000
0!
0'
#147800000000
1!
b1001 %
1'
b1001 +
#147810000000
0!
0'
#147820000000
1!
b0 %
1'
b0 +
#147830000000
0!
0'
#147840000000
1!
1$
b1 %
1'
1*
b1 +
#147850000000
0!
0'
#147860000000
1!
b10 %
1'
b10 +
#147870000000
0!
0'
#147880000000
1!
b11 %
1'
b11 +
#147890000000
0!
0'
#147900000000
1!
b100 %
1'
b100 +
#147910000000
0!
0'
#147920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#147930000000
0!
0'
#147940000000
1!
0$
b110 %
1'
0*
b110 +
#147950000000
0!
0'
#147960000000
1!
b111 %
1'
b111 +
#147970000000
0!
0'
#147980000000
1!
b1000 %
1'
b1000 +
#147990000000
0!
0'
#148000000000
1!
b1001 %
1'
b1001 +
#148010000000
0!
0'
#148020000000
1!
b0 %
1'
b0 +
#148030000000
0!
0'
#148040000000
1!
1$
b1 %
1'
1*
b1 +
#148050000000
0!
0'
#148060000000
1!
b10 %
1'
b10 +
#148070000000
0!
0'
#148080000000
1!
b11 %
1'
b11 +
#148090000000
0!
0'
#148100000000
1!
b100 %
1'
b100 +
#148110000000
0!
0'
#148120000000
1!
b101 %
1'
b101 +
#148130000000
1"
1(
#148140000000
0!
0"
b100 &
0'
0(
b100 ,
#148150000000
1!
b110 %
1'
b110 +
#148160000000
0!
0'
#148170000000
1!
b111 %
1'
b111 +
#148180000000
0!
0'
#148190000000
1!
0$
b1000 %
1'
0*
b1000 +
#148200000000
0!
0'
#148210000000
1!
b1001 %
1'
b1001 +
#148220000000
0!
0'
#148230000000
1!
b0 %
1'
b0 +
#148240000000
0!
0'
#148250000000
1!
1$
b1 %
1'
1*
b1 +
#148260000000
0!
0'
#148270000000
1!
b10 %
1'
b10 +
#148280000000
0!
0'
#148290000000
1!
b11 %
1'
b11 +
#148300000000
0!
0'
#148310000000
1!
b100 %
1'
b100 +
#148320000000
0!
0'
#148330000000
1!
b101 %
1'
b101 +
#148340000000
0!
0'
#148350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#148360000000
0!
0'
#148370000000
1!
b111 %
1'
b111 +
#148380000000
0!
0'
#148390000000
1!
b1000 %
1'
b1000 +
#148400000000
0!
0'
#148410000000
1!
b1001 %
1'
b1001 +
#148420000000
0!
0'
#148430000000
1!
b0 %
1'
b0 +
#148440000000
0!
0'
#148450000000
1!
1$
b1 %
1'
1*
b1 +
#148460000000
0!
0'
#148470000000
1!
b10 %
1'
b10 +
#148480000000
0!
0'
#148490000000
1!
b11 %
1'
b11 +
#148500000000
0!
0'
#148510000000
1!
b100 %
1'
b100 +
#148520000000
0!
0'
#148530000000
1!
b101 %
1'
b101 +
#148540000000
0!
0'
#148550000000
1!
0$
b110 %
1'
0*
b110 +
#148560000000
1"
1(
#148570000000
0!
0"
b100 &
0'
0(
b100 ,
#148580000000
1!
1$
b111 %
1'
1*
b111 +
#148590000000
0!
0'
#148600000000
1!
0$
b1000 %
1'
0*
b1000 +
#148610000000
0!
0'
#148620000000
1!
b1001 %
1'
b1001 +
#148630000000
0!
0'
#148640000000
1!
b0 %
1'
b0 +
#148650000000
0!
0'
#148660000000
1!
1$
b1 %
1'
1*
b1 +
#148670000000
0!
0'
#148680000000
1!
b10 %
1'
b10 +
#148690000000
0!
0'
#148700000000
1!
b11 %
1'
b11 +
#148710000000
0!
0'
#148720000000
1!
b100 %
1'
b100 +
#148730000000
0!
0'
#148740000000
1!
b101 %
1'
b101 +
#148750000000
0!
0'
#148760000000
1!
b110 %
1'
b110 +
#148770000000
0!
0'
#148780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#148790000000
0!
0'
#148800000000
1!
b1000 %
1'
b1000 +
#148810000000
0!
0'
#148820000000
1!
b1001 %
1'
b1001 +
#148830000000
0!
0'
#148840000000
1!
b0 %
1'
b0 +
#148850000000
0!
0'
#148860000000
1!
1$
b1 %
1'
1*
b1 +
#148870000000
0!
0'
#148880000000
1!
b10 %
1'
b10 +
#148890000000
0!
0'
#148900000000
1!
b11 %
1'
b11 +
#148910000000
0!
0'
#148920000000
1!
b100 %
1'
b100 +
#148930000000
0!
0'
#148940000000
1!
b101 %
1'
b101 +
#148950000000
0!
0'
#148960000000
1!
0$
b110 %
1'
0*
b110 +
#148970000000
0!
0'
#148980000000
1!
b111 %
1'
b111 +
#148990000000
1"
1(
#149000000000
0!
0"
b100 &
0'
0(
b100 ,
#149010000000
1!
b1000 %
1'
b1000 +
#149020000000
0!
0'
#149030000000
1!
b1001 %
1'
b1001 +
#149040000000
0!
0'
#149050000000
1!
b0 %
1'
b0 +
#149060000000
0!
0'
#149070000000
1!
1$
b1 %
1'
1*
b1 +
#149080000000
0!
0'
#149090000000
1!
b10 %
1'
b10 +
#149100000000
0!
0'
#149110000000
1!
b11 %
1'
b11 +
#149120000000
0!
0'
#149130000000
1!
b100 %
1'
b100 +
#149140000000
0!
0'
#149150000000
1!
b101 %
1'
b101 +
#149160000000
0!
0'
#149170000000
1!
b110 %
1'
b110 +
#149180000000
0!
0'
#149190000000
1!
b111 %
1'
b111 +
#149200000000
0!
0'
#149210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#149220000000
0!
0'
#149230000000
1!
b1001 %
1'
b1001 +
#149240000000
0!
0'
#149250000000
1!
b0 %
1'
b0 +
#149260000000
0!
0'
#149270000000
1!
1$
b1 %
1'
1*
b1 +
#149280000000
0!
0'
#149290000000
1!
b10 %
1'
b10 +
#149300000000
0!
0'
#149310000000
1!
b11 %
1'
b11 +
#149320000000
0!
0'
#149330000000
1!
b100 %
1'
b100 +
#149340000000
0!
0'
#149350000000
1!
b101 %
1'
b101 +
#149360000000
0!
0'
#149370000000
1!
0$
b110 %
1'
0*
b110 +
#149380000000
0!
0'
#149390000000
1!
b111 %
1'
b111 +
#149400000000
0!
0'
#149410000000
1!
b1000 %
1'
b1000 +
#149420000000
1"
1(
#149430000000
0!
0"
b100 &
0'
0(
b100 ,
#149440000000
1!
b1001 %
1'
b1001 +
#149450000000
0!
0'
#149460000000
1!
b0 %
1'
b0 +
#149470000000
0!
0'
#149480000000
1!
1$
b1 %
1'
1*
b1 +
#149490000000
0!
0'
#149500000000
1!
b10 %
1'
b10 +
#149510000000
0!
0'
#149520000000
1!
b11 %
1'
b11 +
#149530000000
0!
0'
#149540000000
1!
b100 %
1'
b100 +
#149550000000
0!
0'
#149560000000
1!
b101 %
1'
b101 +
#149570000000
0!
0'
#149580000000
1!
b110 %
1'
b110 +
#149590000000
0!
0'
#149600000000
1!
b111 %
1'
b111 +
#149610000000
0!
0'
#149620000000
1!
0$
b1000 %
1'
0*
b1000 +
#149630000000
0!
0'
#149640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#149650000000
0!
0'
#149660000000
1!
b0 %
1'
b0 +
#149670000000
0!
0'
#149680000000
1!
1$
b1 %
1'
1*
b1 +
#149690000000
0!
0'
#149700000000
1!
b10 %
1'
b10 +
#149710000000
0!
0'
#149720000000
1!
b11 %
1'
b11 +
#149730000000
0!
0'
#149740000000
1!
b100 %
1'
b100 +
#149750000000
0!
0'
#149760000000
1!
b101 %
1'
b101 +
#149770000000
0!
0'
#149780000000
1!
0$
b110 %
1'
0*
b110 +
#149790000000
0!
0'
#149800000000
1!
b111 %
1'
b111 +
#149810000000
0!
0'
#149820000000
1!
b1000 %
1'
b1000 +
#149830000000
0!
0'
#149840000000
1!
b1001 %
1'
b1001 +
#149850000000
1"
1(
#149860000000
0!
0"
b100 &
0'
0(
b100 ,
#149870000000
1!
b0 %
1'
b0 +
#149880000000
0!
0'
#149890000000
1!
1$
b1 %
1'
1*
b1 +
#149900000000
0!
0'
#149910000000
1!
b10 %
1'
b10 +
#149920000000
0!
0'
#149930000000
1!
b11 %
1'
b11 +
#149940000000
0!
0'
#149950000000
1!
b100 %
1'
b100 +
#149960000000
0!
0'
#149970000000
1!
b101 %
1'
b101 +
#149980000000
0!
0'
#149990000000
1!
b110 %
1'
b110 +
#150000000000
0!
0'
#150010000000
1!
b111 %
1'
b111 +
#150020000000
0!
0'
#150030000000
1!
0$
b1000 %
1'
0*
b1000 +
#150040000000
0!
0'
#150050000000
1!
b1001 %
1'
b1001 +
#150060000000
0!
0'
#150070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#150080000000
0!
0'
#150090000000
1!
1$
b1 %
1'
1*
b1 +
#150100000000
0!
0'
#150110000000
1!
b10 %
1'
b10 +
#150120000000
0!
0'
#150130000000
1!
b11 %
1'
b11 +
#150140000000
0!
0'
#150150000000
1!
b100 %
1'
b100 +
#150160000000
0!
0'
#150170000000
1!
b101 %
1'
b101 +
#150180000000
0!
0'
#150190000000
1!
0$
b110 %
1'
0*
b110 +
#150200000000
0!
0'
#150210000000
1!
b111 %
1'
b111 +
#150220000000
0!
0'
#150230000000
1!
b1000 %
1'
b1000 +
#150240000000
0!
0'
#150250000000
1!
b1001 %
1'
b1001 +
#150260000000
0!
0'
#150270000000
1!
b0 %
1'
b0 +
#150280000000
1"
1(
#150290000000
0!
0"
b100 &
0'
0(
b100 ,
#150300000000
1!
1$
b1 %
1'
1*
b1 +
#150310000000
0!
0'
#150320000000
1!
b10 %
1'
b10 +
#150330000000
0!
0'
#150340000000
1!
b11 %
1'
b11 +
#150350000000
0!
0'
#150360000000
1!
b100 %
1'
b100 +
#150370000000
0!
0'
#150380000000
1!
b101 %
1'
b101 +
#150390000000
0!
0'
#150400000000
1!
b110 %
1'
b110 +
#150410000000
0!
0'
#150420000000
1!
b111 %
1'
b111 +
#150430000000
0!
0'
#150440000000
1!
0$
b1000 %
1'
0*
b1000 +
#150450000000
0!
0'
#150460000000
1!
b1001 %
1'
b1001 +
#150470000000
0!
0'
#150480000000
1!
b0 %
1'
b0 +
#150490000000
0!
0'
#150500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#150510000000
0!
0'
#150520000000
1!
b10 %
1'
b10 +
#150530000000
0!
0'
#150540000000
1!
b11 %
1'
b11 +
#150550000000
0!
0'
#150560000000
1!
b100 %
1'
b100 +
#150570000000
0!
0'
#150580000000
1!
b101 %
1'
b101 +
#150590000000
0!
0'
#150600000000
1!
0$
b110 %
1'
0*
b110 +
#150610000000
0!
0'
#150620000000
1!
b111 %
1'
b111 +
#150630000000
0!
0'
#150640000000
1!
b1000 %
1'
b1000 +
#150650000000
0!
0'
#150660000000
1!
b1001 %
1'
b1001 +
#150670000000
0!
0'
#150680000000
1!
b0 %
1'
b0 +
#150690000000
0!
0'
#150700000000
1!
1$
b1 %
1'
1*
b1 +
#150710000000
1"
1(
#150720000000
0!
0"
b100 &
0'
0(
b100 ,
#150730000000
1!
b10 %
1'
b10 +
#150740000000
0!
0'
#150750000000
1!
b11 %
1'
b11 +
#150760000000
0!
0'
#150770000000
1!
b100 %
1'
b100 +
#150780000000
0!
0'
#150790000000
1!
b101 %
1'
b101 +
#150800000000
0!
0'
#150810000000
1!
b110 %
1'
b110 +
#150820000000
0!
0'
#150830000000
1!
b111 %
1'
b111 +
#150840000000
0!
0'
#150850000000
1!
0$
b1000 %
1'
0*
b1000 +
#150860000000
0!
0'
#150870000000
1!
b1001 %
1'
b1001 +
#150880000000
0!
0'
#150890000000
1!
b0 %
1'
b0 +
#150900000000
0!
0'
#150910000000
1!
1$
b1 %
1'
1*
b1 +
#150920000000
0!
0'
#150930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#150940000000
0!
0'
#150950000000
1!
b11 %
1'
b11 +
#150960000000
0!
0'
#150970000000
1!
b100 %
1'
b100 +
#150980000000
0!
0'
#150990000000
1!
b101 %
1'
b101 +
#151000000000
0!
0'
#151010000000
1!
0$
b110 %
1'
0*
b110 +
#151020000000
0!
0'
#151030000000
1!
b111 %
1'
b111 +
#151040000000
0!
0'
#151050000000
1!
b1000 %
1'
b1000 +
#151060000000
0!
0'
#151070000000
1!
b1001 %
1'
b1001 +
#151080000000
0!
0'
#151090000000
1!
b0 %
1'
b0 +
#151100000000
0!
0'
#151110000000
1!
1$
b1 %
1'
1*
b1 +
#151120000000
0!
0'
#151130000000
1!
b10 %
1'
b10 +
#151140000000
1"
1(
#151150000000
0!
0"
b100 &
0'
0(
b100 ,
#151160000000
1!
b11 %
1'
b11 +
#151170000000
0!
0'
#151180000000
1!
b100 %
1'
b100 +
#151190000000
0!
0'
#151200000000
1!
b101 %
1'
b101 +
#151210000000
0!
0'
#151220000000
1!
b110 %
1'
b110 +
#151230000000
0!
0'
#151240000000
1!
b111 %
1'
b111 +
#151250000000
0!
0'
#151260000000
1!
0$
b1000 %
1'
0*
b1000 +
#151270000000
0!
0'
#151280000000
1!
b1001 %
1'
b1001 +
#151290000000
0!
0'
#151300000000
1!
b0 %
1'
b0 +
#151310000000
0!
0'
#151320000000
1!
1$
b1 %
1'
1*
b1 +
#151330000000
0!
0'
#151340000000
1!
b10 %
1'
b10 +
#151350000000
0!
0'
#151360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#151370000000
0!
0'
#151380000000
1!
b100 %
1'
b100 +
#151390000000
0!
0'
#151400000000
1!
b101 %
1'
b101 +
#151410000000
0!
0'
#151420000000
1!
0$
b110 %
1'
0*
b110 +
#151430000000
0!
0'
#151440000000
1!
b111 %
1'
b111 +
#151450000000
0!
0'
#151460000000
1!
b1000 %
1'
b1000 +
#151470000000
0!
0'
#151480000000
1!
b1001 %
1'
b1001 +
#151490000000
0!
0'
#151500000000
1!
b0 %
1'
b0 +
#151510000000
0!
0'
#151520000000
1!
1$
b1 %
1'
1*
b1 +
#151530000000
0!
0'
#151540000000
1!
b10 %
1'
b10 +
#151550000000
0!
0'
#151560000000
1!
b11 %
1'
b11 +
#151570000000
1"
1(
#151580000000
0!
0"
b100 &
0'
0(
b100 ,
#151590000000
1!
b100 %
1'
b100 +
#151600000000
0!
0'
#151610000000
1!
b101 %
1'
b101 +
#151620000000
0!
0'
#151630000000
1!
b110 %
1'
b110 +
#151640000000
0!
0'
#151650000000
1!
b111 %
1'
b111 +
#151660000000
0!
0'
#151670000000
1!
0$
b1000 %
1'
0*
b1000 +
#151680000000
0!
0'
#151690000000
1!
b1001 %
1'
b1001 +
#151700000000
0!
0'
#151710000000
1!
b0 %
1'
b0 +
#151720000000
0!
0'
#151730000000
1!
1$
b1 %
1'
1*
b1 +
#151740000000
0!
0'
#151750000000
1!
b10 %
1'
b10 +
#151760000000
0!
0'
#151770000000
1!
b11 %
1'
b11 +
#151780000000
0!
0'
#151790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#151800000000
0!
0'
#151810000000
1!
b101 %
1'
b101 +
#151820000000
0!
0'
#151830000000
1!
0$
b110 %
1'
0*
b110 +
#151840000000
0!
0'
#151850000000
1!
b111 %
1'
b111 +
#151860000000
0!
0'
#151870000000
1!
b1000 %
1'
b1000 +
#151880000000
0!
0'
#151890000000
1!
b1001 %
1'
b1001 +
#151900000000
0!
0'
#151910000000
1!
b0 %
1'
b0 +
#151920000000
0!
0'
#151930000000
1!
1$
b1 %
1'
1*
b1 +
#151940000000
0!
0'
#151950000000
1!
b10 %
1'
b10 +
#151960000000
0!
0'
#151970000000
1!
b11 %
1'
b11 +
#151980000000
0!
0'
#151990000000
1!
b100 %
1'
b100 +
#152000000000
1"
1(
#152010000000
0!
0"
b100 &
0'
0(
b100 ,
#152020000000
1!
b101 %
1'
b101 +
#152030000000
0!
0'
#152040000000
1!
b110 %
1'
b110 +
#152050000000
0!
0'
#152060000000
1!
b111 %
1'
b111 +
#152070000000
0!
0'
#152080000000
1!
0$
b1000 %
1'
0*
b1000 +
#152090000000
0!
0'
#152100000000
1!
b1001 %
1'
b1001 +
#152110000000
0!
0'
#152120000000
1!
b0 %
1'
b0 +
#152130000000
0!
0'
#152140000000
1!
1$
b1 %
1'
1*
b1 +
#152150000000
0!
0'
#152160000000
1!
b10 %
1'
b10 +
#152170000000
0!
0'
#152180000000
1!
b11 %
1'
b11 +
#152190000000
0!
0'
#152200000000
1!
b100 %
1'
b100 +
#152210000000
0!
0'
#152220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#152230000000
0!
0'
#152240000000
1!
0$
b110 %
1'
0*
b110 +
#152250000000
0!
0'
#152260000000
1!
b111 %
1'
b111 +
#152270000000
0!
0'
#152280000000
1!
b1000 %
1'
b1000 +
#152290000000
0!
0'
#152300000000
1!
b1001 %
1'
b1001 +
#152310000000
0!
0'
#152320000000
1!
b0 %
1'
b0 +
#152330000000
0!
0'
#152340000000
1!
1$
b1 %
1'
1*
b1 +
#152350000000
0!
0'
#152360000000
1!
b10 %
1'
b10 +
#152370000000
0!
0'
#152380000000
1!
b11 %
1'
b11 +
#152390000000
0!
0'
#152400000000
1!
b100 %
1'
b100 +
#152410000000
0!
0'
#152420000000
1!
b101 %
1'
b101 +
#152430000000
1"
1(
#152440000000
0!
0"
b100 &
0'
0(
b100 ,
#152450000000
1!
b110 %
1'
b110 +
#152460000000
0!
0'
#152470000000
1!
b111 %
1'
b111 +
#152480000000
0!
0'
#152490000000
1!
0$
b1000 %
1'
0*
b1000 +
#152500000000
0!
0'
#152510000000
1!
b1001 %
1'
b1001 +
#152520000000
0!
0'
#152530000000
1!
b0 %
1'
b0 +
#152540000000
0!
0'
#152550000000
1!
1$
b1 %
1'
1*
b1 +
#152560000000
0!
0'
#152570000000
1!
b10 %
1'
b10 +
#152580000000
0!
0'
#152590000000
1!
b11 %
1'
b11 +
#152600000000
0!
0'
#152610000000
1!
b100 %
1'
b100 +
#152620000000
0!
0'
#152630000000
1!
b101 %
1'
b101 +
#152640000000
0!
0'
#152650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#152660000000
0!
0'
#152670000000
1!
b111 %
1'
b111 +
#152680000000
0!
0'
#152690000000
1!
b1000 %
1'
b1000 +
#152700000000
0!
0'
#152710000000
1!
b1001 %
1'
b1001 +
#152720000000
0!
0'
#152730000000
1!
b0 %
1'
b0 +
#152740000000
0!
0'
#152750000000
1!
1$
b1 %
1'
1*
b1 +
#152760000000
0!
0'
#152770000000
1!
b10 %
1'
b10 +
#152780000000
0!
0'
#152790000000
1!
b11 %
1'
b11 +
#152800000000
0!
0'
#152810000000
1!
b100 %
1'
b100 +
#152820000000
0!
0'
#152830000000
1!
b101 %
1'
b101 +
#152840000000
0!
0'
#152850000000
1!
0$
b110 %
1'
0*
b110 +
#152860000000
1"
1(
#152870000000
0!
0"
b100 &
0'
0(
b100 ,
#152880000000
1!
1$
b111 %
1'
1*
b111 +
#152890000000
0!
0'
#152900000000
1!
0$
b1000 %
1'
0*
b1000 +
#152910000000
0!
0'
#152920000000
1!
b1001 %
1'
b1001 +
#152930000000
0!
0'
#152940000000
1!
b0 %
1'
b0 +
#152950000000
0!
0'
#152960000000
1!
1$
b1 %
1'
1*
b1 +
#152970000000
0!
0'
#152980000000
1!
b10 %
1'
b10 +
#152990000000
0!
0'
#153000000000
1!
b11 %
1'
b11 +
#153010000000
0!
0'
#153020000000
1!
b100 %
1'
b100 +
#153030000000
0!
0'
#153040000000
1!
b101 %
1'
b101 +
#153050000000
0!
0'
#153060000000
1!
b110 %
1'
b110 +
#153070000000
0!
0'
#153080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#153090000000
0!
0'
#153100000000
1!
b1000 %
1'
b1000 +
#153110000000
0!
0'
#153120000000
1!
b1001 %
1'
b1001 +
#153130000000
0!
0'
#153140000000
1!
b0 %
1'
b0 +
#153150000000
0!
0'
#153160000000
1!
1$
b1 %
1'
1*
b1 +
#153170000000
0!
0'
#153180000000
1!
b10 %
1'
b10 +
#153190000000
0!
0'
#153200000000
1!
b11 %
1'
b11 +
#153210000000
0!
0'
#153220000000
1!
b100 %
1'
b100 +
#153230000000
0!
0'
#153240000000
1!
b101 %
1'
b101 +
#153250000000
0!
0'
#153260000000
1!
0$
b110 %
1'
0*
b110 +
#153270000000
0!
0'
#153280000000
1!
b111 %
1'
b111 +
#153290000000
1"
1(
#153300000000
0!
0"
b100 &
0'
0(
b100 ,
#153310000000
1!
b1000 %
1'
b1000 +
#153320000000
0!
0'
#153330000000
1!
b1001 %
1'
b1001 +
#153340000000
0!
0'
#153350000000
1!
b0 %
1'
b0 +
#153360000000
0!
0'
#153370000000
1!
1$
b1 %
1'
1*
b1 +
#153380000000
0!
0'
#153390000000
1!
b10 %
1'
b10 +
#153400000000
0!
0'
#153410000000
1!
b11 %
1'
b11 +
#153420000000
0!
0'
#153430000000
1!
b100 %
1'
b100 +
#153440000000
0!
0'
#153450000000
1!
b101 %
1'
b101 +
#153460000000
0!
0'
#153470000000
1!
b110 %
1'
b110 +
#153480000000
0!
0'
#153490000000
1!
b111 %
1'
b111 +
#153500000000
0!
0'
#153510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#153520000000
0!
0'
#153530000000
1!
b1001 %
1'
b1001 +
#153540000000
0!
0'
#153550000000
1!
b0 %
1'
b0 +
#153560000000
0!
0'
#153570000000
1!
1$
b1 %
1'
1*
b1 +
#153580000000
0!
0'
#153590000000
1!
b10 %
1'
b10 +
#153600000000
0!
0'
#153610000000
1!
b11 %
1'
b11 +
#153620000000
0!
0'
#153630000000
1!
b100 %
1'
b100 +
#153640000000
0!
0'
#153650000000
1!
b101 %
1'
b101 +
#153660000000
0!
0'
#153670000000
1!
0$
b110 %
1'
0*
b110 +
#153680000000
0!
0'
#153690000000
1!
b111 %
1'
b111 +
#153700000000
0!
0'
#153710000000
1!
b1000 %
1'
b1000 +
#153720000000
1"
1(
#153730000000
0!
0"
b100 &
0'
0(
b100 ,
#153740000000
1!
b1001 %
1'
b1001 +
#153750000000
0!
0'
#153760000000
1!
b0 %
1'
b0 +
#153770000000
0!
0'
#153780000000
1!
1$
b1 %
1'
1*
b1 +
#153790000000
0!
0'
#153800000000
1!
b10 %
1'
b10 +
#153810000000
0!
0'
#153820000000
1!
b11 %
1'
b11 +
#153830000000
0!
0'
#153840000000
1!
b100 %
1'
b100 +
#153850000000
0!
0'
#153860000000
1!
b101 %
1'
b101 +
#153870000000
0!
0'
#153880000000
1!
b110 %
1'
b110 +
#153890000000
0!
0'
#153900000000
1!
b111 %
1'
b111 +
#153910000000
0!
0'
#153920000000
1!
0$
b1000 %
1'
0*
b1000 +
#153930000000
0!
0'
#153940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#153950000000
0!
0'
#153960000000
1!
b0 %
1'
b0 +
#153970000000
0!
0'
#153980000000
1!
1$
b1 %
1'
1*
b1 +
#153990000000
0!
0'
#154000000000
1!
b10 %
1'
b10 +
#154010000000
0!
0'
#154020000000
1!
b11 %
1'
b11 +
#154030000000
0!
0'
#154040000000
1!
b100 %
1'
b100 +
#154050000000
0!
0'
#154060000000
1!
b101 %
1'
b101 +
#154070000000
0!
0'
#154080000000
1!
0$
b110 %
1'
0*
b110 +
#154090000000
0!
0'
#154100000000
1!
b111 %
1'
b111 +
#154110000000
0!
0'
#154120000000
1!
b1000 %
1'
b1000 +
#154130000000
0!
0'
#154140000000
1!
b1001 %
1'
b1001 +
#154150000000
1"
1(
#154160000000
0!
0"
b100 &
0'
0(
b100 ,
#154170000000
1!
b0 %
1'
b0 +
#154180000000
0!
0'
#154190000000
1!
1$
b1 %
1'
1*
b1 +
#154200000000
0!
0'
#154210000000
1!
b10 %
1'
b10 +
#154220000000
0!
0'
#154230000000
1!
b11 %
1'
b11 +
#154240000000
0!
0'
#154250000000
1!
b100 %
1'
b100 +
#154260000000
0!
0'
#154270000000
1!
b101 %
1'
b101 +
#154280000000
0!
0'
#154290000000
1!
b110 %
1'
b110 +
#154300000000
0!
0'
#154310000000
1!
b111 %
1'
b111 +
#154320000000
0!
0'
#154330000000
1!
0$
b1000 %
1'
0*
b1000 +
#154340000000
0!
0'
#154350000000
1!
b1001 %
1'
b1001 +
#154360000000
0!
0'
#154370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#154380000000
0!
0'
#154390000000
1!
1$
b1 %
1'
1*
b1 +
#154400000000
0!
0'
#154410000000
1!
b10 %
1'
b10 +
#154420000000
0!
0'
#154430000000
1!
b11 %
1'
b11 +
#154440000000
0!
0'
#154450000000
1!
b100 %
1'
b100 +
#154460000000
0!
0'
#154470000000
1!
b101 %
1'
b101 +
#154480000000
0!
0'
#154490000000
1!
0$
b110 %
1'
0*
b110 +
#154500000000
0!
0'
#154510000000
1!
b111 %
1'
b111 +
#154520000000
0!
0'
#154530000000
1!
b1000 %
1'
b1000 +
#154540000000
0!
0'
#154550000000
1!
b1001 %
1'
b1001 +
#154560000000
0!
0'
#154570000000
1!
b0 %
1'
b0 +
#154580000000
1"
1(
#154590000000
0!
0"
b100 &
0'
0(
b100 ,
#154600000000
1!
1$
b1 %
1'
1*
b1 +
#154610000000
0!
0'
#154620000000
1!
b10 %
1'
b10 +
#154630000000
0!
0'
#154640000000
1!
b11 %
1'
b11 +
#154650000000
0!
0'
#154660000000
1!
b100 %
1'
b100 +
#154670000000
0!
0'
#154680000000
1!
b101 %
1'
b101 +
#154690000000
0!
0'
#154700000000
1!
b110 %
1'
b110 +
#154710000000
0!
0'
#154720000000
1!
b111 %
1'
b111 +
#154730000000
0!
0'
#154740000000
1!
0$
b1000 %
1'
0*
b1000 +
#154750000000
0!
0'
#154760000000
1!
b1001 %
1'
b1001 +
#154770000000
0!
0'
#154780000000
1!
b0 %
1'
b0 +
#154790000000
0!
0'
#154800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#154810000000
0!
0'
#154820000000
1!
b10 %
1'
b10 +
#154830000000
0!
0'
#154840000000
1!
b11 %
1'
b11 +
#154850000000
0!
0'
#154860000000
1!
b100 %
1'
b100 +
#154870000000
0!
0'
#154880000000
1!
b101 %
1'
b101 +
#154890000000
0!
0'
#154900000000
1!
0$
b110 %
1'
0*
b110 +
#154910000000
0!
0'
#154920000000
1!
b111 %
1'
b111 +
#154930000000
0!
0'
#154940000000
1!
b1000 %
1'
b1000 +
#154950000000
0!
0'
#154960000000
1!
b1001 %
1'
b1001 +
#154970000000
0!
0'
#154980000000
1!
b0 %
1'
b0 +
#154990000000
0!
0'
#155000000000
1!
1$
b1 %
1'
1*
b1 +
#155010000000
1"
1(
#155020000000
0!
0"
b100 &
0'
0(
b100 ,
#155030000000
1!
b10 %
1'
b10 +
#155040000000
0!
0'
#155050000000
1!
b11 %
1'
b11 +
#155060000000
0!
0'
#155070000000
1!
b100 %
1'
b100 +
#155080000000
0!
0'
#155090000000
1!
b101 %
1'
b101 +
#155100000000
0!
0'
#155110000000
1!
b110 %
1'
b110 +
#155120000000
0!
0'
#155130000000
1!
b111 %
1'
b111 +
#155140000000
0!
0'
#155150000000
1!
0$
b1000 %
1'
0*
b1000 +
#155160000000
0!
0'
#155170000000
1!
b1001 %
1'
b1001 +
#155180000000
0!
0'
#155190000000
1!
b0 %
1'
b0 +
#155200000000
0!
0'
#155210000000
1!
1$
b1 %
1'
1*
b1 +
#155220000000
0!
0'
#155230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#155240000000
0!
0'
#155250000000
1!
b11 %
1'
b11 +
#155260000000
0!
0'
#155270000000
1!
b100 %
1'
b100 +
#155280000000
0!
0'
#155290000000
1!
b101 %
1'
b101 +
#155300000000
0!
0'
#155310000000
1!
0$
b110 %
1'
0*
b110 +
#155320000000
0!
0'
#155330000000
1!
b111 %
1'
b111 +
#155340000000
0!
0'
#155350000000
1!
b1000 %
1'
b1000 +
#155360000000
0!
0'
#155370000000
1!
b1001 %
1'
b1001 +
#155380000000
0!
0'
#155390000000
1!
b0 %
1'
b0 +
#155400000000
0!
0'
#155410000000
1!
1$
b1 %
1'
1*
b1 +
#155420000000
0!
0'
#155430000000
1!
b10 %
1'
b10 +
#155440000000
1"
1(
#155450000000
0!
0"
b100 &
0'
0(
b100 ,
#155460000000
1!
b11 %
1'
b11 +
#155470000000
0!
0'
#155480000000
1!
b100 %
1'
b100 +
#155490000000
0!
0'
#155500000000
1!
b101 %
1'
b101 +
#155510000000
0!
0'
#155520000000
1!
b110 %
1'
b110 +
#155530000000
0!
0'
#155540000000
1!
b111 %
1'
b111 +
#155550000000
0!
0'
#155560000000
1!
0$
b1000 %
1'
0*
b1000 +
#155570000000
0!
0'
#155580000000
1!
b1001 %
1'
b1001 +
#155590000000
0!
0'
#155600000000
1!
b0 %
1'
b0 +
#155610000000
0!
0'
#155620000000
1!
1$
b1 %
1'
1*
b1 +
#155630000000
0!
0'
#155640000000
1!
b10 %
1'
b10 +
#155650000000
0!
0'
#155660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#155670000000
0!
0'
#155680000000
1!
b100 %
1'
b100 +
#155690000000
0!
0'
#155700000000
1!
b101 %
1'
b101 +
#155710000000
0!
0'
#155720000000
1!
0$
b110 %
1'
0*
b110 +
#155730000000
0!
0'
#155740000000
1!
b111 %
1'
b111 +
#155750000000
0!
0'
#155760000000
1!
b1000 %
1'
b1000 +
#155770000000
0!
0'
#155780000000
1!
b1001 %
1'
b1001 +
#155790000000
0!
0'
#155800000000
1!
b0 %
1'
b0 +
#155810000000
0!
0'
#155820000000
1!
1$
b1 %
1'
1*
b1 +
#155830000000
0!
0'
#155840000000
1!
b10 %
1'
b10 +
#155850000000
0!
0'
#155860000000
1!
b11 %
1'
b11 +
#155870000000
1"
1(
#155880000000
0!
0"
b100 &
0'
0(
b100 ,
#155890000000
1!
b100 %
1'
b100 +
#155900000000
0!
0'
#155910000000
1!
b101 %
1'
b101 +
#155920000000
0!
0'
#155930000000
1!
b110 %
1'
b110 +
#155940000000
0!
0'
#155950000000
1!
b111 %
1'
b111 +
#155960000000
0!
0'
#155970000000
1!
0$
b1000 %
1'
0*
b1000 +
#155980000000
0!
0'
#155990000000
1!
b1001 %
1'
b1001 +
#156000000000
0!
0'
#156010000000
1!
b0 %
1'
b0 +
#156020000000
0!
0'
#156030000000
1!
1$
b1 %
1'
1*
b1 +
#156040000000
0!
0'
#156050000000
1!
b10 %
1'
b10 +
#156060000000
0!
0'
#156070000000
1!
b11 %
1'
b11 +
#156080000000
0!
0'
#156090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#156100000000
0!
0'
#156110000000
1!
b101 %
1'
b101 +
#156120000000
0!
0'
#156130000000
1!
0$
b110 %
1'
0*
b110 +
#156140000000
0!
0'
#156150000000
1!
b111 %
1'
b111 +
#156160000000
0!
0'
#156170000000
1!
b1000 %
1'
b1000 +
#156180000000
0!
0'
#156190000000
1!
b1001 %
1'
b1001 +
#156200000000
0!
0'
#156210000000
1!
b0 %
1'
b0 +
#156220000000
0!
0'
#156230000000
1!
1$
b1 %
1'
1*
b1 +
#156240000000
0!
0'
#156250000000
1!
b10 %
1'
b10 +
#156260000000
0!
0'
#156270000000
1!
b11 %
1'
b11 +
#156280000000
0!
0'
#156290000000
1!
b100 %
1'
b100 +
#156300000000
1"
1(
#156310000000
0!
0"
b100 &
0'
0(
b100 ,
#156320000000
1!
b101 %
1'
b101 +
#156330000000
0!
0'
#156340000000
1!
b110 %
1'
b110 +
#156350000000
0!
0'
#156360000000
1!
b111 %
1'
b111 +
#156370000000
0!
0'
#156380000000
1!
0$
b1000 %
1'
0*
b1000 +
#156390000000
0!
0'
#156400000000
1!
b1001 %
1'
b1001 +
#156410000000
0!
0'
#156420000000
1!
b0 %
1'
b0 +
#156430000000
0!
0'
#156440000000
1!
1$
b1 %
1'
1*
b1 +
#156450000000
0!
0'
#156460000000
1!
b10 %
1'
b10 +
#156470000000
0!
0'
#156480000000
1!
b11 %
1'
b11 +
#156490000000
0!
0'
#156500000000
1!
b100 %
1'
b100 +
#156510000000
0!
0'
#156520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#156530000000
0!
0'
#156540000000
1!
0$
b110 %
1'
0*
b110 +
#156550000000
0!
0'
#156560000000
1!
b111 %
1'
b111 +
#156570000000
0!
0'
#156580000000
1!
b1000 %
1'
b1000 +
#156590000000
0!
0'
#156600000000
1!
b1001 %
1'
b1001 +
#156610000000
0!
0'
#156620000000
1!
b0 %
1'
b0 +
#156630000000
0!
0'
#156640000000
1!
1$
b1 %
1'
1*
b1 +
#156650000000
0!
0'
#156660000000
1!
b10 %
1'
b10 +
#156670000000
0!
0'
#156680000000
1!
b11 %
1'
b11 +
#156690000000
0!
0'
#156700000000
1!
b100 %
1'
b100 +
#156710000000
0!
0'
#156720000000
1!
b101 %
1'
b101 +
#156730000000
1"
1(
#156740000000
0!
0"
b100 &
0'
0(
b100 ,
#156750000000
1!
b110 %
1'
b110 +
#156760000000
0!
0'
#156770000000
1!
b111 %
1'
b111 +
#156780000000
0!
0'
#156790000000
1!
0$
b1000 %
1'
0*
b1000 +
#156800000000
0!
0'
#156810000000
1!
b1001 %
1'
b1001 +
#156820000000
0!
0'
#156830000000
1!
b0 %
1'
b0 +
#156840000000
0!
0'
#156850000000
1!
1$
b1 %
1'
1*
b1 +
#156860000000
0!
0'
#156870000000
1!
b10 %
1'
b10 +
#156880000000
0!
0'
#156890000000
1!
b11 %
1'
b11 +
#156900000000
0!
0'
#156910000000
1!
b100 %
1'
b100 +
#156920000000
0!
0'
#156930000000
1!
b101 %
1'
b101 +
#156940000000
0!
0'
#156950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#156960000000
0!
0'
#156970000000
1!
b111 %
1'
b111 +
#156980000000
0!
0'
#156990000000
1!
b1000 %
1'
b1000 +
#157000000000
0!
0'
#157010000000
1!
b1001 %
1'
b1001 +
#157020000000
0!
0'
#157030000000
1!
b0 %
1'
b0 +
#157040000000
0!
0'
#157050000000
1!
1$
b1 %
1'
1*
b1 +
#157060000000
0!
0'
#157070000000
1!
b10 %
1'
b10 +
#157080000000
0!
0'
#157090000000
1!
b11 %
1'
b11 +
#157100000000
0!
0'
#157110000000
1!
b100 %
1'
b100 +
#157120000000
0!
0'
#157130000000
1!
b101 %
1'
b101 +
#157140000000
0!
0'
#157150000000
1!
0$
b110 %
1'
0*
b110 +
#157160000000
1"
1(
#157170000000
0!
0"
b100 &
0'
0(
b100 ,
#157180000000
1!
1$
b111 %
1'
1*
b111 +
#157190000000
0!
0'
#157200000000
1!
0$
b1000 %
1'
0*
b1000 +
#157210000000
0!
0'
#157220000000
1!
b1001 %
1'
b1001 +
#157230000000
0!
0'
#157240000000
1!
b0 %
1'
b0 +
#157250000000
0!
0'
#157260000000
1!
1$
b1 %
1'
1*
b1 +
#157270000000
0!
0'
#157280000000
1!
b10 %
1'
b10 +
#157290000000
0!
0'
#157300000000
1!
b11 %
1'
b11 +
#157310000000
0!
0'
#157320000000
1!
b100 %
1'
b100 +
#157330000000
0!
0'
#157340000000
1!
b101 %
1'
b101 +
#157350000000
0!
0'
#157360000000
1!
b110 %
1'
b110 +
#157370000000
0!
0'
#157380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#157390000000
0!
0'
#157400000000
1!
b1000 %
1'
b1000 +
#157410000000
0!
0'
#157420000000
1!
b1001 %
1'
b1001 +
#157430000000
0!
0'
#157440000000
1!
b0 %
1'
b0 +
#157450000000
0!
0'
#157460000000
1!
1$
b1 %
1'
1*
b1 +
#157470000000
0!
0'
#157480000000
1!
b10 %
1'
b10 +
#157490000000
0!
0'
#157500000000
1!
b11 %
1'
b11 +
#157510000000
0!
0'
#157520000000
1!
b100 %
1'
b100 +
#157530000000
0!
0'
#157540000000
1!
b101 %
1'
b101 +
#157550000000
0!
0'
#157560000000
1!
0$
b110 %
1'
0*
b110 +
#157570000000
0!
0'
#157580000000
1!
b111 %
1'
b111 +
#157590000000
1"
1(
#157600000000
0!
0"
b100 &
0'
0(
b100 ,
#157610000000
1!
b1000 %
1'
b1000 +
#157620000000
0!
0'
#157630000000
1!
b1001 %
1'
b1001 +
#157640000000
0!
0'
#157650000000
1!
b0 %
1'
b0 +
#157660000000
0!
0'
#157670000000
1!
1$
b1 %
1'
1*
b1 +
#157680000000
0!
0'
#157690000000
1!
b10 %
1'
b10 +
#157700000000
0!
0'
#157710000000
1!
b11 %
1'
b11 +
#157720000000
0!
0'
#157730000000
1!
b100 %
1'
b100 +
#157740000000
0!
0'
#157750000000
1!
b101 %
1'
b101 +
#157760000000
0!
0'
#157770000000
1!
b110 %
1'
b110 +
#157780000000
0!
0'
#157790000000
1!
b111 %
1'
b111 +
#157800000000
0!
0'
#157810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#157820000000
0!
0'
#157830000000
1!
b1001 %
1'
b1001 +
#157840000000
0!
0'
#157850000000
1!
b0 %
1'
b0 +
#157860000000
0!
0'
#157870000000
1!
1$
b1 %
1'
1*
b1 +
#157880000000
0!
0'
#157890000000
1!
b10 %
1'
b10 +
#157900000000
0!
0'
#157910000000
1!
b11 %
1'
b11 +
#157920000000
0!
0'
#157930000000
1!
b100 %
1'
b100 +
#157940000000
0!
0'
#157950000000
1!
b101 %
1'
b101 +
#157960000000
0!
0'
#157970000000
1!
0$
b110 %
1'
0*
b110 +
#157980000000
0!
0'
#157990000000
1!
b111 %
1'
b111 +
#158000000000
0!
0'
#158010000000
1!
b1000 %
1'
b1000 +
#158020000000
1"
1(
#158030000000
0!
0"
b100 &
0'
0(
b100 ,
#158040000000
1!
b1001 %
1'
b1001 +
#158050000000
0!
0'
#158060000000
1!
b0 %
1'
b0 +
#158070000000
0!
0'
#158080000000
1!
1$
b1 %
1'
1*
b1 +
#158090000000
0!
0'
#158100000000
1!
b10 %
1'
b10 +
#158110000000
0!
0'
#158120000000
1!
b11 %
1'
b11 +
#158130000000
0!
0'
#158140000000
1!
b100 %
1'
b100 +
#158150000000
0!
0'
#158160000000
1!
b101 %
1'
b101 +
#158170000000
0!
0'
#158180000000
1!
b110 %
1'
b110 +
#158190000000
0!
0'
#158200000000
1!
b111 %
1'
b111 +
#158210000000
0!
0'
#158220000000
1!
0$
b1000 %
1'
0*
b1000 +
#158230000000
0!
0'
#158240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#158250000000
0!
0'
#158260000000
1!
b0 %
1'
b0 +
#158270000000
0!
0'
#158280000000
1!
1$
b1 %
1'
1*
b1 +
#158290000000
0!
0'
#158300000000
1!
b10 %
1'
b10 +
#158310000000
0!
0'
#158320000000
1!
b11 %
1'
b11 +
#158330000000
0!
0'
#158340000000
1!
b100 %
1'
b100 +
#158350000000
0!
0'
#158360000000
1!
b101 %
1'
b101 +
#158370000000
0!
0'
#158380000000
1!
0$
b110 %
1'
0*
b110 +
#158390000000
0!
0'
#158400000000
1!
b111 %
1'
b111 +
#158410000000
0!
0'
#158420000000
1!
b1000 %
1'
b1000 +
#158430000000
0!
0'
#158440000000
1!
b1001 %
1'
b1001 +
#158450000000
1"
1(
#158460000000
0!
0"
b100 &
0'
0(
b100 ,
#158470000000
1!
b0 %
1'
b0 +
#158480000000
0!
0'
#158490000000
1!
1$
b1 %
1'
1*
b1 +
#158500000000
0!
0'
#158510000000
1!
b10 %
1'
b10 +
#158520000000
0!
0'
#158530000000
1!
b11 %
1'
b11 +
#158540000000
0!
0'
#158550000000
1!
b100 %
1'
b100 +
#158560000000
0!
0'
#158570000000
1!
b101 %
1'
b101 +
#158580000000
0!
0'
#158590000000
1!
b110 %
1'
b110 +
#158600000000
0!
0'
#158610000000
1!
b111 %
1'
b111 +
#158620000000
0!
0'
#158630000000
1!
0$
b1000 %
1'
0*
b1000 +
#158640000000
0!
0'
#158650000000
1!
b1001 %
1'
b1001 +
#158660000000
0!
0'
#158670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#158680000000
0!
0'
#158690000000
1!
1$
b1 %
1'
1*
b1 +
#158700000000
0!
0'
#158710000000
1!
b10 %
1'
b10 +
#158720000000
0!
0'
#158730000000
1!
b11 %
1'
b11 +
#158740000000
0!
0'
#158750000000
1!
b100 %
1'
b100 +
#158760000000
0!
0'
#158770000000
1!
b101 %
1'
b101 +
#158780000000
0!
0'
#158790000000
1!
0$
b110 %
1'
0*
b110 +
#158800000000
0!
0'
#158810000000
1!
b111 %
1'
b111 +
#158820000000
0!
0'
#158830000000
1!
b1000 %
1'
b1000 +
#158840000000
0!
0'
#158850000000
1!
b1001 %
1'
b1001 +
#158860000000
0!
0'
#158870000000
1!
b0 %
1'
b0 +
#158880000000
1"
1(
#158890000000
0!
0"
b100 &
0'
0(
b100 ,
#158900000000
1!
1$
b1 %
1'
1*
b1 +
#158910000000
0!
0'
#158920000000
1!
b10 %
1'
b10 +
#158930000000
0!
0'
#158940000000
1!
b11 %
1'
b11 +
#158950000000
0!
0'
#158960000000
1!
b100 %
1'
b100 +
#158970000000
0!
0'
#158980000000
1!
b101 %
1'
b101 +
#158990000000
0!
0'
#159000000000
1!
b110 %
1'
b110 +
#159010000000
0!
0'
#159020000000
1!
b111 %
1'
b111 +
#159030000000
0!
0'
#159040000000
1!
0$
b1000 %
1'
0*
b1000 +
#159050000000
0!
0'
#159060000000
1!
b1001 %
1'
b1001 +
#159070000000
0!
0'
#159080000000
1!
b0 %
1'
b0 +
#159090000000
0!
0'
#159100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#159110000000
0!
0'
#159120000000
1!
b10 %
1'
b10 +
#159130000000
0!
0'
#159140000000
1!
b11 %
1'
b11 +
#159150000000
0!
0'
#159160000000
1!
b100 %
1'
b100 +
#159170000000
0!
0'
#159180000000
1!
b101 %
1'
b101 +
#159190000000
0!
0'
#159200000000
1!
0$
b110 %
1'
0*
b110 +
#159210000000
0!
0'
#159220000000
1!
b111 %
1'
b111 +
#159230000000
0!
0'
#159240000000
1!
b1000 %
1'
b1000 +
#159250000000
0!
0'
#159260000000
1!
b1001 %
1'
b1001 +
#159270000000
0!
0'
#159280000000
1!
b0 %
1'
b0 +
#159290000000
0!
0'
#159300000000
1!
1$
b1 %
1'
1*
b1 +
#159310000000
1"
1(
#159320000000
0!
0"
b100 &
0'
0(
b100 ,
#159330000000
1!
b10 %
1'
b10 +
#159340000000
0!
0'
#159350000000
1!
b11 %
1'
b11 +
#159360000000
0!
0'
#159370000000
1!
b100 %
1'
b100 +
#159380000000
0!
0'
#159390000000
1!
b101 %
1'
b101 +
#159400000000
0!
0'
#159410000000
1!
b110 %
1'
b110 +
#159420000000
0!
0'
#159430000000
1!
b111 %
1'
b111 +
#159440000000
0!
0'
#159450000000
1!
0$
b1000 %
1'
0*
b1000 +
#159460000000
0!
0'
#159470000000
1!
b1001 %
1'
b1001 +
#159480000000
0!
0'
#159490000000
1!
b0 %
1'
b0 +
#159500000000
0!
0'
#159510000000
1!
1$
b1 %
1'
1*
b1 +
#159520000000
0!
0'
#159530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#159540000000
0!
0'
#159550000000
1!
b11 %
1'
b11 +
#159560000000
0!
0'
#159570000000
1!
b100 %
1'
b100 +
#159580000000
0!
0'
#159590000000
1!
b101 %
1'
b101 +
#159600000000
0!
0'
#159610000000
1!
0$
b110 %
1'
0*
b110 +
#159620000000
0!
0'
#159630000000
1!
b111 %
1'
b111 +
#159640000000
0!
0'
#159650000000
1!
b1000 %
1'
b1000 +
#159660000000
0!
0'
#159670000000
1!
b1001 %
1'
b1001 +
#159680000000
0!
0'
#159690000000
1!
b0 %
1'
b0 +
#159700000000
0!
0'
#159710000000
1!
1$
b1 %
1'
1*
b1 +
#159720000000
0!
0'
#159730000000
1!
b10 %
1'
b10 +
#159740000000
1"
1(
#159750000000
0!
0"
b100 &
0'
0(
b100 ,
#159760000000
1!
b11 %
1'
b11 +
#159770000000
0!
0'
#159780000000
1!
b100 %
1'
b100 +
#159790000000
0!
0'
#159800000000
1!
b101 %
1'
b101 +
#159810000000
0!
0'
#159820000000
1!
b110 %
1'
b110 +
#159830000000
0!
0'
#159840000000
1!
b111 %
1'
b111 +
#159850000000
0!
0'
#159860000000
1!
0$
b1000 %
1'
0*
b1000 +
#159870000000
0!
0'
#159880000000
1!
b1001 %
1'
b1001 +
#159890000000
0!
0'
#159900000000
1!
b0 %
1'
b0 +
#159910000000
0!
0'
#159920000000
1!
1$
b1 %
1'
1*
b1 +
#159930000000
0!
0'
#159940000000
1!
b10 %
1'
b10 +
#159950000000
0!
0'
#159960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#159970000000
0!
0'
#159980000000
1!
b100 %
1'
b100 +
#159990000000
0!
0'
#160000000000
1!
b101 %
1'
b101 +
#160010000000
0!
0'
#160020000000
1!
0$
b110 %
1'
0*
b110 +
#160030000000
0!
0'
#160040000000
1!
b111 %
1'
b111 +
#160050000000
0!
0'
#160060000000
1!
b1000 %
1'
b1000 +
#160070000000
0!
0'
#160080000000
1!
b1001 %
1'
b1001 +
#160090000000
0!
0'
#160100000000
1!
b0 %
1'
b0 +
#160110000000
0!
0'
#160120000000
1!
1$
b1 %
1'
1*
b1 +
#160130000000
0!
0'
#160140000000
1!
b10 %
1'
b10 +
#160150000000
0!
0'
#160160000000
1!
b11 %
1'
b11 +
#160170000000
1"
1(
#160180000000
0!
0"
b100 &
0'
0(
b100 ,
#160190000000
1!
b100 %
1'
b100 +
#160200000000
0!
0'
#160210000000
1!
b101 %
1'
b101 +
#160220000000
0!
0'
#160230000000
1!
b110 %
1'
b110 +
#160240000000
0!
0'
#160250000000
1!
b111 %
1'
b111 +
#160260000000
0!
0'
#160270000000
1!
0$
b1000 %
1'
0*
b1000 +
#160280000000
0!
0'
#160290000000
1!
b1001 %
1'
b1001 +
#160300000000
0!
0'
#160310000000
1!
b0 %
1'
b0 +
#160320000000
0!
0'
#160330000000
1!
1$
b1 %
1'
1*
b1 +
#160340000000
0!
0'
#160350000000
1!
b10 %
1'
b10 +
#160360000000
0!
0'
#160370000000
1!
b11 %
1'
b11 +
#160380000000
0!
0'
#160390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#160400000000
0!
0'
#160410000000
1!
b101 %
1'
b101 +
#160420000000
0!
0'
#160430000000
1!
0$
b110 %
1'
0*
b110 +
#160440000000
0!
0'
#160450000000
1!
b111 %
1'
b111 +
#160460000000
0!
0'
#160470000000
1!
b1000 %
1'
b1000 +
#160480000000
0!
0'
#160490000000
1!
b1001 %
1'
b1001 +
#160500000000
0!
0'
#160510000000
1!
b0 %
1'
b0 +
#160520000000
0!
0'
#160530000000
1!
1$
b1 %
1'
1*
b1 +
#160540000000
0!
0'
#160550000000
1!
b10 %
1'
b10 +
#160560000000
0!
0'
#160570000000
1!
b11 %
1'
b11 +
#160580000000
0!
0'
#160590000000
1!
b100 %
1'
b100 +
#160600000000
1"
1(
#160610000000
0!
0"
b100 &
0'
0(
b100 ,
#160620000000
1!
b101 %
1'
b101 +
#160630000000
0!
0'
#160640000000
1!
b110 %
1'
b110 +
#160650000000
0!
0'
#160660000000
1!
b111 %
1'
b111 +
#160670000000
0!
0'
#160680000000
1!
0$
b1000 %
1'
0*
b1000 +
#160690000000
0!
0'
#160700000000
1!
b1001 %
1'
b1001 +
#160710000000
0!
0'
#160720000000
1!
b0 %
1'
b0 +
#160730000000
0!
0'
#160740000000
1!
1$
b1 %
1'
1*
b1 +
#160750000000
0!
0'
#160760000000
1!
b10 %
1'
b10 +
#160770000000
0!
0'
#160780000000
1!
b11 %
1'
b11 +
#160790000000
0!
0'
#160800000000
1!
b100 %
1'
b100 +
#160810000000
0!
0'
#160820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#160830000000
0!
0'
#160840000000
1!
0$
b110 %
1'
0*
b110 +
#160850000000
0!
0'
#160860000000
1!
b111 %
1'
b111 +
#160870000000
0!
0'
#160880000000
1!
b1000 %
1'
b1000 +
#160890000000
0!
0'
#160900000000
1!
b1001 %
1'
b1001 +
#160910000000
0!
0'
#160920000000
1!
b0 %
1'
b0 +
#160930000000
0!
0'
#160940000000
1!
1$
b1 %
1'
1*
b1 +
#160950000000
0!
0'
#160960000000
1!
b10 %
1'
b10 +
#160970000000
0!
0'
#160980000000
1!
b11 %
1'
b11 +
#160990000000
0!
0'
#161000000000
1!
b100 %
1'
b100 +
#161010000000
0!
0'
#161020000000
1!
b101 %
1'
b101 +
#161030000000
1"
1(
#161040000000
0!
0"
b100 &
0'
0(
b100 ,
#161050000000
1!
b110 %
1'
b110 +
#161060000000
0!
0'
#161070000000
1!
b111 %
1'
b111 +
#161080000000
0!
0'
#161090000000
1!
0$
b1000 %
1'
0*
b1000 +
#161100000000
0!
0'
#161110000000
1!
b1001 %
1'
b1001 +
#161120000000
0!
0'
#161130000000
1!
b0 %
1'
b0 +
#161140000000
0!
0'
#161150000000
1!
1$
b1 %
1'
1*
b1 +
#161160000000
0!
0'
#161170000000
1!
b10 %
1'
b10 +
#161180000000
0!
0'
#161190000000
1!
b11 %
1'
b11 +
#161200000000
0!
0'
#161210000000
1!
b100 %
1'
b100 +
#161220000000
0!
0'
#161230000000
1!
b101 %
1'
b101 +
#161240000000
0!
0'
#161250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#161260000000
0!
0'
#161270000000
1!
b111 %
1'
b111 +
#161280000000
0!
0'
#161290000000
1!
b1000 %
1'
b1000 +
#161300000000
0!
0'
#161310000000
1!
b1001 %
1'
b1001 +
#161320000000
0!
0'
#161330000000
1!
b0 %
1'
b0 +
#161340000000
0!
0'
#161350000000
1!
1$
b1 %
1'
1*
b1 +
#161360000000
0!
0'
#161370000000
1!
b10 %
1'
b10 +
#161380000000
0!
0'
#161390000000
1!
b11 %
1'
b11 +
#161400000000
0!
0'
#161410000000
1!
b100 %
1'
b100 +
#161420000000
0!
0'
#161430000000
1!
b101 %
1'
b101 +
#161440000000
0!
0'
#161450000000
1!
0$
b110 %
1'
0*
b110 +
#161460000000
1"
1(
#161470000000
0!
0"
b100 &
0'
0(
b100 ,
#161480000000
1!
1$
b111 %
1'
1*
b111 +
#161490000000
0!
0'
#161500000000
1!
0$
b1000 %
1'
0*
b1000 +
#161510000000
0!
0'
#161520000000
1!
b1001 %
1'
b1001 +
#161530000000
0!
0'
#161540000000
1!
b0 %
1'
b0 +
#161550000000
0!
0'
#161560000000
1!
1$
b1 %
1'
1*
b1 +
#161570000000
0!
0'
#161580000000
1!
b10 %
1'
b10 +
#161590000000
0!
0'
#161600000000
1!
b11 %
1'
b11 +
#161610000000
0!
0'
#161620000000
1!
b100 %
1'
b100 +
#161630000000
0!
0'
#161640000000
1!
b101 %
1'
b101 +
#161650000000
0!
0'
#161660000000
1!
b110 %
1'
b110 +
#161670000000
0!
0'
#161680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#161690000000
0!
0'
#161700000000
1!
b1000 %
1'
b1000 +
#161710000000
0!
0'
#161720000000
1!
b1001 %
1'
b1001 +
#161730000000
0!
0'
#161740000000
1!
b0 %
1'
b0 +
#161750000000
0!
0'
#161760000000
1!
1$
b1 %
1'
1*
b1 +
#161770000000
0!
0'
#161780000000
1!
b10 %
1'
b10 +
#161790000000
0!
0'
#161800000000
1!
b11 %
1'
b11 +
#161810000000
0!
0'
#161820000000
1!
b100 %
1'
b100 +
#161830000000
0!
0'
#161840000000
1!
b101 %
1'
b101 +
#161850000000
0!
0'
#161860000000
1!
0$
b110 %
1'
0*
b110 +
#161870000000
0!
0'
#161880000000
1!
b111 %
1'
b111 +
#161890000000
1"
1(
#161900000000
0!
0"
b100 &
0'
0(
b100 ,
#161910000000
1!
b1000 %
1'
b1000 +
#161920000000
0!
0'
#161930000000
1!
b1001 %
1'
b1001 +
#161940000000
0!
0'
#161950000000
1!
b0 %
1'
b0 +
#161960000000
0!
0'
#161970000000
1!
1$
b1 %
1'
1*
b1 +
#161980000000
0!
0'
#161990000000
1!
b10 %
1'
b10 +
#162000000000
0!
0'
#162010000000
1!
b11 %
1'
b11 +
#162020000000
0!
0'
#162030000000
1!
b100 %
1'
b100 +
#162040000000
0!
0'
#162050000000
1!
b101 %
1'
b101 +
#162060000000
0!
0'
#162070000000
1!
b110 %
1'
b110 +
#162080000000
0!
0'
#162090000000
1!
b111 %
1'
b111 +
#162100000000
0!
0'
#162110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#162120000000
0!
0'
#162130000000
1!
b1001 %
1'
b1001 +
#162140000000
0!
0'
#162150000000
1!
b0 %
1'
b0 +
#162160000000
0!
0'
#162170000000
1!
1$
b1 %
1'
1*
b1 +
#162180000000
0!
0'
#162190000000
1!
b10 %
1'
b10 +
#162200000000
0!
0'
#162210000000
1!
b11 %
1'
b11 +
#162220000000
0!
0'
#162230000000
1!
b100 %
1'
b100 +
#162240000000
0!
0'
#162250000000
1!
b101 %
1'
b101 +
#162260000000
0!
0'
#162270000000
1!
0$
b110 %
1'
0*
b110 +
#162280000000
0!
0'
#162290000000
1!
b111 %
1'
b111 +
#162300000000
0!
0'
#162310000000
1!
b1000 %
1'
b1000 +
#162320000000
1"
1(
#162330000000
0!
0"
b100 &
0'
0(
b100 ,
#162340000000
1!
b1001 %
1'
b1001 +
#162350000000
0!
0'
#162360000000
1!
b0 %
1'
b0 +
#162370000000
0!
0'
#162380000000
1!
1$
b1 %
1'
1*
b1 +
#162390000000
0!
0'
#162400000000
1!
b10 %
1'
b10 +
#162410000000
0!
0'
#162420000000
1!
b11 %
1'
b11 +
#162430000000
0!
0'
#162440000000
1!
b100 %
1'
b100 +
#162450000000
0!
0'
#162460000000
1!
b101 %
1'
b101 +
#162470000000
0!
0'
#162480000000
1!
b110 %
1'
b110 +
#162490000000
0!
0'
#162500000000
1!
b111 %
1'
b111 +
#162510000000
0!
0'
#162520000000
1!
0$
b1000 %
1'
0*
b1000 +
#162530000000
0!
0'
#162540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#162550000000
0!
0'
#162560000000
1!
b0 %
1'
b0 +
#162570000000
0!
0'
#162580000000
1!
1$
b1 %
1'
1*
b1 +
#162590000000
0!
0'
#162600000000
1!
b10 %
1'
b10 +
#162610000000
0!
0'
#162620000000
1!
b11 %
1'
b11 +
#162630000000
0!
0'
#162640000000
1!
b100 %
1'
b100 +
#162650000000
0!
0'
#162660000000
1!
b101 %
1'
b101 +
#162670000000
0!
0'
#162680000000
1!
0$
b110 %
1'
0*
b110 +
#162690000000
0!
0'
#162700000000
1!
b111 %
1'
b111 +
#162710000000
0!
0'
#162720000000
1!
b1000 %
1'
b1000 +
#162730000000
0!
0'
#162740000000
1!
b1001 %
1'
b1001 +
#162750000000
1"
1(
#162760000000
0!
0"
b100 &
0'
0(
b100 ,
#162770000000
1!
b0 %
1'
b0 +
#162780000000
0!
0'
#162790000000
1!
1$
b1 %
1'
1*
b1 +
#162800000000
0!
0'
#162810000000
1!
b10 %
1'
b10 +
#162820000000
0!
0'
#162830000000
1!
b11 %
1'
b11 +
#162840000000
0!
0'
#162850000000
1!
b100 %
1'
b100 +
#162860000000
0!
0'
#162870000000
1!
b101 %
1'
b101 +
#162880000000
0!
0'
#162890000000
1!
b110 %
1'
b110 +
#162900000000
0!
0'
#162910000000
1!
b111 %
1'
b111 +
#162920000000
0!
0'
#162930000000
1!
0$
b1000 %
1'
0*
b1000 +
#162940000000
0!
0'
#162950000000
1!
b1001 %
1'
b1001 +
#162960000000
0!
0'
#162970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#162980000000
0!
0'
#162990000000
1!
1$
b1 %
1'
1*
b1 +
#163000000000
0!
0'
#163010000000
1!
b10 %
1'
b10 +
#163020000000
0!
0'
#163030000000
1!
b11 %
1'
b11 +
#163040000000
0!
0'
#163050000000
1!
b100 %
1'
b100 +
#163060000000
0!
0'
#163070000000
1!
b101 %
1'
b101 +
#163080000000
0!
0'
#163090000000
1!
0$
b110 %
1'
0*
b110 +
#163100000000
0!
0'
#163110000000
1!
b111 %
1'
b111 +
#163120000000
0!
0'
#163130000000
1!
b1000 %
1'
b1000 +
#163140000000
0!
0'
#163150000000
1!
b1001 %
1'
b1001 +
#163160000000
0!
0'
#163170000000
1!
b0 %
1'
b0 +
#163180000000
1"
1(
#163190000000
0!
0"
b100 &
0'
0(
b100 ,
#163200000000
1!
1$
b1 %
1'
1*
b1 +
#163210000000
0!
0'
#163220000000
1!
b10 %
1'
b10 +
#163230000000
0!
0'
#163240000000
1!
b11 %
1'
b11 +
#163250000000
0!
0'
#163260000000
1!
b100 %
1'
b100 +
#163270000000
0!
0'
#163280000000
1!
b101 %
1'
b101 +
#163290000000
0!
0'
#163300000000
1!
b110 %
1'
b110 +
#163310000000
0!
0'
#163320000000
1!
b111 %
1'
b111 +
#163330000000
0!
0'
#163340000000
1!
0$
b1000 %
1'
0*
b1000 +
#163350000000
0!
0'
#163360000000
1!
b1001 %
1'
b1001 +
#163370000000
0!
0'
#163380000000
1!
b0 %
1'
b0 +
#163390000000
0!
0'
#163400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#163410000000
0!
0'
#163420000000
1!
b10 %
1'
b10 +
#163430000000
0!
0'
#163440000000
1!
b11 %
1'
b11 +
#163450000000
0!
0'
#163460000000
1!
b100 %
1'
b100 +
#163470000000
0!
0'
#163480000000
1!
b101 %
1'
b101 +
#163490000000
0!
0'
#163500000000
1!
0$
b110 %
1'
0*
b110 +
#163510000000
0!
0'
#163520000000
1!
b111 %
1'
b111 +
#163530000000
0!
0'
#163540000000
1!
b1000 %
1'
b1000 +
#163550000000
0!
0'
#163560000000
1!
b1001 %
1'
b1001 +
#163570000000
0!
0'
#163580000000
1!
b0 %
1'
b0 +
#163590000000
0!
0'
#163600000000
1!
1$
b1 %
1'
1*
b1 +
#163610000000
1"
1(
#163620000000
0!
0"
b100 &
0'
0(
b100 ,
#163630000000
1!
b10 %
1'
b10 +
#163640000000
0!
0'
#163650000000
1!
b11 %
1'
b11 +
#163660000000
0!
0'
#163670000000
1!
b100 %
1'
b100 +
#163680000000
0!
0'
#163690000000
1!
b101 %
1'
b101 +
#163700000000
0!
0'
#163710000000
1!
b110 %
1'
b110 +
#163720000000
0!
0'
#163730000000
1!
b111 %
1'
b111 +
#163740000000
0!
0'
#163750000000
1!
0$
b1000 %
1'
0*
b1000 +
#163760000000
0!
0'
#163770000000
1!
b1001 %
1'
b1001 +
#163780000000
0!
0'
#163790000000
1!
b0 %
1'
b0 +
#163800000000
0!
0'
#163810000000
1!
1$
b1 %
1'
1*
b1 +
#163820000000
0!
0'
#163830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#163840000000
0!
0'
#163850000000
1!
b11 %
1'
b11 +
#163860000000
0!
0'
#163870000000
1!
b100 %
1'
b100 +
#163880000000
0!
0'
#163890000000
1!
b101 %
1'
b101 +
#163900000000
0!
0'
#163910000000
1!
0$
b110 %
1'
0*
b110 +
#163920000000
0!
0'
#163930000000
1!
b111 %
1'
b111 +
#163940000000
0!
0'
#163950000000
1!
b1000 %
1'
b1000 +
#163960000000
0!
0'
#163970000000
1!
b1001 %
1'
b1001 +
#163980000000
0!
0'
#163990000000
1!
b0 %
1'
b0 +
#164000000000
0!
0'
#164010000000
1!
1$
b1 %
1'
1*
b1 +
#164020000000
0!
0'
#164030000000
1!
b10 %
1'
b10 +
#164040000000
1"
1(
#164050000000
0!
0"
b100 &
0'
0(
b100 ,
#164060000000
1!
b11 %
1'
b11 +
#164070000000
0!
0'
#164080000000
1!
b100 %
1'
b100 +
#164090000000
0!
0'
#164100000000
1!
b101 %
1'
b101 +
#164110000000
0!
0'
#164120000000
1!
b110 %
1'
b110 +
#164130000000
0!
0'
#164140000000
1!
b111 %
1'
b111 +
#164150000000
0!
0'
#164160000000
1!
0$
b1000 %
1'
0*
b1000 +
#164170000000
0!
0'
#164180000000
1!
b1001 %
1'
b1001 +
#164190000000
0!
0'
#164200000000
1!
b0 %
1'
b0 +
#164210000000
0!
0'
#164220000000
1!
1$
b1 %
1'
1*
b1 +
#164230000000
0!
0'
#164240000000
1!
b10 %
1'
b10 +
#164250000000
0!
0'
#164260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#164270000000
0!
0'
#164280000000
1!
b100 %
1'
b100 +
#164290000000
0!
0'
#164300000000
1!
b101 %
1'
b101 +
#164310000000
0!
0'
#164320000000
1!
0$
b110 %
1'
0*
b110 +
#164330000000
0!
0'
#164340000000
1!
b111 %
1'
b111 +
#164350000000
0!
0'
#164360000000
1!
b1000 %
1'
b1000 +
#164370000000
0!
0'
#164380000000
1!
b1001 %
1'
b1001 +
#164390000000
0!
0'
#164400000000
1!
b0 %
1'
b0 +
#164410000000
0!
0'
#164420000000
1!
1$
b1 %
1'
1*
b1 +
#164430000000
0!
0'
#164440000000
1!
b10 %
1'
b10 +
#164450000000
0!
0'
#164460000000
1!
b11 %
1'
b11 +
#164470000000
1"
1(
#164480000000
0!
0"
b100 &
0'
0(
b100 ,
#164490000000
1!
b100 %
1'
b100 +
#164500000000
0!
0'
#164510000000
1!
b101 %
1'
b101 +
#164520000000
0!
0'
#164530000000
1!
b110 %
1'
b110 +
#164540000000
0!
0'
#164550000000
1!
b111 %
1'
b111 +
#164560000000
0!
0'
#164570000000
1!
0$
b1000 %
1'
0*
b1000 +
#164580000000
0!
0'
#164590000000
1!
b1001 %
1'
b1001 +
#164600000000
0!
0'
#164610000000
1!
b0 %
1'
b0 +
#164620000000
0!
0'
#164630000000
1!
1$
b1 %
1'
1*
b1 +
#164640000000
0!
0'
#164650000000
1!
b10 %
1'
b10 +
#164660000000
0!
0'
#164670000000
1!
b11 %
1'
b11 +
#164680000000
0!
0'
#164690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#164700000000
0!
0'
#164710000000
1!
b101 %
1'
b101 +
#164720000000
0!
0'
#164730000000
1!
0$
b110 %
1'
0*
b110 +
#164740000000
0!
0'
#164750000000
1!
b111 %
1'
b111 +
#164760000000
0!
0'
#164770000000
1!
b1000 %
1'
b1000 +
#164780000000
0!
0'
#164790000000
1!
b1001 %
1'
b1001 +
#164800000000
0!
0'
#164810000000
1!
b0 %
1'
b0 +
#164820000000
0!
0'
#164830000000
1!
1$
b1 %
1'
1*
b1 +
#164840000000
0!
0'
#164850000000
1!
b10 %
1'
b10 +
#164860000000
0!
0'
#164870000000
1!
b11 %
1'
b11 +
#164880000000
0!
0'
#164890000000
1!
b100 %
1'
b100 +
#164900000000
1"
1(
#164910000000
0!
0"
b100 &
0'
0(
b100 ,
#164920000000
1!
b101 %
1'
b101 +
#164930000000
0!
0'
#164940000000
1!
b110 %
1'
b110 +
#164950000000
0!
0'
#164960000000
1!
b111 %
1'
b111 +
#164970000000
0!
0'
#164980000000
1!
0$
b1000 %
1'
0*
b1000 +
#164990000000
0!
0'
#165000000000
1!
b1001 %
1'
b1001 +
#165010000000
0!
0'
#165020000000
1!
b0 %
1'
b0 +
#165030000000
0!
0'
#165040000000
1!
1$
b1 %
1'
1*
b1 +
#165050000000
0!
0'
#165060000000
1!
b10 %
1'
b10 +
#165070000000
0!
0'
#165080000000
1!
b11 %
1'
b11 +
#165090000000
0!
0'
#165100000000
1!
b100 %
1'
b100 +
#165110000000
0!
0'
#165120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#165130000000
0!
0'
#165140000000
1!
0$
b110 %
1'
0*
b110 +
#165150000000
0!
0'
#165160000000
1!
b111 %
1'
b111 +
#165170000000
0!
0'
#165180000000
1!
b1000 %
1'
b1000 +
#165190000000
0!
0'
#165200000000
1!
b1001 %
1'
b1001 +
#165210000000
0!
0'
#165220000000
1!
b0 %
1'
b0 +
#165230000000
0!
0'
#165240000000
1!
1$
b1 %
1'
1*
b1 +
#165250000000
0!
0'
#165260000000
1!
b10 %
1'
b10 +
#165270000000
0!
0'
#165280000000
1!
b11 %
1'
b11 +
#165290000000
0!
0'
#165300000000
1!
b100 %
1'
b100 +
#165310000000
0!
0'
#165320000000
1!
b101 %
1'
b101 +
#165330000000
1"
1(
#165340000000
0!
0"
b100 &
0'
0(
b100 ,
#165350000000
1!
b110 %
1'
b110 +
#165360000000
0!
0'
#165370000000
1!
b111 %
1'
b111 +
#165380000000
0!
0'
#165390000000
1!
0$
b1000 %
1'
0*
b1000 +
#165400000000
0!
0'
#165410000000
1!
b1001 %
1'
b1001 +
#165420000000
0!
0'
#165430000000
1!
b0 %
1'
b0 +
#165440000000
0!
0'
#165450000000
1!
1$
b1 %
1'
1*
b1 +
#165460000000
0!
0'
#165470000000
1!
b10 %
1'
b10 +
#165480000000
0!
0'
#165490000000
1!
b11 %
1'
b11 +
#165500000000
0!
0'
#165510000000
1!
b100 %
1'
b100 +
#165520000000
0!
0'
#165530000000
1!
b101 %
1'
b101 +
#165540000000
0!
0'
#165550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#165560000000
0!
0'
#165570000000
1!
b111 %
1'
b111 +
#165580000000
0!
0'
#165590000000
1!
b1000 %
1'
b1000 +
#165600000000
0!
0'
#165610000000
1!
b1001 %
1'
b1001 +
#165620000000
0!
0'
#165630000000
1!
b0 %
1'
b0 +
#165640000000
0!
0'
#165650000000
1!
1$
b1 %
1'
1*
b1 +
#165660000000
0!
0'
#165670000000
1!
b10 %
1'
b10 +
#165680000000
0!
0'
#165690000000
1!
b11 %
1'
b11 +
#165700000000
0!
0'
#165710000000
1!
b100 %
1'
b100 +
#165720000000
0!
0'
#165730000000
1!
b101 %
1'
b101 +
#165740000000
0!
0'
#165750000000
1!
0$
b110 %
1'
0*
b110 +
#165760000000
1"
1(
#165770000000
0!
0"
b100 &
0'
0(
b100 ,
#165780000000
1!
1$
b111 %
1'
1*
b111 +
#165790000000
0!
0'
#165800000000
1!
0$
b1000 %
1'
0*
b1000 +
#165810000000
0!
0'
#165820000000
1!
b1001 %
1'
b1001 +
#165830000000
0!
0'
#165840000000
1!
b0 %
1'
b0 +
#165850000000
0!
0'
#165860000000
1!
1$
b1 %
1'
1*
b1 +
#165870000000
0!
0'
#165880000000
1!
b10 %
1'
b10 +
#165890000000
0!
0'
#165900000000
1!
b11 %
1'
b11 +
#165910000000
0!
0'
#165920000000
1!
b100 %
1'
b100 +
#165930000000
0!
0'
#165940000000
1!
b101 %
1'
b101 +
#165950000000
0!
0'
#165960000000
1!
b110 %
1'
b110 +
#165970000000
0!
0'
#165980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#165990000000
0!
0'
#166000000000
1!
b1000 %
1'
b1000 +
#166010000000
0!
0'
#166020000000
1!
b1001 %
1'
b1001 +
#166030000000
0!
0'
#166040000000
1!
b0 %
1'
b0 +
#166050000000
0!
0'
#166060000000
1!
1$
b1 %
1'
1*
b1 +
#166070000000
0!
0'
#166080000000
1!
b10 %
1'
b10 +
#166090000000
0!
0'
#166100000000
1!
b11 %
1'
b11 +
#166110000000
0!
0'
#166120000000
1!
b100 %
1'
b100 +
#166130000000
0!
0'
#166140000000
1!
b101 %
1'
b101 +
#166150000000
0!
0'
#166160000000
1!
0$
b110 %
1'
0*
b110 +
#166170000000
0!
0'
#166180000000
1!
b111 %
1'
b111 +
#166190000000
1"
1(
#166200000000
0!
0"
b100 &
0'
0(
b100 ,
#166210000000
1!
b1000 %
1'
b1000 +
#166220000000
0!
0'
#166230000000
1!
b1001 %
1'
b1001 +
#166240000000
0!
0'
#166250000000
1!
b0 %
1'
b0 +
#166260000000
0!
0'
#166270000000
1!
1$
b1 %
1'
1*
b1 +
#166280000000
0!
0'
#166290000000
1!
b10 %
1'
b10 +
#166300000000
0!
0'
#166310000000
1!
b11 %
1'
b11 +
#166320000000
0!
0'
#166330000000
1!
b100 %
1'
b100 +
#166340000000
0!
0'
#166350000000
1!
b101 %
1'
b101 +
#166360000000
0!
0'
#166370000000
1!
b110 %
1'
b110 +
#166380000000
0!
0'
#166390000000
1!
b111 %
1'
b111 +
#166400000000
0!
0'
#166410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#166420000000
0!
0'
#166430000000
1!
b1001 %
1'
b1001 +
#166440000000
0!
0'
#166450000000
1!
b0 %
1'
b0 +
#166460000000
0!
0'
#166470000000
1!
1$
b1 %
1'
1*
b1 +
#166480000000
0!
0'
#166490000000
1!
b10 %
1'
b10 +
#166500000000
0!
0'
#166510000000
1!
b11 %
1'
b11 +
#166520000000
0!
0'
#166530000000
1!
b100 %
1'
b100 +
#166540000000
0!
0'
#166550000000
1!
b101 %
1'
b101 +
#166560000000
0!
0'
#166570000000
1!
0$
b110 %
1'
0*
b110 +
#166580000000
0!
0'
#166590000000
1!
b111 %
1'
b111 +
#166600000000
0!
0'
#166610000000
1!
b1000 %
1'
b1000 +
#166620000000
1"
1(
#166630000000
0!
0"
b100 &
0'
0(
b100 ,
#166640000000
1!
b1001 %
1'
b1001 +
#166650000000
0!
0'
#166660000000
1!
b0 %
1'
b0 +
#166670000000
0!
0'
#166680000000
1!
1$
b1 %
1'
1*
b1 +
#166690000000
0!
0'
#166700000000
1!
b10 %
1'
b10 +
#166710000000
0!
0'
#166720000000
1!
b11 %
1'
b11 +
#166730000000
0!
0'
#166740000000
1!
b100 %
1'
b100 +
#166750000000
0!
0'
#166760000000
1!
b101 %
1'
b101 +
#166770000000
0!
0'
#166780000000
1!
b110 %
1'
b110 +
#166790000000
0!
0'
#166800000000
1!
b111 %
1'
b111 +
#166810000000
0!
0'
#166820000000
1!
0$
b1000 %
1'
0*
b1000 +
#166830000000
0!
0'
#166840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#166850000000
0!
0'
#166860000000
1!
b0 %
1'
b0 +
#166870000000
0!
0'
#166880000000
1!
1$
b1 %
1'
1*
b1 +
#166890000000
0!
0'
#166900000000
1!
b10 %
1'
b10 +
#166910000000
0!
0'
#166920000000
1!
b11 %
1'
b11 +
#166930000000
0!
0'
#166940000000
1!
b100 %
1'
b100 +
#166950000000
0!
0'
#166960000000
1!
b101 %
1'
b101 +
#166970000000
0!
0'
#166980000000
1!
0$
b110 %
1'
0*
b110 +
#166990000000
0!
0'
#167000000000
1!
b111 %
1'
b111 +
#167010000000
0!
0'
#167020000000
1!
b1000 %
1'
b1000 +
#167030000000
0!
0'
#167040000000
1!
b1001 %
1'
b1001 +
#167050000000
1"
1(
#167060000000
0!
0"
b100 &
0'
0(
b100 ,
#167070000000
1!
b0 %
1'
b0 +
#167080000000
0!
0'
#167090000000
1!
1$
b1 %
1'
1*
b1 +
#167100000000
0!
0'
#167110000000
1!
b10 %
1'
b10 +
#167120000000
0!
0'
#167130000000
1!
b11 %
1'
b11 +
#167140000000
0!
0'
#167150000000
1!
b100 %
1'
b100 +
#167160000000
0!
0'
#167170000000
1!
b101 %
1'
b101 +
#167180000000
0!
0'
#167190000000
1!
b110 %
1'
b110 +
#167200000000
0!
0'
#167210000000
1!
b111 %
1'
b111 +
#167220000000
0!
0'
#167230000000
1!
0$
b1000 %
1'
0*
b1000 +
#167240000000
0!
0'
#167250000000
1!
b1001 %
1'
b1001 +
#167260000000
0!
0'
#167270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#167280000000
0!
0'
#167290000000
1!
1$
b1 %
1'
1*
b1 +
#167300000000
0!
0'
#167310000000
1!
b10 %
1'
b10 +
#167320000000
0!
0'
#167330000000
1!
b11 %
1'
b11 +
#167340000000
0!
0'
#167350000000
1!
b100 %
1'
b100 +
#167360000000
0!
0'
#167370000000
1!
b101 %
1'
b101 +
#167380000000
0!
0'
#167390000000
1!
0$
b110 %
1'
0*
b110 +
#167400000000
0!
0'
#167410000000
1!
b111 %
1'
b111 +
#167420000000
0!
0'
#167430000000
1!
b1000 %
1'
b1000 +
#167440000000
0!
0'
#167450000000
1!
b1001 %
1'
b1001 +
#167460000000
0!
0'
#167470000000
1!
b0 %
1'
b0 +
#167480000000
1"
1(
#167490000000
0!
0"
b100 &
0'
0(
b100 ,
#167500000000
1!
1$
b1 %
1'
1*
b1 +
#167510000000
0!
0'
#167520000000
1!
b10 %
1'
b10 +
#167530000000
0!
0'
#167540000000
1!
b11 %
1'
b11 +
#167550000000
0!
0'
#167560000000
1!
b100 %
1'
b100 +
#167570000000
0!
0'
#167580000000
1!
b101 %
1'
b101 +
#167590000000
0!
0'
#167600000000
1!
b110 %
1'
b110 +
#167610000000
0!
0'
#167620000000
1!
b111 %
1'
b111 +
#167630000000
0!
0'
#167640000000
1!
0$
b1000 %
1'
0*
b1000 +
#167650000000
0!
0'
#167660000000
1!
b1001 %
1'
b1001 +
#167670000000
0!
0'
#167680000000
1!
b0 %
1'
b0 +
#167690000000
0!
0'
#167700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#167710000000
0!
0'
#167720000000
1!
b10 %
1'
b10 +
#167730000000
0!
0'
#167740000000
1!
b11 %
1'
b11 +
#167750000000
0!
0'
#167760000000
1!
b100 %
1'
b100 +
#167770000000
0!
0'
#167780000000
1!
b101 %
1'
b101 +
#167790000000
0!
0'
#167800000000
1!
0$
b110 %
1'
0*
b110 +
#167810000000
0!
0'
#167820000000
1!
b111 %
1'
b111 +
#167830000000
0!
0'
#167840000000
1!
b1000 %
1'
b1000 +
#167850000000
0!
0'
#167860000000
1!
b1001 %
1'
b1001 +
#167870000000
0!
0'
#167880000000
1!
b0 %
1'
b0 +
#167890000000
0!
0'
#167900000000
1!
1$
b1 %
1'
1*
b1 +
#167910000000
1"
1(
#167920000000
0!
0"
b100 &
0'
0(
b100 ,
#167930000000
1!
b10 %
1'
b10 +
#167940000000
0!
0'
#167950000000
1!
b11 %
1'
b11 +
#167960000000
0!
0'
#167970000000
1!
b100 %
1'
b100 +
#167980000000
0!
0'
#167990000000
1!
b101 %
1'
b101 +
#168000000000
0!
0'
#168010000000
1!
b110 %
1'
b110 +
#168020000000
0!
0'
#168030000000
1!
b111 %
1'
b111 +
#168040000000
0!
0'
#168050000000
1!
0$
b1000 %
1'
0*
b1000 +
#168060000000
0!
0'
#168070000000
1!
b1001 %
1'
b1001 +
#168080000000
0!
0'
#168090000000
1!
b0 %
1'
b0 +
#168100000000
0!
0'
#168110000000
1!
1$
b1 %
1'
1*
b1 +
#168120000000
0!
0'
#168130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#168140000000
0!
0'
#168150000000
1!
b11 %
1'
b11 +
#168160000000
0!
0'
#168170000000
1!
b100 %
1'
b100 +
#168180000000
0!
0'
#168190000000
1!
b101 %
1'
b101 +
#168200000000
0!
0'
#168210000000
1!
0$
b110 %
1'
0*
b110 +
#168220000000
0!
0'
#168230000000
1!
b111 %
1'
b111 +
#168240000000
0!
0'
#168250000000
1!
b1000 %
1'
b1000 +
#168260000000
0!
0'
#168270000000
1!
b1001 %
1'
b1001 +
#168280000000
0!
0'
#168290000000
1!
b0 %
1'
b0 +
#168300000000
0!
0'
#168310000000
1!
1$
b1 %
1'
1*
b1 +
#168320000000
0!
0'
#168330000000
1!
b10 %
1'
b10 +
#168340000000
1"
1(
#168350000000
0!
0"
b100 &
0'
0(
b100 ,
#168360000000
1!
b11 %
1'
b11 +
#168370000000
0!
0'
#168380000000
1!
b100 %
1'
b100 +
#168390000000
0!
0'
#168400000000
1!
b101 %
1'
b101 +
#168410000000
0!
0'
#168420000000
1!
b110 %
1'
b110 +
#168430000000
0!
0'
#168440000000
1!
b111 %
1'
b111 +
#168450000000
0!
0'
#168460000000
1!
0$
b1000 %
1'
0*
b1000 +
#168470000000
0!
0'
#168480000000
1!
b1001 %
1'
b1001 +
#168490000000
0!
0'
#168500000000
1!
b0 %
1'
b0 +
#168510000000
0!
0'
#168520000000
1!
1$
b1 %
1'
1*
b1 +
#168530000000
0!
0'
#168540000000
1!
b10 %
1'
b10 +
#168550000000
0!
0'
#168560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#168570000000
0!
0'
#168580000000
1!
b100 %
1'
b100 +
#168590000000
0!
0'
#168600000000
1!
b101 %
1'
b101 +
#168610000000
0!
0'
#168620000000
1!
0$
b110 %
1'
0*
b110 +
#168630000000
0!
0'
#168640000000
1!
b111 %
1'
b111 +
#168650000000
0!
0'
#168660000000
1!
b1000 %
1'
b1000 +
#168670000000
0!
0'
#168680000000
1!
b1001 %
1'
b1001 +
#168690000000
0!
0'
#168700000000
1!
b0 %
1'
b0 +
#168710000000
0!
0'
#168720000000
1!
1$
b1 %
1'
1*
b1 +
#168730000000
0!
0'
#168740000000
1!
b10 %
1'
b10 +
#168750000000
0!
0'
#168760000000
1!
b11 %
1'
b11 +
#168770000000
1"
1(
#168780000000
0!
0"
b100 &
0'
0(
b100 ,
#168790000000
1!
b100 %
1'
b100 +
#168800000000
0!
0'
#168810000000
1!
b101 %
1'
b101 +
#168820000000
0!
0'
#168830000000
1!
b110 %
1'
b110 +
#168840000000
0!
0'
#168850000000
1!
b111 %
1'
b111 +
#168860000000
0!
0'
#168870000000
1!
0$
b1000 %
1'
0*
b1000 +
#168880000000
0!
0'
#168890000000
1!
b1001 %
1'
b1001 +
#168900000000
0!
0'
#168910000000
1!
b0 %
1'
b0 +
#168920000000
0!
0'
#168930000000
1!
1$
b1 %
1'
1*
b1 +
#168940000000
0!
0'
#168950000000
1!
b10 %
1'
b10 +
#168960000000
0!
0'
#168970000000
1!
b11 %
1'
b11 +
#168980000000
0!
0'
#168990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#169000000000
0!
0'
#169010000000
1!
b101 %
1'
b101 +
#169020000000
0!
0'
#169030000000
1!
0$
b110 %
1'
0*
b110 +
#169040000000
0!
0'
#169050000000
1!
b111 %
1'
b111 +
#169060000000
0!
0'
#169070000000
1!
b1000 %
1'
b1000 +
#169080000000
0!
0'
#169090000000
1!
b1001 %
1'
b1001 +
#169100000000
0!
0'
#169110000000
1!
b0 %
1'
b0 +
#169120000000
0!
0'
#169130000000
1!
1$
b1 %
1'
1*
b1 +
#169140000000
0!
0'
#169150000000
1!
b10 %
1'
b10 +
#169160000000
0!
0'
#169170000000
1!
b11 %
1'
b11 +
#169180000000
0!
0'
#169190000000
1!
b100 %
1'
b100 +
#169200000000
1"
1(
#169210000000
0!
0"
b100 &
0'
0(
b100 ,
#169220000000
1!
b101 %
1'
b101 +
#169230000000
0!
0'
#169240000000
1!
b110 %
1'
b110 +
#169250000000
0!
0'
#169260000000
1!
b111 %
1'
b111 +
#169270000000
0!
0'
#169280000000
1!
0$
b1000 %
1'
0*
b1000 +
#169290000000
0!
0'
#169300000000
1!
b1001 %
1'
b1001 +
#169310000000
0!
0'
#169320000000
1!
b0 %
1'
b0 +
#169330000000
0!
0'
#169340000000
1!
1$
b1 %
1'
1*
b1 +
#169350000000
0!
0'
#169360000000
1!
b10 %
1'
b10 +
#169370000000
0!
0'
#169380000000
1!
b11 %
1'
b11 +
#169390000000
0!
0'
#169400000000
1!
b100 %
1'
b100 +
#169410000000
0!
0'
#169420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#169430000000
0!
0'
#169440000000
1!
0$
b110 %
1'
0*
b110 +
#169450000000
0!
0'
#169460000000
1!
b111 %
1'
b111 +
#169470000000
0!
0'
#169480000000
1!
b1000 %
1'
b1000 +
#169490000000
0!
0'
#169500000000
1!
b1001 %
1'
b1001 +
#169510000000
0!
0'
#169520000000
1!
b0 %
1'
b0 +
#169530000000
0!
0'
#169540000000
1!
1$
b1 %
1'
1*
b1 +
#169550000000
0!
0'
#169560000000
1!
b10 %
1'
b10 +
#169570000000
0!
0'
#169580000000
1!
b11 %
1'
b11 +
#169590000000
0!
0'
#169600000000
1!
b100 %
1'
b100 +
#169610000000
0!
0'
#169620000000
1!
b101 %
1'
b101 +
#169630000000
1"
1(
#169640000000
0!
0"
b100 &
0'
0(
b100 ,
#169650000000
1!
b110 %
1'
b110 +
#169660000000
0!
0'
#169670000000
1!
b111 %
1'
b111 +
#169680000000
0!
0'
#169690000000
1!
0$
b1000 %
1'
0*
b1000 +
#169700000000
0!
0'
#169710000000
1!
b1001 %
1'
b1001 +
#169720000000
0!
0'
#169730000000
1!
b0 %
1'
b0 +
#169740000000
0!
0'
#169750000000
1!
1$
b1 %
1'
1*
b1 +
#169760000000
0!
0'
#169770000000
1!
b10 %
1'
b10 +
#169780000000
0!
0'
#169790000000
1!
b11 %
1'
b11 +
#169800000000
0!
0'
#169810000000
1!
b100 %
1'
b100 +
#169820000000
0!
0'
#169830000000
1!
b101 %
1'
b101 +
#169840000000
0!
0'
#169850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#169860000000
0!
0'
#169870000000
1!
b111 %
1'
b111 +
#169880000000
0!
0'
#169890000000
1!
b1000 %
1'
b1000 +
#169900000000
0!
0'
#169910000000
1!
b1001 %
1'
b1001 +
#169920000000
0!
0'
#169930000000
1!
b0 %
1'
b0 +
#169940000000
0!
0'
#169950000000
1!
1$
b1 %
1'
1*
b1 +
#169960000000
0!
0'
#169970000000
1!
b10 %
1'
b10 +
#169980000000
0!
0'
#169990000000
1!
b11 %
1'
b11 +
#170000000000
0!
0'
#170010000000
1!
b100 %
1'
b100 +
#170020000000
0!
0'
#170030000000
1!
b101 %
1'
b101 +
#170040000000
0!
0'
#170050000000
1!
0$
b110 %
1'
0*
b110 +
#170060000000
1"
1(
#170070000000
0!
0"
b100 &
0'
0(
b100 ,
#170080000000
1!
1$
b111 %
1'
1*
b111 +
#170090000000
0!
0'
#170100000000
1!
0$
b1000 %
1'
0*
b1000 +
#170110000000
0!
0'
#170120000000
1!
b1001 %
1'
b1001 +
#170130000000
0!
0'
#170140000000
1!
b0 %
1'
b0 +
#170150000000
0!
0'
#170160000000
1!
1$
b1 %
1'
1*
b1 +
#170170000000
0!
0'
#170180000000
1!
b10 %
1'
b10 +
#170190000000
0!
0'
#170200000000
1!
b11 %
1'
b11 +
#170210000000
0!
0'
#170220000000
1!
b100 %
1'
b100 +
#170230000000
0!
0'
#170240000000
1!
b101 %
1'
b101 +
#170250000000
0!
0'
#170260000000
1!
b110 %
1'
b110 +
#170270000000
0!
0'
#170280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#170290000000
0!
0'
#170300000000
1!
b1000 %
1'
b1000 +
#170310000000
0!
0'
#170320000000
1!
b1001 %
1'
b1001 +
#170330000000
0!
0'
#170340000000
1!
b0 %
1'
b0 +
#170350000000
0!
0'
#170360000000
1!
1$
b1 %
1'
1*
b1 +
#170370000000
0!
0'
#170380000000
1!
b10 %
1'
b10 +
#170390000000
0!
0'
#170400000000
1!
b11 %
1'
b11 +
#170410000000
0!
0'
#170420000000
1!
b100 %
1'
b100 +
#170430000000
0!
0'
#170440000000
1!
b101 %
1'
b101 +
#170450000000
0!
0'
#170460000000
1!
0$
b110 %
1'
0*
b110 +
#170470000000
0!
0'
#170480000000
1!
b111 %
1'
b111 +
#170490000000
1"
1(
#170500000000
0!
0"
b100 &
0'
0(
b100 ,
#170510000000
1!
b1000 %
1'
b1000 +
#170520000000
0!
0'
#170530000000
1!
b1001 %
1'
b1001 +
#170540000000
0!
0'
#170550000000
1!
b0 %
1'
b0 +
#170560000000
0!
0'
#170570000000
1!
1$
b1 %
1'
1*
b1 +
#170580000000
0!
0'
#170590000000
1!
b10 %
1'
b10 +
#170600000000
0!
0'
#170610000000
1!
b11 %
1'
b11 +
#170620000000
0!
0'
#170630000000
1!
b100 %
1'
b100 +
#170640000000
0!
0'
#170650000000
1!
b101 %
1'
b101 +
#170660000000
0!
0'
#170670000000
1!
b110 %
1'
b110 +
#170680000000
0!
0'
#170690000000
1!
b111 %
1'
b111 +
#170700000000
0!
0'
#170710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#170720000000
0!
0'
#170730000000
1!
b1001 %
1'
b1001 +
#170740000000
0!
0'
#170750000000
1!
b0 %
1'
b0 +
#170760000000
0!
0'
#170770000000
1!
1$
b1 %
1'
1*
b1 +
#170780000000
0!
0'
#170790000000
1!
b10 %
1'
b10 +
#170800000000
0!
0'
#170810000000
1!
b11 %
1'
b11 +
#170820000000
0!
0'
#170830000000
1!
b100 %
1'
b100 +
#170840000000
0!
0'
#170850000000
1!
b101 %
1'
b101 +
#170860000000
0!
0'
#170870000000
1!
0$
b110 %
1'
0*
b110 +
#170880000000
0!
0'
#170890000000
1!
b111 %
1'
b111 +
#170900000000
0!
0'
#170910000000
1!
b1000 %
1'
b1000 +
#170920000000
1"
1(
#170930000000
0!
0"
b100 &
0'
0(
b100 ,
#170940000000
1!
b1001 %
1'
b1001 +
#170950000000
0!
0'
#170960000000
1!
b0 %
1'
b0 +
#170970000000
0!
0'
#170980000000
1!
1$
b1 %
1'
1*
b1 +
#170990000000
0!
0'
#171000000000
1!
b10 %
1'
b10 +
#171010000000
0!
0'
#171020000000
1!
b11 %
1'
b11 +
#171030000000
0!
0'
#171040000000
1!
b100 %
1'
b100 +
#171050000000
0!
0'
#171060000000
1!
b101 %
1'
b101 +
#171070000000
0!
0'
#171080000000
1!
b110 %
1'
b110 +
#171090000000
0!
0'
#171100000000
1!
b111 %
1'
b111 +
#171110000000
0!
0'
#171120000000
1!
0$
b1000 %
1'
0*
b1000 +
#171130000000
0!
0'
#171140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#171150000000
0!
0'
#171160000000
1!
b0 %
1'
b0 +
#171170000000
0!
0'
#171180000000
1!
1$
b1 %
1'
1*
b1 +
#171190000000
0!
0'
#171200000000
1!
b10 %
1'
b10 +
#171210000000
0!
0'
#171220000000
1!
b11 %
1'
b11 +
#171230000000
0!
0'
#171240000000
1!
b100 %
1'
b100 +
#171250000000
0!
0'
#171260000000
1!
b101 %
1'
b101 +
#171270000000
0!
0'
#171280000000
1!
0$
b110 %
1'
0*
b110 +
#171290000000
0!
0'
#171300000000
1!
b111 %
1'
b111 +
#171310000000
0!
0'
#171320000000
1!
b1000 %
1'
b1000 +
#171330000000
0!
0'
#171340000000
1!
b1001 %
1'
b1001 +
#171350000000
1"
1(
#171360000000
0!
0"
b100 &
0'
0(
b100 ,
#171370000000
1!
b0 %
1'
b0 +
#171380000000
0!
0'
#171390000000
1!
1$
b1 %
1'
1*
b1 +
#171400000000
0!
0'
#171410000000
1!
b10 %
1'
b10 +
#171420000000
0!
0'
#171430000000
1!
b11 %
1'
b11 +
#171440000000
0!
0'
#171450000000
1!
b100 %
1'
b100 +
#171460000000
0!
0'
#171470000000
1!
b101 %
1'
b101 +
#171480000000
0!
0'
#171490000000
1!
b110 %
1'
b110 +
#171500000000
0!
0'
#171510000000
1!
b111 %
1'
b111 +
#171520000000
0!
0'
#171530000000
1!
0$
b1000 %
1'
0*
b1000 +
#171540000000
0!
0'
#171550000000
1!
b1001 %
1'
b1001 +
#171560000000
0!
0'
#171570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#171580000000
0!
0'
#171590000000
1!
1$
b1 %
1'
1*
b1 +
#171600000000
0!
0'
#171610000000
1!
b10 %
1'
b10 +
#171620000000
0!
0'
#171630000000
1!
b11 %
1'
b11 +
#171640000000
0!
0'
#171650000000
1!
b100 %
1'
b100 +
#171660000000
0!
0'
#171670000000
1!
b101 %
1'
b101 +
#171680000000
0!
0'
#171690000000
1!
0$
b110 %
1'
0*
b110 +
#171700000000
0!
0'
#171710000000
1!
b111 %
1'
b111 +
#171720000000
0!
0'
#171730000000
1!
b1000 %
1'
b1000 +
#171740000000
0!
0'
#171750000000
1!
b1001 %
1'
b1001 +
#171760000000
0!
0'
#171770000000
1!
b0 %
1'
b0 +
#171780000000
1"
1(
#171790000000
0!
0"
b100 &
0'
0(
b100 ,
#171800000000
1!
1$
b1 %
1'
1*
b1 +
#171810000000
0!
0'
#171820000000
1!
b10 %
1'
b10 +
#171830000000
0!
0'
#171840000000
1!
b11 %
1'
b11 +
#171850000000
0!
0'
#171860000000
1!
b100 %
1'
b100 +
#171870000000
0!
0'
#171880000000
1!
b101 %
1'
b101 +
#171890000000
0!
0'
#171900000000
1!
b110 %
1'
b110 +
#171910000000
0!
0'
#171920000000
1!
b111 %
1'
b111 +
#171930000000
0!
0'
#171940000000
1!
0$
b1000 %
1'
0*
b1000 +
#171950000000
0!
0'
#171960000000
1!
b1001 %
1'
b1001 +
#171970000000
0!
0'
#171980000000
1!
b0 %
1'
b0 +
#171990000000
0!
0'
#172000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#172010000000
0!
0'
#172020000000
1!
b10 %
1'
b10 +
#172030000000
0!
0'
#172040000000
1!
b11 %
1'
b11 +
#172050000000
0!
0'
#172060000000
1!
b100 %
1'
b100 +
#172070000000
0!
0'
#172080000000
1!
b101 %
1'
b101 +
#172090000000
0!
0'
#172100000000
1!
0$
b110 %
1'
0*
b110 +
#172110000000
0!
0'
#172120000000
1!
b111 %
1'
b111 +
#172130000000
0!
0'
#172140000000
1!
b1000 %
1'
b1000 +
#172150000000
0!
0'
#172160000000
1!
b1001 %
1'
b1001 +
#172170000000
0!
0'
#172180000000
1!
b0 %
1'
b0 +
#172190000000
0!
0'
#172200000000
1!
1$
b1 %
1'
1*
b1 +
#172210000000
1"
1(
#172220000000
0!
0"
b100 &
0'
0(
b100 ,
#172230000000
1!
b10 %
1'
b10 +
#172240000000
0!
0'
#172250000000
1!
b11 %
1'
b11 +
#172260000000
0!
0'
#172270000000
1!
b100 %
1'
b100 +
#172280000000
0!
0'
#172290000000
1!
b101 %
1'
b101 +
#172300000000
0!
0'
#172310000000
1!
b110 %
1'
b110 +
#172320000000
0!
0'
#172330000000
1!
b111 %
1'
b111 +
#172340000000
0!
0'
#172350000000
1!
0$
b1000 %
1'
0*
b1000 +
#172360000000
0!
0'
#172370000000
1!
b1001 %
1'
b1001 +
#172380000000
0!
0'
#172390000000
1!
b0 %
1'
b0 +
#172400000000
0!
0'
#172410000000
1!
1$
b1 %
1'
1*
b1 +
#172420000000
0!
0'
#172430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#172440000000
0!
0'
#172450000000
1!
b11 %
1'
b11 +
#172460000000
0!
0'
#172470000000
1!
b100 %
1'
b100 +
#172480000000
0!
0'
#172490000000
1!
b101 %
1'
b101 +
#172500000000
0!
0'
#172510000000
1!
0$
b110 %
1'
0*
b110 +
#172520000000
0!
0'
#172530000000
1!
b111 %
1'
b111 +
#172540000000
0!
0'
#172550000000
1!
b1000 %
1'
b1000 +
#172560000000
0!
0'
#172570000000
1!
b1001 %
1'
b1001 +
#172580000000
0!
0'
#172590000000
1!
b0 %
1'
b0 +
#172600000000
0!
0'
#172610000000
1!
1$
b1 %
1'
1*
b1 +
#172620000000
0!
0'
#172630000000
1!
b10 %
1'
b10 +
#172640000000
1"
1(
#172650000000
0!
0"
b100 &
0'
0(
b100 ,
#172660000000
1!
b11 %
1'
b11 +
#172670000000
0!
0'
#172680000000
1!
b100 %
1'
b100 +
#172690000000
0!
0'
#172700000000
1!
b101 %
1'
b101 +
#172710000000
0!
0'
#172720000000
1!
b110 %
1'
b110 +
#172730000000
0!
0'
#172740000000
1!
b111 %
1'
b111 +
#172750000000
0!
0'
#172760000000
1!
0$
b1000 %
1'
0*
b1000 +
#172770000000
0!
0'
#172780000000
1!
b1001 %
1'
b1001 +
#172790000000
0!
0'
#172800000000
1!
b0 %
1'
b0 +
#172810000000
0!
0'
#172820000000
1!
1$
b1 %
1'
1*
b1 +
#172830000000
0!
0'
#172840000000
1!
b10 %
1'
b10 +
#172850000000
0!
0'
#172860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#172870000000
0!
0'
#172880000000
1!
b100 %
1'
b100 +
#172890000000
0!
0'
#172900000000
1!
b101 %
1'
b101 +
#172910000000
0!
0'
#172920000000
1!
0$
b110 %
1'
0*
b110 +
#172930000000
0!
0'
#172940000000
1!
b111 %
1'
b111 +
#172950000000
0!
0'
#172960000000
1!
b1000 %
1'
b1000 +
#172970000000
0!
0'
#172980000000
1!
b1001 %
1'
b1001 +
#172990000000
0!
0'
#173000000000
1!
b0 %
1'
b0 +
#173010000000
0!
0'
#173020000000
1!
1$
b1 %
1'
1*
b1 +
#173030000000
0!
0'
#173040000000
1!
b10 %
1'
b10 +
#173050000000
0!
0'
#173060000000
1!
b11 %
1'
b11 +
#173070000000
1"
1(
#173080000000
0!
0"
b100 &
0'
0(
b100 ,
#173090000000
1!
b100 %
1'
b100 +
#173100000000
0!
0'
#173110000000
1!
b101 %
1'
b101 +
#173120000000
0!
0'
#173130000000
1!
b110 %
1'
b110 +
#173140000000
0!
0'
#173150000000
1!
b111 %
1'
b111 +
#173160000000
0!
0'
#173170000000
1!
0$
b1000 %
1'
0*
b1000 +
#173180000000
0!
0'
#173190000000
1!
b1001 %
1'
b1001 +
#173200000000
0!
0'
#173210000000
1!
b0 %
1'
b0 +
#173220000000
0!
0'
#173230000000
1!
1$
b1 %
1'
1*
b1 +
#173240000000
0!
0'
#173250000000
1!
b10 %
1'
b10 +
#173260000000
0!
0'
#173270000000
1!
b11 %
1'
b11 +
#173280000000
0!
0'
#173290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#173300000000
0!
0'
#173310000000
1!
b101 %
1'
b101 +
#173320000000
0!
0'
#173330000000
1!
0$
b110 %
1'
0*
b110 +
#173340000000
0!
0'
#173350000000
1!
b111 %
1'
b111 +
#173360000000
0!
0'
#173370000000
1!
b1000 %
1'
b1000 +
#173380000000
0!
0'
#173390000000
1!
b1001 %
1'
b1001 +
#173400000000
0!
0'
#173410000000
1!
b0 %
1'
b0 +
#173420000000
0!
0'
#173430000000
1!
1$
b1 %
1'
1*
b1 +
#173440000000
0!
0'
#173450000000
1!
b10 %
1'
b10 +
#173460000000
0!
0'
#173470000000
1!
b11 %
1'
b11 +
#173480000000
0!
0'
#173490000000
1!
b100 %
1'
b100 +
#173500000000
1"
1(
#173510000000
0!
0"
b100 &
0'
0(
b100 ,
#173520000000
1!
b101 %
1'
b101 +
#173530000000
0!
0'
#173540000000
1!
b110 %
1'
b110 +
#173550000000
0!
0'
#173560000000
1!
b111 %
1'
b111 +
#173570000000
0!
0'
#173580000000
1!
0$
b1000 %
1'
0*
b1000 +
#173590000000
0!
0'
#173600000000
1!
b1001 %
1'
b1001 +
#173610000000
0!
0'
#173620000000
1!
b0 %
1'
b0 +
#173630000000
0!
0'
#173640000000
1!
1$
b1 %
1'
1*
b1 +
#173650000000
0!
0'
#173660000000
1!
b10 %
1'
b10 +
#173670000000
0!
0'
#173680000000
1!
b11 %
1'
b11 +
#173690000000
0!
0'
#173700000000
1!
b100 %
1'
b100 +
#173710000000
0!
0'
#173720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#173730000000
0!
0'
#173740000000
1!
0$
b110 %
1'
0*
b110 +
#173750000000
0!
0'
#173760000000
1!
b111 %
1'
b111 +
#173770000000
0!
0'
#173780000000
1!
b1000 %
1'
b1000 +
#173790000000
0!
0'
#173800000000
1!
b1001 %
1'
b1001 +
#173810000000
0!
0'
#173820000000
1!
b0 %
1'
b0 +
#173830000000
0!
0'
#173840000000
1!
1$
b1 %
1'
1*
b1 +
#173850000000
0!
0'
#173860000000
1!
b10 %
1'
b10 +
#173870000000
0!
0'
#173880000000
1!
b11 %
1'
b11 +
#173890000000
0!
0'
#173900000000
1!
b100 %
1'
b100 +
#173910000000
0!
0'
#173920000000
1!
b101 %
1'
b101 +
#173930000000
1"
1(
#173940000000
0!
0"
b100 &
0'
0(
b100 ,
#173950000000
1!
b110 %
1'
b110 +
#173960000000
0!
0'
#173970000000
1!
b111 %
1'
b111 +
#173980000000
0!
0'
#173990000000
1!
0$
b1000 %
1'
0*
b1000 +
#174000000000
0!
0'
#174010000000
1!
b1001 %
1'
b1001 +
#174020000000
0!
0'
#174030000000
1!
b0 %
1'
b0 +
#174040000000
0!
0'
#174050000000
1!
1$
b1 %
1'
1*
b1 +
#174060000000
0!
0'
#174070000000
1!
b10 %
1'
b10 +
#174080000000
0!
0'
#174090000000
1!
b11 %
1'
b11 +
#174100000000
0!
0'
#174110000000
1!
b100 %
1'
b100 +
#174120000000
0!
0'
#174130000000
1!
b101 %
1'
b101 +
#174140000000
0!
0'
#174150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#174160000000
0!
0'
#174170000000
1!
b111 %
1'
b111 +
#174180000000
0!
0'
#174190000000
1!
b1000 %
1'
b1000 +
#174200000000
0!
0'
#174210000000
1!
b1001 %
1'
b1001 +
#174220000000
0!
0'
#174230000000
1!
b0 %
1'
b0 +
#174240000000
0!
0'
#174250000000
1!
1$
b1 %
1'
1*
b1 +
#174260000000
0!
0'
#174270000000
1!
b10 %
1'
b10 +
#174280000000
0!
0'
#174290000000
1!
b11 %
1'
b11 +
#174300000000
0!
0'
#174310000000
1!
b100 %
1'
b100 +
#174320000000
0!
0'
#174330000000
1!
b101 %
1'
b101 +
#174340000000
0!
0'
#174350000000
1!
0$
b110 %
1'
0*
b110 +
#174360000000
1"
1(
#174370000000
0!
0"
b100 &
0'
0(
b100 ,
#174380000000
1!
1$
b111 %
1'
1*
b111 +
#174390000000
0!
0'
#174400000000
1!
0$
b1000 %
1'
0*
b1000 +
#174410000000
0!
0'
#174420000000
1!
b1001 %
1'
b1001 +
#174430000000
0!
0'
#174440000000
1!
b0 %
1'
b0 +
#174450000000
0!
0'
#174460000000
1!
1$
b1 %
1'
1*
b1 +
#174470000000
0!
0'
#174480000000
1!
b10 %
1'
b10 +
#174490000000
0!
0'
#174500000000
1!
b11 %
1'
b11 +
#174510000000
0!
0'
#174520000000
1!
b100 %
1'
b100 +
#174530000000
0!
0'
#174540000000
1!
b101 %
1'
b101 +
#174550000000
0!
0'
#174560000000
1!
b110 %
1'
b110 +
#174570000000
0!
0'
#174580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#174590000000
0!
0'
#174600000000
1!
b1000 %
1'
b1000 +
#174610000000
0!
0'
#174620000000
1!
b1001 %
1'
b1001 +
#174630000000
0!
0'
#174640000000
1!
b0 %
1'
b0 +
#174650000000
0!
0'
#174660000000
1!
1$
b1 %
1'
1*
b1 +
#174670000000
0!
0'
#174680000000
1!
b10 %
1'
b10 +
#174690000000
0!
0'
#174700000000
1!
b11 %
1'
b11 +
#174710000000
0!
0'
#174720000000
1!
b100 %
1'
b100 +
#174730000000
0!
0'
#174740000000
1!
b101 %
1'
b101 +
#174750000000
0!
0'
#174760000000
1!
0$
b110 %
1'
0*
b110 +
#174770000000
0!
0'
#174780000000
1!
b111 %
1'
b111 +
#174790000000
1"
1(
#174800000000
0!
0"
b100 &
0'
0(
b100 ,
#174810000000
1!
b1000 %
1'
b1000 +
#174820000000
0!
0'
#174830000000
1!
b1001 %
1'
b1001 +
#174840000000
0!
0'
#174850000000
1!
b0 %
1'
b0 +
#174860000000
0!
0'
#174870000000
1!
1$
b1 %
1'
1*
b1 +
#174880000000
0!
0'
#174890000000
1!
b10 %
1'
b10 +
#174900000000
0!
0'
#174910000000
1!
b11 %
1'
b11 +
#174920000000
0!
0'
#174930000000
1!
b100 %
1'
b100 +
#174940000000
0!
0'
#174950000000
1!
b101 %
1'
b101 +
#174960000000
0!
0'
#174970000000
1!
b110 %
1'
b110 +
#174980000000
0!
0'
#174990000000
1!
b111 %
1'
b111 +
#175000000000
0!
0'
#175010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#175020000000
0!
0'
#175030000000
1!
b1001 %
1'
b1001 +
#175040000000
0!
0'
#175050000000
1!
b0 %
1'
b0 +
#175060000000
0!
0'
#175070000000
1!
1$
b1 %
1'
1*
b1 +
#175080000000
0!
0'
#175090000000
1!
b10 %
1'
b10 +
#175100000000
0!
0'
#175110000000
1!
b11 %
1'
b11 +
#175120000000
0!
0'
#175130000000
1!
b100 %
1'
b100 +
#175140000000
0!
0'
#175150000000
1!
b101 %
1'
b101 +
#175160000000
0!
0'
#175170000000
1!
0$
b110 %
1'
0*
b110 +
#175180000000
0!
0'
#175190000000
1!
b111 %
1'
b111 +
#175200000000
0!
0'
#175210000000
1!
b1000 %
1'
b1000 +
#175220000000
1"
1(
#175230000000
0!
0"
b100 &
0'
0(
b100 ,
#175240000000
1!
b1001 %
1'
b1001 +
#175250000000
0!
0'
#175260000000
1!
b0 %
1'
b0 +
#175270000000
0!
0'
#175280000000
1!
1$
b1 %
1'
1*
b1 +
#175290000000
0!
0'
#175300000000
1!
b10 %
1'
b10 +
#175310000000
0!
0'
#175320000000
1!
b11 %
1'
b11 +
#175330000000
0!
0'
#175340000000
1!
b100 %
1'
b100 +
#175350000000
0!
0'
#175360000000
1!
b101 %
1'
b101 +
#175370000000
0!
0'
#175380000000
1!
b110 %
1'
b110 +
#175390000000
0!
0'
#175400000000
1!
b111 %
1'
b111 +
#175410000000
0!
0'
#175420000000
1!
0$
b1000 %
1'
0*
b1000 +
#175430000000
0!
0'
#175440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#175450000000
0!
0'
#175460000000
1!
b0 %
1'
b0 +
#175470000000
0!
0'
#175480000000
1!
1$
b1 %
1'
1*
b1 +
#175490000000
0!
0'
#175500000000
1!
b10 %
1'
b10 +
#175510000000
0!
0'
#175520000000
1!
b11 %
1'
b11 +
#175530000000
0!
0'
#175540000000
1!
b100 %
1'
b100 +
#175550000000
0!
0'
#175560000000
1!
b101 %
1'
b101 +
#175570000000
0!
0'
#175580000000
1!
0$
b110 %
1'
0*
b110 +
#175590000000
0!
0'
#175600000000
1!
b111 %
1'
b111 +
#175610000000
0!
0'
#175620000000
1!
b1000 %
1'
b1000 +
#175630000000
0!
0'
#175640000000
1!
b1001 %
1'
b1001 +
#175650000000
1"
1(
#175660000000
0!
0"
b100 &
0'
0(
b100 ,
#175670000000
1!
b0 %
1'
b0 +
#175680000000
0!
0'
#175690000000
1!
1$
b1 %
1'
1*
b1 +
#175700000000
0!
0'
#175710000000
1!
b10 %
1'
b10 +
#175720000000
0!
0'
#175730000000
1!
b11 %
1'
b11 +
#175740000000
0!
0'
#175750000000
1!
b100 %
1'
b100 +
#175760000000
0!
0'
#175770000000
1!
b101 %
1'
b101 +
#175780000000
0!
0'
#175790000000
1!
b110 %
1'
b110 +
#175800000000
0!
0'
#175810000000
1!
b111 %
1'
b111 +
#175820000000
0!
0'
#175830000000
1!
0$
b1000 %
1'
0*
b1000 +
#175840000000
0!
0'
#175850000000
1!
b1001 %
1'
b1001 +
#175860000000
0!
0'
#175870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#175880000000
0!
0'
#175890000000
1!
1$
b1 %
1'
1*
b1 +
#175900000000
0!
0'
#175910000000
1!
b10 %
1'
b10 +
#175920000000
0!
0'
#175930000000
1!
b11 %
1'
b11 +
#175940000000
0!
0'
#175950000000
1!
b100 %
1'
b100 +
#175960000000
0!
0'
#175970000000
1!
b101 %
1'
b101 +
#175980000000
0!
0'
#175990000000
1!
0$
b110 %
1'
0*
b110 +
#176000000000
0!
0'
#176010000000
1!
b111 %
1'
b111 +
#176020000000
0!
0'
#176030000000
1!
b1000 %
1'
b1000 +
#176040000000
0!
0'
#176050000000
1!
b1001 %
1'
b1001 +
#176060000000
0!
0'
#176070000000
1!
b0 %
1'
b0 +
#176080000000
1"
1(
#176090000000
0!
0"
b100 &
0'
0(
b100 ,
#176100000000
1!
1$
b1 %
1'
1*
b1 +
#176110000000
0!
0'
#176120000000
1!
b10 %
1'
b10 +
#176130000000
0!
0'
#176140000000
1!
b11 %
1'
b11 +
#176150000000
0!
0'
#176160000000
1!
b100 %
1'
b100 +
#176170000000
0!
0'
#176180000000
1!
b101 %
1'
b101 +
#176190000000
0!
0'
#176200000000
1!
b110 %
1'
b110 +
#176210000000
0!
0'
#176220000000
1!
b111 %
1'
b111 +
#176230000000
0!
0'
#176240000000
1!
0$
b1000 %
1'
0*
b1000 +
#176250000000
0!
0'
#176260000000
1!
b1001 %
1'
b1001 +
#176270000000
0!
0'
#176280000000
1!
b0 %
1'
b0 +
#176290000000
0!
0'
#176300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#176310000000
0!
0'
#176320000000
1!
b10 %
1'
b10 +
#176330000000
0!
0'
#176340000000
1!
b11 %
1'
b11 +
#176350000000
0!
0'
#176360000000
1!
b100 %
1'
b100 +
#176370000000
0!
0'
#176380000000
1!
b101 %
1'
b101 +
#176390000000
0!
0'
#176400000000
1!
0$
b110 %
1'
0*
b110 +
#176410000000
0!
0'
#176420000000
1!
b111 %
1'
b111 +
#176430000000
0!
0'
#176440000000
1!
b1000 %
1'
b1000 +
#176450000000
0!
0'
#176460000000
1!
b1001 %
1'
b1001 +
#176470000000
0!
0'
#176480000000
1!
b0 %
1'
b0 +
#176490000000
0!
0'
#176500000000
1!
1$
b1 %
1'
1*
b1 +
#176510000000
1"
1(
#176520000000
0!
0"
b100 &
0'
0(
b100 ,
#176530000000
1!
b10 %
1'
b10 +
#176540000000
0!
0'
#176550000000
1!
b11 %
1'
b11 +
#176560000000
0!
0'
#176570000000
1!
b100 %
1'
b100 +
#176580000000
0!
0'
#176590000000
1!
b101 %
1'
b101 +
#176600000000
0!
0'
#176610000000
1!
b110 %
1'
b110 +
#176620000000
0!
0'
#176630000000
1!
b111 %
1'
b111 +
#176640000000
0!
0'
#176650000000
1!
0$
b1000 %
1'
0*
b1000 +
#176660000000
0!
0'
#176670000000
1!
b1001 %
1'
b1001 +
#176680000000
0!
0'
#176690000000
1!
b0 %
1'
b0 +
#176700000000
0!
0'
#176710000000
1!
1$
b1 %
1'
1*
b1 +
#176720000000
0!
0'
#176730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#176740000000
0!
0'
#176750000000
1!
b11 %
1'
b11 +
#176760000000
0!
0'
#176770000000
1!
b100 %
1'
b100 +
#176780000000
0!
0'
#176790000000
1!
b101 %
1'
b101 +
#176800000000
0!
0'
#176810000000
1!
0$
b110 %
1'
0*
b110 +
#176820000000
0!
0'
#176830000000
1!
b111 %
1'
b111 +
#176840000000
0!
0'
#176850000000
1!
b1000 %
1'
b1000 +
#176860000000
0!
0'
#176870000000
1!
b1001 %
1'
b1001 +
#176880000000
0!
0'
#176890000000
1!
b0 %
1'
b0 +
#176900000000
0!
0'
#176910000000
1!
1$
b1 %
1'
1*
b1 +
#176920000000
0!
0'
#176930000000
1!
b10 %
1'
b10 +
#176940000000
1"
1(
#176950000000
0!
0"
b100 &
0'
0(
b100 ,
#176960000000
1!
b11 %
1'
b11 +
#176970000000
0!
0'
#176980000000
1!
b100 %
1'
b100 +
#176990000000
0!
0'
#177000000000
1!
b101 %
1'
b101 +
#177010000000
0!
0'
#177020000000
1!
b110 %
1'
b110 +
#177030000000
0!
0'
#177040000000
1!
b111 %
1'
b111 +
#177050000000
0!
0'
#177060000000
1!
0$
b1000 %
1'
0*
b1000 +
#177070000000
0!
0'
#177080000000
1!
b1001 %
1'
b1001 +
#177090000000
0!
0'
#177100000000
1!
b0 %
1'
b0 +
#177110000000
0!
0'
#177120000000
1!
1$
b1 %
1'
1*
b1 +
#177130000000
0!
0'
#177140000000
1!
b10 %
1'
b10 +
#177150000000
0!
0'
#177160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#177170000000
0!
0'
#177180000000
1!
b100 %
1'
b100 +
#177190000000
0!
0'
#177200000000
1!
b101 %
1'
b101 +
#177210000000
0!
0'
#177220000000
1!
0$
b110 %
1'
0*
b110 +
#177230000000
0!
0'
#177240000000
1!
b111 %
1'
b111 +
#177250000000
0!
0'
#177260000000
1!
b1000 %
1'
b1000 +
#177270000000
0!
0'
#177280000000
1!
b1001 %
1'
b1001 +
#177290000000
0!
0'
#177300000000
1!
b0 %
1'
b0 +
#177310000000
0!
0'
#177320000000
1!
1$
b1 %
1'
1*
b1 +
#177330000000
0!
0'
#177340000000
1!
b10 %
1'
b10 +
#177350000000
0!
0'
#177360000000
1!
b11 %
1'
b11 +
#177370000000
1"
1(
#177380000000
0!
0"
b100 &
0'
0(
b100 ,
#177390000000
1!
b100 %
1'
b100 +
#177400000000
0!
0'
#177410000000
1!
b101 %
1'
b101 +
#177420000000
0!
0'
#177430000000
1!
b110 %
1'
b110 +
#177440000000
0!
0'
#177450000000
1!
b111 %
1'
b111 +
#177460000000
0!
0'
#177470000000
1!
0$
b1000 %
1'
0*
b1000 +
#177480000000
0!
0'
#177490000000
1!
b1001 %
1'
b1001 +
#177500000000
0!
0'
#177510000000
1!
b0 %
1'
b0 +
#177520000000
0!
0'
#177530000000
1!
1$
b1 %
1'
1*
b1 +
#177540000000
0!
0'
#177550000000
1!
b10 %
1'
b10 +
#177560000000
0!
0'
#177570000000
1!
b11 %
1'
b11 +
#177580000000
0!
0'
#177590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#177600000000
0!
0'
#177610000000
1!
b101 %
1'
b101 +
#177620000000
0!
0'
#177630000000
1!
0$
b110 %
1'
0*
b110 +
#177640000000
0!
0'
#177650000000
1!
b111 %
1'
b111 +
#177660000000
0!
0'
#177670000000
1!
b1000 %
1'
b1000 +
#177680000000
0!
0'
#177690000000
1!
b1001 %
1'
b1001 +
#177700000000
0!
0'
#177710000000
1!
b0 %
1'
b0 +
#177720000000
0!
0'
#177730000000
1!
1$
b1 %
1'
1*
b1 +
#177740000000
0!
0'
#177750000000
1!
b10 %
1'
b10 +
#177760000000
0!
0'
#177770000000
1!
b11 %
1'
b11 +
#177780000000
0!
0'
#177790000000
1!
b100 %
1'
b100 +
#177800000000
1"
1(
#177810000000
0!
0"
b100 &
0'
0(
b100 ,
#177820000000
1!
b101 %
1'
b101 +
#177830000000
0!
0'
#177840000000
1!
b110 %
1'
b110 +
#177850000000
0!
0'
#177860000000
1!
b111 %
1'
b111 +
#177870000000
0!
0'
#177880000000
1!
0$
b1000 %
1'
0*
b1000 +
#177890000000
0!
0'
#177900000000
1!
b1001 %
1'
b1001 +
#177910000000
0!
0'
#177920000000
1!
b0 %
1'
b0 +
#177930000000
0!
0'
#177940000000
1!
1$
b1 %
1'
1*
b1 +
#177950000000
0!
0'
#177960000000
1!
b10 %
1'
b10 +
#177970000000
0!
0'
#177980000000
1!
b11 %
1'
b11 +
#177990000000
0!
0'
#178000000000
1!
b100 %
1'
b100 +
#178010000000
0!
0'
#178020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#178030000000
0!
0'
#178040000000
1!
0$
b110 %
1'
0*
b110 +
#178050000000
0!
0'
#178060000000
1!
b111 %
1'
b111 +
#178070000000
0!
0'
#178080000000
1!
b1000 %
1'
b1000 +
#178090000000
0!
0'
#178100000000
1!
b1001 %
1'
b1001 +
#178110000000
0!
0'
#178120000000
1!
b0 %
1'
b0 +
#178130000000
0!
0'
#178140000000
1!
1$
b1 %
1'
1*
b1 +
#178150000000
0!
0'
#178160000000
1!
b10 %
1'
b10 +
#178170000000
0!
0'
#178180000000
1!
b11 %
1'
b11 +
#178190000000
0!
0'
#178200000000
1!
b100 %
1'
b100 +
#178210000000
0!
0'
#178220000000
1!
b101 %
1'
b101 +
#178230000000
1"
1(
#178240000000
0!
0"
b100 &
0'
0(
b100 ,
#178250000000
1!
b110 %
1'
b110 +
#178260000000
0!
0'
#178270000000
1!
b111 %
1'
b111 +
#178280000000
0!
0'
#178290000000
1!
0$
b1000 %
1'
0*
b1000 +
#178300000000
0!
0'
#178310000000
1!
b1001 %
1'
b1001 +
#178320000000
0!
0'
#178330000000
1!
b0 %
1'
b0 +
#178340000000
0!
0'
#178350000000
1!
1$
b1 %
1'
1*
b1 +
#178360000000
0!
0'
#178370000000
1!
b10 %
1'
b10 +
#178380000000
0!
0'
#178390000000
1!
b11 %
1'
b11 +
#178400000000
0!
0'
#178410000000
1!
b100 %
1'
b100 +
#178420000000
0!
0'
#178430000000
1!
b101 %
1'
b101 +
#178440000000
0!
0'
#178450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#178460000000
0!
0'
#178470000000
1!
b111 %
1'
b111 +
#178480000000
0!
0'
#178490000000
1!
b1000 %
1'
b1000 +
#178500000000
0!
0'
#178510000000
1!
b1001 %
1'
b1001 +
#178520000000
0!
0'
#178530000000
1!
b0 %
1'
b0 +
#178540000000
0!
0'
#178550000000
1!
1$
b1 %
1'
1*
b1 +
#178560000000
0!
0'
#178570000000
1!
b10 %
1'
b10 +
#178580000000
0!
0'
#178590000000
1!
b11 %
1'
b11 +
#178600000000
0!
0'
#178610000000
1!
b100 %
1'
b100 +
#178620000000
0!
0'
#178630000000
1!
b101 %
1'
b101 +
#178640000000
0!
0'
#178650000000
1!
0$
b110 %
1'
0*
b110 +
#178660000000
1"
1(
#178670000000
0!
0"
b100 &
0'
0(
b100 ,
#178680000000
1!
1$
b111 %
1'
1*
b111 +
#178690000000
0!
0'
#178700000000
1!
0$
b1000 %
1'
0*
b1000 +
#178710000000
0!
0'
#178720000000
1!
b1001 %
1'
b1001 +
#178730000000
0!
0'
#178740000000
1!
b0 %
1'
b0 +
#178750000000
0!
0'
#178760000000
1!
1$
b1 %
1'
1*
b1 +
#178770000000
0!
0'
#178780000000
1!
b10 %
1'
b10 +
#178790000000
0!
0'
#178800000000
1!
b11 %
1'
b11 +
#178810000000
0!
0'
#178820000000
1!
b100 %
1'
b100 +
#178830000000
0!
0'
#178840000000
1!
b101 %
1'
b101 +
#178850000000
0!
0'
#178860000000
1!
b110 %
1'
b110 +
#178870000000
0!
0'
#178880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#178890000000
0!
0'
#178900000000
1!
b1000 %
1'
b1000 +
#178910000000
0!
0'
#178920000000
1!
b1001 %
1'
b1001 +
#178930000000
0!
0'
#178940000000
1!
b0 %
1'
b0 +
#178950000000
0!
0'
#178960000000
1!
1$
b1 %
1'
1*
b1 +
#178970000000
0!
0'
#178980000000
1!
b10 %
1'
b10 +
#178990000000
0!
0'
#179000000000
1!
b11 %
1'
b11 +
#179010000000
0!
0'
#179020000000
1!
b100 %
1'
b100 +
#179030000000
0!
0'
#179040000000
1!
b101 %
1'
b101 +
#179050000000
0!
0'
#179060000000
1!
0$
b110 %
1'
0*
b110 +
#179070000000
0!
0'
#179080000000
1!
b111 %
1'
b111 +
#179090000000
1"
1(
#179100000000
0!
0"
b100 &
0'
0(
b100 ,
#179110000000
1!
b1000 %
1'
b1000 +
#179120000000
0!
0'
#179130000000
1!
b1001 %
1'
b1001 +
#179140000000
0!
0'
#179150000000
1!
b0 %
1'
b0 +
#179160000000
0!
0'
#179170000000
1!
1$
b1 %
1'
1*
b1 +
#179180000000
0!
0'
#179190000000
1!
b10 %
1'
b10 +
#179200000000
0!
0'
#179210000000
1!
b11 %
1'
b11 +
#179220000000
0!
0'
#179230000000
1!
b100 %
1'
b100 +
#179240000000
0!
0'
#179250000000
1!
b101 %
1'
b101 +
#179260000000
0!
0'
#179270000000
1!
b110 %
1'
b110 +
#179280000000
0!
0'
#179290000000
1!
b111 %
1'
b111 +
#179300000000
0!
0'
#179310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#179320000000
0!
0'
#179330000000
1!
b1001 %
1'
b1001 +
#179340000000
0!
0'
#179350000000
1!
b0 %
1'
b0 +
#179360000000
0!
0'
#179370000000
1!
1$
b1 %
1'
1*
b1 +
#179380000000
0!
0'
#179390000000
1!
b10 %
1'
b10 +
#179400000000
0!
0'
#179410000000
1!
b11 %
1'
b11 +
#179420000000
0!
0'
#179430000000
1!
b100 %
1'
b100 +
#179440000000
0!
0'
#179450000000
1!
b101 %
1'
b101 +
#179460000000
0!
0'
#179470000000
1!
0$
b110 %
1'
0*
b110 +
#179480000000
0!
0'
#179490000000
1!
b111 %
1'
b111 +
#179500000000
0!
0'
#179510000000
1!
b1000 %
1'
b1000 +
#179520000000
1"
1(
#179530000000
0!
0"
b100 &
0'
0(
b100 ,
#179540000000
1!
b1001 %
1'
b1001 +
#179550000000
0!
0'
#179560000000
1!
b0 %
1'
b0 +
#179570000000
0!
0'
#179580000000
1!
1$
b1 %
1'
1*
b1 +
#179590000000
0!
0'
#179600000000
1!
b10 %
1'
b10 +
#179610000000
0!
0'
#179620000000
1!
b11 %
1'
b11 +
#179630000000
0!
0'
#179640000000
1!
b100 %
1'
b100 +
#179650000000
0!
0'
#179660000000
1!
b101 %
1'
b101 +
#179670000000
0!
0'
#179680000000
1!
b110 %
1'
b110 +
#179690000000
0!
0'
#179700000000
1!
b111 %
1'
b111 +
#179710000000
0!
0'
#179720000000
1!
0$
b1000 %
1'
0*
b1000 +
#179730000000
0!
0'
#179740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#179750000000
0!
0'
#179760000000
1!
b0 %
1'
b0 +
#179770000000
0!
0'
#179780000000
1!
1$
b1 %
1'
1*
b1 +
#179790000000
0!
0'
#179800000000
1!
b10 %
1'
b10 +
#179810000000
0!
0'
#179820000000
1!
b11 %
1'
b11 +
#179830000000
0!
0'
#179840000000
1!
b100 %
1'
b100 +
#179850000000
0!
0'
#179860000000
1!
b101 %
1'
b101 +
#179870000000
0!
0'
#179880000000
1!
0$
b110 %
1'
0*
b110 +
#179890000000
0!
0'
#179900000000
1!
b111 %
1'
b111 +
#179910000000
0!
0'
#179920000000
1!
b1000 %
1'
b1000 +
#179930000000
0!
0'
#179940000000
1!
b1001 %
1'
b1001 +
#179950000000
1"
1(
#179960000000
0!
0"
b100 &
0'
0(
b100 ,
#179970000000
1!
b0 %
1'
b0 +
#179980000000
0!
0'
#179990000000
1!
1$
b1 %
1'
1*
b1 +
#180000000000
0!
0'
#180010000000
1!
b10 %
1'
b10 +
#180020000000
0!
0'
#180030000000
1!
b11 %
1'
b11 +
#180040000000
0!
0'
#180050000000
1!
b100 %
1'
b100 +
#180060000000
0!
0'
#180070000000
1!
b101 %
1'
b101 +
#180080000000
0!
0'
#180090000000
1!
b110 %
1'
b110 +
#180100000000
0!
0'
#180110000000
1!
b111 %
1'
b111 +
#180120000000
0!
0'
#180130000000
1!
0$
b1000 %
1'
0*
b1000 +
#180140000000
0!
0'
#180150000000
1!
b1001 %
1'
b1001 +
#180160000000
0!
0'
#180170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#180180000000
0!
0'
#180190000000
1!
1$
b1 %
1'
1*
b1 +
#180200000000
0!
0'
#180210000000
1!
b10 %
1'
b10 +
#180220000000
0!
0'
#180230000000
1!
b11 %
1'
b11 +
#180240000000
0!
0'
#180250000000
1!
b100 %
1'
b100 +
#180260000000
0!
0'
#180270000000
1!
b101 %
1'
b101 +
#180280000000
0!
0'
#180290000000
1!
0$
b110 %
1'
0*
b110 +
#180300000000
0!
0'
#180310000000
1!
b111 %
1'
b111 +
#180320000000
0!
0'
#180330000000
1!
b1000 %
1'
b1000 +
#180340000000
0!
0'
#180350000000
1!
b1001 %
1'
b1001 +
#180360000000
0!
0'
#180370000000
1!
b0 %
1'
b0 +
#180380000000
1"
1(
#180390000000
0!
0"
b100 &
0'
0(
b100 ,
#180400000000
1!
1$
b1 %
1'
1*
b1 +
#180410000000
0!
0'
#180420000000
1!
b10 %
1'
b10 +
#180430000000
0!
0'
#180440000000
1!
b11 %
1'
b11 +
#180450000000
0!
0'
#180460000000
1!
b100 %
1'
b100 +
#180470000000
0!
0'
#180480000000
1!
b101 %
1'
b101 +
#180490000000
0!
0'
#180500000000
1!
b110 %
1'
b110 +
#180510000000
0!
0'
#180520000000
1!
b111 %
1'
b111 +
#180530000000
0!
0'
#180540000000
1!
0$
b1000 %
1'
0*
b1000 +
#180550000000
0!
0'
#180560000000
1!
b1001 %
1'
b1001 +
#180570000000
0!
0'
#180580000000
1!
b0 %
1'
b0 +
#180590000000
0!
0'
#180600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#180610000000
0!
0'
#180620000000
1!
b10 %
1'
b10 +
#180630000000
0!
0'
#180640000000
1!
b11 %
1'
b11 +
#180650000000
0!
0'
#180660000000
1!
b100 %
1'
b100 +
#180670000000
0!
0'
#180680000000
1!
b101 %
1'
b101 +
#180690000000
0!
0'
#180700000000
1!
0$
b110 %
1'
0*
b110 +
#180710000000
0!
0'
#180720000000
1!
b111 %
1'
b111 +
#180730000000
0!
0'
#180740000000
1!
b1000 %
1'
b1000 +
#180750000000
0!
0'
#180760000000
1!
b1001 %
1'
b1001 +
#180770000000
0!
0'
#180780000000
1!
b0 %
1'
b0 +
#180790000000
0!
0'
#180800000000
1!
1$
b1 %
1'
1*
b1 +
#180810000000
1"
1(
#180820000000
0!
0"
b100 &
0'
0(
b100 ,
#180830000000
1!
b10 %
1'
b10 +
#180840000000
0!
0'
#180850000000
1!
b11 %
1'
b11 +
#180860000000
0!
0'
#180870000000
1!
b100 %
1'
b100 +
#180880000000
0!
0'
#180890000000
1!
b101 %
1'
b101 +
#180900000000
0!
0'
#180910000000
1!
b110 %
1'
b110 +
#180920000000
0!
0'
#180930000000
1!
b111 %
1'
b111 +
#180940000000
0!
0'
#180950000000
1!
0$
b1000 %
1'
0*
b1000 +
#180960000000
0!
0'
#180970000000
1!
b1001 %
1'
b1001 +
#180980000000
0!
0'
#180990000000
1!
b0 %
1'
b0 +
#181000000000
0!
0'
#181010000000
1!
1$
b1 %
1'
1*
b1 +
#181020000000
0!
0'
#181030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#181040000000
0!
0'
#181050000000
1!
b11 %
1'
b11 +
#181060000000
0!
0'
#181070000000
1!
b100 %
1'
b100 +
#181080000000
0!
0'
#181090000000
1!
b101 %
1'
b101 +
#181100000000
0!
0'
#181110000000
1!
0$
b110 %
1'
0*
b110 +
#181120000000
0!
0'
#181130000000
1!
b111 %
1'
b111 +
#181140000000
0!
0'
#181150000000
1!
b1000 %
1'
b1000 +
#181160000000
0!
0'
#181170000000
1!
b1001 %
1'
b1001 +
#181180000000
0!
0'
#181190000000
1!
b0 %
1'
b0 +
#181200000000
0!
0'
#181210000000
1!
1$
b1 %
1'
1*
b1 +
#181220000000
0!
0'
#181230000000
1!
b10 %
1'
b10 +
#181240000000
1"
1(
#181250000000
0!
0"
b100 &
0'
0(
b100 ,
#181260000000
1!
b11 %
1'
b11 +
#181270000000
0!
0'
#181280000000
1!
b100 %
1'
b100 +
#181290000000
0!
0'
#181300000000
1!
b101 %
1'
b101 +
#181310000000
0!
0'
#181320000000
1!
b110 %
1'
b110 +
#181330000000
0!
0'
#181340000000
1!
b111 %
1'
b111 +
#181350000000
0!
0'
#181360000000
1!
0$
b1000 %
1'
0*
b1000 +
#181370000000
0!
0'
#181380000000
1!
b1001 %
1'
b1001 +
#181390000000
0!
0'
#181400000000
1!
b0 %
1'
b0 +
#181410000000
0!
0'
#181420000000
1!
1$
b1 %
1'
1*
b1 +
#181430000000
0!
0'
#181440000000
1!
b10 %
1'
b10 +
#181450000000
0!
0'
#181460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#181470000000
0!
0'
#181480000000
1!
b100 %
1'
b100 +
#181490000000
0!
0'
#181500000000
1!
b101 %
1'
b101 +
#181510000000
0!
0'
#181520000000
1!
0$
b110 %
1'
0*
b110 +
#181530000000
0!
0'
#181540000000
1!
b111 %
1'
b111 +
#181550000000
0!
0'
#181560000000
1!
b1000 %
1'
b1000 +
#181570000000
0!
0'
#181580000000
1!
b1001 %
1'
b1001 +
#181590000000
0!
0'
#181600000000
1!
b0 %
1'
b0 +
#181610000000
0!
0'
#181620000000
1!
1$
b1 %
1'
1*
b1 +
#181630000000
0!
0'
#181640000000
1!
b10 %
1'
b10 +
#181650000000
0!
0'
#181660000000
1!
b11 %
1'
b11 +
#181670000000
1"
1(
#181680000000
0!
0"
b100 &
0'
0(
b100 ,
#181690000000
1!
b100 %
1'
b100 +
#181700000000
0!
0'
#181710000000
1!
b101 %
1'
b101 +
#181720000000
0!
0'
#181730000000
1!
b110 %
1'
b110 +
#181740000000
0!
0'
#181750000000
1!
b111 %
1'
b111 +
#181760000000
0!
0'
#181770000000
1!
0$
b1000 %
1'
0*
b1000 +
#181780000000
0!
0'
#181790000000
1!
b1001 %
1'
b1001 +
#181800000000
0!
0'
#181810000000
1!
b0 %
1'
b0 +
#181820000000
0!
0'
#181830000000
1!
1$
b1 %
1'
1*
b1 +
#181840000000
0!
0'
#181850000000
1!
b10 %
1'
b10 +
#181860000000
0!
0'
#181870000000
1!
b11 %
1'
b11 +
#181880000000
0!
0'
#181890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#181900000000
0!
0'
#181910000000
1!
b101 %
1'
b101 +
#181920000000
0!
0'
#181930000000
1!
0$
b110 %
1'
0*
b110 +
#181940000000
0!
0'
#181950000000
1!
b111 %
1'
b111 +
#181960000000
0!
0'
#181970000000
1!
b1000 %
1'
b1000 +
#181980000000
0!
0'
#181990000000
1!
b1001 %
1'
b1001 +
#182000000000
0!
0'
#182010000000
1!
b0 %
1'
b0 +
#182020000000
0!
0'
#182030000000
1!
1$
b1 %
1'
1*
b1 +
#182040000000
0!
0'
#182050000000
1!
b10 %
1'
b10 +
#182060000000
0!
0'
#182070000000
1!
b11 %
1'
b11 +
#182080000000
0!
0'
#182090000000
1!
b100 %
1'
b100 +
#182100000000
1"
1(
#182110000000
0!
0"
b100 &
0'
0(
b100 ,
#182120000000
1!
b101 %
1'
b101 +
#182130000000
0!
0'
#182140000000
1!
b110 %
1'
b110 +
#182150000000
0!
0'
#182160000000
1!
b111 %
1'
b111 +
#182170000000
0!
0'
#182180000000
1!
0$
b1000 %
1'
0*
b1000 +
#182190000000
0!
0'
#182200000000
1!
b1001 %
1'
b1001 +
#182210000000
0!
0'
#182220000000
1!
b0 %
1'
b0 +
#182230000000
0!
0'
#182240000000
1!
1$
b1 %
1'
1*
b1 +
#182250000000
0!
0'
#182260000000
1!
b10 %
1'
b10 +
#182270000000
0!
0'
#182280000000
1!
b11 %
1'
b11 +
#182290000000
0!
0'
#182300000000
1!
b100 %
1'
b100 +
#182310000000
0!
0'
#182320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#182330000000
0!
0'
#182340000000
1!
0$
b110 %
1'
0*
b110 +
#182350000000
0!
0'
#182360000000
1!
b111 %
1'
b111 +
#182370000000
0!
0'
#182380000000
1!
b1000 %
1'
b1000 +
#182390000000
0!
0'
#182400000000
1!
b1001 %
1'
b1001 +
#182410000000
0!
0'
#182420000000
1!
b0 %
1'
b0 +
#182430000000
0!
0'
#182440000000
1!
1$
b1 %
1'
1*
b1 +
#182450000000
0!
0'
#182460000000
1!
b10 %
1'
b10 +
#182470000000
0!
0'
#182480000000
1!
b11 %
1'
b11 +
#182490000000
0!
0'
#182500000000
1!
b100 %
1'
b100 +
#182510000000
0!
0'
#182520000000
1!
b101 %
1'
b101 +
#182530000000
1"
1(
#182540000000
0!
0"
b100 &
0'
0(
b100 ,
#182550000000
1!
b110 %
1'
b110 +
#182560000000
0!
0'
#182570000000
1!
b111 %
1'
b111 +
#182580000000
0!
0'
#182590000000
1!
0$
b1000 %
1'
0*
b1000 +
#182600000000
0!
0'
#182610000000
1!
b1001 %
1'
b1001 +
#182620000000
0!
0'
#182630000000
1!
b0 %
1'
b0 +
#182640000000
0!
0'
#182650000000
1!
1$
b1 %
1'
1*
b1 +
#182660000000
0!
0'
#182670000000
1!
b10 %
1'
b10 +
#182680000000
0!
0'
#182690000000
1!
b11 %
1'
b11 +
#182700000000
0!
0'
#182710000000
1!
b100 %
1'
b100 +
#182720000000
0!
0'
#182730000000
1!
b101 %
1'
b101 +
#182740000000
0!
0'
#182750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#182760000000
0!
0'
#182770000000
1!
b111 %
1'
b111 +
#182780000000
0!
0'
#182790000000
1!
b1000 %
1'
b1000 +
#182800000000
0!
0'
#182810000000
1!
b1001 %
1'
b1001 +
#182820000000
0!
0'
#182830000000
1!
b0 %
1'
b0 +
#182840000000
0!
0'
#182850000000
1!
1$
b1 %
1'
1*
b1 +
#182860000000
0!
0'
#182870000000
1!
b10 %
1'
b10 +
#182880000000
0!
0'
#182890000000
1!
b11 %
1'
b11 +
#182900000000
0!
0'
#182910000000
1!
b100 %
1'
b100 +
#182920000000
0!
0'
#182930000000
1!
b101 %
1'
b101 +
#182940000000
0!
0'
#182950000000
1!
0$
b110 %
1'
0*
b110 +
#182960000000
1"
1(
#182970000000
0!
0"
b100 &
0'
0(
b100 ,
#182980000000
1!
1$
b111 %
1'
1*
b111 +
#182990000000
0!
0'
#183000000000
1!
0$
b1000 %
1'
0*
b1000 +
#183010000000
0!
0'
#183020000000
1!
b1001 %
1'
b1001 +
#183030000000
0!
0'
#183040000000
1!
b0 %
1'
b0 +
#183050000000
0!
0'
#183060000000
1!
1$
b1 %
1'
1*
b1 +
#183070000000
0!
0'
#183080000000
1!
b10 %
1'
b10 +
#183090000000
0!
0'
#183100000000
1!
b11 %
1'
b11 +
#183110000000
0!
0'
#183120000000
1!
b100 %
1'
b100 +
#183130000000
0!
0'
#183140000000
1!
b101 %
1'
b101 +
#183150000000
0!
0'
#183160000000
1!
b110 %
1'
b110 +
#183170000000
0!
0'
#183180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#183190000000
0!
0'
#183200000000
1!
b1000 %
1'
b1000 +
#183210000000
0!
0'
#183220000000
1!
b1001 %
1'
b1001 +
#183230000000
0!
0'
#183240000000
1!
b0 %
1'
b0 +
#183250000000
0!
0'
#183260000000
1!
1$
b1 %
1'
1*
b1 +
#183270000000
0!
0'
#183280000000
1!
b10 %
1'
b10 +
#183290000000
0!
0'
#183300000000
1!
b11 %
1'
b11 +
#183310000000
0!
0'
#183320000000
1!
b100 %
1'
b100 +
#183330000000
0!
0'
#183340000000
1!
b101 %
1'
b101 +
#183350000000
0!
0'
#183360000000
1!
0$
b110 %
1'
0*
b110 +
#183370000000
0!
0'
#183380000000
1!
b111 %
1'
b111 +
#183390000000
1"
1(
#183400000000
0!
0"
b100 &
0'
0(
b100 ,
#183410000000
1!
b1000 %
1'
b1000 +
#183420000000
0!
0'
#183430000000
1!
b1001 %
1'
b1001 +
#183440000000
0!
0'
#183450000000
1!
b0 %
1'
b0 +
#183460000000
0!
0'
#183470000000
1!
1$
b1 %
1'
1*
b1 +
#183480000000
0!
0'
#183490000000
1!
b10 %
1'
b10 +
#183500000000
0!
0'
#183510000000
1!
b11 %
1'
b11 +
#183520000000
0!
0'
#183530000000
1!
b100 %
1'
b100 +
#183540000000
0!
0'
#183550000000
1!
b101 %
1'
b101 +
#183560000000
0!
0'
#183570000000
1!
b110 %
1'
b110 +
#183580000000
0!
0'
#183590000000
1!
b111 %
1'
b111 +
#183600000000
0!
0'
#183610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#183620000000
0!
0'
#183630000000
1!
b1001 %
1'
b1001 +
#183640000000
0!
0'
#183650000000
1!
b0 %
1'
b0 +
#183660000000
0!
0'
#183670000000
1!
1$
b1 %
1'
1*
b1 +
#183680000000
0!
0'
#183690000000
1!
b10 %
1'
b10 +
#183700000000
0!
0'
#183710000000
1!
b11 %
1'
b11 +
#183720000000
0!
0'
#183730000000
1!
b100 %
1'
b100 +
#183740000000
0!
0'
#183750000000
1!
b101 %
1'
b101 +
#183760000000
0!
0'
#183770000000
1!
0$
b110 %
1'
0*
b110 +
#183780000000
0!
0'
#183790000000
1!
b111 %
1'
b111 +
#183800000000
0!
0'
#183810000000
1!
b1000 %
1'
b1000 +
#183820000000
1"
1(
#183830000000
0!
0"
b100 &
0'
0(
b100 ,
#183840000000
1!
b1001 %
1'
b1001 +
#183850000000
0!
0'
#183860000000
1!
b0 %
1'
b0 +
#183870000000
0!
0'
#183880000000
1!
1$
b1 %
1'
1*
b1 +
#183890000000
0!
0'
#183900000000
1!
b10 %
1'
b10 +
#183910000000
0!
0'
#183920000000
1!
b11 %
1'
b11 +
#183930000000
0!
0'
#183940000000
1!
b100 %
1'
b100 +
#183950000000
0!
0'
#183960000000
1!
b101 %
1'
b101 +
#183970000000
0!
0'
#183980000000
1!
b110 %
1'
b110 +
#183990000000
0!
0'
#184000000000
1!
b111 %
1'
b111 +
#184010000000
0!
0'
#184020000000
1!
0$
b1000 %
1'
0*
b1000 +
#184030000000
0!
0'
#184040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#184050000000
0!
0'
#184060000000
1!
b0 %
1'
b0 +
#184070000000
0!
0'
#184080000000
1!
1$
b1 %
1'
1*
b1 +
#184090000000
0!
0'
#184100000000
1!
b10 %
1'
b10 +
#184110000000
0!
0'
#184120000000
1!
b11 %
1'
b11 +
#184130000000
0!
0'
#184140000000
1!
b100 %
1'
b100 +
#184150000000
0!
0'
#184160000000
1!
b101 %
1'
b101 +
#184170000000
0!
0'
#184180000000
1!
0$
b110 %
1'
0*
b110 +
#184190000000
0!
0'
#184200000000
1!
b111 %
1'
b111 +
#184210000000
0!
0'
#184220000000
1!
b1000 %
1'
b1000 +
#184230000000
0!
0'
#184240000000
1!
b1001 %
1'
b1001 +
#184250000000
1"
1(
#184260000000
0!
0"
b100 &
0'
0(
b100 ,
#184270000000
1!
b0 %
1'
b0 +
#184280000000
0!
0'
#184290000000
1!
1$
b1 %
1'
1*
b1 +
#184300000000
0!
0'
#184310000000
1!
b10 %
1'
b10 +
#184320000000
0!
0'
#184330000000
1!
b11 %
1'
b11 +
#184340000000
0!
0'
#184350000000
1!
b100 %
1'
b100 +
#184360000000
0!
0'
#184370000000
1!
b101 %
1'
b101 +
#184380000000
0!
0'
#184390000000
1!
b110 %
1'
b110 +
#184400000000
0!
0'
#184410000000
1!
b111 %
1'
b111 +
#184420000000
0!
0'
#184430000000
1!
0$
b1000 %
1'
0*
b1000 +
#184440000000
0!
0'
#184450000000
1!
b1001 %
1'
b1001 +
#184460000000
0!
0'
#184470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#184480000000
0!
0'
#184490000000
1!
1$
b1 %
1'
1*
b1 +
#184500000000
0!
0'
#184510000000
1!
b10 %
1'
b10 +
#184520000000
0!
0'
#184530000000
1!
b11 %
1'
b11 +
#184540000000
0!
0'
#184550000000
1!
b100 %
1'
b100 +
#184560000000
0!
0'
#184570000000
1!
b101 %
1'
b101 +
#184580000000
0!
0'
#184590000000
1!
0$
b110 %
1'
0*
b110 +
#184600000000
0!
0'
#184610000000
1!
b111 %
1'
b111 +
#184620000000
0!
0'
#184630000000
1!
b1000 %
1'
b1000 +
#184640000000
0!
0'
#184650000000
1!
b1001 %
1'
b1001 +
#184660000000
0!
0'
#184670000000
1!
b0 %
1'
b0 +
#184680000000
1"
1(
#184690000000
0!
0"
b100 &
0'
0(
b100 ,
#184700000000
1!
1$
b1 %
1'
1*
b1 +
#184710000000
0!
0'
#184720000000
1!
b10 %
1'
b10 +
#184730000000
0!
0'
#184740000000
1!
b11 %
1'
b11 +
#184750000000
0!
0'
#184760000000
1!
b100 %
1'
b100 +
#184770000000
0!
0'
#184780000000
1!
b101 %
1'
b101 +
#184790000000
0!
0'
#184800000000
1!
b110 %
1'
b110 +
#184810000000
0!
0'
#184820000000
1!
b111 %
1'
b111 +
#184830000000
0!
0'
#184840000000
1!
0$
b1000 %
1'
0*
b1000 +
#184850000000
0!
0'
#184860000000
1!
b1001 %
1'
b1001 +
#184870000000
0!
0'
#184880000000
1!
b0 %
1'
b0 +
#184890000000
0!
0'
#184900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#184910000000
0!
0'
#184920000000
1!
b10 %
1'
b10 +
#184930000000
0!
0'
#184940000000
1!
b11 %
1'
b11 +
#184950000000
0!
0'
#184960000000
1!
b100 %
1'
b100 +
#184970000000
0!
0'
#184980000000
1!
b101 %
1'
b101 +
#184990000000
0!
0'
#185000000000
1!
0$
b110 %
1'
0*
b110 +
#185010000000
0!
0'
#185020000000
1!
b111 %
1'
b111 +
#185030000000
0!
0'
#185040000000
1!
b1000 %
1'
b1000 +
#185050000000
0!
0'
#185060000000
1!
b1001 %
1'
b1001 +
#185070000000
0!
0'
#185080000000
1!
b0 %
1'
b0 +
#185090000000
0!
0'
#185100000000
1!
1$
b1 %
1'
1*
b1 +
#185110000000
1"
1(
#185120000000
0!
0"
b100 &
0'
0(
b100 ,
#185130000000
1!
b10 %
1'
b10 +
#185140000000
0!
0'
#185150000000
1!
b11 %
1'
b11 +
#185160000000
0!
0'
#185170000000
1!
b100 %
1'
b100 +
#185180000000
0!
0'
#185190000000
1!
b101 %
1'
b101 +
#185200000000
0!
0'
#185210000000
1!
b110 %
1'
b110 +
#185220000000
0!
0'
#185230000000
1!
b111 %
1'
b111 +
#185240000000
0!
0'
#185250000000
1!
0$
b1000 %
1'
0*
b1000 +
#185260000000
0!
0'
#185270000000
1!
b1001 %
1'
b1001 +
#185280000000
0!
0'
#185290000000
1!
b0 %
1'
b0 +
#185300000000
0!
0'
#185310000000
1!
1$
b1 %
1'
1*
b1 +
#185320000000
0!
0'
#185330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#185340000000
0!
0'
#185350000000
1!
b11 %
1'
b11 +
#185360000000
0!
0'
#185370000000
1!
b100 %
1'
b100 +
#185380000000
0!
0'
#185390000000
1!
b101 %
1'
b101 +
#185400000000
0!
0'
#185410000000
1!
0$
b110 %
1'
0*
b110 +
#185420000000
0!
0'
#185430000000
1!
b111 %
1'
b111 +
#185440000000
0!
0'
#185450000000
1!
b1000 %
1'
b1000 +
#185460000000
0!
0'
#185470000000
1!
b1001 %
1'
b1001 +
#185480000000
0!
0'
#185490000000
1!
b0 %
1'
b0 +
#185500000000
0!
0'
#185510000000
1!
1$
b1 %
1'
1*
b1 +
#185520000000
0!
0'
#185530000000
1!
b10 %
1'
b10 +
#185540000000
1"
1(
#185550000000
0!
0"
b100 &
0'
0(
b100 ,
#185560000000
1!
b11 %
1'
b11 +
#185570000000
0!
0'
#185580000000
1!
b100 %
1'
b100 +
#185590000000
0!
0'
#185600000000
1!
b101 %
1'
b101 +
#185610000000
0!
0'
#185620000000
1!
b110 %
1'
b110 +
#185630000000
0!
0'
#185640000000
1!
b111 %
1'
b111 +
#185650000000
0!
0'
#185660000000
1!
0$
b1000 %
1'
0*
b1000 +
#185670000000
0!
0'
#185680000000
1!
b1001 %
1'
b1001 +
#185690000000
0!
0'
#185700000000
1!
b0 %
1'
b0 +
#185710000000
0!
0'
#185720000000
1!
1$
b1 %
1'
1*
b1 +
#185730000000
0!
0'
#185740000000
1!
b10 %
1'
b10 +
#185750000000
0!
0'
#185760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#185770000000
0!
0'
#185780000000
1!
b100 %
1'
b100 +
#185790000000
0!
0'
#185800000000
1!
b101 %
1'
b101 +
#185810000000
0!
0'
#185820000000
1!
0$
b110 %
1'
0*
b110 +
#185830000000
0!
0'
#185840000000
1!
b111 %
1'
b111 +
#185850000000
0!
0'
#185860000000
1!
b1000 %
1'
b1000 +
#185870000000
0!
0'
#185880000000
1!
b1001 %
1'
b1001 +
#185890000000
0!
0'
#185900000000
1!
b0 %
1'
b0 +
#185910000000
0!
0'
#185920000000
1!
1$
b1 %
1'
1*
b1 +
#185930000000
0!
0'
#185940000000
1!
b10 %
1'
b10 +
#185950000000
0!
0'
#185960000000
1!
b11 %
1'
b11 +
#185970000000
1"
1(
#185980000000
0!
0"
b100 &
0'
0(
b100 ,
#185990000000
1!
b100 %
1'
b100 +
#186000000000
0!
0'
#186010000000
1!
b101 %
1'
b101 +
#186020000000
0!
0'
#186030000000
1!
b110 %
1'
b110 +
#186040000000
0!
0'
#186050000000
1!
b111 %
1'
b111 +
#186060000000
0!
0'
#186070000000
1!
0$
b1000 %
1'
0*
b1000 +
#186080000000
0!
0'
#186090000000
1!
b1001 %
1'
b1001 +
#186100000000
0!
0'
#186110000000
1!
b0 %
1'
b0 +
#186120000000
0!
0'
#186130000000
1!
1$
b1 %
1'
1*
b1 +
#186140000000
0!
0'
#186150000000
1!
b10 %
1'
b10 +
#186160000000
0!
0'
#186170000000
1!
b11 %
1'
b11 +
#186180000000
0!
0'
#186190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#186200000000
0!
0'
#186210000000
1!
b101 %
1'
b101 +
#186220000000
0!
0'
#186230000000
1!
0$
b110 %
1'
0*
b110 +
#186240000000
0!
0'
#186250000000
1!
b111 %
1'
b111 +
#186260000000
0!
0'
#186270000000
1!
b1000 %
1'
b1000 +
#186280000000
0!
0'
#186290000000
1!
b1001 %
1'
b1001 +
#186300000000
0!
0'
#186310000000
1!
b0 %
1'
b0 +
#186320000000
0!
0'
#186330000000
1!
1$
b1 %
1'
1*
b1 +
#186340000000
0!
0'
#186350000000
1!
b10 %
1'
b10 +
#186360000000
0!
0'
#186370000000
1!
b11 %
1'
b11 +
#186380000000
0!
0'
#186390000000
1!
b100 %
1'
b100 +
#186400000000
1"
1(
#186410000000
0!
0"
b100 &
0'
0(
b100 ,
#186420000000
1!
b101 %
1'
b101 +
#186430000000
0!
0'
#186440000000
1!
b110 %
1'
b110 +
#186450000000
0!
0'
#186460000000
1!
b111 %
1'
b111 +
#186470000000
0!
0'
#186480000000
1!
0$
b1000 %
1'
0*
b1000 +
#186490000000
0!
0'
#186500000000
1!
b1001 %
1'
b1001 +
#186510000000
0!
0'
#186520000000
1!
b0 %
1'
b0 +
#186530000000
0!
0'
#186540000000
1!
1$
b1 %
1'
1*
b1 +
#186550000000
0!
0'
#186560000000
1!
b10 %
1'
b10 +
#186570000000
0!
0'
#186580000000
1!
b11 %
1'
b11 +
#186590000000
0!
0'
#186600000000
1!
b100 %
1'
b100 +
#186610000000
0!
0'
#186620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#186630000000
0!
0'
#186640000000
1!
0$
b110 %
1'
0*
b110 +
#186650000000
0!
0'
#186660000000
1!
b111 %
1'
b111 +
#186670000000
0!
0'
#186680000000
1!
b1000 %
1'
b1000 +
#186690000000
0!
0'
#186700000000
1!
b1001 %
1'
b1001 +
#186710000000
0!
0'
#186720000000
1!
b0 %
1'
b0 +
#186730000000
0!
0'
#186740000000
1!
1$
b1 %
1'
1*
b1 +
#186750000000
0!
0'
#186760000000
1!
b10 %
1'
b10 +
#186770000000
0!
0'
#186780000000
1!
b11 %
1'
b11 +
#186790000000
0!
0'
#186800000000
1!
b100 %
1'
b100 +
#186810000000
0!
0'
#186820000000
1!
b101 %
1'
b101 +
#186830000000
1"
1(
#186840000000
0!
0"
b100 &
0'
0(
b100 ,
#186850000000
1!
b110 %
1'
b110 +
#186860000000
0!
0'
#186870000000
1!
b111 %
1'
b111 +
#186880000000
0!
0'
#186890000000
1!
0$
b1000 %
1'
0*
b1000 +
#186900000000
0!
0'
#186910000000
1!
b1001 %
1'
b1001 +
#186920000000
0!
0'
#186930000000
1!
b0 %
1'
b0 +
#186940000000
0!
0'
#186950000000
1!
1$
b1 %
1'
1*
b1 +
#186960000000
0!
0'
#186970000000
1!
b10 %
1'
b10 +
#186980000000
0!
0'
#186990000000
1!
b11 %
1'
b11 +
#187000000000
0!
0'
#187010000000
1!
b100 %
1'
b100 +
#187020000000
0!
0'
#187030000000
1!
b101 %
1'
b101 +
#187040000000
0!
0'
#187050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#187060000000
0!
0'
#187070000000
1!
b111 %
1'
b111 +
#187080000000
0!
0'
#187090000000
1!
b1000 %
1'
b1000 +
#187100000000
0!
0'
#187110000000
1!
b1001 %
1'
b1001 +
#187120000000
0!
0'
#187130000000
1!
b0 %
1'
b0 +
#187140000000
0!
0'
#187150000000
1!
1$
b1 %
1'
1*
b1 +
#187160000000
0!
0'
#187170000000
1!
b10 %
1'
b10 +
#187180000000
0!
0'
#187190000000
1!
b11 %
1'
b11 +
#187200000000
0!
0'
#187210000000
1!
b100 %
1'
b100 +
#187220000000
0!
0'
#187230000000
1!
b101 %
1'
b101 +
#187240000000
0!
0'
#187250000000
1!
0$
b110 %
1'
0*
b110 +
#187260000000
1"
1(
#187270000000
0!
0"
b100 &
0'
0(
b100 ,
#187280000000
1!
1$
b111 %
1'
1*
b111 +
#187290000000
0!
0'
#187300000000
1!
0$
b1000 %
1'
0*
b1000 +
#187310000000
0!
0'
#187320000000
1!
b1001 %
1'
b1001 +
#187330000000
0!
0'
#187340000000
1!
b0 %
1'
b0 +
#187350000000
0!
0'
#187360000000
1!
1$
b1 %
1'
1*
b1 +
#187370000000
0!
0'
#187380000000
1!
b10 %
1'
b10 +
#187390000000
0!
0'
#187400000000
1!
b11 %
1'
b11 +
#187410000000
0!
0'
#187420000000
1!
b100 %
1'
b100 +
#187430000000
0!
0'
#187440000000
1!
b101 %
1'
b101 +
#187450000000
0!
0'
#187460000000
1!
b110 %
1'
b110 +
#187470000000
0!
0'
#187480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#187490000000
0!
0'
#187500000000
1!
b1000 %
1'
b1000 +
#187510000000
0!
0'
#187520000000
1!
b1001 %
1'
b1001 +
#187530000000
0!
0'
#187540000000
1!
b0 %
1'
b0 +
#187550000000
0!
0'
#187560000000
1!
1$
b1 %
1'
1*
b1 +
#187570000000
0!
0'
#187580000000
1!
b10 %
1'
b10 +
#187590000000
0!
0'
#187600000000
1!
b11 %
1'
b11 +
#187610000000
0!
0'
#187620000000
1!
b100 %
1'
b100 +
#187630000000
0!
0'
#187640000000
1!
b101 %
1'
b101 +
#187650000000
0!
0'
#187660000000
1!
0$
b110 %
1'
0*
b110 +
#187670000000
0!
0'
#187680000000
1!
b111 %
1'
b111 +
#187690000000
1"
1(
#187700000000
0!
0"
b100 &
0'
0(
b100 ,
#187710000000
1!
b1000 %
1'
b1000 +
#187720000000
0!
0'
#187730000000
1!
b1001 %
1'
b1001 +
#187740000000
0!
0'
#187750000000
1!
b0 %
1'
b0 +
#187760000000
0!
0'
#187770000000
1!
1$
b1 %
1'
1*
b1 +
#187780000000
0!
0'
#187790000000
1!
b10 %
1'
b10 +
#187800000000
0!
0'
#187810000000
1!
b11 %
1'
b11 +
#187820000000
0!
0'
#187830000000
1!
b100 %
1'
b100 +
#187840000000
0!
0'
#187850000000
1!
b101 %
1'
b101 +
#187860000000
0!
0'
#187870000000
1!
b110 %
1'
b110 +
#187880000000
0!
0'
#187890000000
1!
b111 %
1'
b111 +
#187900000000
0!
0'
#187910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#187920000000
0!
0'
#187930000000
1!
b1001 %
1'
b1001 +
#187940000000
0!
0'
#187950000000
1!
b0 %
1'
b0 +
#187960000000
0!
0'
#187970000000
1!
1$
b1 %
1'
1*
b1 +
#187980000000
0!
0'
#187990000000
1!
b10 %
1'
b10 +
#188000000000
0!
0'
#188010000000
1!
b11 %
1'
b11 +
#188020000000
0!
0'
#188030000000
1!
b100 %
1'
b100 +
#188040000000
0!
0'
#188050000000
1!
b101 %
1'
b101 +
#188060000000
0!
0'
#188070000000
1!
0$
b110 %
1'
0*
b110 +
#188080000000
0!
0'
#188090000000
1!
b111 %
1'
b111 +
#188100000000
0!
0'
#188110000000
1!
b1000 %
1'
b1000 +
#188120000000
1"
1(
#188130000000
0!
0"
b100 &
0'
0(
b100 ,
#188140000000
1!
b1001 %
1'
b1001 +
#188150000000
0!
0'
#188160000000
1!
b0 %
1'
b0 +
#188170000000
0!
0'
#188180000000
1!
1$
b1 %
1'
1*
b1 +
#188190000000
0!
0'
#188200000000
1!
b10 %
1'
b10 +
#188210000000
0!
0'
#188220000000
1!
b11 %
1'
b11 +
#188230000000
0!
0'
#188240000000
1!
b100 %
1'
b100 +
#188250000000
0!
0'
#188260000000
1!
b101 %
1'
b101 +
#188270000000
0!
0'
#188280000000
1!
b110 %
1'
b110 +
#188290000000
0!
0'
#188300000000
1!
b111 %
1'
b111 +
#188310000000
0!
0'
#188320000000
1!
0$
b1000 %
1'
0*
b1000 +
#188330000000
0!
0'
#188340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#188350000000
0!
0'
#188360000000
1!
b0 %
1'
b0 +
#188370000000
0!
0'
#188380000000
1!
1$
b1 %
1'
1*
b1 +
#188390000000
0!
0'
#188400000000
1!
b10 %
1'
b10 +
#188410000000
0!
0'
#188420000000
1!
b11 %
1'
b11 +
#188430000000
0!
0'
#188440000000
1!
b100 %
1'
b100 +
#188450000000
0!
0'
#188460000000
1!
b101 %
1'
b101 +
#188470000000
0!
0'
#188480000000
1!
0$
b110 %
1'
0*
b110 +
#188490000000
0!
0'
#188500000000
1!
b111 %
1'
b111 +
#188510000000
0!
0'
#188520000000
1!
b1000 %
1'
b1000 +
#188530000000
0!
0'
#188540000000
1!
b1001 %
1'
b1001 +
#188550000000
1"
1(
#188560000000
0!
0"
b100 &
0'
0(
b100 ,
#188570000000
1!
b0 %
1'
b0 +
#188580000000
0!
0'
#188590000000
1!
1$
b1 %
1'
1*
b1 +
#188600000000
0!
0'
#188610000000
1!
b10 %
1'
b10 +
#188620000000
0!
0'
#188630000000
1!
b11 %
1'
b11 +
#188640000000
0!
0'
#188650000000
1!
b100 %
1'
b100 +
#188660000000
0!
0'
#188670000000
1!
b101 %
1'
b101 +
#188680000000
0!
0'
#188690000000
1!
b110 %
1'
b110 +
#188700000000
0!
0'
#188710000000
1!
b111 %
1'
b111 +
#188720000000
0!
0'
#188730000000
1!
0$
b1000 %
1'
0*
b1000 +
#188740000000
0!
0'
#188750000000
1!
b1001 %
1'
b1001 +
#188760000000
0!
0'
#188770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#188780000000
0!
0'
#188790000000
1!
1$
b1 %
1'
1*
b1 +
#188800000000
0!
0'
#188810000000
1!
b10 %
1'
b10 +
#188820000000
0!
0'
#188830000000
1!
b11 %
1'
b11 +
#188840000000
0!
0'
#188850000000
1!
b100 %
1'
b100 +
#188860000000
0!
0'
#188870000000
1!
b101 %
1'
b101 +
#188880000000
0!
0'
#188890000000
1!
0$
b110 %
1'
0*
b110 +
#188900000000
0!
0'
#188910000000
1!
b111 %
1'
b111 +
#188920000000
0!
0'
#188930000000
1!
b1000 %
1'
b1000 +
#188940000000
0!
0'
#188950000000
1!
b1001 %
1'
b1001 +
#188960000000
0!
0'
#188970000000
1!
b0 %
1'
b0 +
#188980000000
1"
1(
#188990000000
0!
0"
b100 &
0'
0(
b100 ,
#189000000000
1!
1$
b1 %
1'
1*
b1 +
#189010000000
0!
0'
#189020000000
1!
b10 %
1'
b10 +
#189030000000
0!
0'
#189040000000
1!
b11 %
1'
b11 +
#189050000000
0!
0'
#189060000000
1!
b100 %
1'
b100 +
#189070000000
0!
0'
#189080000000
1!
b101 %
1'
b101 +
#189090000000
0!
0'
#189100000000
1!
b110 %
1'
b110 +
#189110000000
0!
0'
#189120000000
1!
b111 %
1'
b111 +
#189130000000
0!
0'
#189140000000
1!
0$
b1000 %
1'
0*
b1000 +
#189150000000
0!
0'
#189160000000
1!
b1001 %
1'
b1001 +
#189170000000
0!
0'
#189180000000
1!
b0 %
1'
b0 +
#189190000000
0!
0'
#189200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#189210000000
0!
0'
#189220000000
1!
b10 %
1'
b10 +
#189230000000
0!
0'
#189240000000
1!
b11 %
1'
b11 +
#189250000000
0!
0'
#189260000000
1!
b100 %
1'
b100 +
#189270000000
0!
0'
#189280000000
1!
b101 %
1'
b101 +
#189290000000
0!
0'
#189300000000
1!
0$
b110 %
1'
0*
b110 +
#189310000000
0!
0'
#189320000000
1!
b111 %
1'
b111 +
#189330000000
0!
0'
#189340000000
1!
b1000 %
1'
b1000 +
#189350000000
0!
0'
#189360000000
1!
b1001 %
1'
b1001 +
#189370000000
0!
0'
#189380000000
1!
b0 %
1'
b0 +
#189390000000
0!
0'
#189400000000
1!
1$
b1 %
1'
1*
b1 +
#189410000000
1"
1(
#189420000000
0!
0"
b100 &
0'
0(
b100 ,
#189430000000
1!
b10 %
1'
b10 +
#189440000000
0!
0'
#189450000000
1!
b11 %
1'
b11 +
#189460000000
0!
0'
#189470000000
1!
b100 %
1'
b100 +
#189480000000
0!
0'
#189490000000
1!
b101 %
1'
b101 +
#189500000000
0!
0'
#189510000000
1!
b110 %
1'
b110 +
#189520000000
0!
0'
#189530000000
1!
b111 %
1'
b111 +
#189540000000
0!
0'
#189550000000
1!
0$
b1000 %
1'
0*
b1000 +
#189560000000
0!
0'
#189570000000
1!
b1001 %
1'
b1001 +
#189580000000
0!
0'
#189590000000
1!
b0 %
1'
b0 +
#189600000000
0!
0'
#189610000000
1!
1$
b1 %
1'
1*
b1 +
#189620000000
0!
0'
#189630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#189640000000
0!
0'
#189650000000
1!
b11 %
1'
b11 +
#189660000000
0!
0'
#189670000000
1!
b100 %
1'
b100 +
#189680000000
0!
0'
#189690000000
1!
b101 %
1'
b101 +
#189700000000
0!
0'
#189710000000
1!
0$
b110 %
1'
0*
b110 +
#189720000000
0!
0'
#189730000000
1!
b111 %
1'
b111 +
#189740000000
0!
0'
#189750000000
1!
b1000 %
1'
b1000 +
#189760000000
0!
0'
#189770000000
1!
b1001 %
1'
b1001 +
#189780000000
0!
0'
#189790000000
1!
b0 %
1'
b0 +
#189800000000
0!
0'
#189810000000
1!
1$
b1 %
1'
1*
b1 +
#189820000000
0!
0'
#189830000000
1!
b10 %
1'
b10 +
#189840000000
1"
1(
#189850000000
0!
0"
b100 &
0'
0(
b100 ,
#189860000000
1!
b11 %
1'
b11 +
#189870000000
0!
0'
#189880000000
1!
b100 %
1'
b100 +
#189890000000
0!
0'
#189900000000
1!
b101 %
1'
b101 +
#189910000000
0!
0'
#189920000000
1!
b110 %
1'
b110 +
#189930000000
0!
0'
#189940000000
1!
b111 %
1'
b111 +
#189950000000
0!
0'
#189960000000
1!
0$
b1000 %
1'
0*
b1000 +
#189970000000
0!
0'
#189980000000
1!
b1001 %
1'
b1001 +
#189990000000
0!
0'
#190000000000
1!
b0 %
1'
b0 +
#190010000000
0!
0'
#190020000000
1!
1$
b1 %
1'
1*
b1 +
#190030000000
0!
0'
#190040000000
1!
b10 %
1'
b10 +
#190050000000
0!
0'
#190060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#190070000000
0!
0'
#190080000000
1!
b100 %
1'
b100 +
#190090000000
0!
0'
#190100000000
1!
b101 %
1'
b101 +
#190110000000
0!
0'
#190120000000
1!
0$
b110 %
1'
0*
b110 +
#190130000000
0!
0'
#190140000000
1!
b111 %
1'
b111 +
#190150000000
0!
0'
#190160000000
1!
b1000 %
1'
b1000 +
#190170000000
0!
0'
#190180000000
1!
b1001 %
1'
b1001 +
#190190000000
0!
0'
#190200000000
1!
b0 %
1'
b0 +
#190210000000
0!
0'
#190220000000
1!
1$
b1 %
1'
1*
b1 +
#190230000000
0!
0'
#190240000000
1!
b10 %
1'
b10 +
#190250000000
0!
0'
#190260000000
1!
b11 %
1'
b11 +
#190270000000
1"
1(
#190280000000
0!
0"
b100 &
0'
0(
b100 ,
#190290000000
1!
b100 %
1'
b100 +
#190300000000
0!
0'
#190310000000
1!
b101 %
1'
b101 +
#190320000000
0!
0'
#190330000000
1!
b110 %
1'
b110 +
#190340000000
0!
0'
#190350000000
1!
b111 %
1'
b111 +
#190360000000
0!
0'
#190370000000
1!
0$
b1000 %
1'
0*
b1000 +
#190380000000
0!
0'
#190390000000
1!
b1001 %
1'
b1001 +
#190400000000
0!
0'
#190410000000
1!
b0 %
1'
b0 +
#190420000000
0!
0'
#190430000000
1!
1$
b1 %
1'
1*
b1 +
#190440000000
0!
0'
#190450000000
1!
b10 %
1'
b10 +
#190460000000
0!
0'
#190470000000
1!
b11 %
1'
b11 +
#190480000000
0!
0'
#190490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#190500000000
0!
0'
#190510000000
1!
b101 %
1'
b101 +
#190520000000
0!
0'
#190530000000
1!
0$
b110 %
1'
0*
b110 +
#190540000000
0!
0'
#190550000000
1!
b111 %
1'
b111 +
#190560000000
0!
0'
#190570000000
1!
b1000 %
1'
b1000 +
#190580000000
0!
0'
#190590000000
1!
b1001 %
1'
b1001 +
#190600000000
0!
0'
#190610000000
1!
b0 %
1'
b0 +
#190620000000
0!
0'
#190630000000
1!
1$
b1 %
1'
1*
b1 +
#190640000000
0!
0'
#190650000000
1!
b10 %
1'
b10 +
#190660000000
0!
0'
#190670000000
1!
b11 %
1'
b11 +
#190680000000
0!
0'
#190690000000
1!
b100 %
1'
b100 +
#190700000000
1"
1(
#190710000000
0!
0"
b100 &
0'
0(
b100 ,
#190720000000
1!
b101 %
1'
b101 +
#190730000000
0!
0'
#190740000000
1!
b110 %
1'
b110 +
#190750000000
0!
0'
#190760000000
1!
b111 %
1'
b111 +
#190770000000
0!
0'
#190780000000
1!
0$
b1000 %
1'
0*
b1000 +
#190790000000
0!
0'
#190800000000
1!
b1001 %
1'
b1001 +
#190810000000
0!
0'
#190820000000
1!
b0 %
1'
b0 +
#190830000000
0!
0'
#190840000000
1!
1$
b1 %
1'
1*
b1 +
#190850000000
0!
0'
#190860000000
1!
b10 %
1'
b10 +
#190870000000
0!
0'
#190880000000
1!
b11 %
1'
b11 +
#190890000000
0!
0'
#190900000000
1!
b100 %
1'
b100 +
#190910000000
0!
0'
#190920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#190930000000
0!
0'
#190940000000
1!
0$
b110 %
1'
0*
b110 +
#190950000000
0!
0'
#190960000000
1!
b111 %
1'
b111 +
#190970000000
0!
0'
#190980000000
1!
b1000 %
1'
b1000 +
#190990000000
0!
0'
#191000000000
1!
b1001 %
1'
b1001 +
#191010000000
0!
0'
#191020000000
1!
b0 %
1'
b0 +
#191030000000
0!
0'
#191040000000
1!
1$
b1 %
1'
1*
b1 +
#191050000000
0!
0'
#191060000000
1!
b10 %
1'
b10 +
#191070000000
0!
0'
#191080000000
1!
b11 %
1'
b11 +
#191090000000
0!
0'
#191100000000
1!
b100 %
1'
b100 +
#191110000000
0!
0'
#191120000000
1!
b101 %
1'
b101 +
#191130000000
1"
1(
#191140000000
0!
0"
b100 &
0'
0(
b100 ,
#191150000000
1!
b110 %
1'
b110 +
#191160000000
0!
0'
#191170000000
1!
b111 %
1'
b111 +
#191180000000
0!
0'
#191190000000
1!
0$
b1000 %
1'
0*
b1000 +
#191200000000
0!
0'
#191210000000
1!
b1001 %
1'
b1001 +
#191220000000
0!
0'
#191230000000
1!
b0 %
1'
b0 +
#191240000000
0!
0'
#191250000000
1!
1$
b1 %
1'
1*
b1 +
#191260000000
0!
0'
#191270000000
1!
b10 %
1'
b10 +
#191280000000
0!
0'
#191290000000
1!
b11 %
1'
b11 +
#191300000000
0!
0'
#191310000000
1!
b100 %
1'
b100 +
#191320000000
0!
0'
#191330000000
1!
b101 %
1'
b101 +
#191340000000
0!
0'
#191350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#191360000000
0!
0'
#191370000000
1!
b111 %
1'
b111 +
#191380000000
0!
0'
#191390000000
1!
b1000 %
1'
b1000 +
#191400000000
0!
0'
#191410000000
1!
b1001 %
1'
b1001 +
#191420000000
0!
0'
#191430000000
1!
b0 %
1'
b0 +
#191440000000
0!
0'
#191450000000
1!
1$
b1 %
1'
1*
b1 +
#191460000000
0!
0'
#191470000000
1!
b10 %
1'
b10 +
#191480000000
0!
0'
#191490000000
1!
b11 %
1'
b11 +
#191500000000
0!
0'
#191510000000
1!
b100 %
1'
b100 +
#191520000000
0!
0'
#191530000000
1!
b101 %
1'
b101 +
#191540000000
0!
0'
#191550000000
1!
0$
b110 %
1'
0*
b110 +
#191560000000
1"
1(
#191570000000
0!
0"
b100 &
0'
0(
b100 ,
#191580000000
1!
1$
b111 %
1'
1*
b111 +
#191590000000
0!
0'
#191600000000
1!
0$
b1000 %
1'
0*
b1000 +
#191610000000
0!
0'
#191620000000
1!
b1001 %
1'
b1001 +
#191630000000
0!
0'
#191640000000
1!
b0 %
1'
b0 +
#191650000000
0!
0'
#191660000000
1!
1$
b1 %
1'
1*
b1 +
#191670000000
0!
0'
#191680000000
1!
b10 %
1'
b10 +
#191690000000
0!
0'
#191700000000
1!
b11 %
1'
b11 +
#191710000000
0!
0'
#191720000000
1!
b100 %
1'
b100 +
#191730000000
0!
0'
#191740000000
1!
b101 %
1'
b101 +
#191750000000
0!
0'
#191760000000
1!
b110 %
1'
b110 +
#191770000000
0!
0'
#191780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#191790000000
0!
0'
#191800000000
1!
b1000 %
1'
b1000 +
#191810000000
0!
0'
#191820000000
1!
b1001 %
1'
b1001 +
#191830000000
0!
0'
#191840000000
1!
b0 %
1'
b0 +
#191850000000
0!
0'
#191860000000
1!
1$
b1 %
1'
1*
b1 +
#191870000000
0!
0'
#191880000000
1!
b10 %
1'
b10 +
#191890000000
0!
0'
#191900000000
1!
b11 %
1'
b11 +
#191910000000
0!
0'
#191920000000
1!
b100 %
1'
b100 +
#191930000000
0!
0'
#191940000000
1!
b101 %
1'
b101 +
#191950000000
0!
0'
#191960000000
1!
0$
b110 %
1'
0*
b110 +
#191970000000
0!
0'
#191980000000
1!
b111 %
1'
b111 +
#191990000000
1"
1(
#192000000000
0!
0"
b100 &
0'
0(
b100 ,
#192010000000
1!
b1000 %
1'
b1000 +
#192020000000
0!
0'
#192030000000
1!
b1001 %
1'
b1001 +
#192040000000
0!
0'
#192050000000
1!
b0 %
1'
b0 +
#192060000000
0!
0'
#192070000000
1!
1$
b1 %
1'
1*
b1 +
#192080000000
0!
0'
#192090000000
1!
b10 %
1'
b10 +
#192100000000
0!
0'
#192110000000
1!
b11 %
1'
b11 +
#192120000000
0!
0'
#192130000000
1!
b100 %
1'
b100 +
#192140000000
0!
0'
#192150000000
1!
b101 %
1'
b101 +
#192160000000
0!
0'
#192170000000
1!
b110 %
1'
b110 +
#192180000000
0!
0'
#192190000000
1!
b111 %
1'
b111 +
#192200000000
0!
0'
#192210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#192220000000
0!
0'
#192230000000
1!
b1001 %
1'
b1001 +
#192240000000
0!
0'
#192250000000
1!
b0 %
1'
b0 +
#192260000000
0!
0'
#192270000000
1!
1$
b1 %
1'
1*
b1 +
#192280000000
0!
0'
#192290000000
1!
b10 %
1'
b10 +
#192300000000
0!
0'
#192310000000
1!
b11 %
1'
b11 +
#192320000000
0!
0'
#192330000000
1!
b100 %
1'
b100 +
#192340000000
0!
0'
#192350000000
1!
b101 %
1'
b101 +
#192360000000
0!
0'
#192370000000
1!
0$
b110 %
1'
0*
b110 +
#192380000000
0!
0'
#192390000000
1!
b111 %
1'
b111 +
#192400000000
0!
0'
#192410000000
1!
b1000 %
1'
b1000 +
#192420000000
1"
1(
#192430000000
0!
0"
b100 &
0'
0(
b100 ,
#192440000000
1!
b1001 %
1'
b1001 +
#192450000000
0!
0'
#192460000000
1!
b0 %
1'
b0 +
#192470000000
0!
0'
#192480000000
1!
1$
b1 %
1'
1*
b1 +
#192490000000
0!
0'
#192500000000
1!
b10 %
1'
b10 +
#192510000000
0!
0'
#192520000000
1!
b11 %
1'
b11 +
#192530000000
0!
0'
#192540000000
1!
b100 %
1'
b100 +
#192550000000
0!
0'
#192560000000
1!
b101 %
1'
b101 +
#192570000000
0!
0'
#192580000000
1!
b110 %
1'
b110 +
#192590000000
0!
0'
#192600000000
1!
b111 %
1'
b111 +
#192610000000
0!
0'
#192620000000
1!
0$
b1000 %
1'
0*
b1000 +
#192630000000
0!
0'
#192640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#192650000000
0!
0'
#192660000000
1!
b0 %
1'
b0 +
#192670000000
0!
0'
#192680000000
1!
1$
b1 %
1'
1*
b1 +
#192690000000
0!
0'
#192700000000
1!
b10 %
1'
b10 +
#192710000000
0!
0'
#192720000000
1!
b11 %
1'
b11 +
#192730000000
0!
0'
#192740000000
1!
b100 %
1'
b100 +
#192750000000
0!
0'
#192760000000
1!
b101 %
1'
b101 +
#192770000000
0!
0'
#192780000000
1!
0$
b110 %
1'
0*
b110 +
#192790000000
0!
0'
#192800000000
1!
b111 %
1'
b111 +
#192810000000
0!
0'
#192820000000
1!
b1000 %
1'
b1000 +
#192830000000
0!
0'
#192840000000
1!
b1001 %
1'
b1001 +
#192850000000
1"
1(
#192860000000
0!
0"
b100 &
0'
0(
b100 ,
#192870000000
1!
b0 %
1'
b0 +
#192880000000
0!
0'
#192890000000
1!
1$
b1 %
1'
1*
b1 +
#192900000000
0!
0'
#192910000000
1!
b10 %
1'
b10 +
#192920000000
0!
0'
#192930000000
1!
b11 %
1'
b11 +
#192940000000
0!
0'
#192950000000
1!
b100 %
1'
b100 +
#192960000000
0!
0'
#192970000000
1!
b101 %
1'
b101 +
#192980000000
0!
0'
#192990000000
1!
b110 %
1'
b110 +
#193000000000
0!
0'
#193010000000
1!
b111 %
1'
b111 +
#193020000000
0!
0'
#193030000000
1!
0$
b1000 %
1'
0*
b1000 +
#193040000000
0!
0'
#193050000000
1!
b1001 %
1'
b1001 +
#193060000000
0!
0'
#193070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#193080000000
0!
0'
#193090000000
1!
1$
b1 %
1'
1*
b1 +
#193100000000
0!
0'
#193110000000
1!
b10 %
1'
b10 +
#193120000000
0!
0'
#193130000000
1!
b11 %
1'
b11 +
#193140000000
0!
0'
#193150000000
1!
b100 %
1'
b100 +
#193160000000
0!
0'
#193170000000
1!
b101 %
1'
b101 +
#193180000000
0!
0'
#193190000000
1!
0$
b110 %
1'
0*
b110 +
#193200000000
0!
0'
#193210000000
1!
b111 %
1'
b111 +
#193220000000
0!
0'
#193230000000
1!
b1000 %
1'
b1000 +
#193240000000
0!
0'
#193250000000
1!
b1001 %
1'
b1001 +
#193260000000
0!
0'
#193270000000
1!
b0 %
1'
b0 +
#193280000000
1"
1(
#193290000000
0!
0"
b100 &
0'
0(
b100 ,
#193300000000
1!
1$
b1 %
1'
1*
b1 +
#193310000000
0!
0'
#193320000000
1!
b10 %
1'
b10 +
#193330000000
0!
0'
#193340000000
1!
b11 %
1'
b11 +
#193350000000
0!
0'
#193360000000
1!
b100 %
1'
b100 +
#193370000000
0!
0'
#193380000000
1!
b101 %
1'
b101 +
#193390000000
0!
0'
#193400000000
1!
b110 %
1'
b110 +
#193410000000
0!
0'
#193420000000
1!
b111 %
1'
b111 +
#193430000000
0!
0'
#193440000000
1!
0$
b1000 %
1'
0*
b1000 +
#193450000000
0!
0'
#193460000000
1!
b1001 %
1'
b1001 +
#193470000000
0!
0'
#193480000000
1!
b0 %
1'
b0 +
#193490000000
0!
0'
#193500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#193510000000
0!
0'
#193520000000
1!
b10 %
1'
b10 +
#193530000000
0!
0'
#193540000000
1!
b11 %
1'
b11 +
#193550000000
0!
0'
#193560000000
1!
b100 %
1'
b100 +
#193570000000
0!
0'
#193580000000
1!
b101 %
1'
b101 +
#193590000000
0!
0'
#193600000000
1!
0$
b110 %
1'
0*
b110 +
#193610000000
0!
0'
#193620000000
1!
b111 %
1'
b111 +
#193630000000
0!
0'
#193640000000
1!
b1000 %
1'
b1000 +
#193650000000
0!
0'
#193660000000
1!
b1001 %
1'
b1001 +
#193670000000
0!
0'
#193680000000
1!
b0 %
1'
b0 +
#193690000000
0!
0'
#193700000000
1!
1$
b1 %
1'
1*
b1 +
#193710000000
1"
1(
#193720000000
0!
0"
b100 &
0'
0(
b100 ,
#193730000000
1!
b10 %
1'
b10 +
#193740000000
0!
0'
#193750000000
1!
b11 %
1'
b11 +
#193760000000
0!
0'
#193770000000
1!
b100 %
1'
b100 +
#193780000000
0!
0'
#193790000000
1!
b101 %
1'
b101 +
#193800000000
0!
0'
#193810000000
1!
b110 %
1'
b110 +
#193820000000
0!
0'
#193830000000
1!
b111 %
1'
b111 +
#193840000000
0!
0'
#193850000000
1!
0$
b1000 %
1'
0*
b1000 +
#193860000000
0!
0'
#193870000000
1!
b1001 %
1'
b1001 +
#193880000000
0!
0'
#193890000000
1!
b0 %
1'
b0 +
#193900000000
0!
0'
#193910000000
1!
1$
b1 %
1'
1*
b1 +
#193920000000
0!
0'
#193930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#193940000000
0!
0'
#193950000000
1!
b11 %
1'
b11 +
#193960000000
0!
0'
#193970000000
1!
b100 %
1'
b100 +
#193980000000
0!
0'
#193990000000
1!
b101 %
1'
b101 +
#194000000000
0!
0'
#194010000000
1!
0$
b110 %
1'
0*
b110 +
#194020000000
0!
0'
#194030000000
1!
b111 %
1'
b111 +
#194040000000
0!
0'
#194050000000
1!
b1000 %
1'
b1000 +
#194060000000
0!
0'
#194070000000
1!
b1001 %
1'
b1001 +
#194080000000
0!
0'
#194090000000
1!
b0 %
1'
b0 +
#194100000000
0!
0'
#194110000000
1!
1$
b1 %
1'
1*
b1 +
#194120000000
0!
0'
#194130000000
1!
b10 %
1'
b10 +
#194140000000
1"
1(
#194150000000
0!
0"
b100 &
0'
0(
b100 ,
#194160000000
1!
b11 %
1'
b11 +
#194170000000
0!
0'
#194180000000
1!
b100 %
1'
b100 +
#194190000000
0!
0'
#194200000000
1!
b101 %
1'
b101 +
#194210000000
0!
0'
#194220000000
1!
b110 %
1'
b110 +
#194230000000
0!
0'
#194240000000
1!
b111 %
1'
b111 +
#194250000000
0!
0'
#194260000000
1!
0$
b1000 %
1'
0*
b1000 +
#194270000000
0!
0'
#194280000000
1!
b1001 %
1'
b1001 +
#194290000000
0!
0'
#194300000000
1!
b0 %
1'
b0 +
#194310000000
0!
0'
#194320000000
1!
1$
b1 %
1'
1*
b1 +
#194330000000
0!
0'
#194340000000
1!
b10 %
1'
b10 +
#194350000000
0!
0'
#194360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#194370000000
0!
0'
#194380000000
1!
b100 %
1'
b100 +
#194390000000
0!
0'
#194400000000
1!
b101 %
1'
b101 +
#194410000000
0!
0'
#194420000000
1!
0$
b110 %
1'
0*
b110 +
#194430000000
0!
0'
#194440000000
1!
b111 %
1'
b111 +
#194450000000
0!
0'
#194460000000
1!
b1000 %
1'
b1000 +
#194470000000
0!
0'
#194480000000
1!
b1001 %
1'
b1001 +
#194490000000
0!
0'
#194500000000
1!
b0 %
1'
b0 +
#194510000000
0!
0'
#194520000000
1!
1$
b1 %
1'
1*
b1 +
#194530000000
0!
0'
#194540000000
1!
b10 %
1'
b10 +
#194550000000
0!
0'
#194560000000
1!
b11 %
1'
b11 +
#194570000000
1"
1(
#194580000000
0!
0"
b100 &
0'
0(
b100 ,
#194590000000
1!
b100 %
1'
b100 +
#194600000000
0!
0'
#194610000000
1!
b101 %
1'
b101 +
#194620000000
0!
0'
#194630000000
1!
b110 %
1'
b110 +
#194640000000
0!
0'
#194650000000
1!
b111 %
1'
b111 +
#194660000000
0!
0'
#194670000000
1!
0$
b1000 %
1'
0*
b1000 +
#194680000000
0!
0'
#194690000000
1!
b1001 %
1'
b1001 +
#194700000000
0!
0'
#194710000000
1!
b0 %
1'
b0 +
#194720000000
0!
0'
#194730000000
1!
1$
b1 %
1'
1*
b1 +
#194740000000
0!
0'
#194750000000
1!
b10 %
1'
b10 +
#194760000000
0!
0'
#194770000000
1!
b11 %
1'
b11 +
#194780000000
0!
0'
#194790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#194800000000
0!
0'
#194810000000
1!
b101 %
1'
b101 +
#194820000000
0!
0'
#194830000000
1!
0$
b110 %
1'
0*
b110 +
#194840000000
0!
0'
#194850000000
1!
b111 %
1'
b111 +
#194860000000
0!
0'
#194870000000
1!
b1000 %
1'
b1000 +
#194880000000
0!
0'
#194890000000
1!
b1001 %
1'
b1001 +
#194900000000
0!
0'
#194910000000
1!
b0 %
1'
b0 +
#194920000000
0!
0'
#194930000000
1!
1$
b1 %
1'
1*
b1 +
#194940000000
0!
0'
#194950000000
1!
b10 %
1'
b10 +
#194960000000
0!
0'
#194970000000
1!
b11 %
1'
b11 +
#194980000000
0!
0'
#194990000000
1!
b100 %
1'
b100 +
#195000000000
1"
1(
#195010000000
0!
0"
b100 &
0'
0(
b100 ,
#195020000000
1!
b101 %
1'
b101 +
#195030000000
0!
0'
#195040000000
1!
b110 %
1'
b110 +
#195050000000
0!
0'
#195060000000
1!
b111 %
1'
b111 +
#195070000000
0!
0'
#195080000000
1!
0$
b1000 %
1'
0*
b1000 +
#195090000000
0!
0'
#195100000000
1!
b1001 %
1'
b1001 +
#195110000000
0!
0'
#195120000000
1!
b0 %
1'
b0 +
#195130000000
0!
0'
#195140000000
1!
1$
b1 %
1'
1*
b1 +
#195150000000
0!
0'
#195160000000
1!
b10 %
1'
b10 +
#195170000000
0!
0'
#195180000000
1!
b11 %
1'
b11 +
#195190000000
0!
0'
#195200000000
1!
b100 %
1'
b100 +
#195210000000
0!
0'
#195220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#195230000000
0!
0'
#195240000000
1!
0$
b110 %
1'
0*
b110 +
#195250000000
0!
0'
#195260000000
1!
b111 %
1'
b111 +
#195270000000
0!
0'
#195280000000
1!
b1000 %
1'
b1000 +
#195290000000
0!
0'
#195300000000
1!
b1001 %
1'
b1001 +
#195310000000
0!
0'
#195320000000
1!
b0 %
1'
b0 +
#195330000000
0!
0'
#195340000000
1!
1$
b1 %
1'
1*
b1 +
#195350000000
0!
0'
#195360000000
1!
b10 %
1'
b10 +
#195370000000
0!
0'
#195380000000
1!
b11 %
1'
b11 +
#195390000000
0!
0'
#195400000000
1!
b100 %
1'
b100 +
#195410000000
0!
0'
#195420000000
1!
b101 %
1'
b101 +
#195430000000
1"
1(
#195440000000
0!
0"
b100 &
0'
0(
b100 ,
#195450000000
1!
b110 %
1'
b110 +
#195460000000
0!
0'
#195470000000
1!
b111 %
1'
b111 +
#195480000000
0!
0'
#195490000000
1!
0$
b1000 %
1'
0*
b1000 +
#195500000000
0!
0'
#195510000000
1!
b1001 %
1'
b1001 +
#195520000000
0!
0'
#195530000000
1!
b0 %
1'
b0 +
#195540000000
0!
0'
#195550000000
1!
1$
b1 %
1'
1*
b1 +
#195560000000
0!
0'
#195570000000
1!
b10 %
1'
b10 +
#195580000000
0!
0'
#195590000000
1!
b11 %
1'
b11 +
#195600000000
0!
0'
#195610000000
1!
b100 %
1'
b100 +
#195620000000
0!
0'
#195630000000
1!
b101 %
1'
b101 +
#195640000000
0!
0'
#195650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#195660000000
0!
0'
#195670000000
1!
b111 %
1'
b111 +
#195680000000
0!
0'
#195690000000
1!
b1000 %
1'
b1000 +
#195700000000
0!
0'
#195710000000
1!
b1001 %
1'
b1001 +
#195720000000
0!
0'
#195730000000
1!
b0 %
1'
b0 +
#195740000000
0!
0'
#195750000000
1!
1$
b1 %
1'
1*
b1 +
#195760000000
0!
0'
#195770000000
1!
b10 %
1'
b10 +
#195780000000
0!
0'
#195790000000
1!
b11 %
1'
b11 +
#195800000000
0!
0'
#195810000000
1!
b100 %
1'
b100 +
#195820000000
0!
0'
#195830000000
1!
b101 %
1'
b101 +
#195840000000
0!
0'
#195850000000
1!
0$
b110 %
1'
0*
b110 +
#195860000000
1"
1(
#195870000000
0!
0"
b100 &
0'
0(
b100 ,
#195880000000
1!
1$
b111 %
1'
1*
b111 +
#195890000000
0!
0'
#195900000000
1!
0$
b1000 %
1'
0*
b1000 +
#195910000000
0!
0'
#195920000000
1!
b1001 %
1'
b1001 +
#195930000000
0!
0'
#195940000000
1!
b0 %
1'
b0 +
#195950000000
0!
0'
#195960000000
1!
1$
b1 %
1'
1*
b1 +
#195970000000
0!
0'
#195980000000
1!
b10 %
1'
b10 +
#195990000000
0!
0'
#196000000000
1!
b11 %
1'
b11 +
#196010000000
0!
0'
#196020000000
1!
b100 %
1'
b100 +
#196030000000
0!
0'
#196040000000
1!
b101 %
1'
b101 +
#196050000000
0!
0'
#196060000000
1!
b110 %
1'
b110 +
#196070000000
0!
0'
#196080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#196090000000
0!
0'
#196100000000
1!
b1000 %
1'
b1000 +
#196110000000
0!
0'
#196120000000
1!
b1001 %
1'
b1001 +
#196130000000
0!
0'
#196140000000
1!
b0 %
1'
b0 +
#196150000000
0!
0'
#196160000000
1!
1$
b1 %
1'
1*
b1 +
#196170000000
0!
0'
#196180000000
1!
b10 %
1'
b10 +
#196190000000
0!
0'
#196200000000
1!
b11 %
1'
b11 +
#196210000000
0!
0'
#196220000000
1!
b100 %
1'
b100 +
#196230000000
0!
0'
#196240000000
1!
b101 %
1'
b101 +
#196250000000
0!
0'
#196260000000
1!
0$
b110 %
1'
0*
b110 +
#196270000000
0!
0'
#196280000000
1!
b111 %
1'
b111 +
#196290000000
1"
1(
#196300000000
0!
0"
b100 &
0'
0(
b100 ,
#196310000000
1!
b1000 %
1'
b1000 +
#196320000000
0!
0'
#196330000000
1!
b1001 %
1'
b1001 +
#196340000000
0!
0'
#196350000000
1!
b0 %
1'
b0 +
#196360000000
0!
0'
#196370000000
1!
1$
b1 %
1'
1*
b1 +
#196380000000
0!
0'
#196390000000
1!
b10 %
1'
b10 +
#196400000000
0!
0'
#196410000000
1!
b11 %
1'
b11 +
#196420000000
0!
0'
#196430000000
1!
b100 %
1'
b100 +
#196440000000
0!
0'
#196450000000
1!
b101 %
1'
b101 +
#196460000000
0!
0'
#196470000000
1!
b110 %
1'
b110 +
#196480000000
0!
0'
#196490000000
1!
b111 %
1'
b111 +
#196500000000
0!
0'
#196510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#196520000000
0!
0'
#196530000000
1!
b1001 %
1'
b1001 +
#196540000000
0!
0'
#196550000000
1!
b0 %
1'
b0 +
#196560000000
0!
0'
#196570000000
1!
1$
b1 %
1'
1*
b1 +
#196580000000
0!
0'
#196590000000
1!
b10 %
1'
b10 +
#196600000000
0!
0'
#196610000000
1!
b11 %
1'
b11 +
#196620000000
0!
0'
#196630000000
1!
b100 %
1'
b100 +
#196640000000
0!
0'
#196650000000
1!
b101 %
1'
b101 +
#196660000000
0!
0'
#196670000000
1!
0$
b110 %
1'
0*
b110 +
#196680000000
0!
0'
#196690000000
1!
b111 %
1'
b111 +
#196700000000
0!
0'
#196710000000
1!
b1000 %
1'
b1000 +
#196720000000
1"
1(
#196730000000
0!
0"
b100 &
0'
0(
b100 ,
#196740000000
1!
b1001 %
1'
b1001 +
#196750000000
0!
0'
#196760000000
1!
b0 %
1'
b0 +
#196770000000
0!
0'
#196780000000
1!
1$
b1 %
1'
1*
b1 +
#196790000000
0!
0'
#196800000000
1!
b10 %
1'
b10 +
#196810000000
0!
0'
#196820000000
1!
b11 %
1'
b11 +
#196830000000
0!
0'
#196840000000
1!
b100 %
1'
b100 +
#196850000000
0!
0'
#196860000000
1!
b101 %
1'
b101 +
#196870000000
0!
0'
#196880000000
1!
b110 %
1'
b110 +
#196890000000
0!
0'
#196900000000
1!
b111 %
1'
b111 +
#196910000000
0!
0'
#196920000000
1!
0$
b1000 %
1'
0*
b1000 +
#196930000000
0!
0'
#196940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#196950000000
0!
0'
#196960000000
1!
b0 %
1'
b0 +
#196970000000
0!
0'
#196980000000
1!
1$
b1 %
1'
1*
b1 +
#196990000000
0!
0'
#197000000000
1!
b10 %
1'
b10 +
#197010000000
0!
0'
#197020000000
1!
b11 %
1'
b11 +
#197030000000
0!
0'
#197040000000
1!
b100 %
1'
b100 +
#197050000000
0!
0'
#197060000000
1!
b101 %
1'
b101 +
#197070000000
0!
0'
#197080000000
1!
0$
b110 %
1'
0*
b110 +
#197090000000
0!
0'
#197100000000
1!
b111 %
1'
b111 +
#197110000000
0!
0'
#197120000000
1!
b1000 %
1'
b1000 +
#197130000000
0!
0'
#197140000000
1!
b1001 %
1'
b1001 +
#197150000000
1"
1(
#197160000000
0!
0"
b100 &
0'
0(
b100 ,
#197170000000
1!
b0 %
1'
b0 +
#197180000000
0!
0'
#197190000000
1!
1$
b1 %
1'
1*
b1 +
#197200000000
0!
0'
#197210000000
1!
b10 %
1'
b10 +
#197220000000
0!
0'
#197230000000
1!
b11 %
1'
b11 +
#197240000000
0!
0'
#197250000000
1!
b100 %
1'
b100 +
#197260000000
0!
0'
#197270000000
1!
b101 %
1'
b101 +
#197280000000
0!
0'
#197290000000
1!
b110 %
1'
b110 +
#197300000000
0!
0'
#197310000000
1!
b111 %
1'
b111 +
#197320000000
0!
0'
#197330000000
1!
0$
b1000 %
1'
0*
b1000 +
#197340000000
0!
0'
#197350000000
1!
b1001 %
1'
b1001 +
#197360000000
0!
0'
#197370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#197380000000
0!
0'
#197390000000
1!
1$
b1 %
1'
1*
b1 +
#197400000000
0!
0'
#197410000000
1!
b10 %
1'
b10 +
#197420000000
0!
0'
#197430000000
1!
b11 %
1'
b11 +
#197440000000
0!
0'
#197450000000
1!
b100 %
1'
b100 +
#197460000000
0!
0'
#197470000000
1!
b101 %
1'
b101 +
#197480000000
0!
0'
#197490000000
1!
0$
b110 %
1'
0*
b110 +
#197500000000
0!
0'
#197510000000
1!
b111 %
1'
b111 +
#197520000000
0!
0'
#197530000000
1!
b1000 %
1'
b1000 +
#197540000000
0!
0'
#197550000000
1!
b1001 %
1'
b1001 +
#197560000000
0!
0'
#197570000000
1!
b0 %
1'
b0 +
#197580000000
1"
1(
#197590000000
0!
0"
b100 &
0'
0(
b100 ,
#197600000000
1!
1$
b1 %
1'
1*
b1 +
#197610000000
0!
0'
#197620000000
1!
b10 %
1'
b10 +
#197630000000
0!
0'
#197640000000
1!
b11 %
1'
b11 +
#197650000000
0!
0'
#197660000000
1!
b100 %
1'
b100 +
#197670000000
0!
0'
#197680000000
1!
b101 %
1'
b101 +
#197690000000
0!
0'
#197700000000
1!
b110 %
1'
b110 +
#197710000000
0!
0'
#197720000000
1!
b111 %
1'
b111 +
#197730000000
0!
0'
#197740000000
1!
0$
b1000 %
1'
0*
b1000 +
#197750000000
0!
0'
#197760000000
1!
b1001 %
1'
b1001 +
#197770000000
0!
0'
#197780000000
1!
b0 %
1'
b0 +
#197790000000
0!
0'
#197800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#197810000000
0!
0'
#197820000000
1!
b10 %
1'
b10 +
#197830000000
0!
0'
#197840000000
1!
b11 %
1'
b11 +
#197850000000
0!
0'
#197860000000
1!
b100 %
1'
b100 +
#197870000000
0!
0'
#197880000000
1!
b101 %
1'
b101 +
#197890000000
0!
0'
#197900000000
1!
0$
b110 %
1'
0*
b110 +
#197910000000
0!
0'
#197920000000
1!
b111 %
1'
b111 +
#197930000000
0!
0'
#197940000000
1!
b1000 %
1'
b1000 +
#197950000000
0!
0'
#197960000000
1!
b1001 %
1'
b1001 +
#197970000000
0!
0'
#197980000000
1!
b0 %
1'
b0 +
#197990000000
0!
0'
#198000000000
1!
1$
b1 %
1'
1*
b1 +
#198010000000
1"
1(
#198020000000
0!
0"
b100 &
0'
0(
b100 ,
#198030000000
1!
b10 %
1'
b10 +
#198040000000
0!
0'
#198050000000
1!
b11 %
1'
b11 +
#198060000000
0!
0'
#198070000000
1!
b100 %
1'
b100 +
#198080000000
0!
0'
#198090000000
1!
b101 %
1'
b101 +
#198100000000
0!
0'
#198110000000
1!
b110 %
1'
b110 +
#198120000000
0!
0'
#198130000000
1!
b111 %
1'
b111 +
#198140000000
0!
0'
#198150000000
1!
0$
b1000 %
1'
0*
b1000 +
#198160000000
0!
0'
#198170000000
1!
b1001 %
1'
b1001 +
#198180000000
0!
0'
#198190000000
1!
b0 %
1'
b0 +
#198200000000
0!
0'
#198210000000
1!
1$
b1 %
1'
1*
b1 +
#198220000000
0!
0'
#198230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#198240000000
0!
0'
#198250000000
1!
b11 %
1'
b11 +
#198260000000
0!
0'
#198270000000
1!
b100 %
1'
b100 +
#198280000000
0!
0'
#198290000000
1!
b101 %
1'
b101 +
#198300000000
0!
0'
#198310000000
1!
0$
b110 %
1'
0*
b110 +
#198320000000
0!
0'
#198330000000
1!
b111 %
1'
b111 +
#198340000000
0!
0'
#198350000000
1!
b1000 %
1'
b1000 +
#198360000000
0!
0'
#198370000000
1!
b1001 %
1'
b1001 +
#198380000000
0!
0'
#198390000000
1!
b0 %
1'
b0 +
#198400000000
0!
0'
#198410000000
1!
1$
b1 %
1'
1*
b1 +
#198420000000
0!
0'
#198430000000
1!
b10 %
1'
b10 +
#198440000000
1"
1(
#198450000000
0!
0"
b100 &
0'
0(
b100 ,
#198460000000
1!
b11 %
1'
b11 +
#198470000000
0!
0'
#198480000000
1!
b100 %
1'
b100 +
#198490000000
0!
0'
#198500000000
1!
b101 %
1'
b101 +
#198510000000
0!
0'
#198520000000
1!
b110 %
1'
b110 +
#198530000000
0!
0'
#198540000000
1!
b111 %
1'
b111 +
#198550000000
0!
0'
#198560000000
1!
0$
b1000 %
1'
0*
b1000 +
#198570000000
0!
0'
#198580000000
1!
b1001 %
1'
b1001 +
#198590000000
0!
0'
#198600000000
1!
b0 %
1'
b0 +
#198610000000
0!
0'
#198620000000
1!
1$
b1 %
1'
1*
b1 +
#198630000000
0!
0'
#198640000000
1!
b10 %
1'
b10 +
#198650000000
0!
0'
#198660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#198670000000
0!
0'
#198680000000
1!
b100 %
1'
b100 +
#198690000000
0!
0'
#198700000000
1!
b101 %
1'
b101 +
#198710000000
0!
0'
#198720000000
1!
0$
b110 %
1'
0*
b110 +
#198730000000
0!
0'
#198740000000
1!
b111 %
1'
b111 +
#198750000000
0!
0'
#198760000000
1!
b1000 %
1'
b1000 +
#198770000000
0!
0'
#198780000000
1!
b1001 %
1'
b1001 +
#198790000000
0!
0'
#198800000000
1!
b0 %
1'
b0 +
#198810000000
0!
0'
#198820000000
1!
1$
b1 %
1'
1*
b1 +
#198830000000
0!
0'
#198840000000
1!
b10 %
1'
b10 +
#198850000000
0!
0'
#198860000000
1!
b11 %
1'
b11 +
#198870000000
1"
1(
#198880000000
0!
0"
b100 &
0'
0(
b100 ,
#198890000000
1!
b100 %
1'
b100 +
#198900000000
0!
0'
#198910000000
1!
b101 %
1'
b101 +
#198920000000
0!
0'
#198930000000
1!
b110 %
1'
b110 +
#198940000000
0!
0'
#198950000000
1!
b111 %
1'
b111 +
#198960000000
0!
0'
#198970000000
1!
0$
b1000 %
1'
0*
b1000 +
#198980000000
0!
0'
#198990000000
1!
b1001 %
1'
b1001 +
#199000000000
0!
0'
#199010000000
1!
b0 %
1'
b0 +
#199020000000
0!
0'
#199030000000
1!
1$
b1 %
1'
1*
b1 +
#199040000000
0!
0'
#199050000000
1!
b10 %
1'
b10 +
#199060000000
0!
0'
#199070000000
1!
b11 %
1'
b11 +
#199080000000
0!
0'
#199090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#199100000000
0!
0'
#199110000000
1!
b101 %
1'
b101 +
#199120000000
0!
0'
#199130000000
1!
0$
b110 %
1'
0*
b110 +
#199140000000
0!
0'
#199150000000
1!
b111 %
1'
b111 +
#199160000000
0!
0'
#199170000000
1!
b1000 %
1'
b1000 +
#199180000000
0!
0'
#199190000000
1!
b1001 %
1'
b1001 +
#199200000000
0!
0'
#199210000000
1!
b0 %
1'
b0 +
#199220000000
0!
0'
#199230000000
1!
1$
b1 %
1'
1*
b1 +
#199240000000
0!
0'
#199250000000
1!
b10 %
1'
b10 +
#199260000000
0!
0'
#199270000000
1!
b11 %
1'
b11 +
#199280000000
0!
0'
#199290000000
1!
b100 %
1'
b100 +
#199300000000
1"
1(
#199310000000
0!
0"
b100 &
0'
0(
b100 ,
#199320000000
1!
b101 %
1'
b101 +
#199330000000
0!
0'
#199340000000
1!
b110 %
1'
b110 +
#199350000000
0!
0'
#199360000000
1!
b111 %
1'
b111 +
#199370000000
0!
0'
#199380000000
1!
0$
b1000 %
1'
0*
b1000 +
#199390000000
0!
0'
#199400000000
1!
b1001 %
1'
b1001 +
#199410000000
0!
0'
#199420000000
1!
b0 %
1'
b0 +
#199430000000
0!
0'
#199440000000
1!
1$
b1 %
1'
1*
b1 +
#199450000000
0!
0'
#199460000000
1!
b10 %
1'
b10 +
#199470000000
0!
0'
#199480000000
1!
b11 %
1'
b11 +
#199490000000
0!
0'
#199500000000
1!
b100 %
1'
b100 +
#199510000000
0!
0'
#199520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#199530000000
0!
0'
#199540000000
1!
0$
b110 %
1'
0*
b110 +
#199550000000
0!
0'
#199560000000
1!
b111 %
1'
b111 +
#199570000000
0!
0'
#199580000000
1!
b1000 %
1'
b1000 +
#199590000000
0!
0'
#199600000000
1!
b1001 %
1'
b1001 +
#199610000000
0!
0'
#199620000000
1!
b0 %
1'
b0 +
#199630000000
0!
0'
#199640000000
1!
1$
b1 %
1'
1*
b1 +
#199650000000
0!
0'
#199660000000
1!
b10 %
1'
b10 +
#199670000000
0!
0'
#199680000000
1!
b11 %
1'
b11 +
#199690000000
0!
0'
#199700000000
1!
b100 %
1'
b100 +
#199710000000
0!
0'
#199720000000
1!
b101 %
1'
b101 +
#199730000000
1"
1(
#199740000000
0!
0"
b100 &
0'
0(
b100 ,
#199750000000
1!
b110 %
1'
b110 +
#199760000000
0!
0'
#199770000000
1!
b111 %
1'
b111 +
#199780000000
0!
0'
#199790000000
1!
0$
b1000 %
1'
0*
b1000 +
#199800000000
0!
0'
#199810000000
1!
b1001 %
1'
b1001 +
#199820000000
0!
0'
#199830000000
1!
b0 %
1'
b0 +
#199840000000
0!
0'
#199850000000
1!
1$
b1 %
1'
1*
b1 +
#199860000000
0!
0'
#199870000000
1!
b10 %
1'
b10 +
#199880000000
0!
0'
#199890000000
1!
b11 %
1'
b11 +
#199900000000
0!
0'
#199910000000
1!
b100 %
1'
b100 +
#199920000000
0!
0'
#199930000000
1!
b101 %
1'
b101 +
#199940000000
0!
0'
#199950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#199960000000
0!
0'
#199970000000
1!
b111 %
1'
b111 +
#199980000000
0!
0'
#199990000000
1!
b1000 %
1'
b1000 +
#200000000000
0!
0'
#200010000000
1!
b1001 %
1'
b1001 +
#200020000000
0!
0'
#200030000000
1!
b0 %
1'
b0 +
#200040000000
0!
0'
#200050000000
1!
1$
b1 %
1'
1*
b1 +
#200060000000
0!
0'
#200070000000
1!
b10 %
1'
b10 +
#200080000000
0!
0'
#200090000000
1!
b11 %
1'
b11 +
#200100000000
0!
0'
#200110000000
1!
b100 %
1'
b100 +
#200120000000
0!
0'
#200130000000
1!
b101 %
1'
b101 +
#200140000000
0!
0'
#200150000000
1!
0$
b110 %
1'
0*
b110 +
#200160000000
1"
1(
#200170000000
0!
0"
b100 &
0'
0(
b100 ,
#200180000000
1!
1$
b111 %
1'
1*
b111 +
#200190000000
0!
0'
#200200000000
1!
0$
b1000 %
1'
0*
b1000 +
#200210000000
0!
0'
#200220000000
1!
b1001 %
1'
b1001 +
#200230000000
0!
0'
#200240000000
1!
b0 %
1'
b0 +
#200250000000
0!
0'
#200260000000
1!
1$
b1 %
1'
1*
b1 +
#200270000000
0!
0'
#200280000000
1!
b10 %
1'
b10 +
#200290000000
0!
0'
#200300000000
1!
b11 %
1'
b11 +
#200310000000
0!
0'
#200320000000
1!
b100 %
1'
b100 +
#200330000000
0!
0'
#200340000000
1!
b101 %
1'
b101 +
#200350000000
0!
0'
#200360000000
1!
b110 %
1'
b110 +
#200370000000
0!
0'
#200380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#200390000000
0!
0'
#200400000000
1!
b1000 %
1'
b1000 +
#200410000000
0!
0'
#200420000000
1!
b1001 %
1'
b1001 +
#200430000000
0!
0'
#200440000000
1!
b0 %
1'
b0 +
#200450000000
0!
0'
#200460000000
1!
1$
b1 %
1'
1*
b1 +
#200470000000
0!
0'
#200480000000
1!
b10 %
1'
b10 +
#200490000000
0!
0'
#200500000000
1!
b11 %
1'
b11 +
#200510000000
0!
0'
#200520000000
1!
b100 %
1'
b100 +
#200530000000
0!
0'
#200540000000
1!
b101 %
1'
b101 +
#200550000000
0!
0'
#200560000000
1!
0$
b110 %
1'
0*
b110 +
#200570000000
0!
0'
#200580000000
1!
b111 %
1'
b111 +
#200590000000
1"
1(
#200600000000
0!
0"
b100 &
0'
0(
b100 ,
#200610000000
1!
b1000 %
1'
b1000 +
#200620000000
0!
0'
#200630000000
1!
b1001 %
1'
b1001 +
#200640000000
0!
0'
#200650000000
1!
b0 %
1'
b0 +
#200660000000
0!
0'
#200670000000
1!
1$
b1 %
1'
1*
b1 +
#200680000000
0!
0'
#200690000000
1!
b10 %
1'
b10 +
#200700000000
0!
0'
#200710000000
1!
b11 %
1'
b11 +
#200720000000
0!
0'
#200730000000
1!
b100 %
1'
b100 +
#200740000000
0!
0'
#200750000000
1!
b101 %
1'
b101 +
#200760000000
0!
0'
#200770000000
1!
b110 %
1'
b110 +
#200780000000
0!
0'
#200790000000
1!
b111 %
1'
b111 +
#200800000000
0!
0'
#200810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#200820000000
0!
0'
#200830000000
1!
b1001 %
1'
b1001 +
#200840000000
0!
0'
#200850000000
1!
b0 %
1'
b0 +
#200860000000
0!
0'
#200870000000
1!
1$
b1 %
1'
1*
b1 +
#200880000000
0!
0'
#200890000000
1!
b10 %
1'
b10 +
#200900000000
0!
0'
#200910000000
1!
b11 %
1'
b11 +
#200920000000
0!
0'
#200930000000
1!
b100 %
1'
b100 +
#200940000000
0!
0'
#200950000000
1!
b101 %
1'
b101 +
#200960000000
0!
0'
#200970000000
1!
0$
b110 %
1'
0*
b110 +
#200980000000
0!
0'
#200990000000
1!
b111 %
1'
b111 +
#201000000000
0!
0'
#201010000000
1!
b1000 %
1'
b1000 +
#201020000000
1"
1(
#201030000000
0!
0"
b100 &
0'
0(
b100 ,
#201040000000
1!
b1001 %
1'
b1001 +
#201050000000
0!
0'
#201060000000
1!
b0 %
1'
b0 +
#201070000000
0!
0'
#201080000000
1!
1$
b1 %
1'
1*
b1 +
#201090000000
0!
0'
#201100000000
1!
b10 %
1'
b10 +
#201110000000
0!
0'
#201120000000
1!
b11 %
1'
b11 +
#201130000000
0!
0'
#201140000000
1!
b100 %
1'
b100 +
#201150000000
0!
0'
#201160000000
1!
b101 %
1'
b101 +
#201170000000
0!
0'
#201180000000
1!
b110 %
1'
b110 +
#201190000000
0!
0'
#201200000000
1!
b111 %
1'
b111 +
#201210000000
0!
0'
#201220000000
1!
0$
b1000 %
1'
0*
b1000 +
#201230000000
0!
0'
#201240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#201250000000
0!
0'
#201260000000
1!
b0 %
1'
b0 +
#201270000000
0!
0'
#201280000000
1!
1$
b1 %
1'
1*
b1 +
#201290000000
0!
0'
#201300000000
1!
b10 %
1'
b10 +
#201310000000
0!
0'
#201320000000
1!
b11 %
1'
b11 +
#201330000000
0!
0'
#201340000000
1!
b100 %
1'
b100 +
#201350000000
0!
0'
#201360000000
1!
b101 %
1'
b101 +
#201370000000
0!
0'
#201380000000
1!
0$
b110 %
1'
0*
b110 +
#201390000000
0!
0'
#201400000000
1!
b111 %
1'
b111 +
#201410000000
0!
0'
#201420000000
1!
b1000 %
1'
b1000 +
#201430000000
0!
0'
#201440000000
1!
b1001 %
1'
b1001 +
#201450000000
1"
1(
#201460000000
0!
0"
b100 &
0'
0(
b100 ,
#201470000000
1!
b0 %
1'
b0 +
#201480000000
0!
0'
#201490000000
1!
1$
b1 %
1'
1*
b1 +
#201500000000
0!
0'
#201510000000
1!
b10 %
1'
b10 +
#201520000000
0!
0'
#201530000000
1!
b11 %
1'
b11 +
#201540000000
0!
0'
#201550000000
1!
b100 %
1'
b100 +
#201560000000
0!
0'
#201570000000
1!
b101 %
1'
b101 +
#201580000000
0!
0'
#201590000000
1!
b110 %
1'
b110 +
#201600000000
0!
0'
#201610000000
1!
b111 %
1'
b111 +
#201620000000
0!
0'
#201630000000
1!
0$
b1000 %
1'
0*
b1000 +
#201640000000
0!
0'
#201650000000
1!
b1001 %
1'
b1001 +
#201660000000
0!
0'
#201670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#201680000000
0!
0'
#201690000000
1!
1$
b1 %
1'
1*
b1 +
#201700000000
0!
0'
#201710000000
1!
b10 %
1'
b10 +
#201720000000
0!
0'
#201730000000
1!
b11 %
1'
b11 +
#201740000000
0!
0'
#201750000000
1!
b100 %
1'
b100 +
#201760000000
0!
0'
#201770000000
1!
b101 %
1'
b101 +
#201780000000
0!
0'
#201790000000
1!
0$
b110 %
1'
0*
b110 +
#201800000000
0!
0'
#201810000000
1!
b111 %
1'
b111 +
#201820000000
0!
0'
#201830000000
1!
b1000 %
1'
b1000 +
#201840000000
0!
0'
#201850000000
1!
b1001 %
1'
b1001 +
#201860000000
0!
0'
#201870000000
1!
b0 %
1'
b0 +
#201880000000
1"
1(
#201890000000
0!
0"
b100 &
0'
0(
b100 ,
#201900000000
1!
1$
b1 %
1'
1*
b1 +
#201910000000
0!
0'
#201920000000
1!
b10 %
1'
b10 +
#201930000000
0!
0'
#201940000000
1!
b11 %
1'
b11 +
#201950000000
0!
0'
#201960000000
1!
b100 %
1'
b100 +
#201970000000
0!
0'
#201980000000
1!
b101 %
1'
b101 +
#201990000000
0!
0'
#202000000000
1!
b110 %
1'
b110 +
#202010000000
0!
0'
#202020000000
1!
b111 %
1'
b111 +
#202030000000
0!
0'
#202040000000
1!
0$
b1000 %
1'
0*
b1000 +
#202050000000
0!
0'
#202060000000
1!
b1001 %
1'
b1001 +
#202070000000
0!
0'
#202080000000
1!
b0 %
1'
b0 +
#202090000000
0!
0'
#202100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#202110000000
0!
0'
#202120000000
1!
b10 %
1'
b10 +
#202130000000
0!
0'
#202140000000
1!
b11 %
1'
b11 +
#202150000000
0!
0'
#202160000000
1!
b100 %
1'
b100 +
#202170000000
0!
0'
#202180000000
1!
b101 %
1'
b101 +
#202190000000
0!
0'
#202200000000
1!
0$
b110 %
1'
0*
b110 +
#202210000000
0!
0'
#202220000000
1!
b111 %
1'
b111 +
#202230000000
0!
0'
#202240000000
1!
b1000 %
1'
b1000 +
#202250000000
0!
0'
#202260000000
1!
b1001 %
1'
b1001 +
#202270000000
0!
0'
#202280000000
1!
b0 %
1'
b0 +
#202290000000
0!
0'
#202300000000
1!
1$
b1 %
1'
1*
b1 +
#202310000000
1"
1(
#202320000000
0!
0"
b100 &
0'
0(
b100 ,
#202330000000
1!
b10 %
1'
b10 +
#202340000000
0!
0'
#202350000000
1!
b11 %
1'
b11 +
#202360000000
0!
0'
#202370000000
1!
b100 %
1'
b100 +
#202380000000
0!
0'
#202390000000
1!
b101 %
1'
b101 +
#202400000000
0!
0'
#202410000000
1!
b110 %
1'
b110 +
#202420000000
0!
0'
#202430000000
1!
b111 %
1'
b111 +
#202440000000
0!
0'
#202450000000
1!
0$
b1000 %
1'
0*
b1000 +
#202460000000
0!
0'
#202470000000
1!
b1001 %
1'
b1001 +
#202480000000
0!
0'
#202490000000
1!
b0 %
1'
b0 +
#202500000000
0!
0'
#202510000000
1!
1$
b1 %
1'
1*
b1 +
#202520000000
0!
0'
#202530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#202540000000
0!
0'
#202550000000
1!
b11 %
1'
b11 +
#202560000000
0!
0'
#202570000000
1!
b100 %
1'
b100 +
#202580000000
0!
0'
#202590000000
1!
b101 %
1'
b101 +
#202600000000
0!
0'
#202610000000
1!
0$
b110 %
1'
0*
b110 +
#202620000000
0!
0'
#202630000000
1!
b111 %
1'
b111 +
#202640000000
0!
0'
#202650000000
1!
b1000 %
1'
b1000 +
#202660000000
0!
0'
#202670000000
1!
b1001 %
1'
b1001 +
#202680000000
0!
0'
#202690000000
1!
b0 %
1'
b0 +
#202700000000
0!
0'
#202710000000
1!
1$
b1 %
1'
1*
b1 +
#202720000000
0!
0'
#202730000000
1!
b10 %
1'
b10 +
#202740000000
1"
1(
#202750000000
0!
0"
b100 &
0'
0(
b100 ,
#202760000000
1!
b11 %
1'
b11 +
#202770000000
0!
0'
#202780000000
1!
b100 %
1'
b100 +
#202790000000
0!
0'
#202800000000
1!
b101 %
1'
b101 +
#202810000000
0!
0'
#202820000000
1!
b110 %
1'
b110 +
#202830000000
0!
0'
#202840000000
1!
b111 %
1'
b111 +
#202850000000
0!
0'
#202860000000
1!
0$
b1000 %
1'
0*
b1000 +
#202870000000
0!
0'
#202880000000
1!
b1001 %
1'
b1001 +
#202890000000
0!
0'
#202900000000
1!
b0 %
1'
b0 +
#202910000000
0!
0'
#202920000000
1!
1$
b1 %
1'
1*
b1 +
#202930000000
0!
0'
#202940000000
1!
b10 %
1'
b10 +
#202950000000
0!
0'
#202960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#202970000000
0!
0'
#202980000000
1!
b100 %
1'
b100 +
#202990000000
0!
0'
#203000000000
1!
b101 %
1'
b101 +
#203010000000
0!
0'
#203020000000
1!
0$
b110 %
1'
0*
b110 +
#203030000000
0!
0'
#203040000000
1!
b111 %
1'
b111 +
#203050000000
0!
0'
#203060000000
1!
b1000 %
1'
b1000 +
#203070000000
0!
0'
#203080000000
1!
b1001 %
1'
b1001 +
#203090000000
0!
0'
#203100000000
1!
b0 %
1'
b0 +
#203110000000
0!
0'
#203120000000
1!
1$
b1 %
1'
1*
b1 +
#203130000000
0!
0'
#203140000000
1!
b10 %
1'
b10 +
#203150000000
0!
0'
#203160000000
1!
b11 %
1'
b11 +
#203170000000
1"
1(
#203180000000
0!
0"
b100 &
0'
0(
b100 ,
#203190000000
1!
b100 %
1'
b100 +
#203200000000
0!
0'
#203210000000
1!
b101 %
1'
b101 +
#203220000000
0!
0'
#203230000000
1!
b110 %
1'
b110 +
#203240000000
0!
0'
#203250000000
1!
b111 %
1'
b111 +
#203260000000
0!
0'
#203270000000
1!
0$
b1000 %
1'
0*
b1000 +
#203280000000
0!
0'
#203290000000
1!
b1001 %
1'
b1001 +
#203300000000
0!
0'
#203310000000
1!
b0 %
1'
b0 +
#203320000000
0!
0'
#203330000000
1!
1$
b1 %
1'
1*
b1 +
#203340000000
0!
0'
#203350000000
1!
b10 %
1'
b10 +
#203360000000
0!
0'
#203370000000
1!
b11 %
1'
b11 +
#203380000000
0!
0'
#203390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#203400000000
0!
0'
#203410000000
1!
b101 %
1'
b101 +
#203420000000
0!
0'
#203430000000
1!
0$
b110 %
1'
0*
b110 +
#203440000000
0!
0'
#203450000000
1!
b111 %
1'
b111 +
#203460000000
0!
0'
#203470000000
1!
b1000 %
1'
b1000 +
#203480000000
0!
0'
#203490000000
1!
b1001 %
1'
b1001 +
#203500000000
0!
0'
#203510000000
1!
b0 %
1'
b0 +
#203520000000
0!
0'
#203530000000
1!
1$
b1 %
1'
1*
b1 +
#203540000000
0!
0'
#203550000000
1!
b10 %
1'
b10 +
#203560000000
0!
0'
#203570000000
1!
b11 %
1'
b11 +
#203580000000
0!
0'
#203590000000
1!
b100 %
1'
b100 +
#203600000000
1"
1(
#203610000000
0!
0"
b100 &
0'
0(
b100 ,
#203620000000
1!
b101 %
1'
b101 +
#203630000000
0!
0'
#203640000000
1!
b110 %
1'
b110 +
#203650000000
0!
0'
#203660000000
1!
b111 %
1'
b111 +
#203670000000
0!
0'
#203680000000
1!
0$
b1000 %
1'
0*
b1000 +
#203690000000
0!
0'
#203700000000
1!
b1001 %
1'
b1001 +
#203710000000
0!
0'
#203720000000
1!
b0 %
1'
b0 +
#203730000000
0!
0'
#203740000000
1!
1$
b1 %
1'
1*
b1 +
#203750000000
0!
0'
#203760000000
1!
b10 %
1'
b10 +
#203770000000
0!
0'
#203780000000
1!
b11 %
1'
b11 +
#203790000000
0!
0'
#203800000000
1!
b100 %
1'
b100 +
#203810000000
0!
0'
#203820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#203830000000
0!
0'
#203840000000
1!
0$
b110 %
1'
0*
b110 +
#203850000000
0!
0'
#203860000000
1!
b111 %
1'
b111 +
#203870000000
0!
0'
#203880000000
1!
b1000 %
1'
b1000 +
#203890000000
0!
0'
#203900000000
1!
b1001 %
1'
b1001 +
#203910000000
0!
0'
#203920000000
1!
b0 %
1'
b0 +
#203930000000
0!
0'
#203940000000
1!
1$
b1 %
1'
1*
b1 +
#203950000000
0!
0'
#203960000000
1!
b10 %
1'
b10 +
#203970000000
0!
0'
#203980000000
1!
b11 %
1'
b11 +
#203990000000
0!
0'
#204000000000
1!
b100 %
1'
b100 +
#204010000000
0!
0'
#204020000000
1!
b101 %
1'
b101 +
#204030000000
1"
1(
#204040000000
0!
0"
b100 &
0'
0(
b100 ,
#204050000000
1!
b110 %
1'
b110 +
#204060000000
0!
0'
#204070000000
1!
b111 %
1'
b111 +
#204080000000
0!
0'
#204090000000
1!
0$
b1000 %
1'
0*
b1000 +
#204100000000
0!
0'
#204110000000
1!
b1001 %
1'
b1001 +
#204120000000
0!
0'
#204130000000
1!
b0 %
1'
b0 +
#204140000000
0!
0'
#204150000000
1!
1$
b1 %
1'
1*
b1 +
#204160000000
0!
0'
#204170000000
1!
b10 %
1'
b10 +
#204180000000
0!
0'
#204190000000
1!
b11 %
1'
b11 +
#204200000000
0!
0'
#204210000000
1!
b100 %
1'
b100 +
#204220000000
0!
0'
#204230000000
1!
b101 %
1'
b101 +
#204240000000
0!
0'
#204250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#204260000000
0!
0'
#204270000000
1!
b111 %
1'
b111 +
#204280000000
0!
0'
#204290000000
1!
b1000 %
1'
b1000 +
#204300000000
0!
0'
#204310000000
1!
b1001 %
1'
b1001 +
#204320000000
0!
0'
#204330000000
1!
b0 %
1'
b0 +
#204340000000
0!
0'
#204350000000
1!
1$
b1 %
1'
1*
b1 +
#204360000000
0!
0'
#204370000000
1!
b10 %
1'
b10 +
#204380000000
0!
0'
#204390000000
1!
b11 %
1'
b11 +
#204400000000
0!
0'
#204410000000
1!
b100 %
1'
b100 +
#204420000000
0!
0'
#204430000000
1!
b101 %
1'
b101 +
#204440000000
0!
0'
#204450000000
1!
0$
b110 %
1'
0*
b110 +
#204460000000
1"
1(
#204470000000
0!
0"
b100 &
0'
0(
b100 ,
#204480000000
1!
1$
b111 %
1'
1*
b111 +
#204490000000
0!
0'
#204500000000
1!
0$
b1000 %
1'
0*
b1000 +
#204510000000
0!
0'
#204520000000
1!
b1001 %
1'
b1001 +
#204530000000
0!
0'
#204540000000
1!
b0 %
1'
b0 +
#204550000000
0!
0'
#204560000000
1!
1$
b1 %
1'
1*
b1 +
#204570000000
0!
0'
#204580000000
1!
b10 %
1'
b10 +
#204590000000
0!
0'
#204600000000
1!
b11 %
1'
b11 +
#204610000000
0!
0'
#204620000000
1!
b100 %
1'
b100 +
#204630000000
0!
0'
#204640000000
1!
b101 %
1'
b101 +
#204650000000
0!
0'
#204660000000
1!
b110 %
1'
b110 +
#204670000000
0!
0'
#204680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#204690000000
0!
0'
#204700000000
1!
b1000 %
1'
b1000 +
#204710000000
0!
0'
#204720000000
1!
b1001 %
1'
b1001 +
#204730000000
0!
0'
#204740000000
1!
b0 %
1'
b0 +
#204750000000
0!
0'
#204760000000
1!
1$
b1 %
1'
1*
b1 +
#204770000000
0!
0'
#204780000000
1!
b10 %
1'
b10 +
#204790000000
0!
0'
#204800000000
1!
b11 %
1'
b11 +
#204810000000
0!
0'
#204820000000
1!
b100 %
1'
b100 +
#204830000000
0!
0'
#204840000000
1!
b101 %
1'
b101 +
#204850000000
0!
0'
#204860000000
1!
0$
b110 %
1'
0*
b110 +
#204870000000
0!
0'
#204880000000
1!
b111 %
1'
b111 +
#204890000000
1"
1(
#204900000000
0!
0"
b100 &
0'
0(
b100 ,
#204910000000
1!
b1000 %
1'
b1000 +
#204920000000
0!
0'
#204930000000
1!
b1001 %
1'
b1001 +
#204940000000
0!
0'
#204950000000
1!
b0 %
1'
b0 +
#204960000000
0!
0'
#204970000000
1!
1$
b1 %
1'
1*
b1 +
#204980000000
0!
0'
#204990000000
1!
b10 %
1'
b10 +
#205000000000
0!
0'
#205010000000
1!
b11 %
1'
b11 +
#205020000000
0!
0'
#205030000000
1!
b100 %
1'
b100 +
#205040000000
0!
0'
#205050000000
1!
b101 %
1'
b101 +
#205060000000
0!
0'
#205070000000
1!
b110 %
1'
b110 +
#205080000000
0!
0'
#205090000000
1!
b111 %
1'
b111 +
#205100000000
0!
0'
#205110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#205120000000
0!
0'
#205130000000
1!
b1001 %
1'
b1001 +
#205140000000
0!
0'
#205150000000
1!
b0 %
1'
b0 +
#205160000000
0!
0'
#205170000000
1!
1$
b1 %
1'
1*
b1 +
#205180000000
0!
0'
#205190000000
1!
b10 %
1'
b10 +
#205200000000
0!
0'
#205210000000
1!
b11 %
1'
b11 +
#205220000000
0!
0'
#205230000000
1!
b100 %
1'
b100 +
#205240000000
0!
0'
#205250000000
1!
b101 %
1'
b101 +
#205260000000
0!
0'
#205270000000
1!
0$
b110 %
1'
0*
b110 +
#205280000000
0!
0'
#205290000000
1!
b111 %
1'
b111 +
#205300000000
0!
0'
#205310000000
1!
b1000 %
1'
b1000 +
#205320000000
1"
1(
#205330000000
0!
0"
b100 &
0'
0(
b100 ,
#205340000000
1!
b1001 %
1'
b1001 +
#205350000000
0!
0'
#205360000000
1!
b0 %
1'
b0 +
#205370000000
0!
0'
#205380000000
1!
1$
b1 %
1'
1*
b1 +
#205390000000
0!
0'
#205400000000
1!
b10 %
1'
b10 +
#205410000000
0!
0'
#205420000000
1!
b11 %
1'
b11 +
#205430000000
0!
0'
#205440000000
1!
b100 %
1'
b100 +
#205450000000
0!
0'
#205460000000
1!
b101 %
1'
b101 +
#205470000000
0!
0'
#205480000000
1!
b110 %
1'
b110 +
#205490000000
0!
0'
#205500000000
1!
b111 %
1'
b111 +
#205510000000
0!
0'
#205520000000
1!
0$
b1000 %
1'
0*
b1000 +
#205530000000
0!
0'
#205540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#205550000000
0!
0'
#205560000000
1!
b0 %
1'
b0 +
#205570000000
0!
0'
#205580000000
1!
1$
b1 %
1'
1*
b1 +
#205590000000
0!
0'
#205600000000
1!
b10 %
1'
b10 +
#205610000000
0!
0'
#205620000000
1!
b11 %
1'
b11 +
#205630000000
0!
0'
#205640000000
1!
b100 %
1'
b100 +
#205650000000
0!
0'
#205660000000
1!
b101 %
1'
b101 +
#205670000000
0!
0'
#205680000000
1!
0$
b110 %
1'
0*
b110 +
#205690000000
0!
0'
#205700000000
1!
b111 %
1'
b111 +
#205710000000
0!
0'
#205720000000
1!
b1000 %
1'
b1000 +
#205730000000
0!
0'
#205740000000
1!
b1001 %
1'
b1001 +
#205750000000
1"
1(
#205760000000
0!
0"
b100 &
0'
0(
b100 ,
#205770000000
1!
b0 %
1'
b0 +
#205780000000
0!
0'
#205790000000
1!
1$
b1 %
1'
1*
b1 +
#205800000000
0!
0'
#205810000000
1!
b10 %
1'
b10 +
#205820000000
0!
0'
#205830000000
1!
b11 %
1'
b11 +
#205840000000
0!
0'
#205850000000
1!
b100 %
1'
b100 +
#205860000000
0!
0'
#205870000000
1!
b101 %
1'
b101 +
#205880000000
0!
0'
#205890000000
1!
b110 %
1'
b110 +
#205900000000
0!
0'
#205910000000
1!
b111 %
1'
b111 +
#205920000000
0!
0'
#205930000000
1!
0$
b1000 %
1'
0*
b1000 +
#205940000000
0!
0'
#205950000000
1!
b1001 %
1'
b1001 +
#205960000000
0!
0'
#205970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#205980000000
0!
0'
#205990000000
1!
1$
b1 %
1'
1*
b1 +
#206000000000
0!
0'
#206010000000
1!
b10 %
1'
b10 +
#206020000000
0!
0'
#206030000000
1!
b11 %
1'
b11 +
#206040000000
0!
0'
#206050000000
1!
b100 %
1'
b100 +
#206060000000
0!
0'
#206070000000
1!
b101 %
1'
b101 +
#206080000000
0!
0'
#206090000000
1!
0$
b110 %
1'
0*
b110 +
#206100000000
0!
0'
#206110000000
1!
b111 %
1'
b111 +
#206120000000
0!
0'
#206130000000
1!
b1000 %
1'
b1000 +
#206140000000
0!
0'
#206150000000
1!
b1001 %
1'
b1001 +
#206160000000
0!
0'
#206170000000
1!
b0 %
1'
b0 +
#206180000000
1"
1(
#206190000000
0!
0"
b100 &
0'
0(
b100 ,
#206200000000
1!
1$
b1 %
1'
1*
b1 +
#206210000000
0!
0'
#206220000000
1!
b10 %
1'
b10 +
#206230000000
0!
0'
#206240000000
1!
b11 %
1'
b11 +
#206250000000
0!
0'
#206260000000
1!
b100 %
1'
b100 +
#206270000000
0!
0'
#206280000000
1!
b101 %
1'
b101 +
#206290000000
0!
0'
#206300000000
1!
b110 %
1'
b110 +
#206310000000
0!
0'
#206320000000
1!
b111 %
1'
b111 +
#206330000000
0!
0'
#206340000000
1!
0$
b1000 %
1'
0*
b1000 +
#206350000000
0!
0'
#206360000000
1!
b1001 %
1'
b1001 +
#206370000000
0!
0'
#206380000000
1!
b0 %
1'
b0 +
#206390000000
0!
0'
#206400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#206410000000
0!
0'
#206420000000
1!
b10 %
1'
b10 +
#206430000000
0!
0'
#206440000000
1!
b11 %
1'
b11 +
#206450000000
0!
0'
#206460000000
1!
b100 %
1'
b100 +
#206470000000
0!
0'
#206480000000
1!
b101 %
1'
b101 +
#206490000000
0!
0'
#206500000000
1!
0$
b110 %
1'
0*
b110 +
#206510000000
0!
0'
#206520000000
1!
b111 %
1'
b111 +
#206530000000
0!
0'
#206540000000
1!
b1000 %
1'
b1000 +
#206550000000
0!
0'
#206560000000
1!
b1001 %
1'
b1001 +
#206570000000
0!
0'
#206580000000
1!
b0 %
1'
b0 +
#206590000000
0!
0'
#206600000000
1!
1$
b1 %
1'
1*
b1 +
#206610000000
1"
1(
#206620000000
0!
0"
b100 &
0'
0(
b100 ,
#206630000000
1!
b10 %
1'
b10 +
#206640000000
0!
0'
#206650000000
1!
b11 %
1'
b11 +
#206660000000
0!
0'
#206670000000
1!
b100 %
1'
b100 +
#206680000000
0!
0'
#206690000000
1!
b101 %
1'
b101 +
#206700000000
0!
0'
#206710000000
1!
b110 %
1'
b110 +
#206720000000
0!
0'
#206730000000
1!
b111 %
1'
b111 +
#206740000000
0!
0'
#206750000000
1!
0$
b1000 %
1'
0*
b1000 +
#206760000000
0!
0'
#206770000000
1!
b1001 %
1'
b1001 +
#206780000000
0!
0'
#206790000000
1!
b0 %
1'
b0 +
#206800000000
0!
0'
#206810000000
1!
1$
b1 %
1'
1*
b1 +
#206820000000
0!
0'
#206830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#206840000000
0!
0'
#206850000000
1!
b11 %
1'
b11 +
#206860000000
0!
0'
#206870000000
1!
b100 %
1'
b100 +
#206880000000
0!
0'
#206890000000
1!
b101 %
1'
b101 +
#206900000000
0!
0'
#206910000000
1!
0$
b110 %
1'
0*
b110 +
#206920000000
0!
0'
#206930000000
1!
b111 %
1'
b111 +
#206940000000
0!
0'
#206950000000
1!
b1000 %
1'
b1000 +
#206960000000
0!
0'
#206970000000
1!
b1001 %
1'
b1001 +
#206980000000
0!
0'
#206990000000
1!
b0 %
1'
b0 +
#207000000000
0!
0'
#207010000000
1!
1$
b1 %
1'
1*
b1 +
#207020000000
0!
0'
#207030000000
1!
b10 %
1'
b10 +
#207040000000
1"
1(
#207050000000
0!
0"
b100 &
0'
0(
b100 ,
#207060000000
1!
b11 %
1'
b11 +
#207070000000
0!
0'
#207080000000
1!
b100 %
1'
b100 +
#207090000000
0!
0'
#207100000000
1!
b101 %
1'
b101 +
#207110000000
0!
0'
#207120000000
1!
b110 %
1'
b110 +
#207130000000
0!
0'
#207140000000
1!
b111 %
1'
b111 +
#207150000000
0!
0'
#207160000000
1!
0$
b1000 %
1'
0*
b1000 +
#207170000000
0!
0'
#207180000000
1!
b1001 %
1'
b1001 +
#207190000000
0!
0'
#207200000000
1!
b0 %
1'
b0 +
#207210000000
0!
0'
#207220000000
1!
1$
b1 %
1'
1*
b1 +
#207230000000
0!
0'
#207240000000
1!
b10 %
1'
b10 +
#207250000000
0!
0'
#207260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#207270000000
0!
0'
#207280000000
1!
b100 %
1'
b100 +
#207290000000
0!
0'
#207300000000
1!
b101 %
1'
b101 +
#207310000000
0!
0'
#207320000000
1!
0$
b110 %
1'
0*
b110 +
#207330000000
0!
0'
#207340000000
1!
b111 %
1'
b111 +
#207350000000
0!
0'
#207360000000
1!
b1000 %
1'
b1000 +
#207370000000
0!
0'
#207380000000
1!
b1001 %
1'
b1001 +
#207390000000
0!
0'
#207400000000
1!
b0 %
1'
b0 +
#207410000000
0!
0'
#207420000000
1!
1$
b1 %
1'
1*
b1 +
#207430000000
0!
0'
#207440000000
1!
b10 %
1'
b10 +
#207450000000
0!
0'
#207460000000
1!
b11 %
1'
b11 +
#207470000000
1"
1(
#207480000000
0!
0"
b100 &
0'
0(
b100 ,
#207490000000
1!
b100 %
1'
b100 +
#207500000000
0!
0'
#207510000000
1!
b101 %
1'
b101 +
#207520000000
0!
0'
#207530000000
1!
b110 %
1'
b110 +
#207540000000
0!
0'
#207550000000
1!
b111 %
1'
b111 +
#207560000000
0!
0'
#207570000000
1!
0$
b1000 %
1'
0*
b1000 +
#207580000000
0!
0'
#207590000000
1!
b1001 %
1'
b1001 +
#207600000000
0!
0'
#207610000000
1!
b0 %
1'
b0 +
#207620000000
0!
0'
#207630000000
1!
1$
b1 %
1'
1*
b1 +
#207640000000
0!
0'
#207650000000
1!
b10 %
1'
b10 +
#207660000000
0!
0'
#207670000000
1!
b11 %
1'
b11 +
#207680000000
0!
0'
#207690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#207700000000
0!
0'
#207710000000
1!
b101 %
1'
b101 +
#207720000000
0!
0'
#207730000000
1!
0$
b110 %
1'
0*
b110 +
#207740000000
0!
0'
#207750000000
1!
b111 %
1'
b111 +
#207760000000
0!
0'
#207770000000
1!
b1000 %
1'
b1000 +
#207780000000
0!
0'
#207790000000
1!
b1001 %
1'
b1001 +
#207800000000
0!
0'
#207810000000
1!
b0 %
1'
b0 +
#207820000000
0!
0'
#207830000000
1!
1$
b1 %
1'
1*
b1 +
#207840000000
0!
0'
#207850000000
1!
b10 %
1'
b10 +
#207860000000
0!
0'
#207870000000
1!
b11 %
1'
b11 +
#207880000000
0!
0'
#207890000000
1!
b100 %
1'
b100 +
#207900000000
1"
1(
#207910000000
0!
0"
b100 &
0'
0(
b100 ,
#207920000000
1!
b101 %
1'
b101 +
#207930000000
0!
0'
#207940000000
1!
b110 %
1'
b110 +
#207950000000
0!
0'
#207960000000
1!
b111 %
1'
b111 +
#207970000000
0!
0'
#207980000000
1!
0$
b1000 %
1'
0*
b1000 +
#207990000000
0!
0'
#208000000000
1!
b1001 %
1'
b1001 +
#208010000000
0!
0'
#208020000000
1!
b0 %
1'
b0 +
#208030000000
0!
0'
#208040000000
1!
1$
b1 %
1'
1*
b1 +
#208050000000
0!
0'
#208060000000
1!
b10 %
1'
b10 +
#208070000000
0!
0'
#208080000000
1!
b11 %
1'
b11 +
#208090000000
0!
0'
#208100000000
1!
b100 %
1'
b100 +
#208110000000
0!
0'
#208120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#208130000000
0!
0'
#208140000000
1!
0$
b110 %
1'
0*
b110 +
#208150000000
0!
0'
#208160000000
1!
b111 %
1'
b111 +
#208170000000
0!
0'
#208180000000
1!
b1000 %
1'
b1000 +
#208190000000
0!
0'
#208200000000
1!
b1001 %
1'
b1001 +
#208210000000
0!
0'
#208220000000
1!
b0 %
1'
b0 +
#208230000000
0!
0'
#208240000000
1!
1$
b1 %
1'
1*
b1 +
#208250000000
0!
0'
#208260000000
1!
b10 %
1'
b10 +
#208270000000
0!
0'
#208280000000
1!
b11 %
1'
b11 +
#208290000000
0!
0'
#208300000000
1!
b100 %
1'
b100 +
#208310000000
0!
0'
#208320000000
1!
b101 %
1'
b101 +
#208330000000
1"
1(
#208340000000
0!
0"
b100 &
0'
0(
b100 ,
#208350000000
1!
b110 %
1'
b110 +
#208360000000
0!
0'
#208370000000
1!
b111 %
1'
b111 +
#208380000000
0!
0'
#208390000000
1!
0$
b1000 %
1'
0*
b1000 +
#208400000000
0!
0'
#208410000000
1!
b1001 %
1'
b1001 +
#208420000000
0!
0'
#208430000000
1!
b0 %
1'
b0 +
#208440000000
0!
0'
#208450000000
1!
1$
b1 %
1'
1*
b1 +
#208460000000
0!
0'
#208470000000
1!
b10 %
1'
b10 +
#208480000000
0!
0'
#208490000000
1!
b11 %
1'
b11 +
#208500000000
0!
0'
#208510000000
1!
b100 %
1'
b100 +
#208520000000
0!
0'
#208530000000
1!
b101 %
1'
b101 +
#208540000000
0!
0'
#208550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#208560000000
0!
0'
#208570000000
1!
b111 %
1'
b111 +
#208580000000
0!
0'
#208590000000
1!
b1000 %
1'
b1000 +
#208600000000
0!
0'
#208610000000
1!
b1001 %
1'
b1001 +
#208620000000
0!
0'
#208630000000
1!
b0 %
1'
b0 +
#208640000000
0!
0'
#208650000000
1!
1$
b1 %
1'
1*
b1 +
#208660000000
0!
0'
#208670000000
1!
b10 %
1'
b10 +
#208680000000
0!
0'
#208690000000
1!
b11 %
1'
b11 +
#208700000000
0!
0'
#208710000000
1!
b100 %
1'
b100 +
#208720000000
0!
0'
#208730000000
1!
b101 %
1'
b101 +
#208740000000
0!
0'
#208750000000
1!
0$
b110 %
1'
0*
b110 +
#208760000000
1"
1(
#208770000000
0!
0"
b100 &
0'
0(
b100 ,
#208780000000
1!
1$
b111 %
1'
1*
b111 +
#208790000000
0!
0'
#208800000000
1!
0$
b1000 %
1'
0*
b1000 +
#208810000000
0!
0'
#208820000000
1!
b1001 %
1'
b1001 +
#208830000000
0!
0'
#208840000000
1!
b0 %
1'
b0 +
#208850000000
0!
0'
#208860000000
1!
1$
b1 %
1'
1*
b1 +
#208870000000
0!
0'
#208880000000
1!
b10 %
1'
b10 +
#208890000000
0!
0'
#208900000000
1!
b11 %
1'
b11 +
#208910000000
0!
0'
#208920000000
1!
b100 %
1'
b100 +
#208930000000
0!
0'
#208940000000
1!
b101 %
1'
b101 +
#208950000000
0!
0'
#208960000000
1!
b110 %
1'
b110 +
#208970000000
0!
0'
#208980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#208990000000
0!
0'
#209000000000
1!
b1000 %
1'
b1000 +
#209010000000
0!
0'
#209020000000
1!
b1001 %
1'
b1001 +
#209030000000
0!
0'
#209040000000
1!
b0 %
1'
b0 +
#209050000000
0!
0'
#209060000000
1!
1$
b1 %
1'
1*
b1 +
#209070000000
0!
0'
#209080000000
1!
b10 %
1'
b10 +
#209090000000
0!
0'
#209100000000
1!
b11 %
1'
b11 +
#209110000000
0!
0'
#209120000000
1!
b100 %
1'
b100 +
#209130000000
0!
0'
#209140000000
1!
b101 %
1'
b101 +
#209150000000
0!
0'
#209160000000
1!
0$
b110 %
1'
0*
b110 +
#209170000000
0!
0'
#209180000000
1!
b111 %
1'
b111 +
#209190000000
1"
1(
#209200000000
0!
0"
b100 &
0'
0(
b100 ,
#209210000000
1!
b1000 %
1'
b1000 +
#209220000000
0!
0'
#209230000000
1!
b1001 %
1'
b1001 +
#209240000000
0!
0'
#209250000000
1!
b0 %
1'
b0 +
#209260000000
0!
0'
#209270000000
1!
1$
b1 %
1'
1*
b1 +
#209280000000
0!
0'
#209290000000
1!
b10 %
1'
b10 +
#209300000000
0!
0'
#209310000000
1!
b11 %
1'
b11 +
#209320000000
0!
0'
#209330000000
1!
b100 %
1'
b100 +
#209340000000
0!
0'
#209350000000
1!
b101 %
1'
b101 +
#209360000000
0!
0'
#209370000000
1!
b110 %
1'
b110 +
#209380000000
0!
0'
#209390000000
1!
b111 %
1'
b111 +
#209400000000
0!
0'
#209410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#209420000000
0!
0'
#209430000000
1!
b1001 %
1'
b1001 +
#209440000000
0!
0'
#209450000000
1!
b0 %
1'
b0 +
#209460000000
0!
0'
#209470000000
1!
1$
b1 %
1'
1*
b1 +
#209480000000
0!
0'
#209490000000
1!
b10 %
1'
b10 +
#209500000000
0!
0'
#209510000000
1!
b11 %
1'
b11 +
#209520000000
0!
0'
#209530000000
1!
b100 %
1'
b100 +
#209540000000
0!
0'
#209550000000
1!
b101 %
1'
b101 +
#209560000000
0!
0'
#209570000000
1!
0$
b110 %
1'
0*
b110 +
#209580000000
0!
0'
#209590000000
1!
b111 %
1'
b111 +
#209600000000
0!
0'
#209610000000
1!
b1000 %
1'
b1000 +
#209620000000
1"
1(
#209630000000
0!
0"
b100 &
0'
0(
b100 ,
#209640000000
1!
b1001 %
1'
b1001 +
#209650000000
0!
0'
#209660000000
1!
b0 %
1'
b0 +
#209670000000
0!
0'
#209680000000
1!
1$
b1 %
1'
1*
b1 +
#209690000000
0!
0'
#209700000000
1!
b10 %
1'
b10 +
#209710000000
0!
0'
#209720000000
1!
b11 %
1'
b11 +
#209730000000
0!
0'
#209740000000
1!
b100 %
1'
b100 +
#209750000000
0!
0'
#209760000000
1!
b101 %
1'
b101 +
#209770000000
0!
0'
#209780000000
1!
b110 %
1'
b110 +
#209790000000
0!
0'
#209800000000
1!
b111 %
1'
b111 +
#209810000000
0!
0'
#209820000000
1!
0$
b1000 %
1'
0*
b1000 +
#209830000000
0!
0'
#209840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#209850000000
0!
0'
#209860000000
1!
b0 %
1'
b0 +
#209870000000
0!
0'
#209880000000
1!
1$
b1 %
1'
1*
b1 +
#209890000000
0!
0'
#209900000000
1!
b10 %
1'
b10 +
#209910000000
0!
0'
#209920000000
1!
b11 %
1'
b11 +
#209930000000
0!
0'
#209940000000
1!
b100 %
1'
b100 +
#209950000000
0!
0'
#209960000000
1!
b101 %
1'
b101 +
#209970000000
0!
0'
#209980000000
1!
0$
b110 %
1'
0*
b110 +
#209990000000
0!
0'
#210000000000
1!
b111 %
1'
b111 +
#210010000000
0!
0'
#210020000000
1!
b1000 %
1'
b1000 +
#210030000000
0!
0'
#210040000000
1!
b1001 %
1'
b1001 +
#210050000000
1"
1(
#210060000000
0!
0"
b100 &
0'
0(
b100 ,
#210070000000
1!
b0 %
1'
b0 +
#210080000000
0!
0'
#210090000000
1!
1$
b1 %
1'
1*
b1 +
#210100000000
0!
0'
#210110000000
1!
b10 %
1'
b10 +
#210120000000
0!
0'
#210130000000
1!
b11 %
1'
b11 +
#210140000000
0!
0'
#210150000000
1!
b100 %
1'
b100 +
#210160000000
0!
0'
#210170000000
1!
b101 %
1'
b101 +
#210180000000
0!
0'
#210190000000
1!
b110 %
1'
b110 +
#210200000000
0!
0'
#210210000000
1!
b111 %
1'
b111 +
#210220000000
0!
0'
#210230000000
1!
0$
b1000 %
1'
0*
b1000 +
#210240000000
0!
0'
#210250000000
1!
b1001 %
1'
b1001 +
#210260000000
0!
0'
#210270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#210280000000
0!
0'
#210290000000
1!
1$
b1 %
1'
1*
b1 +
#210300000000
0!
0'
#210310000000
1!
b10 %
1'
b10 +
#210320000000
0!
0'
#210330000000
1!
b11 %
1'
b11 +
#210340000000
0!
0'
#210350000000
1!
b100 %
1'
b100 +
#210360000000
0!
0'
#210370000000
1!
b101 %
1'
b101 +
#210380000000
0!
0'
#210390000000
1!
0$
b110 %
1'
0*
b110 +
#210400000000
0!
0'
#210410000000
1!
b111 %
1'
b111 +
#210420000000
0!
0'
#210430000000
1!
b1000 %
1'
b1000 +
#210440000000
0!
0'
#210450000000
1!
b1001 %
1'
b1001 +
#210460000000
0!
0'
#210470000000
1!
b0 %
1'
b0 +
#210480000000
1"
1(
#210490000000
0!
0"
b100 &
0'
0(
b100 ,
#210500000000
1!
1$
b1 %
1'
1*
b1 +
#210510000000
0!
0'
#210520000000
1!
b10 %
1'
b10 +
#210530000000
0!
0'
#210540000000
1!
b11 %
1'
b11 +
#210550000000
0!
0'
#210560000000
1!
b100 %
1'
b100 +
#210570000000
0!
0'
#210580000000
1!
b101 %
1'
b101 +
#210590000000
0!
0'
#210600000000
1!
b110 %
1'
b110 +
#210610000000
0!
0'
#210620000000
1!
b111 %
1'
b111 +
#210630000000
0!
0'
#210640000000
1!
0$
b1000 %
1'
0*
b1000 +
#210650000000
0!
0'
#210660000000
1!
b1001 %
1'
b1001 +
#210670000000
0!
0'
#210680000000
1!
b0 %
1'
b0 +
#210690000000
0!
0'
#210700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#210710000000
0!
0'
#210720000000
1!
b10 %
1'
b10 +
#210730000000
0!
0'
#210740000000
1!
b11 %
1'
b11 +
#210750000000
0!
0'
#210760000000
1!
b100 %
1'
b100 +
#210770000000
0!
0'
#210780000000
1!
b101 %
1'
b101 +
#210790000000
0!
0'
#210800000000
1!
0$
b110 %
1'
0*
b110 +
#210810000000
0!
0'
#210820000000
1!
b111 %
1'
b111 +
#210830000000
0!
0'
#210840000000
1!
b1000 %
1'
b1000 +
#210850000000
0!
0'
#210860000000
1!
b1001 %
1'
b1001 +
#210870000000
0!
0'
#210880000000
1!
b0 %
1'
b0 +
#210890000000
0!
0'
#210900000000
1!
1$
b1 %
1'
1*
b1 +
#210910000000
1"
1(
#210920000000
0!
0"
b100 &
0'
0(
b100 ,
#210930000000
1!
b10 %
1'
b10 +
#210940000000
0!
0'
#210950000000
1!
b11 %
1'
b11 +
#210960000000
0!
0'
#210970000000
1!
b100 %
1'
b100 +
#210980000000
0!
0'
#210990000000
1!
b101 %
1'
b101 +
#211000000000
0!
0'
#211010000000
1!
b110 %
1'
b110 +
#211020000000
0!
0'
#211030000000
1!
b111 %
1'
b111 +
#211040000000
0!
0'
#211050000000
1!
0$
b1000 %
1'
0*
b1000 +
#211060000000
0!
0'
#211070000000
1!
b1001 %
1'
b1001 +
#211080000000
0!
0'
#211090000000
1!
b0 %
1'
b0 +
#211100000000
0!
0'
#211110000000
1!
1$
b1 %
1'
1*
b1 +
#211120000000
0!
0'
#211130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#211140000000
0!
0'
#211150000000
1!
b11 %
1'
b11 +
#211160000000
0!
0'
#211170000000
1!
b100 %
1'
b100 +
#211180000000
0!
0'
#211190000000
1!
b101 %
1'
b101 +
#211200000000
0!
0'
#211210000000
1!
0$
b110 %
1'
0*
b110 +
#211220000000
0!
0'
#211230000000
1!
b111 %
1'
b111 +
#211240000000
0!
0'
#211250000000
1!
b1000 %
1'
b1000 +
#211260000000
0!
0'
#211270000000
1!
b1001 %
1'
b1001 +
#211280000000
0!
0'
#211290000000
1!
b0 %
1'
b0 +
#211300000000
0!
0'
#211310000000
1!
1$
b1 %
1'
1*
b1 +
#211320000000
0!
0'
#211330000000
1!
b10 %
1'
b10 +
#211340000000
1"
1(
#211350000000
0!
0"
b100 &
0'
0(
b100 ,
#211360000000
1!
b11 %
1'
b11 +
#211370000000
0!
0'
#211380000000
1!
b100 %
1'
b100 +
#211390000000
0!
0'
#211400000000
1!
b101 %
1'
b101 +
#211410000000
0!
0'
#211420000000
1!
b110 %
1'
b110 +
#211430000000
0!
0'
#211440000000
1!
b111 %
1'
b111 +
#211450000000
0!
0'
#211460000000
1!
0$
b1000 %
1'
0*
b1000 +
#211470000000
0!
0'
#211480000000
1!
b1001 %
1'
b1001 +
#211490000000
0!
0'
#211500000000
1!
b0 %
1'
b0 +
#211510000000
0!
0'
#211520000000
1!
1$
b1 %
1'
1*
b1 +
#211530000000
0!
0'
#211540000000
1!
b10 %
1'
b10 +
#211550000000
0!
0'
#211560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#211570000000
0!
0'
#211580000000
1!
b100 %
1'
b100 +
#211590000000
0!
0'
#211600000000
1!
b101 %
1'
b101 +
#211610000000
0!
0'
#211620000000
1!
0$
b110 %
1'
0*
b110 +
#211630000000
0!
0'
#211640000000
1!
b111 %
1'
b111 +
#211650000000
0!
0'
#211660000000
1!
b1000 %
1'
b1000 +
#211670000000
0!
0'
#211680000000
1!
b1001 %
1'
b1001 +
#211690000000
0!
0'
#211700000000
1!
b0 %
1'
b0 +
#211710000000
0!
0'
#211720000000
1!
1$
b1 %
1'
1*
b1 +
#211730000000
0!
0'
#211740000000
1!
b10 %
1'
b10 +
#211750000000
0!
0'
#211760000000
1!
b11 %
1'
b11 +
#211770000000
1"
1(
#211780000000
0!
0"
b100 &
0'
0(
b100 ,
#211790000000
1!
b100 %
1'
b100 +
#211800000000
0!
0'
#211810000000
1!
b101 %
1'
b101 +
#211820000000
0!
0'
#211830000000
1!
b110 %
1'
b110 +
#211840000000
0!
0'
#211850000000
1!
b111 %
1'
b111 +
#211860000000
0!
0'
#211870000000
1!
0$
b1000 %
1'
0*
b1000 +
#211880000000
0!
0'
#211890000000
1!
b1001 %
1'
b1001 +
#211900000000
0!
0'
#211910000000
1!
b0 %
1'
b0 +
#211920000000
0!
0'
#211930000000
1!
1$
b1 %
1'
1*
b1 +
#211940000000
0!
0'
#211950000000
1!
b10 %
1'
b10 +
#211960000000
0!
0'
#211970000000
1!
b11 %
1'
b11 +
#211980000000
0!
0'
#211990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#212000000000
0!
0'
#212010000000
1!
b101 %
1'
b101 +
#212020000000
0!
0'
#212030000000
1!
0$
b110 %
1'
0*
b110 +
#212040000000
0!
0'
#212050000000
1!
b111 %
1'
b111 +
#212060000000
0!
0'
#212070000000
1!
b1000 %
1'
b1000 +
#212080000000
0!
0'
#212090000000
1!
b1001 %
1'
b1001 +
#212100000000
0!
0'
#212110000000
1!
b0 %
1'
b0 +
#212120000000
0!
0'
#212130000000
1!
1$
b1 %
1'
1*
b1 +
#212140000000
0!
0'
#212150000000
1!
b10 %
1'
b10 +
#212160000000
0!
0'
#212170000000
1!
b11 %
1'
b11 +
#212180000000
0!
0'
#212190000000
1!
b100 %
1'
b100 +
#212200000000
1"
1(
#212210000000
0!
0"
b100 &
0'
0(
b100 ,
#212220000000
1!
b101 %
1'
b101 +
#212230000000
0!
0'
#212240000000
1!
b110 %
1'
b110 +
#212250000000
0!
0'
#212260000000
1!
b111 %
1'
b111 +
#212270000000
0!
0'
#212280000000
1!
0$
b1000 %
1'
0*
b1000 +
#212290000000
0!
0'
#212300000000
1!
b1001 %
1'
b1001 +
#212310000000
0!
0'
#212320000000
1!
b0 %
1'
b0 +
#212330000000
0!
0'
#212340000000
1!
1$
b1 %
1'
1*
b1 +
#212350000000
0!
0'
#212360000000
1!
b10 %
1'
b10 +
#212370000000
0!
0'
#212380000000
1!
b11 %
1'
b11 +
#212390000000
0!
0'
#212400000000
1!
b100 %
1'
b100 +
#212410000000
0!
0'
#212420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#212430000000
0!
0'
#212440000000
1!
0$
b110 %
1'
0*
b110 +
#212450000000
0!
0'
#212460000000
1!
b111 %
1'
b111 +
#212470000000
0!
0'
#212480000000
1!
b1000 %
1'
b1000 +
#212490000000
0!
0'
#212500000000
1!
b1001 %
1'
b1001 +
#212510000000
0!
0'
#212520000000
1!
b0 %
1'
b0 +
#212530000000
0!
0'
#212540000000
1!
1$
b1 %
1'
1*
b1 +
#212550000000
0!
0'
#212560000000
1!
b10 %
1'
b10 +
#212570000000
0!
0'
#212580000000
1!
b11 %
1'
b11 +
#212590000000
0!
0'
#212600000000
1!
b100 %
1'
b100 +
#212610000000
0!
0'
#212620000000
1!
b101 %
1'
b101 +
#212630000000
1"
1(
#212640000000
0!
0"
b100 &
0'
0(
b100 ,
#212650000000
1!
b110 %
1'
b110 +
#212660000000
0!
0'
#212670000000
1!
b111 %
1'
b111 +
#212680000000
0!
0'
#212690000000
1!
0$
b1000 %
1'
0*
b1000 +
#212700000000
0!
0'
#212710000000
1!
b1001 %
1'
b1001 +
#212720000000
0!
0'
#212730000000
1!
b0 %
1'
b0 +
#212740000000
0!
0'
#212750000000
1!
1$
b1 %
1'
1*
b1 +
#212760000000
0!
0'
#212770000000
1!
b10 %
1'
b10 +
#212780000000
0!
0'
#212790000000
1!
b11 %
1'
b11 +
#212800000000
0!
0'
#212810000000
1!
b100 %
1'
b100 +
#212820000000
0!
0'
#212830000000
1!
b101 %
1'
b101 +
#212840000000
0!
0'
#212850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#212860000000
0!
0'
#212870000000
1!
b111 %
1'
b111 +
#212880000000
0!
0'
#212890000000
1!
b1000 %
1'
b1000 +
#212900000000
0!
0'
#212910000000
1!
b1001 %
1'
b1001 +
#212920000000
0!
0'
#212930000000
1!
b0 %
1'
b0 +
#212940000000
0!
0'
#212950000000
1!
1$
b1 %
1'
1*
b1 +
#212960000000
0!
0'
#212970000000
1!
b10 %
1'
b10 +
#212980000000
0!
0'
#212990000000
1!
b11 %
1'
b11 +
#213000000000
0!
0'
#213010000000
1!
b100 %
1'
b100 +
#213020000000
0!
0'
#213030000000
1!
b101 %
1'
b101 +
#213040000000
0!
0'
#213050000000
1!
0$
b110 %
1'
0*
b110 +
#213060000000
1"
1(
#213070000000
0!
0"
b100 &
0'
0(
b100 ,
#213080000000
1!
1$
b111 %
1'
1*
b111 +
#213090000000
0!
0'
#213100000000
1!
0$
b1000 %
1'
0*
b1000 +
#213110000000
0!
0'
#213120000000
1!
b1001 %
1'
b1001 +
#213130000000
0!
0'
#213140000000
1!
b0 %
1'
b0 +
#213150000000
0!
0'
#213160000000
1!
1$
b1 %
1'
1*
b1 +
#213170000000
0!
0'
#213180000000
1!
b10 %
1'
b10 +
#213190000000
0!
0'
#213200000000
1!
b11 %
1'
b11 +
#213210000000
0!
0'
#213220000000
1!
b100 %
1'
b100 +
#213230000000
0!
0'
#213240000000
1!
b101 %
1'
b101 +
#213250000000
0!
0'
#213260000000
1!
b110 %
1'
b110 +
#213270000000
0!
0'
#213280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#213290000000
0!
0'
#213300000000
1!
b1000 %
1'
b1000 +
#213310000000
0!
0'
#213320000000
1!
b1001 %
1'
b1001 +
#213330000000
0!
0'
#213340000000
1!
b0 %
1'
b0 +
#213350000000
0!
0'
#213360000000
1!
1$
b1 %
1'
1*
b1 +
#213370000000
0!
0'
#213380000000
1!
b10 %
1'
b10 +
#213390000000
0!
0'
#213400000000
1!
b11 %
1'
b11 +
#213410000000
0!
0'
#213420000000
1!
b100 %
1'
b100 +
#213430000000
0!
0'
#213440000000
1!
b101 %
1'
b101 +
#213450000000
0!
0'
#213460000000
1!
0$
b110 %
1'
0*
b110 +
#213470000000
0!
0'
#213480000000
1!
b111 %
1'
b111 +
#213490000000
1"
1(
#213500000000
0!
0"
b100 &
0'
0(
b100 ,
#213510000000
1!
b1000 %
1'
b1000 +
#213520000000
0!
0'
#213530000000
1!
b1001 %
1'
b1001 +
#213540000000
0!
0'
#213550000000
1!
b0 %
1'
b0 +
#213560000000
0!
0'
#213570000000
1!
1$
b1 %
1'
1*
b1 +
#213580000000
0!
0'
#213590000000
1!
b10 %
1'
b10 +
#213600000000
0!
0'
#213610000000
1!
b11 %
1'
b11 +
#213620000000
0!
0'
#213630000000
1!
b100 %
1'
b100 +
#213640000000
0!
0'
#213650000000
1!
b101 %
1'
b101 +
#213660000000
0!
0'
#213670000000
1!
b110 %
1'
b110 +
#213680000000
0!
0'
#213690000000
1!
b111 %
1'
b111 +
#213700000000
0!
0'
#213710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#213720000000
0!
0'
#213730000000
1!
b1001 %
1'
b1001 +
#213740000000
0!
0'
#213750000000
1!
b0 %
1'
b0 +
#213760000000
0!
0'
#213770000000
1!
1$
b1 %
1'
1*
b1 +
#213780000000
0!
0'
#213790000000
1!
b10 %
1'
b10 +
#213800000000
0!
0'
#213810000000
1!
b11 %
1'
b11 +
#213820000000
0!
0'
#213830000000
1!
b100 %
1'
b100 +
#213840000000
0!
0'
#213850000000
1!
b101 %
1'
b101 +
#213860000000
0!
0'
#213870000000
1!
0$
b110 %
1'
0*
b110 +
#213880000000
0!
0'
#213890000000
1!
b111 %
1'
b111 +
#213900000000
0!
0'
#213910000000
1!
b1000 %
1'
b1000 +
#213920000000
1"
1(
#213930000000
0!
0"
b100 &
0'
0(
b100 ,
#213940000000
1!
b1001 %
1'
b1001 +
#213950000000
0!
0'
#213960000000
1!
b0 %
1'
b0 +
#213970000000
0!
0'
#213980000000
1!
1$
b1 %
1'
1*
b1 +
#213990000000
0!
0'
#214000000000
1!
b10 %
1'
b10 +
#214010000000
0!
0'
#214020000000
1!
b11 %
1'
b11 +
#214030000000
0!
0'
#214040000000
1!
b100 %
1'
b100 +
#214050000000
0!
0'
#214060000000
1!
b101 %
1'
b101 +
#214070000000
0!
0'
#214080000000
1!
b110 %
1'
b110 +
#214090000000
0!
0'
#214100000000
1!
b111 %
1'
b111 +
#214110000000
0!
0'
#214120000000
1!
0$
b1000 %
1'
0*
b1000 +
#214130000000
0!
0'
#214140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#214150000000
0!
0'
#214160000000
1!
b0 %
1'
b0 +
#214170000000
0!
0'
#214180000000
1!
1$
b1 %
1'
1*
b1 +
#214190000000
0!
0'
#214200000000
1!
b10 %
1'
b10 +
#214210000000
0!
0'
#214220000000
1!
b11 %
1'
b11 +
#214230000000
0!
0'
#214240000000
1!
b100 %
1'
b100 +
#214250000000
0!
0'
#214260000000
1!
b101 %
1'
b101 +
#214270000000
0!
0'
#214280000000
1!
0$
b110 %
1'
0*
b110 +
#214290000000
0!
0'
#214300000000
1!
b111 %
1'
b111 +
#214310000000
0!
0'
#214320000000
1!
b1000 %
1'
b1000 +
#214330000000
0!
0'
#214340000000
1!
b1001 %
1'
b1001 +
#214350000000
1"
1(
#214360000000
0!
0"
b100 &
0'
0(
b100 ,
#214370000000
1!
b0 %
1'
b0 +
#214380000000
0!
0'
#214390000000
1!
1$
b1 %
1'
1*
b1 +
#214400000000
0!
0'
#214410000000
1!
b10 %
1'
b10 +
#214420000000
0!
0'
#214430000000
1!
b11 %
1'
b11 +
#214440000000
0!
0'
#214450000000
1!
b100 %
1'
b100 +
#214460000000
0!
0'
#214470000000
1!
b101 %
1'
b101 +
#214480000000
0!
0'
#214490000000
1!
b110 %
1'
b110 +
#214500000000
0!
0'
#214510000000
1!
b111 %
1'
b111 +
#214520000000
0!
0'
#214530000000
1!
0$
b1000 %
1'
0*
b1000 +
#214540000000
0!
0'
#214550000000
1!
b1001 %
1'
b1001 +
#214560000000
0!
0'
#214570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#214580000000
0!
0'
#214590000000
1!
1$
b1 %
1'
1*
b1 +
#214600000000
0!
0'
#214610000000
1!
b10 %
1'
b10 +
#214620000000
0!
0'
#214630000000
1!
b11 %
1'
b11 +
#214640000000
0!
0'
#214650000000
1!
b100 %
1'
b100 +
#214660000000
0!
0'
#214670000000
1!
b101 %
1'
b101 +
#214680000000
0!
0'
#214690000000
1!
0$
b110 %
1'
0*
b110 +
#214700000000
0!
0'
#214710000000
1!
b111 %
1'
b111 +
#214720000000
0!
0'
#214730000000
1!
b1000 %
1'
b1000 +
#214740000000
0!
0'
#214750000000
1!
b1001 %
1'
b1001 +
#214760000000
0!
0'
#214770000000
1!
b0 %
1'
b0 +
#214780000000
1"
1(
#214790000000
0!
0"
b100 &
0'
0(
b100 ,
#214800000000
1!
1$
b1 %
1'
1*
b1 +
#214810000000
0!
0'
#214820000000
1!
b10 %
1'
b10 +
#214830000000
0!
0'
#214840000000
1!
b11 %
1'
b11 +
#214850000000
0!
0'
#214860000000
1!
b100 %
1'
b100 +
#214870000000
0!
0'
#214880000000
1!
b101 %
1'
b101 +
#214890000000
0!
0'
#214900000000
1!
b110 %
1'
b110 +
#214910000000
0!
0'
#214920000000
1!
b111 %
1'
b111 +
#214930000000
0!
0'
#214940000000
1!
0$
b1000 %
1'
0*
b1000 +
#214950000000
0!
0'
#214960000000
1!
b1001 %
1'
b1001 +
#214970000000
0!
0'
#214980000000
1!
b0 %
1'
b0 +
#214990000000
0!
0'
#215000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#215010000000
0!
0'
#215020000000
1!
b10 %
1'
b10 +
#215030000000
0!
0'
#215040000000
1!
b11 %
1'
b11 +
#215050000000
0!
0'
#215060000000
1!
b100 %
1'
b100 +
#215070000000
0!
0'
#215080000000
1!
b101 %
1'
b101 +
#215090000000
0!
0'
#215100000000
1!
0$
b110 %
1'
0*
b110 +
#215110000000
0!
0'
#215120000000
1!
b111 %
1'
b111 +
#215130000000
0!
0'
#215140000000
1!
b1000 %
1'
b1000 +
#215150000000
0!
0'
#215160000000
1!
b1001 %
1'
b1001 +
#215170000000
0!
0'
#215180000000
1!
b0 %
1'
b0 +
#215190000000
0!
0'
#215200000000
1!
1$
b1 %
1'
1*
b1 +
#215210000000
1"
1(
#215220000000
0!
0"
b100 &
0'
0(
b100 ,
#215230000000
1!
b10 %
1'
b10 +
#215240000000
0!
0'
#215250000000
1!
b11 %
1'
b11 +
#215260000000
0!
0'
#215270000000
1!
b100 %
1'
b100 +
#215280000000
0!
0'
#215290000000
1!
b101 %
1'
b101 +
#215300000000
0!
0'
#215310000000
1!
b110 %
1'
b110 +
#215320000000
0!
0'
#215330000000
1!
b111 %
1'
b111 +
#215340000000
0!
0'
#215350000000
1!
0$
b1000 %
1'
0*
b1000 +
#215360000000
0!
0'
#215370000000
1!
b1001 %
1'
b1001 +
#215380000000
0!
0'
#215390000000
1!
b0 %
1'
b0 +
#215400000000
0!
0'
#215410000000
1!
1$
b1 %
1'
1*
b1 +
#215420000000
0!
0'
#215430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#215440000000
0!
0'
#215450000000
1!
b11 %
1'
b11 +
#215460000000
0!
0'
#215470000000
1!
b100 %
1'
b100 +
#215480000000
0!
0'
#215490000000
1!
b101 %
1'
b101 +
#215500000000
0!
0'
#215510000000
1!
0$
b110 %
1'
0*
b110 +
#215520000000
0!
0'
#215530000000
1!
b111 %
1'
b111 +
#215540000000
0!
0'
#215550000000
1!
b1000 %
1'
b1000 +
#215560000000
0!
0'
#215570000000
1!
b1001 %
1'
b1001 +
#215580000000
0!
0'
#215590000000
1!
b0 %
1'
b0 +
#215600000000
0!
0'
#215610000000
1!
1$
b1 %
1'
1*
b1 +
#215620000000
0!
0'
#215630000000
1!
b10 %
1'
b10 +
#215640000000
1"
1(
#215650000000
0!
0"
b100 &
0'
0(
b100 ,
#215660000000
1!
b11 %
1'
b11 +
#215670000000
0!
0'
#215680000000
1!
b100 %
1'
b100 +
#215690000000
0!
0'
#215700000000
1!
b101 %
1'
b101 +
#215710000000
0!
0'
#215720000000
1!
b110 %
1'
b110 +
#215730000000
0!
0'
#215740000000
1!
b111 %
1'
b111 +
#215750000000
0!
0'
#215760000000
1!
0$
b1000 %
1'
0*
b1000 +
#215770000000
0!
0'
#215780000000
1!
b1001 %
1'
b1001 +
#215790000000
0!
0'
#215800000000
1!
b0 %
1'
b0 +
#215810000000
0!
0'
#215820000000
1!
1$
b1 %
1'
1*
b1 +
#215830000000
0!
0'
#215840000000
1!
b10 %
1'
b10 +
#215850000000
0!
0'
#215860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#215870000000
0!
0'
#215880000000
1!
b100 %
1'
b100 +
#215890000000
0!
0'
#215900000000
1!
b101 %
1'
b101 +
#215910000000
0!
0'
#215920000000
1!
0$
b110 %
1'
0*
b110 +
#215930000000
0!
0'
#215940000000
1!
b111 %
1'
b111 +
#215950000000
0!
0'
#215960000000
1!
b1000 %
1'
b1000 +
#215970000000
0!
0'
#215980000000
1!
b1001 %
1'
b1001 +
#215990000000
0!
0'
#216000000000
1!
b0 %
1'
b0 +
#216010000000
0!
0'
#216020000000
1!
1$
b1 %
1'
1*
b1 +
#216030000000
0!
0'
#216040000000
1!
b10 %
1'
b10 +
#216050000000
0!
0'
#216060000000
1!
b11 %
1'
b11 +
#216070000000
1"
1(
#216080000000
0!
0"
b100 &
0'
0(
b100 ,
#216090000000
1!
b100 %
1'
b100 +
#216100000000
0!
0'
#216110000000
1!
b101 %
1'
b101 +
#216120000000
0!
0'
#216130000000
1!
b110 %
1'
b110 +
#216140000000
0!
0'
#216150000000
1!
b111 %
1'
b111 +
#216160000000
0!
0'
#216170000000
1!
0$
b1000 %
1'
0*
b1000 +
#216180000000
0!
0'
#216190000000
1!
b1001 %
1'
b1001 +
#216200000000
0!
0'
#216210000000
1!
b0 %
1'
b0 +
#216220000000
0!
0'
#216230000000
1!
1$
b1 %
1'
1*
b1 +
#216240000000
0!
0'
#216250000000
1!
b10 %
1'
b10 +
#216260000000
0!
0'
#216270000000
1!
b11 %
1'
b11 +
#216280000000
0!
0'
#216290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#216300000000
0!
0'
#216310000000
1!
b101 %
1'
b101 +
#216320000000
0!
0'
#216330000000
1!
0$
b110 %
1'
0*
b110 +
#216340000000
0!
0'
#216350000000
1!
b111 %
1'
b111 +
#216360000000
0!
0'
#216370000000
1!
b1000 %
1'
b1000 +
#216380000000
0!
0'
#216390000000
1!
b1001 %
1'
b1001 +
#216400000000
0!
0'
#216410000000
1!
b0 %
1'
b0 +
#216420000000
0!
0'
#216430000000
1!
1$
b1 %
1'
1*
b1 +
#216440000000
0!
0'
#216450000000
1!
b10 %
1'
b10 +
#216460000000
0!
0'
#216470000000
1!
b11 %
1'
b11 +
#216480000000
0!
0'
#216490000000
1!
b100 %
1'
b100 +
#216500000000
1"
1(
#216510000000
0!
0"
b100 &
0'
0(
b100 ,
#216520000000
1!
b101 %
1'
b101 +
#216530000000
0!
0'
#216540000000
1!
b110 %
1'
b110 +
#216550000000
0!
0'
#216560000000
1!
b111 %
1'
b111 +
#216570000000
0!
0'
#216580000000
1!
0$
b1000 %
1'
0*
b1000 +
#216590000000
0!
0'
#216600000000
1!
b1001 %
1'
b1001 +
#216610000000
0!
0'
#216620000000
1!
b0 %
1'
b0 +
#216630000000
0!
0'
#216640000000
1!
1$
b1 %
1'
1*
b1 +
#216650000000
0!
0'
#216660000000
1!
b10 %
1'
b10 +
#216670000000
0!
0'
#216680000000
1!
b11 %
1'
b11 +
#216690000000
0!
0'
#216700000000
1!
b100 %
1'
b100 +
#216710000000
0!
0'
#216720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#216730000000
0!
0'
#216740000000
1!
0$
b110 %
1'
0*
b110 +
#216750000000
0!
0'
#216760000000
1!
b111 %
1'
b111 +
#216770000000
0!
0'
#216780000000
1!
b1000 %
1'
b1000 +
#216790000000
0!
0'
#216800000000
1!
b1001 %
1'
b1001 +
#216810000000
0!
0'
#216820000000
1!
b0 %
1'
b0 +
#216830000000
0!
0'
#216840000000
1!
1$
b1 %
1'
1*
b1 +
#216850000000
0!
0'
#216860000000
1!
b10 %
1'
b10 +
#216870000000
0!
0'
#216880000000
1!
b11 %
1'
b11 +
#216890000000
0!
0'
#216900000000
1!
b100 %
1'
b100 +
#216910000000
0!
0'
#216920000000
1!
b101 %
1'
b101 +
#216930000000
1"
1(
#216940000000
0!
0"
b100 &
0'
0(
b100 ,
#216950000000
1!
b110 %
1'
b110 +
#216960000000
0!
0'
#216970000000
1!
b111 %
1'
b111 +
#216980000000
0!
0'
#216990000000
1!
0$
b1000 %
1'
0*
b1000 +
#217000000000
0!
0'
#217010000000
1!
b1001 %
1'
b1001 +
#217020000000
0!
0'
#217030000000
1!
b0 %
1'
b0 +
#217040000000
0!
0'
#217050000000
1!
1$
b1 %
1'
1*
b1 +
#217060000000
0!
0'
#217070000000
1!
b10 %
1'
b10 +
#217080000000
0!
0'
#217090000000
1!
b11 %
1'
b11 +
#217100000000
0!
0'
#217110000000
1!
b100 %
1'
b100 +
#217120000000
0!
0'
#217130000000
1!
b101 %
1'
b101 +
#217140000000
0!
0'
#217150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#217160000000
0!
0'
#217170000000
1!
b111 %
1'
b111 +
#217180000000
0!
0'
#217190000000
1!
b1000 %
1'
b1000 +
#217200000000
0!
0'
#217210000000
1!
b1001 %
1'
b1001 +
#217220000000
0!
0'
#217230000000
1!
b0 %
1'
b0 +
#217240000000
0!
0'
#217250000000
1!
1$
b1 %
1'
1*
b1 +
#217260000000
0!
0'
#217270000000
1!
b10 %
1'
b10 +
#217280000000
0!
0'
#217290000000
1!
b11 %
1'
b11 +
#217300000000
0!
0'
#217310000000
1!
b100 %
1'
b100 +
#217320000000
0!
0'
#217330000000
1!
b101 %
1'
b101 +
#217340000000
0!
0'
#217350000000
1!
0$
b110 %
1'
0*
b110 +
#217360000000
1"
1(
#217370000000
0!
0"
b100 &
0'
0(
b100 ,
#217380000000
1!
1$
b111 %
1'
1*
b111 +
#217390000000
0!
0'
#217400000000
1!
0$
b1000 %
1'
0*
b1000 +
#217410000000
0!
0'
#217420000000
1!
b1001 %
1'
b1001 +
#217430000000
0!
0'
#217440000000
1!
b0 %
1'
b0 +
#217450000000
0!
0'
#217460000000
1!
1$
b1 %
1'
1*
b1 +
#217470000000
0!
0'
#217480000000
1!
b10 %
1'
b10 +
#217490000000
0!
0'
#217500000000
1!
b11 %
1'
b11 +
#217510000000
0!
0'
#217520000000
1!
b100 %
1'
b100 +
#217530000000
0!
0'
#217540000000
1!
b101 %
1'
b101 +
#217550000000
0!
0'
#217560000000
1!
b110 %
1'
b110 +
#217570000000
0!
0'
#217580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#217590000000
0!
0'
#217600000000
1!
b1000 %
1'
b1000 +
#217610000000
0!
0'
#217620000000
1!
b1001 %
1'
b1001 +
#217630000000
0!
0'
#217640000000
1!
b0 %
1'
b0 +
#217650000000
0!
0'
#217660000000
1!
1$
b1 %
1'
1*
b1 +
#217670000000
0!
0'
#217680000000
1!
b10 %
1'
b10 +
#217690000000
0!
0'
#217700000000
1!
b11 %
1'
b11 +
#217710000000
0!
0'
#217720000000
1!
b100 %
1'
b100 +
#217730000000
0!
0'
#217740000000
1!
b101 %
1'
b101 +
#217750000000
0!
0'
#217760000000
1!
0$
b110 %
1'
0*
b110 +
#217770000000
0!
0'
#217780000000
1!
b111 %
1'
b111 +
#217790000000
1"
1(
#217800000000
0!
0"
b100 &
0'
0(
b100 ,
#217810000000
1!
b1000 %
1'
b1000 +
#217820000000
0!
0'
#217830000000
1!
b1001 %
1'
b1001 +
#217840000000
0!
0'
#217850000000
1!
b0 %
1'
b0 +
#217860000000
0!
0'
#217870000000
1!
1$
b1 %
1'
1*
b1 +
#217880000000
0!
0'
#217890000000
1!
b10 %
1'
b10 +
#217900000000
0!
0'
#217910000000
1!
b11 %
1'
b11 +
#217920000000
0!
0'
#217930000000
1!
b100 %
1'
b100 +
#217940000000
0!
0'
#217950000000
1!
b101 %
1'
b101 +
#217960000000
0!
0'
#217970000000
1!
b110 %
1'
b110 +
#217980000000
0!
0'
#217990000000
1!
b111 %
1'
b111 +
#218000000000
0!
0'
#218010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#218020000000
0!
0'
#218030000000
1!
b1001 %
1'
b1001 +
#218040000000
0!
0'
#218050000000
1!
b0 %
1'
b0 +
#218060000000
0!
0'
#218070000000
1!
1$
b1 %
1'
1*
b1 +
#218080000000
0!
0'
#218090000000
1!
b10 %
1'
b10 +
#218100000000
0!
0'
#218110000000
1!
b11 %
1'
b11 +
#218120000000
0!
0'
#218130000000
1!
b100 %
1'
b100 +
#218140000000
0!
0'
#218150000000
1!
b101 %
1'
b101 +
#218160000000
0!
0'
#218170000000
1!
0$
b110 %
1'
0*
b110 +
#218180000000
0!
0'
#218190000000
1!
b111 %
1'
b111 +
#218200000000
0!
0'
#218210000000
1!
b1000 %
1'
b1000 +
#218220000000
1"
1(
#218230000000
0!
0"
b100 &
0'
0(
b100 ,
#218240000000
1!
b1001 %
1'
b1001 +
#218250000000
0!
0'
#218260000000
1!
b0 %
1'
b0 +
#218270000000
0!
0'
#218280000000
1!
1$
b1 %
1'
1*
b1 +
#218290000000
0!
0'
#218300000000
1!
b10 %
1'
b10 +
#218310000000
0!
0'
#218320000000
1!
b11 %
1'
b11 +
#218330000000
0!
0'
#218340000000
1!
b100 %
1'
b100 +
#218350000000
0!
0'
#218360000000
1!
b101 %
1'
b101 +
#218370000000
0!
0'
#218380000000
1!
b110 %
1'
b110 +
#218390000000
0!
0'
#218400000000
1!
b111 %
1'
b111 +
#218410000000
0!
0'
#218420000000
1!
0$
b1000 %
1'
0*
b1000 +
#218430000000
0!
0'
#218440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#218450000000
0!
0'
#218460000000
1!
b0 %
1'
b0 +
#218470000000
0!
0'
#218480000000
1!
1$
b1 %
1'
1*
b1 +
#218490000000
0!
0'
#218500000000
1!
b10 %
1'
b10 +
#218510000000
0!
0'
#218520000000
1!
b11 %
1'
b11 +
#218530000000
0!
0'
#218540000000
1!
b100 %
1'
b100 +
#218550000000
0!
0'
#218560000000
1!
b101 %
1'
b101 +
#218570000000
0!
0'
#218580000000
1!
0$
b110 %
1'
0*
b110 +
#218590000000
0!
0'
#218600000000
1!
b111 %
1'
b111 +
#218610000000
0!
0'
#218620000000
1!
b1000 %
1'
b1000 +
#218630000000
0!
0'
#218640000000
1!
b1001 %
1'
b1001 +
#218650000000
1"
1(
#218660000000
0!
0"
b100 &
0'
0(
b100 ,
#218670000000
1!
b0 %
1'
b0 +
#218680000000
0!
0'
#218690000000
1!
1$
b1 %
1'
1*
b1 +
#218700000000
0!
0'
#218710000000
1!
b10 %
1'
b10 +
#218720000000
0!
0'
#218730000000
1!
b11 %
1'
b11 +
#218740000000
0!
0'
#218750000000
1!
b100 %
1'
b100 +
#218760000000
0!
0'
#218770000000
1!
b101 %
1'
b101 +
#218780000000
0!
0'
#218790000000
1!
b110 %
1'
b110 +
#218800000000
0!
0'
#218810000000
1!
b111 %
1'
b111 +
#218820000000
0!
0'
#218830000000
1!
0$
b1000 %
1'
0*
b1000 +
#218840000000
0!
0'
#218850000000
1!
b1001 %
1'
b1001 +
#218860000000
0!
0'
#218870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#218880000000
0!
0'
#218890000000
1!
1$
b1 %
1'
1*
b1 +
#218900000000
0!
0'
#218910000000
1!
b10 %
1'
b10 +
#218920000000
0!
0'
#218930000000
1!
b11 %
1'
b11 +
#218940000000
0!
0'
#218950000000
1!
b100 %
1'
b100 +
#218960000000
0!
0'
#218970000000
1!
b101 %
1'
b101 +
#218980000000
0!
0'
#218990000000
1!
0$
b110 %
1'
0*
b110 +
#219000000000
0!
0'
#219010000000
1!
b111 %
1'
b111 +
#219020000000
0!
0'
#219030000000
1!
b1000 %
1'
b1000 +
#219040000000
0!
0'
#219050000000
1!
b1001 %
1'
b1001 +
#219060000000
0!
0'
#219070000000
1!
b0 %
1'
b0 +
#219080000000
1"
1(
#219090000000
0!
0"
b100 &
0'
0(
b100 ,
#219100000000
1!
1$
b1 %
1'
1*
b1 +
#219110000000
0!
0'
#219120000000
1!
b10 %
1'
b10 +
#219130000000
0!
0'
#219140000000
1!
b11 %
1'
b11 +
#219150000000
0!
0'
#219160000000
1!
b100 %
1'
b100 +
#219170000000
0!
0'
#219180000000
1!
b101 %
1'
b101 +
#219190000000
0!
0'
#219200000000
1!
b110 %
1'
b110 +
#219210000000
0!
0'
#219220000000
1!
b111 %
1'
b111 +
#219230000000
0!
0'
#219240000000
1!
0$
b1000 %
1'
0*
b1000 +
#219250000000
0!
0'
#219260000000
1!
b1001 %
1'
b1001 +
#219270000000
0!
0'
#219280000000
1!
b0 %
1'
b0 +
#219290000000
0!
0'
#219300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#219310000000
0!
0'
#219320000000
1!
b10 %
1'
b10 +
#219330000000
0!
0'
#219340000000
1!
b11 %
1'
b11 +
#219350000000
0!
0'
#219360000000
1!
b100 %
1'
b100 +
#219370000000
0!
0'
#219380000000
1!
b101 %
1'
b101 +
#219390000000
0!
0'
#219400000000
1!
0$
b110 %
1'
0*
b110 +
#219410000000
0!
0'
#219420000000
1!
b111 %
1'
b111 +
#219430000000
0!
0'
#219440000000
1!
b1000 %
1'
b1000 +
#219450000000
0!
0'
#219460000000
1!
b1001 %
1'
b1001 +
#219470000000
0!
0'
#219480000000
1!
b0 %
1'
b0 +
#219490000000
0!
0'
#219500000000
1!
1$
b1 %
1'
1*
b1 +
#219510000000
1"
1(
#219520000000
0!
0"
b100 &
0'
0(
b100 ,
#219530000000
1!
b10 %
1'
b10 +
#219540000000
0!
0'
#219550000000
1!
b11 %
1'
b11 +
#219560000000
0!
0'
#219570000000
1!
b100 %
1'
b100 +
#219580000000
0!
0'
#219590000000
1!
b101 %
1'
b101 +
#219600000000
0!
0'
#219610000000
1!
b110 %
1'
b110 +
#219620000000
0!
0'
#219630000000
1!
b111 %
1'
b111 +
#219640000000
0!
0'
#219650000000
1!
0$
b1000 %
1'
0*
b1000 +
#219660000000
0!
0'
#219670000000
1!
b1001 %
1'
b1001 +
#219680000000
0!
0'
#219690000000
1!
b0 %
1'
b0 +
#219700000000
0!
0'
#219710000000
1!
1$
b1 %
1'
1*
b1 +
#219720000000
0!
0'
#219730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#219740000000
0!
0'
#219750000000
1!
b11 %
1'
b11 +
#219760000000
0!
0'
#219770000000
1!
b100 %
1'
b100 +
#219780000000
0!
0'
#219790000000
1!
b101 %
1'
b101 +
#219800000000
0!
0'
#219810000000
1!
0$
b110 %
1'
0*
b110 +
#219820000000
0!
0'
#219830000000
1!
b111 %
1'
b111 +
#219840000000
0!
0'
#219850000000
1!
b1000 %
1'
b1000 +
#219860000000
0!
0'
#219870000000
1!
b1001 %
1'
b1001 +
#219880000000
0!
0'
#219890000000
1!
b0 %
1'
b0 +
#219900000000
0!
0'
#219910000000
1!
1$
b1 %
1'
1*
b1 +
#219920000000
0!
0'
#219930000000
1!
b10 %
1'
b10 +
#219940000000
1"
1(
#219950000000
0!
0"
b100 &
0'
0(
b100 ,
#219960000000
1!
b11 %
1'
b11 +
#219970000000
0!
0'
#219980000000
1!
b100 %
1'
b100 +
#219990000000
0!
0'
#220000000000
1!
b101 %
1'
b101 +
#220010000000
0!
0'
#220020000000
1!
b110 %
1'
b110 +
#220030000000
0!
0'
#220040000000
1!
b111 %
1'
b111 +
#220050000000
0!
0'
#220060000000
1!
0$
b1000 %
1'
0*
b1000 +
#220070000000
0!
0'
#220080000000
1!
b1001 %
1'
b1001 +
#220090000000
0!
0'
#220100000000
1!
b0 %
1'
b0 +
#220110000000
0!
0'
#220120000000
1!
1$
b1 %
1'
1*
b1 +
#220130000000
0!
0'
#220140000000
1!
b10 %
1'
b10 +
#220150000000
0!
0'
#220160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#220170000000
0!
0'
#220180000000
1!
b100 %
1'
b100 +
#220190000000
0!
0'
#220200000000
1!
b101 %
1'
b101 +
#220210000000
0!
0'
#220220000000
1!
0$
b110 %
1'
0*
b110 +
#220230000000
0!
0'
#220240000000
1!
b111 %
1'
b111 +
#220250000000
0!
0'
#220260000000
1!
b1000 %
1'
b1000 +
#220270000000
0!
0'
#220280000000
1!
b1001 %
1'
b1001 +
#220290000000
0!
0'
#220300000000
1!
b0 %
1'
b0 +
#220310000000
0!
0'
#220320000000
1!
1$
b1 %
1'
1*
b1 +
#220330000000
0!
0'
#220340000000
1!
b10 %
1'
b10 +
#220350000000
0!
0'
#220360000000
1!
b11 %
1'
b11 +
#220370000000
1"
1(
#220380000000
0!
0"
b100 &
0'
0(
b100 ,
#220390000000
1!
b100 %
1'
b100 +
#220400000000
0!
0'
#220410000000
1!
b101 %
1'
b101 +
#220420000000
0!
0'
#220430000000
1!
b110 %
1'
b110 +
#220440000000
0!
0'
#220450000000
1!
b111 %
1'
b111 +
#220460000000
0!
0'
#220470000000
1!
0$
b1000 %
1'
0*
b1000 +
#220480000000
0!
0'
#220490000000
1!
b1001 %
1'
b1001 +
#220500000000
0!
0'
#220510000000
1!
b0 %
1'
b0 +
#220520000000
0!
0'
#220530000000
1!
1$
b1 %
1'
1*
b1 +
#220540000000
0!
0'
#220550000000
1!
b10 %
1'
b10 +
#220560000000
0!
0'
#220570000000
1!
b11 %
1'
b11 +
#220580000000
0!
0'
#220590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#220600000000
0!
0'
#220610000000
1!
b101 %
1'
b101 +
#220620000000
0!
0'
#220630000000
1!
0$
b110 %
1'
0*
b110 +
#220640000000
0!
0'
#220650000000
1!
b111 %
1'
b111 +
#220660000000
0!
0'
#220670000000
1!
b1000 %
1'
b1000 +
#220680000000
0!
0'
#220690000000
1!
b1001 %
1'
b1001 +
#220700000000
0!
0'
#220710000000
1!
b0 %
1'
b0 +
#220720000000
0!
0'
#220730000000
1!
1$
b1 %
1'
1*
b1 +
#220740000000
0!
0'
#220750000000
1!
b10 %
1'
b10 +
#220760000000
0!
0'
#220770000000
1!
b11 %
1'
b11 +
#220780000000
0!
0'
#220790000000
1!
b100 %
1'
b100 +
#220800000000
1"
1(
#220810000000
0!
0"
b100 &
0'
0(
b100 ,
#220820000000
1!
b101 %
1'
b101 +
#220830000000
0!
0'
#220840000000
1!
b110 %
1'
b110 +
#220850000000
0!
0'
#220860000000
1!
b111 %
1'
b111 +
#220870000000
0!
0'
#220880000000
1!
0$
b1000 %
1'
0*
b1000 +
#220890000000
0!
0'
#220900000000
1!
b1001 %
1'
b1001 +
#220910000000
0!
0'
#220920000000
1!
b0 %
1'
b0 +
#220930000000
0!
0'
#220940000000
1!
1$
b1 %
1'
1*
b1 +
#220950000000
0!
0'
#220960000000
1!
b10 %
1'
b10 +
#220970000000
0!
0'
#220980000000
1!
b11 %
1'
b11 +
#220990000000
0!
0'
#221000000000
1!
b100 %
1'
b100 +
#221010000000
0!
0'
#221020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#221030000000
0!
0'
#221040000000
1!
0$
b110 %
1'
0*
b110 +
#221050000000
0!
0'
#221060000000
1!
b111 %
1'
b111 +
#221070000000
0!
0'
#221080000000
1!
b1000 %
1'
b1000 +
#221090000000
0!
0'
#221100000000
1!
b1001 %
1'
b1001 +
#221110000000
0!
0'
#221120000000
1!
b0 %
1'
b0 +
#221130000000
0!
0'
#221140000000
1!
1$
b1 %
1'
1*
b1 +
#221150000000
0!
0'
#221160000000
1!
b10 %
1'
b10 +
#221170000000
0!
0'
#221180000000
1!
b11 %
1'
b11 +
#221190000000
0!
0'
#221200000000
1!
b100 %
1'
b100 +
#221210000000
0!
0'
#221220000000
1!
b101 %
1'
b101 +
#221230000000
1"
1(
#221240000000
0!
0"
b100 &
0'
0(
b100 ,
#221250000000
1!
b110 %
1'
b110 +
#221260000000
0!
0'
#221270000000
1!
b111 %
1'
b111 +
#221280000000
0!
0'
#221290000000
1!
0$
b1000 %
1'
0*
b1000 +
#221300000000
0!
0'
#221310000000
1!
b1001 %
1'
b1001 +
#221320000000
0!
0'
#221330000000
1!
b0 %
1'
b0 +
#221340000000
0!
0'
#221350000000
1!
1$
b1 %
1'
1*
b1 +
#221360000000
0!
0'
#221370000000
1!
b10 %
1'
b10 +
#221380000000
0!
0'
#221390000000
1!
b11 %
1'
b11 +
#221400000000
0!
0'
#221410000000
1!
b100 %
1'
b100 +
#221420000000
0!
0'
#221430000000
1!
b101 %
1'
b101 +
#221440000000
0!
0'
#221450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#221460000000
0!
0'
#221470000000
1!
b111 %
1'
b111 +
#221480000000
0!
0'
#221490000000
1!
b1000 %
1'
b1000 +
#221500000000
0!
0'
#221510000000
1!
b1001 %
1'
b1001 +
#221520000000
0!
0'
#221530000000
1!
b0 %
1'
b0 +
#221540000000
0!
0'
#221550000000
1!
1$
b1 %
1'
1*
b1 +
#221560000000
0!
0'
#221570000000
1!
b10 %
1'
b10 +
#221580000000
0!
0'
#221590000000
1!
b11 %
1'
b11 +
#221600000000
0!
0'
#221610000000
1!
b100 %
1'
b100 +
#221620000000
0!
0'
#221630000000
1!
b101 %
1'
b101 +
#221640000000
0!
0'
#221650000000
1!
0$
b110 %
1'
0*
b110 +
#221660000000
1"
1(
#221670000000
0!
0"
b100 &
0'
0(
b100 ,
#221680000000
1!
1$
b111 %
1'
1*
b111 +
#221690000000
0!
0'
#221700000000
1!
0$
b1000 %
1'
0*
b1000 +
#221710000000
0!
0'
#221720000000
1!
b1001 %
1'
b1001 +
#221730000000
0!
0'
#221740000000
1!
b0 %
1'
b0 +
#221750000000
0!
0'
#221760000000
1!
1$
b1 %
1'
1*
b1 +
#221770000000
0!
0'
#221780000000
1!
b10 %
1'
b10 +
#221790000000
0!
0'
#221800000000
1!
b11 %
1'
b11 +
#221810000000
0!
0'
#221820000000
1!
b100 %
1'
b100 +
#221830000000
0!
0'
#221840000000
1!
b101 %
1'
b101 +
#221850000000
0!
0'
#221860000000
1!
b110 %
1'
b110 +
#221870000000
0!
0'
#221880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#221890000000
0!
0'
#221900000000
1!
b1000 %
1'
b1000 +
#221910000000
0!
0'
#221920000000
1!
b1001 %
1'
b1001 +
#221930000000
0!
0'
#221940000000
1!
b0 %
1'
b0 +
#221950000000
0!
0'
#221960000000
1!
1$
b1 %
1'
1*
b1 +
#221970000000
0!
0'
#221980000000
1!
b10 %
1'
b10 +
#221990000000
0!
0'
#222000000000
1!
b11 %
1'
b11 +
#222010000000
0!
0'
#222020000000
1!
b100 %
1'
b100 +
#222030000000
0!
0'
#222040000000
1!
b101 %
1'
b101 +
#222050000000
0!
0'
#222060000000
1!
0$
b110 %
1'
0*
b110 +
#222070000000
0!
0'
#222080000000
1!
b111 %
1'
b111 +
#222090000000
1"
1(
#222100000000
0!
0"
b100 &
0'
0(
b100 ,
#222110000000
1!
b1000 %
1'
b1000 +
#222120000000
0!
0'
#222130000000
1!
b1001 %
1'
b1001 +
#222140000000
0!
0'
#222150000000
1!
b0 %
1'
b0 +
#222160000000
0!
0'
#222170000000
1!
1$
b1 %
1'
1*
b1 +
#222180000000
0!
0'
#222190000000
1!
b10 %
1'
b10 +
#222200000000
0!
0'
#222210000000
1!
b11 %
1'
b11 +
#222220000000
0!
0'
#222230000000
1!
b100 %
1'
b100 +
#222240000000
0!
0'
#222250000000
1!
b101 %
1'
b101 +
#222260000000
0!
0'
#222270000000
1!
b110 %
1'
b110 +
#222280000000
0!
0'
#222290000000
1!
b111 %
1'
b111 +
#222300000000
0!
0'
#222310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#222320000000
0!
0'
#222330000000
1!
b1001 %
1'
b1001 +
#222340000000
0!
0'
#222350000000
1!
b0 %
1'
b0 +
#222360000000
0!
0'
#222370000000
1!
1$
b1 %
1'
1*
b1 +
#222380000000
0!
0'
#222390000000
1!
b10 %
1'
b10 +
#222400000000
0!
0'
#222410000000
1!
b11 %
1'
b11 +
#222420000000
0!
0'
#222430000000
1!
b100 %
1'
b100 +
#222440000000
0!
0'
#222450000000
1!
b101 %
1'
b101 +
#222460000000
0!
0'
#222470000000
1!
0$
b110 %
1'
0*
b110 +
#222480000000
0!
0'
#222490000000
1!
b111 %
1'
b111 +
#222500000000
0!
0'
#222510000000
1!
b1000 %
1'
b1000 +
#222520000000
1"
1(
#222530000000
0!
0"
b100 &
0'
0(
b100 ,
#222540000000
1!
b1001 %
1'
b1001 +
#222550000000
0!
0'
#222560000000
1!
b0 %
1'
b0 +
#222570000000
0!
0'
#222580000000
1!
1$
b1 %
1'
1*
b1 +
#222590000000
0!
0'
#222600000000
1!
b10 %
1'
b10 +
#222610000000
0!
0'
#222620000000
1!
b11 %
1'
b11 +
#222630000000
0!
0'
#222640000000
1!
b100 %
1'
b100 +
#222650000000
0!
0'
#222660000000
1!
b101 %
1'
b101 +
#222670000000
0!
0'
#222680000000
1!
b110 %
1'
b110 +
#222690000000
0!
0'
#222700000000
1!
b111 %
1'
b111 +
#222710000000
0!
0'
#222720000000
1!
0$
b1000 %
1'
0*
b1000 +
#222730000000
0!
0'
#222740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#222750000000
0!
0'
#222760000000
1!
b0 %
1'
b0 +
#222770000000
0!
0'
#222780000000
1!
1$
b1 %
1'
1*
b1 +
#222790000000
0!
0'
#222800000000
1!
b10 %
1'
b10 +
#222810000000
0!
0'
#222820000000
1!
b11 %
1'
b11 +
#222830000000
0!
0'
#222840000000
1!
b100 %
1'
b100 +
#222850000000
0!
0'
#222860000000
1!
b101 %
1'
b101 +
#222870000000
0!
0'
#222880000000
1!
0$
b110 %
1'
0*
b110 +
#222890000000
0!
0'
#222900000000
1!
b111 %
1'
b111 +
#222910000000
0!
0'
#222920000000
1!
b1000 %
1'
b1000 +
#222930000000
0!
0'
#222940000000
1!
b1001 %
1'
b1001 +
#222950000000
1"
1(
#222960000000
0!
0"
b100 &
0'
0(
b100 ,
#222970000000
1!
b0 %
1'
b0 +
#222980000000
0!
0'
#222990000000
1!
1$
b1 %
1'
1*
b1 +
#223000000000
0!
0'
#223010000000
1!
b10 %
1'
b10 +
#223020000000
0!
0'
#223030000000
1!
b11 %
1'
b11 +
#223040000000
0!
0'
#223050000000
1!
b100 %
1'
b100 +
#223060000000
0!
0'
#223070000000
1!
b101 %
1'
b101 +
#223080000000
0!
0'
#223090000000
1!
b110 %
1'
b110 +
#223100000000
0!
0'
#223110000000
1!
b111 %
1'
b111 +
#223120000000
0!
0'
#223130000000
1!
0$
b1000 %
1'
0*
b1000 +
#223140000000
0!
0'
#223150000000
1!
b1001 %
1'
b1001 +
#223160000000
0!
0'
#223170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#223180000000
0!
0'
#223190000000
1!
1$
b1 %
1'
1*
b1 +
#223200000000
0!
0'
#223210000000
1!
b10 %
1'
b10 +
#223220000000
0!
0'
#223230000000
1!
b11 %
1'
b11 +
#223240000000
0!
0'
#223250000000
1!
b100 %
1'
b100 +
#223260000000
0!
0'
#223270000000
1!
b101 %
1'
b101 +
#223280000000
0!
0'
#223290000000
1!
0$
b110 %
1'
0*
b110 +
#223300000000
0!
0'
#223310000000
1!
b111 %
1'
b111 +
#223320000000
0!
0'
#223330000000
1!
b1000 %
1'
b1000 +
#223340000000
0!
0'
#223350000000
1!
b1001 %
1'
b1001 +
#223360000000
0!
0'
#223370000000
1!
b0 %
1'
b0 +
#223380000000
1"
1(
#223390000000
0!
0"
b100 &
0'
0(
b100 ,
#223400000000
1!
1$
b1 %
1'
1*
b1 +
#223410000000
0!
0'
#223420000000
1!
b10 %
1'
b10 +
#223430000000
0!
0'
#223440000000
1!
b11 %
1'
b11 +
#223450000000
0!
0'
#223460000000
1!
b100 %
1'
b100 +
#223470000000
0!
0'
#223480000000
1!
b101 %
1'
b101 +
#223490000000
0!
0'
#223500000000
1!
b110 %
1'
b110 +
#223510000000
0!
0'
#223520000000
1!
b111 %
1'
b111 +
#223530000000
0!
0'
#223540000000
1!
0$
b1000 %
1'
0*
b1000 +
#223550000000
0!
0'
#223560000000
1!
b1001 %
1'
b1001 +
#223570000000
0!
0'
#223580000000
1!
b0 %
1'
b0 +
#223590000000
0!
0'
#223600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#223610000000
0!
0'
#223620000000
1!
b10 %
1'
b10 +
#223630000000
0!
0'
#223640000000
1!
b11 %
1'
b11 +
#223650000000
0!
0'
#223660000000
1!
b100 %
1'
b100 +
#223670000000
0!
0'
#223680000000
1!
b101 %
1'
b101 +
#223690000000
0!
0'
#223700000000
1!
0$
b110 %
1'
0*
b110 +
#223710000000
0!
0'
#223720000000
1!
b111 %
1'
b111 +
#223730000000
0!
0'
#223740000000
1!
b1000 %
1'
b1000 +
#223750000000
0!
0'
#223760000000
1!
b1001 %
1'
b1001 +
#223770000000
0!
0'
#223780000000
1!
b0 %
1'
b0 +
#223790000000
0!
0'
#223800000000
1!
1$
b1 %
1'
1*
b1 +
#223810000000
1"
1(
#223820000000
0!
0"
b100 &
0'
0(
b100 ,
#223830000000
1!
b10 %
1'
b10 +
#223840000000
0!
0'
#223850000000
1!
b11 %
1'
b11 +
#223860000000
0!
0'
#223870000000
1!
b100 %
1'
b100 +
#223880000000
0!
0'
#223890000000
1!
b101 %
1'
b101 +
#223900000000
0!
0'
#223910000000
1!
b110 %
1'
b110 +
#223920000000
0!
0'
#223930000000
1!
b111 %
1'
b111 +
#223940000000
0!
0'
#223950000000
1!
0$
b1000 %
1'
0*
b1000 +
#223960000000
0!
0'
#223970000000
1!
b1001 %
1'
b1001 +
#223980000000
0!
0'
#223990000000
1!
b0 %
1'
b0 +
#224000000000
0!
0'
#224010000000
1!
1$
b1 %
1'
1*
b1 +
#224020000000
0!
0'
#224030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#224040000000
0!
0'
#224050000000
1!
b11 %
1'
b11 +
#224060000000
0!
0'
#224070000000
1!
b100 %
1'
b100 +
#224080000000
0!
0'
#224090000000
1!
b101 %
1'
b101 +
#224100000000
0!
0'
#224110000000
1!
0$
b110 %
1'
0*
b110 +
#224120000000
0!
0'
#224130000000
1!
b111 %
1'
b111 +
#224140000000
0!
0'
#224150000000
1!
b1000 %
1'
b1000 +
#224160000000
0!
0'
#224170000000
1!
b1001 %
1'
b1001 +
#224180000000
0!
0'
#224190000000
1!
b0 %
1'
b0 +
#224200000000
0!
0'
#224210000000
1!
1$
b1 %
1'
1*
b1 +
#224220000000
0!
0'
#224230000000
1!
b10 %
1'
b10 +
#224240000000
1"
1(
#224250000000
0!
0"
b100 &
0'
0(
b100 ,
#224260000000
1!
b11 %
1'
b11 +
#224270000000
0!
0'
#224280000000
1!
b100 %
1'
b100 +
#224290000000
0!
0'
#224300000000
1!
b101 %
1'
b101 +
#224310000000
0!
0'
#224320000000
1!
b110 %
1'
b110 +
#224330000000
0!
0'
#224340000000
1!
b111 %
1'
b111 +
#224350000000
0!
0'
#224360000000
1!
0$
b1000 %
1'
0*
b1000 +
#224370000000
0!
0'
#224380000000
1!
b1001 %
1'
b1001 +
#224390000000
0!
0'
#224400000000
1!
b0 %
1'
b0 +
#224410000000
0!
0'
#224420000000
1!
1$
b1 %
1'
1*
b1 +
#224430000000
0!
0'
#224440000000
1!
b10 %
1'
b10 +
#224450000000
0!
0'
#224460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#224470000000
0!
0'
#224480000000
1!
b100 %
1'
b100 +
#224490000000
0!
0'
#224500000000
1!
b101 %
1'
b101 +
#224510000000
0!
0'
#224520000000
1!
0$
b110 %
1'
0*
b110 +
#224530000000
0!
0'
#224540000000
1!
b111 %
1'
b111 +
#224550000000
0!
0'
#224560000000
1!
b1000 %
1'
b1000 +
#224570000000
0!
0'
#224580000000
1!
b1001 %
1'
b1001 +
#224590000000
0!
0'
#224600000000
1!
b0 %
1'
b0 +
#224610000000
0!
0'
#224620000000
1!
1$
b1 %
1'
1*
b1 +
#224630000000
0!
0'
#224640000000
1!
b10 %
1'
b10 +
#224650000000
0!
0'
#224660000000
1!
b11 %
1'
b11 +
#224670000000
1"
1(
#224680000000
0!
0"
b100 &
0'
0(
b100 ,
#224690000000
1!
b100 %
1'
b100 +
#224700000000
0!
0'
#224710000000
1!
b101 %
1'
b101 +
#224720000000
0!
0'
#224730000000
1!
b110 %
1'
b110 +
#224740000000
0!
0'
#224750000000
1!
b111 %
1'
b111 +
#224760000000
0!
0'
#224770000000
1!
0$
b1000 %
1'
0*
b1000 +
#224780000000
0!
0'
#224790000000
1!
b1001 %
1'
b1001 +
#224800000000
0!
0'
#224810000000
1!
b0 %
1'
b0 +
#224820000000
0!
0'
#224830000000
1!
1$
b1 %
1'
1*
b1 +
#224840000000
0!
0'
#224850000000
1!
b10 %
1'
b10 +
#224860000000
0!
0'
#224870000000
1!
b11 %
1'
b11 +
#224880000000
0!
0'
#224890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#224900000000
0!
0'
#224910000000
1!
b101 %
1'
b101 +
#224920000000
0!
0'
#224930000000
1!
0$
b110 %
1'
0*
b110 +
#224940000000
0!
0'
#224950000000
1!
b111 %
1'
b111 +
#224960000000
0!
0'
#224970000000
1!
b1000 %
1'
b1000 +
#224980000000
0!
0'
#224990000000
1!
b1001 %
1'
b1001 +
#225000000000
0!
0'
#225010000000
1!
b0 %
1'
b0 +
#225020000000
0!
0'
#225030000000
1!
1$
b1 %
1'
1*
b1 +
#225040000000
0!
0'
#225050000000
1!
b10 %
1'
b10 +
#225060000000
0!
0'
#225070000000
1!
b11 %
1'
b11 +
#225080000000
0!
0'
#225090000000
1!
b100 %
1'
b100 +
#225100000000
1"
1(
#225110000000
0!
0"
b100 &
0'
0(
b100 ,
#225120000000
1!
b101 %
1'
b101 +
#225130000000
0!
0'
#225140000000
1!
b110 %
1'
b110 +
#225150000000
0!
0'
#225160000000
1!
b111 %
1'
b111 +
#225170000000
0!
0'
#225180000000
1!
0$
b1000 %
1'
0*
b1000 +
#225190000000
0!
0'
#225200000000
1!
b1001 %
1'
b1001 +
#225210000000
0!
0'
#225220000000
1!
b0 %
1'
b0 +
#225230000000
0!
0'
#225240000000
1!
1$
b1 %
1'
1*
b1 +
#225250000000
0!
0'
#225260000000
1!
b10 %
1'
b10 +
#225270000000
0!
0'
#225280000000
1!
b11 %
1'
b11 +
#225290000000
0!
0'
#225300000000
1!
b100 %
1'
b100 +
#225310000000
0!
0'
#225320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#225330000000
0!
0'
#225340000000
1!
0$
b110 %
1'
0*
b110 +
#225350000000
0!
0'
#225360000000
1!
b111 %
1'
b111 +
#225370000000
0!
0'
#225380000000
1!
b1000 %
1'
b1000 +
#225390000000
0!
0'
#225400000000
1!
b1001 %
1'
b1001 +
#225410000000
0!
0'
#225420000000
1!
b0 %
1'
b0 +
#225430000000
0!
0'
#225440000000
1!
1$
b1 %
1'
1*
b1 +
#225450000000
0!
0'
#225460000000
1!
b10 %
1'
b10 +
#225470000000
0!
0'
#225480000000
1!
b11 %
1'
b11 +
#225490000000
0!
0'
#225500000000
1!
b100 %
1'
b100 +
#225510000000
0!
0'
#225520000000
1!
b101 %
1'
b101 +
#225530000000
1"
1(
#225540000000
0!
0"
b100 &
0'
0(
b100 ,
#225550000000
1!
b110 %
1'
b110 +
#225560000000
0!
0'
#225570000000
1!
b111 %
1'
b111 +
#225580000000
0!
0'
#225590000000
1!
0$
b1000 %
1'
0*
b1000 +
#225600000000
0!
0'
#225610000000
1!
b1001 %
1'
b1001 +
#225620000000
0!
0'
#225630000000
1!
b0 %
1'
b0 +
#225640000000
0!
0'
#225650000000
1!
1$
b1 %
1'
1*
b1 +
#225660000000
0!
0'
#225670000000
1!
b10 %
1'
b10 +
#225680000000
0!
0'
#225690000000
1!
b11 %
1'
b11 +
#225700000000
0!
0'
#225710000000
1!
b100 %
1'
b100 +
#225720000000
0!
0'
#225730000000
1!
b101 %
1'
b101 +
#225740000000
0!
0'
#225750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#225760000000
0!
0'
#225770000000
1!
b111 %
1'
b111 +
#225780000000
0!
0'
#225790000000
1!
b1000 %
1'
b1000 +
#225800000000
0!
0'
#225810000000
1!
b1001 %
1'
b1001 +
#225820000000
0!
0'
#225830000000
1!
b0 %
1'
b0 +
#225840000000
0!
0'
#225850000000
1!
1$
b1 %
1'
1*
b1 +
#225860000000
0!
0'
#225870000000
1!
b10 %
1'
b10 +
#225880000000
0!
0'
#225890000000
1!
b11 %
1'
b11 +
#225900000000
0!
0'
#225910000000
1!
b100 %
1'
b100 +
#225920000000
0!
0'
#225930000000
1!
b101 %
1'
b101 +
#225940000000
0!
0'
#225950000000
1!
0$
b110 %
1'
0*
b110 +
#225960000000
1"
1(
#225970000000
0!
0"
b100 &
0'
0(
b100 ,
#225980000000
1!
1$
b111 %
1'
1*
b111 +
#225990000000
0!
0'
#226000000000
1!
0$
b1000 %
1'
0*
b1000 +
#226010000000
0!
0'
#226020000000
1!
b1001 %
1'
b1001 +
#226030000000
0!
0'
#226040000000
1!
b0 %
1'
b0 +
#226050000000
0!
0'
#226060000000
1!
1$
b1 %
1'
1*
b1 +
#226070000000
0!
0'
#226080000000
1!
b10 %
1'
b10 +
#226090000000
0!
0'
#226100000000
1!
b11 %
1'
b11 +
#226110000000
0!
0'
#226120000000
1!
b100 %
1'
b100 +
#226130000000
0!
0'
#226140000000
1!
b101 %
1'
b101 +
#226150000000
0!
0'
#226160000000
1!
b110 %
1'
b110 +
#226170000000
0!
0'
#226180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#226190000000
0!
0'
#226200000000
1!
b1000 %
1'
b1000 +
#226210000000
0!
0'
#226220000000
1!
b1001 %
1'
b1001 +
#226230000000
0!
0'
#226240000000
1!
b0 %
1'
b0 +
#226250000000
0!
0'
#226260000000
1!
1$
b1 %
1'
1*
b1 +
#226270000000
0!
0'
#226280000000
1!
b10 %
1'
b10 +
#226290000000
0!
0'
#226300000000
1!
b11 %
1'
b11 +
#226310000000
0!
0'
#226320000000
1!
b100 %
1'
b100 +
#226330000000
0!
0'
#226340000000
1!
b101 %
1'
b101 +
#226350000000
0!
0'
#226360000000
1!
0$
b110 %
1'
0*
b110 +
#226370000000
0!
0'
#226380000000
1!
b111 %
1'
b111 +
#226390000000
1"
1(
#226400000000
0!
0"
b100 &
0'
0(
b100 ,
#226410000000
1!
b1000 %
1'
b1000 +
#226420000000
0!
0'
#226430000000
1!
b1001 %
1'
b1001 +
#226440000000
0!
0'
#226450000000
1!
b0 %
1'
b0 +
#226460000000
0!
0'
#226470000000
1!
1$
b1 %
1'
1*
b1 +
#226480000000
0!
0'
#226490000000
1!
b10 %
1'
b10 +
#226500000000
0!
0'
#226510000000
1!
b11 %
1'
b11 +
#226520000000
0!
0'
#226530000000
1!
b100 %
1'
b100 +
#226540000000
0!
0'
#226550000000
1!
b101 %
1'
b101 +
#226560000000
0!
0'
#226570000000
1!
b110 %
1'
b110 +
#226580000000
0!
0'
#226590000000
1!
b111 %
1'
b111 +
#226600000000
0!
0'
#226610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#226620000000
0!
0'
#226630000000
1!
b1001 %
1'
b1001 +
#226640000000
0!
0'
#226650000000
1!
b0 %
1'
b0 +
#226660000000
0!
0'
#226670000000
1!
1$
b1 %
1'
1*
b1 +
#226680000000
0!
0'
#226690000000
1!
b10 %
1'
b10 +
#226700000000
0!
0'
#226710000000
1!
b11 %
1'
b11 +
#226720000000
0!
0'
#226730000000
1!
b100 %
1'
b100 +
#226740000000
0!
0'
#226750000000
1!
b101 %
1'
b101 +
#226760000000
0!
0'
#226770000000
1!
0$
b110 %
1'
0*
b110 +
#226780000000
0!
0'
#226790000000
1!
b111 %
1'
b111 +
#226800000000
0!
0'
#226810000000
1!
b1000 %
1'
b1000 +
#226820000000
1"
1(
#226830000000
0!
0"
b100 &
0'
0(
b100 ,
#226840000000
1!
b1001 %
1'
b1001 +
#226850000000
0!
0'
#226860000000
1!
b0 %
1'
b0 +
#226870000000
0!
0'
#226880000000
1!
1$
b1 %
1'
1*
b1 +
#226890000000
0!
0'
#226900000000
1!
b10 %
1'
b10 +
#226910000000
0!
0'
#226920000000
1!
b11 %
1'
b11 +
#226930000000
0!
0'
#226940000000
1!
b100 %
1'
b100 +
#226950000000
0!
0'
#226960000000
1!
b101 %
1'
b101 +
#226970000000
0!
0'
#226980000000
1!
b110 %
1'
b110 +
#226990000000
0!
0'
#227000000000
1!
b111 %
1'
b111 +
#227010000000
0!
0'
#227020000000
1!
0$
b1000 %
1'
0*
b1000 +
#227030000000
0!
0'
#227040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#227050000000
0!
0'
#227060000000
1!
b0 %
1'
b0 +
#227070000000
0!
0'
#227080000000
1!
1$
b1 %
1'
1*
b1 +
#227090000000
0!
0'
#227100000000
1!
b10 %
1'
b10 +
#227110000000
0!
0'
#227120000000
1!
b11 %
1'
b11 +
#227130000000
0!
0'
#227140000000
1!
b100 %
1'
b100 +
#227150000000
0!
0'
#227160000000
1!
b101 %
1'
b101 +
#227170000000
0!
0'
#227180000000
1!
0$
b110 %
1'
0*
b110 +
#227190000000
0!
0'
#227200000000
1!
b111 %
1'
b111 +
#227210000000
0!
0'
#227220000000
1!
b1000 %
1'
b1000 +
#227230000000
0!
0'
#227240000000
1!
b1001 %
1'
b1001 +
#227250000000
1"
1(
#227260000000
0!
0"
b100 &
0'
0(
b100 ,
#227270000000
1!
b0 %
1'
b0 +
#227280000000
0!
0'
#227290000000
1!
1$
b1 %
1'
1*
b1 +
#227300000000
0!
0'
#227310000000
1!
b10 %
1'
b10 +
#227320000000
0!
0'
#227330000000
1!
b11 %
1'
b11 +
#227340000000
0!
0'
#227350000000
1!
b100 %
1'
b100 +
#227360000000
0!
0'
#227370000000
1!
b101 %
1'
b101 +
#227380000000
0!
0'
#227390000000
1!
b110 %
1'
b110 +
#227400000000
0!
0'
#227410000000
1!
b111 %
1'
b111 +
#227420000000
0!
0'
#227430000000
1!
0$
b1000 %
1'
0*
b1000 +
#227440000000
0!
0'
#227450000000
1!
b1001 %
1'
b1001 +
#227460000000
0!
0'
#227470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#227480000000
0!
0'
#227490000000
1!
1$
b1 %
1'
1*
b1 +
#227500000000
0!
0'
#227510000000
1!
b10 %
1'
b10 +
#227520000000
0!
0'
#227530000000
1!
b11 %
1'
b11 +
#227540000000
0!
0'
#227550000000
1!
b100 %
1'
b100 +
#227560000000
0!
0'
#227570000000
1!
b101 %
1'
b101 +
#227580000000
0!
0'
#227590000000
1!
0$
b110 %
1'
0*
b110 +
#227600000000
0!
0'
#227610000000
1!
b111 %
1'
b111 +
#227620000000
0!
0'
#227630000000
1!
b1000 %
1'
b1000 +
#227640000000
0!
0'
#227650000000
1!
b1001 %
1'
b1001 +
#227660000000
0!
0'
#227670000000
1!
b0 %
1'
b0 +
#227680000000
1"
1(
#227690000000
0!
0"
b100 &
0'
0(
b100 ,
#227700000000
1!
1$
b1 %
1'
1*
b1 +
#227710000000
0!
0'
#227720000000
1!
b10 %
1'
b10 +
#227730000000
0!
0'
#227740000000
1!
b11 %
1'
b11 +
#227750000000
0!
0'
#227760000000
1!
b100 %
1'
b100 +
#227770000000
0!
0'
#227780000000
1!
b101 %
1'
b101 +
#227790000000
0!
0'
#227800000000
1!
b110 %
1'
b110 +
#227810000000
0!
0'
#227820000000
1!
b111 %
1'
b111 +
#227830000000
0!
0'
#227840000000
1!
0$
b1000 %
1'
0*
b1000 +
#227850000000
0!
0'
#227860000000
1!
b1001 %
1'
b1001 +
#227870000000
0!
0'
#227880000000
1!
b0 %
1'
b0 +
#227890000000
0!
0'
#227900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#227910000000
0!
0'
#227920000000
1!
b10 %
1'
b10 +
#227930000000
0!
0'
#227940000000
1!
b11 %
1'
b11 +
#227950000000
0!
0'
#227960000000
1!
b100 %
1'
b100 +
#227970000000
0!
0'
#227980000000
1!
b101 %
1'
b101 +
#227990000000
0!
0'
#228000000000
1!
0$
b110 %
1'
0*
b110 +
#228010000000
0!
0'
#228020000000
1!
b111 %
1'
b111 +
#228030000000
0!
0'
#228040000000
1!
b1000 %
1'
b1000 +
#228050000000
0!
0'
#228060000000
1!
b1001 %
1'
b1001 +
#228070000000
0!
0'
#228080000000
1!
b0 %
1'
b0 +
#228090000000
0!
0'
#228100000000
1!
1$
b1 %
1'
1*
b1 +
#228110000000
1"
1(
#228120000000
0!
0"
b100 &
0'
0(
b100 ,
#228130000000
1!
b10 %
1'
b10 +
#228140000000
0!
0'
#228150000000
1!
b11 %
1'
b11 +
#228160000000
0!
0'
#228170000000
1!
b100 %
1'
b100 +
#228180000000
0!
0'
#228190000000
1!
b101 %
1'
b101 +
#228200000000
0!
0'
#228210000000
1!
b110 %
1'
b110 +
#228220000000
0!
0'
#228230000000
1!
b111 %
1'
b111 +
#228240000000
0!
0'
#228250000000
1!
0$
b1000 %
1'
0*
b1000 +
#228260000000
0!
0'
#228270000000
1!
b1001 %
1'
b1001 +
#228280000000
0!
0'
#228290000000
1!
b0 %
1'
b0 +
#228300000000
0!
0'
#228310000000
1!
1$
b1 %
1'
1*
b1 +
#228320000000
0!
0'
#228330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#228340000000
0!
0'
#228350000000
1!
b11 %
1'
b11 +
#228360000000
0!
0'
#228370000000
1!
b100 %
1'
b100 +
#228380000000
0!
0'
#228390000000
1!
b101 %
1'
b101 +
#228400000000
0!
0'
#228410000000
1!
0$
b110 %
1'
0*
b110 +
#228420000000
0!
0'
#228430000000
1!
b111 %
1'
b111 +
#228440000000
0!
0'
#228450000000
1!
b1000 %
1'
b1000 +
#228460000000
0!
0'
#228470000000
1!
b1001 %
1'
b1001 +
#228480000000
0!
0'
#228490000000
1!
b0 %
1'
b0 +
#228500000000
0!
0'
#228510000000
1!
1$
b1 %
1'
1*
b1 +
#228520000000
0!
0'
#228530000000
1!
b10 %
1'
b10 +
#228540000000
1"
1(
#228550000000
0!
0"
b100 &
0'
0(
b100 ,
#228560000000
1!
b11 %
1'
b11 +
#228570000000
0!
0'
#228580000000
1!
b100 %
1'
b100 +
#228590000000
0!
0'
#228600000000
1!
b101 %
1'
b101 +
#228610000000
0!
0'
#228620000000
1!
b110 %
1'
b110 +
#228630000000
0!
0'
#228640000000
1!
b111 %
1'
b111 +
#228650000000
0!
0'
#228660000000
1!
0$
b1000 %
1'
0*
b1000 +
#228670000000
0!
0'
#228680000000
1!
b1001 %
1'
b1001 +
#228690000000
0!
0'
#228700000000
1!
b0 %
1'
b0 +
#228710000000
0!
0'
#228720000000
1!
1$
b1 %
1'
1*
b1 +
#228730000000
0!
0'
#228740000000
1!
b10 %
1'
b10 +
#228750000000
0!
0'
#228760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#228770000000
0!
0'
#228780000000
1!
b100 %
1'
b100 +
#228790000000
0!
0'
#228800000000
1!
b101 %
1'
b101 +
#228810000000
0!
0'
#228820000000
1!
0$
b110 %
1'
0*
b110 +
#228830000000
0!
0'
#228840000000
1!
b111 %
1'
b111 +
#228850000000
0!
0'
#228860000000
1!
b1000 %
1'
b1000 +
#228870000000
0!
0'
#228880000000
1!
b1001 %
1'
b1001 +
#228890000000
0!
0'
#228900000000
1!
b0 %
1'
b0 +
#228910000000
0!
0'
#228920000000
1!
1$
b1 %
1'
1*
b1 +
#228930000000
0!
0'
#228940000000
1!
b10 %
1'
b10 +
#228950000000
0!
0'
#228960000000
1!
b11 %
1'
b11 +
#228970000000
1"
1(
#228980000000
0!
0"
b100 &
0'
0(
b100 ,
#228990000000
1!
b100 %
1'
b100 +
#229000000000
0!
0'
#229010000000
1!
b101 %
1'
b101 +
#229020000000
0!
0'
#229030000000
1!
b110 %
1'
b110 +
#229040000000
0!
0'
#229050000000
1!
b111 %
1'
b111 +
#229060000000
0!
0'
#229070000000
1!
0$
b1000 %
1'
0*
b1000 +
#229080000000
0!
0'
#229090000000
1!
b1001 %
1'
b1001 +
#229100000000
0!
0'
#229110000000
1!
b0 %
1'
b0 +
#229120000000
0!
0'
#229130000000
1!
1$
b1 %
1'
1*
b1 +
#229140000000
0!
0'
#229150000000
1!
b10 %
1'
b10 +
#229160000000
0!
0'
#229170000000
1!
b11 %
1'
b11 +
#229180000000
0!
0'
#229190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#229200000000
0!
0'
#229210000000
1!
b101 %
1'
b101 +
#229220000000
0!
0'
#229230000000
1!
0$
b110 %
1'
0*
b110 +
#229240000000
0!
0'
#229250000000
1!
b111 %
1'
b111 +
#229260000000
0!
0'
#229270000000
1!
b1000 %
1'
b1000 +
#229280000000
0!
0'
#229290000000
1!
b1001 %
1'
b1001 +
#229300000000
0!
0'
#229310000000
1!
b0 %
1'
b0 +
#229320000000
0!
0'
#229330000000
1!
1$
b1 %
1'
1*
b1 +
#229340000000
0!
0'
#229350000000
1!
b10 %
1'
b10 +
#229360000000
0!
0'
#229370000000
1!
b11 %
1'
b11 +
#229380000000
0!
0'
#229390000000
1!
b100 %
1'
b100 +
#229400000000
1"
1(
#229410000000
0!
0"
b100 &
0'
0(
b100 ,
#229420000000
1!
b101 %
1'
b101 +
#229430000000
0!
0'
#229440000000
1!
b110 %
1'
b110 +
#229450000000
0!
0'
#229460000000
1!
b111 %
1'
b111 +
#229470000000
0!
0'
#229480000000
1!
0$
b1000 %
1'
0*
b1000 +
#229490000000
0!
0'
#229500000000
1!
b1001 %
1'
b1001 +
#229510000000
0!
0'
#229520000000
1!
b0 %
1'
b0 +
#229530000000
0!
0'
#229540000000
1!
1$
b1 %
1'
1*
b1 +
#229550000000
0!
0'
#229560000000
1!
b10 %
1'
b10 +
#229570000000
0!
0'
#229580000000
1!
b11 %
1'
b11 +
#229590000000
0!
0'
#229600000000
1!
b100 %
1'
b100 +
#229610000000
0!
0'
#229620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#229630000000
0!
0'
#229640000000
1!
0$
b110 %
1'
0*
b110 +
#229650000000
0!
0'
#229660000000
1!
b111 %
1'
b111 +
#229670000000
0!
0'
#229680000000
1!
b1000 %
1'
b1000 +
#229690000000
0!
0'
#229700000000
1!
b1001 %
1'
b1001 +
#229710000000
0!
0'
#229720000000
1!
b0 %
1'
b0 +
#229730000000
0!
0'
#229740000000
1!
1$
b1 %
1'
1*
b1 +
#229750000000
0!
0'
#229760000000
1!
b10 %
1'
b10 +
#229770000000
0!
0'
#229780000000
1!
b11 %
1'
b11 +
#229790000000
0!
0'
#229800000000
1!
b100 %
1'
b100 +
#229810000000
0!
0'
#229820000000
1!
b101 %
1'
b101 +
#229830000000
1"
1(
#229840000000
0!
0"
b100 &
0'
0(
b100 ,
#229850000000
1!
b110 %
1'
b110 +
#229860000000
0!
0'
#229870000000
1!
b111 %
1'
b111 +
#229880000000
0!
0'
#229890000000
1!
0$
b1000 %
1'
0*
b1000 +
#229900000000
0!
0'
#229910000000
1!
b1001 %
1'
b1001 +
#229920000000
0!
0'
#229930000000
1!
b0 %
1'
b0 +
#229940000000
0!
0'
#229950000000
1!
1$
b1 %
1'
1*
b1 +
#229960000000
0!
0'
#229970000000
1!
b10 %
1'
b10 +
#229980000000
0!
0'
#229990000000
1!
b11 %
1'
b11 +
#230000000000
0!
0'
#230010000000
1!
b100 %
1'
b100 +
#230020000000
0!
0'
#230030000000
1!
b101 %
1'
b101 +
#230040000000
0!
0'
#230050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#230060000000
0!
0'
#230070000000
1!
b111 %
1'
b111 +
#230080000000
0!
0'
#230090000000
1!
b1000 %
1'
b1000 +
#230100000000
0!
0'
#230110000000
1!
b1001 %
1'
b1001 +
#230120000000
0!
0'
#230130000000
1!
b0 %
1'
b0 +
#230140000000
0!
0'
#230150000000
1!
1$
b1 %
1'
1*
b1 +
#230160000000
0!
0'
#230170000000
1!
b10 %
1'
b10 +
#230180000000
0!
0'
#230190000000
1!
b11 %
1'
b11 +
#230200000000
0!
0'
#230210000000
1!
b100 %
1'
b100 +
#230220000000
0!
0'
#230230000000
1!
b101 %
1'
b101 +
#230240000000
0!
0'
#230250000000
1!
0$
b110 %
1'
0*
b110 +
#230260000000
1"
1(
#230270000000
0!
0"
b100 &
0'
0(
b100 ,
#230280000000
1!
1$
b111 %
1'
1*
b111 +
#230290000000
0!
0'
#230300000000
1!
0$
b1000 %
1'
0*
b1000 +
#230310000000
0!
0'
#230320000000
1!
b1001 %
1'
b1001 +
#230330000000
0!
0'
#230340000000
1!
b0 %
1'
b0 +
#230350000000
0!
0'
#230360000000
1!
1$
b1 %
1'
1*
b1 +
#230370000000
0!
0'
#230380000000
1!
b10 %
1'
b10 +
#230390000000
0!
0'
#230400000000
1!
b11 %
1'
b11 +
#230410000000
0!
0'
#230420000000
1!
b100 %
1'
b100 +
#230430000000
0!
0'
#230440000000
1!
b101 %
1'
b101 +
#230450000000
0!
0'
#230460000000
1!
b110 %
1'
b110 +
#230470000000
0!
0'
#230480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#230490000000
0!
0'
#230500000000
1!
b1000 %
1'
b1000 +
#230510000000
0!
0'
#230520000000
1!
b1001 %
1'
b1001 +
#230530000000
0!
0'
#230540000000
1!
b0 %
1'
b0 +
#230550000000
0!
0'
#230560000000
1!
1$
b1 %
1'
1*
b1 +
#230570000000
0!
0'
#230580000000
1!
b10 %
1'
b10 +
#230590000000
0!
0'
#230600000000
1!
b11 %
1'
b11 +
#230610000000
0!
0'
#230620000000
1!
b100 %
1'
b100 +
#230630000000
0!
0'
#230640000000
1!
b101 %
1'
b101 +
#230650000000
0!
0'
#230660000000
1!
0$
b110 %
1'
0*
b110 +
#230670000000
0!
0'
#230680000000
1!
b111 %
1'
b111 +
#230690000000
1"
1(
#230700000000
0!
0"
b100 &
0'
0(
b100 ,
#230710000000
1!
b1000 %
1'
b1000 +
#230720000000
0!
0'
#230730000000
1!
b1001 %
1'
b1001 +
#230740000000
0!
0'
#230750000000
1!
b0 %
1'
b0 +
#230760000000
0!
0'
#230770000000
1!
1$
b1 %
1'
1*
b1 +
#230780000000
0!
0'
#230790000000
1!
b10 %
1'
b10 +
#230800000000
0!
0'
#230810000000
1!
b11 %
1'
b11 +
#230820000000
0!
0'
#230830000000
1!
b100 %
1'
b100 +
#230840000000
0!
0'
#230850000000
1!
b101 %
1'
b101 +
#230860000000
0!
0'
#230870000000
1!
b110 %
1'
b110 +
#230880000000
0!
0'
#230890000000
1!
b111 %
1'
b111 +
#230900000000
0!
0'
#230910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#230920000000
0!
0'
#230930000000
1!
b1001 %
1'
b1001 +
#230940000000
0!
0'
#230950000000
1!
b0 %
1'
b0 +
#230960000000
0!
0'
#230970000000
1!
1$
b1 %
1'
1*
b1 +
#230980000000
0!
0'
#230990000000
1!
b10 %
1'
b10 +
#231000000000
0!
0'
#231010000000
1!
b11 %
1'
b11 +
#231020000000
0!
0'
#231030000000
1!
b100 %
1'
b100 +
#231040000000
0!
0'
#231050000000
1!
b101 %
1'
b101 +
#231060000000
0!
0'
#231070000000
1!
0$
b110 %
1'
0*
b110 +
#231080000000
0!
0'
#231090000000
1!
b111 %
1'
b111 +
#231100000000
0!
0'
#231110000000
1!
b1000 %
1'
b1000 +
#231120000000
1"
1(
#231130000000
0!
0"
b100 &
0'
0(
b100 ,
#231140000000
1!
b1001 %
1'
b1001 +
#231150000000
0!
0'
#231160000000
1!
b0 %
1'
b0 +
#231170000000
0!
0'
#231180000000
1!
1$
b1 %
1'
1*
b1 +
#231190000000
0!
0'
#231200000000
1!
b10 %
1'
b10 +
#231210000000
0!
0'
#231220000000
1!
b11 %
1'
b11 +
#231230000000
0!
0'
#231240000000
1!
b100 %
1'
b100 +
#231250000000
0!
0'
#231260000000
1!
b101 %
1'
b101 +
#231270000000
0!
0'
#231280000000
1!
b110 %
1'
b110 +
#231290000000
0!
0'
#231300000000
1!
b111 %
1'
b111 +
#231310000000
0!
0'
#231320000000
1!
0$
b1000 %
1'
0*
b1000 +
#231330000000
0!
0'
#231340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#231350000000
0!
0'
#231360000000
1!
b0 %
1'
b0 +
#231370000000
0!
0'
#231380000000
1!
1$
b1 %
1'
1*
b1 +
#231390000000
0!
0'
#231400000000
1!
b10 %
1'
b10 +
#231410000000
0!
0'
#231420000000
1!
b11 %
1'
b11 +
#231430000000
0!
0'
#231440000000
1!
b100 %
1'
b100 +
#231450000000
0!
0'
#231460000000
1!
b101 %
1'
b101 +
#231470000000
0!
0'
#231480000000
1!
0$
b110 %
1'
0*
b110 +
#231490000000
0!
0'
#231500000000
1!
b111 %
1'
b111 +
#231510000000
0!
0'
#231520000000
1!
b1000 %
1'
b1000 +
#231530000000
0!
0'
#231540000000
1!
b1001 %
1'
b1001 +
#231550000000
1"
1(
#231560000000
0!
0"
b100 &
0'
0(
b100 ,
#231570000000
1!
b0 %
1'
b0 +
#231580000000
0!
0'
#231590000000
1!
1$
b1 %
1'
1*
b1 +
#231600000000
0!
0'
#231610000000
1!
b10 %
1'
b10 +
#231620000000
0!
0'
#231630000000
1!
b11 %
1'
b11 +
#231640000000
0!
0'
#231650000000
1!
b100 %
1'
b100 +
#231660000000
0!
0'
#231670000000
1!
b101 %
1'
b101 +
#231680000000
0!
0'
#231690000000
1!
b110 %
1'
b110 +
#231700000000
0!
0'
#231710000000
1!
b111 %
1'
b111 +
#231720000000
0!
0'
#231730000000
1!
0$
b1000 %
1'
0*
b1000 +
#231740000000
0!
0'
#231750000000
1!
b1001 %
1'
b1001 +
#231760000000
0!
0'
#231770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#231780000000
0!
0'
#231790000000
1!
1$
b1 %
1'
1*
b1 +
#231800000000
0!
0'
#231810000000
1!
b10 %
1'
b10 +
#231820000000
0!
0'
#231830000000
1!
b11 %
1'
b11 +
#231840000000
0!
0'
#231850000000
1!
b100 %
1'
b100 +
#231860000000
0!
0'
#231870000000
1!
b101 %
1'
b101 +
#231880000000
0!
0'
#231890000000
1!
0$
b110 %
1'
0*
b110 +
#231900000000
0!
0'
#231910000000
1!
b111 %
1'
b111 +
#231920000000
0!
0'
#231930000000
1!
b1000 %
1'
b1000 +
#231940000000
0!
0'
#231950000000
1!
b1001 %
1'
b1001 +
#231960000000
0!
0'
#231970000000
1!
b0 %
1'
b0 +
#231980000000
1"
1(
#231990000000
0!
0"
b100 &
0'
0(
b100 ,
#232000000000
1!
1$
b1 %
1'
1*
b1 +
#232010000000
0!
0'
#232020000000
1!
b10 %
1'
b10 +
#232030000000
0!
0'
#232040000000
1!
b11 %
1'
b11 +
#232050000000
0!
0'
#232060000000
1!
b100 %
1'
b100 +
#232070000000
0!
0'
#232080000000
1!
b101 %
1'
b101 +
#232090000000
0!
0'
#232100000000
1!
b110 %
1'
b110 +
#232110000000
0!
0'
#232120000000
1!
b111 %
1'
b111 +
#232130000000
0!
0'
#232140000000
1!
0$
b1000 %
1'
0*
b1000 +
#232150000000
0!
0'
#232160000000
1!
b1001 %
1'
b1001 +
#232170000000
0!
0'
#232180000000
1!
b0 %
1'
b0 +
#232190000000
0!
0'
#232200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#232210000000
0!
0'
#232220000000
1!
b10 %
1'
b10 +
#232230000000
0!
0'
#232240000000
1!
b11 %
1'
b11 +
#232250000000
0!
0'
#232260000000
1!
b100 %
1'
b100 +
#232270000000
0!
0'
#232280000000
1!
b101 %
1'
b101 +
#232290000000
0!
0'
#232300000000
1!
0$
b110 %
1'
0*
b110 +
#232310000000
0!
0'
#232320000000
1!
b111 %
1'
b111 +
#232330000000
0!
0'
#232340000000
1!
b1000 %
1'
b1000 +
#232350000000
0!
0'
#232360000000
1!
b1001 %
1'
b1001 +
#232370000000
0!
0'
#232380000000
1!
b0 %
1'
b0 +
#232390000000
0!
0'
#232400000000
1!
1$
b1 %
1'
1*
b1 +
#232410000000
1"
1(
#232420000000
0!
0"
b100 &
0'
0(
b100 ,
#232430000000
1!
b10 %
1'
b10 +
#232440000000
0!
0'
#232450000000
1!
b11 %
1'
b11 +
#232460000000
0!
0'
#232470000000
1!
b100 %
1'
b100 +
#232480000000
0!
0'
#232490000000
1!
b101 %
1'
b101 +
#232500000000
0!
0'
#232510000000
1!
b110 %
1'
b110 +
#232520000000
0!
0'
#232530000000
1!
b111 %
1'
b111 +
#232540000000
0!
0'
#232550000000
1!
0$
b1000 %
1'
0*
b1000 +
#232560000000
0!
0'
#232570000000
1!
b1001 %
1'
b1001 +
#232580000000
0!
0'
#232590000000
1!
b0 %
1'
b0 +
#232600000000
0!
0'
#232610000000
1!
1$
b1 %
1'
1*
b1 +
#232620000000
0!
0'
#232630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#232640000000
0!
0'
#232650000000
1!
b11 %
1'
b11 +
#232660000000
0!
0'
#232670000000
1!
b100 %
1'
b100 +
#232680000000
0!
0'
#232690000000
1!
b101 %
1'
b101 +
#232700000000
0!
0'
#232710000000
1!
0$
b110 %
1'
0*
b110 +
#232720000000
0!
0'
#232730000000
1!
b111 %
1'
b111 +
#232740000000
0!
0'
#232750000000
1!
b1000 %
1'
b1000 +
#232760000000
0!
0'
#232770000000
1!
b1001 %
1'
b1001 +
#232780000000
0!
0'
#232790000000
1!
b0 %
1'
b0 +
#232800000000
0!
0'
#232810000000
1!
1$
b1 %
1'
1*
b1 +
#232820000000
0!
0'
#232830000000
1!
b10 %
1'
b10 +
#232840000000
1"
1(
#232850000000
0!
0"
b100 &
0'
0(
b100 ,
#232860000000
1!
b11 %
1'
b11 +
#232870000000
0!
0'
#232880000000
1!
b100 %
1'
b100 +
#232890000000
0!
0'
#232900000000
1!
b101 %
1'
b101 +
#232910000000
0!
0'
#232920000000
1!
b110 %
1'
b110 +
#232930000000
0!
0'
#232940000000
1!
b111 %
1'
b111 +
#232950000000
0!
0'
#232960000000
1!
0$
b1000 %
1'
0*
b1000 +
#232970000000
0!
0'
#232980000000
1!
b1001 %
1'
b1001 +
#232990000000
0!
0'
#233000000000
1!
b0 %
1'
b0 +
#233010000000
0!
0'
#233020000000
1!
1$
b1 %
1'
1*
b1 +
#233030000000
0!
0'
#233040000000
1!
b10 %
1'
b10 +
#233050000000
0!
0'
#233060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#233070000000
0!
0'
#233080000000
1!
b100 %
1'
b100 +
#233090000000
0!
0'
#233100000000
1!
b101 %
1'
b101 +
#233110000000
0!
0'
#233120000000
1!
0$
b110 %
1'
0*
b110 +
#233130000000
0!
0'
#233140000000
1!
b111 %
1'
b111 +
#233150000000
0!
0'
#233160000000
1!
b1000 %
1'
b1000 +
#233170000000
0!
0'
#233180000000
1!
b1001 %
1'
b1001 +
#233190000000
0!
0'
#233200000000
1!
b0 %
1'
b0 +
#233210000000
0!
0'
#233220000000
1!
1$
b1 %
1'
1*
b1 +
#233230000000
0!
0'
#233240000000
1!
b10 %
1'
b10 +
#233250000000
0!
0'
#233260000000
1!
b11 %
1'
b11 +
#233270000000
1"
1(
#233280000000
0!
0"
b100 &
0'
0(
b100 ,
#233290000000
1!
b100 %
1'
b100 +
#233300000000
0!
0'
#233310000000
1!
b101 %
1'
b101 +
#233320000000
0!
0'
#233330000000
1!
b110 %
1'
b110 +
#233340000000
0!
0'
#233350000000
1!
b111 %
1'
b111 +
#233360000000
0!
0'
#233370000000
1!
0$
b1000 %
1'
0*
b1000 +
#233380000000
0!
0'
#233390000000
1!
b1001 %
1'
b1001 +
#233400000000
0!
0'
#233410000000
1!
b0 %
1'
b0 +
#233420000000
0!
0'
#233430000000
1!
1$
b1 %
1'
1*
b1 +
#233440000000
0!
0'
#233450000000
1!
b10 %
1'
b10 +
#233460000000
0!
0'
#233470000000
1!
b11 %
1'
b11 +
#233480000000
0!
0'
#233490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#233500000000
0!
0'
#233510000000
1!
b101 %
1'
b101 +
#233520000000
0!
0'
#233530000000
1!
0$
b110 %
1'
0*
b110 +
#233540000000
0!
0'
#233550000000
1!
b111 %
1'
b111 +
#233560000000
0!
0'
#233570000000
1!
b1000 %
1'
b1000 +
#233580000000
0!
0'
#233590000000
1!
b1001 %
1'
b1001 +
#233600000000
0!
0'
#233610000000
1!
b0 %
1'
b0 +
#233620000000
0!
0'
#233630000000
1!
1$
b1 %
1'
1*
b1 +
#233640000000
0!
0'
#233650000000
1!
b10 %
1'
b10 +
#233660000000
0!
0'
#233670000000
1!
b11 %
1'
b11 +
#233680000000
0!
0'
#233690000000
1!
b100 %
1'
b100 +
#233700000000
1"
1(
#233710000000
0!
0"
b100 &
0'
0(
b100 ,
#233720000000
1!
b101 %
1'
b101 +
#233730000000
0!
0'
#233740000000
1!
b110 %
1'
b110 +
#233750000000
0!
0'
#233760000000
1!
b111 %
1'
b111 +
#233770000000
0!
0'
#233780000000
1!
0$
b1000 %
1'
0*
b1000 +
#233790000000
0!
0'
#233800000000
1!
b1001 %
1'
b1001 +
#233810000000
0!
0'
#233820000000
1!
b0 %
1'
b0 +
#233830000000
0!
0'
#233840000000
1!
1$
b1 %
1'
1*
b1 +
#233850000000
0!
0'
#233860000000
1!
b10 %
1'
b10 +
#233870000000
0!
0'
#233880000000
1!
b11 %
1'
b11 +
#233890000000
0!
0'
#233900000000
1!
b100 %
1'
b100 +
#233910000000
0!
0'
#233920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#233930000000
0!
0'
#233940000000
1!
0$
b110 %
1'
0*
b110 +
#233950000000
0!
0'
#233960000000
1!
b111 %
1'
b111 +
#233970000000
0!
0'
#233980000000
1!
b1000 %
1'
b1000 +
#233990000000
0!
0'
#234000000000
1!
b1001 %
1'
b1001 +
#234010000000
0!
0'
#234020000000
1!
b0 %
1'
b0 +
#234030000000
0!
0'
#234040000000
1!
1$
b1 %
1'
1*
b1 +
#234050000000
0!
0'
#234060000000
1!
b10 %
1'
b10 +
#234070000000
0!
0'
#234080000000
1!
b11 %
1'
b11 +
#234090000000
0!
0'
#234100000000
1!
b100 %
1'
b100 +
#234110000000
0!
0'
#234120000000
1!
b101 %
1'
b101 +
#234130000000
1"
1(
#234140000000
0!
0"
b100 &
0'
0(
b100 ,
#234150000000
1!
b110 %
1'
b110 +
#234160000000
0!
0'
#234170000000
1!
b111 %
1'
b111 +
#234180000000
0!
0'
#234190000000
1!
0$
b1000 %
1'
0*
b1000 +
#234200000000
0!
0'
#234210000000
1!
b1001 %
1'
b1001 +
#234220000000
0!
0'
#234230000000
1!
b0 %
1'
b0 +
#234240000000
0!
0'
#234250000000
1!
1$
b1 %
1'
1*
b1 +
#234260000000
0!
0'
#234270000000
1!
b10 %
1'
b10 +
#234280000000
0!
0'
#234290000000
1!
b11 %
1'
b11 +
#234300000000
0!
0'
#234310000000
1!
b100 %
1'
b100 +
#234320000000
0!
0'
#234330000000
1!
b101 %
1'
b101 +
#234340000000
0!
0'
#234350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#234360000000
0!
0'
#234370000000
1!
b111 %
1'
b111 +
#234380000000
0!
0'
#234390000000
1!
b1000 %
1'
b1000 +
#234400000000
0!
0'
#234410000000
1!
b1001 %
1'
b1001 +
#234420000000
0!
0'
#234430000000
1!
b0 %
1'
b0 +
#234440000000
0!
0'
#234450000000
1!
1$
b1 %
1'
1*
b1 +
#234460000000
0!
0'
#234470000000
1!
b10 %
1'
b10 +
#234480000000
0!
0'
#234490000000
1!
b11 %
1'
b11 +
#234500000000
0!
0'
#234510000000
1!
b100 %
1'
b100 +
#234520000000
0!
0'
#234530000000
1!
b101 %
1'
b101 +
#234540000000
0!
0'
#234550000000
1!
0$
b110 %
1'
0*
b110 +
#234560000000
1"
1(
#234570000000
0!
0"
b100 &
0'
0(
b100 ,
#234580000000
1!
1$
b111 %
1'
1*
b111 +
#234590000000
0!
0'
#234600000000
1!
0$
b1000 %
1'
0*
b1000 +
#234610000000
0!
0'
#234620000000
1!
b1001 %
1'
b1001 +
#234630000000
0!
0'
#234640000000
1!
b0 %
1'
b0 +
#234650000000
0!
0'
#234660000000
1!
1$
b1 %
1'
1*
b1 +
#234670000000
0!
0'
#234680000000
1!
b10 %
1'
b10 +
#234690000000
0!
0'
#234700000000
1!
b11 %
1'
b11 +
#234710000000
0!
0'
#234720000000
1!
b100 %
1'
b100 +
#234730000000
0!
0'
#234740000000
1!
b101 %
1'
b101 +
#234750000000
0!
0'
#234760000000
1!
b110 %
1'
b110 +
#234770000000
0!
0'
#234780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#234790000000
0!
0'
#234800000000
1!
b1000 %
1'
b1000 +
#234810000000
0!
0'
#234820000000
1!
b1001 %
1'
b1001 +
#234830000000
0!
0'
#234840000000
1!
b0 %
1'
b0 +
#234850000000
0!
0'
#234860000000
1!
1$
b1 %
1'
1*
b1 +
#234870000000
0!
0'
#234880000000
1!
b10 %
1'
b10 +
#234890000000
0!
0'
#234900000000
1!
b11 %
1'
b11 +
#234910000000
0!
0'
#234920000000
1!
b100 %
1'
b100 +
#234930000000
0!
0'
#234940000000
1!
b101 %
1'
b101 +
#234950000000
0!
0'
#234960000000
1!
0$
b110 %
1'
0*
b110 +
#234970000000
0!
0'
#234980000000
1!
b111 %
1'
b111 +
#234990000000
1"
1(
#235000000000
0!
0"
b100 &
0'
0(
b100 ,
#235010000000
1!
b1000 %
1'
b1000 +
#235020000000
0!
0'
#235030000000
1!
b1001 %
1'
b1001 +
#235040000000
0!
0'
#235050000000
1!
b0 %
1'
b0 +
#235060000000
0!
0'
#235070000000
1!
1$
b1 %
1'
1*
b1 +
#235080000000
0!
0'
#235090000000
1!
b10 %
1'
b10 +
#235100000000
0!
0'
#235110000000
1!
b11 %
1'
b11 +
#235120000000
0!
0'
#235130000000
1!
b100 %
1'
b100 +
#235140000000
0!
0'
#235150000000
1!
b101 %
1'
b101 +
#235160000000
0!
0'
#235170000000
1!
b110 %
1'
b110 +
#235180000000
0!
0'
#235190000000
1!
b111 %
1'
b111 +
#235200000000
0!
0'
#235210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#235220000000
0!
0'
#235230000000
1!
b1001 %
1'
b1001 +
#235240000000
0!
0'
#235250000000
1!
b0 %
1'
b0 +
#235260000000
0!
0'
#235270000000
1!
1$
b1 %
1'
1*
b1 +
#235280000000
0!
0'
#235290000000
1!
b10 %
1'
b10 +
#235300000000
0!
0'
#235310000000
1!
b11 %
1'
b11 +
#235320000000
0!
0'
#235330000000
1!
b100 %
1'
b100 +
#235340000000
0!
0'
#235350000000
1!
b101 %
1'
b101 +
#235360000000
0!
0'
#235370000000
1!
0$
b110 %
1'
0*
b110 +
#235380000000
0!
0'
#235390000000
1!
b111 %
1'
b111 +
#235400000000
0!
0'
#235410000000
1!
b1000 %
1'
b1000 +
#235420000000
1"
1(
#235430000000
0!
0"
b100 &
0'
0(
b100 ,
#235440000000
1!
b1001 %
1'
b1001 +
#235450000000
0!
0'
#235460000000
1!
b0 %
1'
b0 +
#235470000000
0!
0'
#235480000000
1!
1$
b1 %
1'
1*
b1 +
#235490000000
0!
0'
#235500000000
1!
b10 %
1'
b10 +
#235510000000
0!
0'
#235520000000
1!
b11 %
1'
b11 +
#235530000000
0!
0'
#235540000000
1!
b100 %
1'
b100 +
#235550000000
0!
0'
#235560000000
1!
b101 %
1'
b101 +
#235570000000
0!
0'
#235580000000
1!
b110 %
1'
b110 +
#235590000000
0!
0'
#235600000000
1!
b111 %
1'
b111 +
#235610000000
0!
0'
#235620000000
1!
0$
b1000 %
1'
0*
b1000 +
#235630000000
0!
0'
#235640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#235650000000
0!
0'
#235660000000
1!
b0 %
1'
b0 +
#235670000000
0!
0'
#235680000000
1!
1$
b1 %
1'
1*
b1 +
#235690000000
0!
0'
#235700000000
1!
b10 %
1'
b10 +
#235710000000
0!
0'
#235720000000
1!
b11 %
1'
b11 +
#235730000000
0!
0'
#235740000000
1!
b100 %
1'
b100 +
#235750000000
0!
0'
#235760000000
1!
b101 %
1'
b101 +
#235770000000
0!
0'
#235780000000
1!
0$
b110 %
1'
0*
b110 +
#235790000000
0!
0'
#235800000000
1!
b111 %
1'
b111 +
#235810000000
0!
0'
#235820000000
1!
b1000 %
1'
b1000 +
#235830000000
0!
0'
#235840000000
1!
b1001 %
1'
b1001 +
#235850000000
1"
1(
#235860000000
0!
0"
b100 &
0'
0(
b100 ,
#235870000000
1!
b0 %
1'
b0 +
#235880000000
0!
0'
#235890000000
1!
1$
b1 %
1'
1*
b1 +
#235900000000
0!
0'
#235910000000
1!
b10 %
1'
b10 +
#235920000000
0!
0'
#235930000000
1!
b11 %
1'
b11 +
#235940000000
0!
0'
#235950000000
1!
b100 %
1'
b100 +
#235960000000
0!
0'
#235970000000
1!
b101 %
1'
b101 +
#235980000000
0!
0'
#235990000000
1!
b110 %
1'
b110 +
#236000000000
0!
0'
#236010000000
1!
b111 %
1'
b111 +
#236020000000
0!
0'
#236030000000
1!
0$
b1000 %
1'
0*
b1000 +
#236040000000
0!
0'
#236050000000
1!
b1001 %
1'
b1001 +
#236060000000
0!
0'
#236070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#236080000000
0!
0'
#236090000000
1!
1$
b1 %
1'
1*
b1 +
#236100000000
0!
0'
#236110000000
1!
b10 %
1'
b10 +
#236120000000
0!
0'
#236130000000
1!
b11 %
1'
b11 +
#236140000000
0!
0'
#236150000000
1!
b100 %
1'
b100 +
#236160000000
0!
0'
#236170000000
1!
b101 %
1'
b101 +
#236180000000
0!
0'
#236190000000
1!
0$
b110 %
1'
0*
b110 +
#236200000000
0!
0'
#236210000000
1!
b111 %
1'
b111 +
#236220000000
0!
0'
#236230000000
1!
b1000 %
1'
b1000 +
#236240000000
0!
0'
#236250000000
1!
b1001 %
1'
b1001 +
#236260000000
0!
0'
#236270000000
1!
b0 %
1'
b0 +
#236280000000
1"
1(
#236290000000
0!
0"
b100 &
0'
0(
b100 ,
#236300000000
1!
1$
b1 %
1'
1*
b1 +
#236310000000
0!
0'
#236320000000
1!
b10 %
1'
b10 +
#236330000000
0!
0'
#236340000000
1!
b11 %
1'
b11 +
#236350000000
0!
0'
#236360000000
1!
b100 %
1'
b100 +
#236370000000
0!
0'
#236380000000
1!
b101 %
1'
b101 +
#236390000000
0!
0'
#236400000000
1!
b110 %
1'
b110 +
#236410000000
0!
0'
#236420000000
1!
b111 %
1'
b111 +
#236430000000
0!
0'
#236440000000
1!
0$
b1000 %
1'
0*
b1000 +
#236450000000
0!
0'
#236460000000
1!
b1001 %
1'
b1001 +
#236470000000
0!
0'
#236480000000
1!
b0 %
1'
b0 +
#236490000000
0!
0'
#236500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#236510000000
0!
0'
#236520000000
1!
b10 %
1'
b10 +
#236530000000
0!
0'
#236540000000
1!
b11 %
1'
b11 +
#236550000000
0!
0'
#236560000000
1!
b100 %
1'
b100 +
#236570000000
0!
0'
#236580000000
1!
b101 %
1'
b101 +
#236590000000
0!
0'
#236600000000
1!
0$
b110 %
1'
0*
b110 +
#236610000000
0!
0'
#236620000000
1!
b111 %
1'
b111 +
#236630000000
0!
0'
#236640000000
1!
b1000 %
1'
b1000 +
#236650000000
0!
0'
#236660000000
1!
b1001 %
1'
b1001 +
#236670000000
0!
0'
#236680000000
1!
b0 %
1'
b0 +
#236690000000
0!
0'
#236700000000
1!
1$
b1 %
1'
1*
b1 +
#236710000000
1"
1(
#236720000000
0!
0"
b100 &
0'
0(
b100 ,
#236730000000
1!
b10 %
1'
b10 +
#236740000000
0!
0'
#236750000000
1!
b11 %
1'
b11 +
#236760000000
0!
0'
#236770000000
1!
b100 %
1'
b100 +
#236780000000
0!
0'
#236790000000
1!
b101 %
1'
b101 +
#236800000000
0!
0'
#236810000000
1!
b110 %
1'
b110 +
#236820000000
0!
0'
#236830000000
1!
b111 %
1'
b111 +
#236840000000
0!
0'
#236850000000
1!
0$
b1000 %
1'
0*
b1000 +
#236860000000
0!
0'
#236870000000
1!
b1001 %
1'
b1001 +
#236880000000
0!
0'
#236890000000
1!
b0 %
1'
b0 +
#236900000000
0!
0'
#236910000000
1!
1$
b1 %
1'
1*
b1 +
#236920000000
0!
0'
#236930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#236940000000
0!
0'
#236950000000
1!
b11 %
1'
b11 +
#236960000000
0!
0'
#236970000000
1!
b100 %
1'
b100 +
#236980000000
0!
0'
#236990000000
1!
b101 %
1'
b101 +
#237000000000
0!
0'
#237010000000
1!
0$
b110 %
1'
0*
b110 +
#237020000000
0!
0'
#237030000000
1!
b111 %
1'
b111 +
#237040000000
0!
0'
#237050000000
1!
b1000 %
1'
b1000 +
#237060000000
0!
0'
#237070000000
1!
b1001 %
1'
b1001 +
#237080000000
0!
0'
#237090000000
1!
b0 %
1'
b0 +
#237100000000
0!
0'
#237110000000
1!
1$
b1 %
1'
1*
b1 +
#237120000000
0!
0'
#237130000000
1!
b10 %
1'
b10 +
#237140000000
1"
1(
#237150000000
0!
0"
b100 &
0'
0(
b100 ,
#237160000000
1!
b11 %
1'
b11 +
#237170000000
0!
0'
#237180000000
1!
b100 %
1'
b100 +
#237190000000
0!
0'
#237200000000
1!
b101 %
1'
b101 +
#237210000000
0!
0'
#237220000000
1!
b110 %
1'
b110 +
#237230000000
0!
0'
#237240000000
1!
b111 %
1'
b111 +
#237250000000
0!
0'
#237260000000
1!
0$
b1000 %
1'
0*
b1000 +
#237270000000
0!
0'
#237280000000
1!
b1001 %
1'
b1001 +
#237290000000
0!
0'
#237300000000
1!
b0 %
1'
b0 +
#237310000000
0!
0'
#237320000000
1!
1$
b1 %
1'
1*
b1 +
#237330000000
0!
0'
#237340000000
1!
b10 %
1'
b10 +
#237350000000
0!
0'
#237360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#237370000000
0!
0'
#237380000000
1!
b100 %
1'
b100 +
#237390000000
0!
0'
#237400000000
1!
b101 %
1'
b101 +
#237410000000
0!
0'
#237420000000
1!
0$
b110 %
1'
0*
b110 +
#237430000000
0!
0'
#237440000000
1!
b111 %
1'
b111 +
#237450000000
0!
0'
#237460000000
1!
b1000 %
1'
b1000 +
#237470000000
0!
0'
#237480000000
1!
b1001 %
1'
b1001 +
#237490000000
0!
0'
#237500000000
1!
b0 %
1'
b0 +
#237510000000
0!
0'
#237520000000
1!
1$
b1 %
1'
1*
b1 +
#237530000000
0!
0'
#237540000000
1!
b10 %
1'
b10 +
#237550000000
0!
0'
#237560000000
1!
b11 %
1'
b11 +
#237570000000
1"
1(
#237580000000
0!
0"
b100 &
0'
0(
b100 ,
#237590000000
1!
b100 %
1'
b100 +
#237600000000
0!
0'
#237610000000
1!
b101 %
1'
b101 +
#237620000000
0!
0'
#237630000000
1!
b110 %
1'
b110 +
#237640000000
0!
0'
#237650000000
1!
b111 %
1'
b111 +
#237660000000
0!
0'
#237670000000
1!
0$
b1000 %
1'
0*
b1000 +
#237680000000
0!
0'
#237690000000
1!
b1001 %
1'
b1001 +
#237700000000
0!
0'
#237710000000
1!
b0 %
1'
b0 +
#237720000000
0!
0'
#237730000000
1!
1$
b1 %
1'
1*
b1 +
#237740000000
0!
0'
#237750000000
1!
b10 %
1'
b10 +
#237760000000
0!
0'
#237770000000
1!
b11 %
1'
b11 +
#237780000000
0!
0'
#237790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#237800000000
0!
0'
#237810000000
1!
b101 %
1'
b101 +
#237820000000
0!
0'
#237830000000
1!
0$
b110 %
1'
0*
b110 +
#237840000000
0!
0'
#237850000000
1!
b111 %
1'
b111 +
#237860000000
0!
0'
#237870000000
1!
b1000 %
1'
b1000 +
#237880000000
0!
0'
#237890000000
1!
b1001 %
1'
b1001 +
#237900000000
0!
0'
#237910000000
1!
b0 %
1'
b0 +
#237920000000
0!
0'
#237930000000
1!
1$
b1 %
1'
1*
b1 +
#237940000000
0!
0'
#237950000000
1!
b10 %
1'
b10 +
#237960000000
0!
0'
#237970000000
1!
b11 %
1'
b11 +
#237980000000
0!
0'
#237990000000
1!
b100 %
1'
b100 +
#238000000000
1"
1(
#238010000000
0!
0"
b100 &
0'
0(
b100 ,
#238020000000
1!
b101 %
1'
b101 +
#238030000000
0!
0'
#238040000000
1!
b110 %
1'
b110 +
#238050000000
0!
0'
#238060000000
1!
b111 %
1'
b111 +
#238070000000
0!
0'
#238080000000
1!
0$
b1000 %
1'
0*
b1000 +
#238090000000
0!
0'
#238100000000
1!
b1001 %
1'
b1001 +
#238110000000
0!
0'
#238120000000
1!
b0 %
1'
b0 +
#238130000000
0!
0'
#238140000000
1!
1$
b1 %
1'
1*
b1 +
#238150000000
0!
0'
#238160000000
1!
b10 %
1'
b10 +
#238170000000
0!
0'
#238180000000
1!
b11 %
1'
b11 +
#238190000000
0!
0'
#238200000000
1!
b100 %
1'
b100 +
#238210000000
0!
0'
#238220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#238230000000
0!
0'
#238240000000
1!
0$
b110 %
1'
0*
b110 +
#238250000000
0!
0'
#238260000000
1!
b111 %
1'
b111 +
#238270000000
0!
0'
#238280000000
1!
b1000 %
1'
b1000 +
#238290000000
0!
0'
#238300000000
1!
b1001 %
1'
b1001 +
#238310000000
0!
0'
#238320000000
1!
b0 %
1'
b0 +
#238330000000
0!
0'
#238340000000
1!
1$
b1 %
1'
1*
b1 +
#238350000000
0!
0'
#238360000000
1!
b10 %
1'
b10 +
#238370000000
0!
0'
#238380000000
1!
b11 %
1'
b11 +
#238390000000
0!
0'
#238400000000
1!
b100 %
1'
b100 +
#238410000000
0!
0'
#238420000000
1!
b101 %
1'
b101 +
#238430000000
1"
1(
#238440000000
0!
0"
b100 &
0'
0(
b100 ,
#238450000000
1!
b110 %
1'
b110 +
#238460000000
0!
0'
#238470000000
1!
b111 %
1'
b111 +
#238480000000
0!
0'
#238490000000
1!
0$
b1000 %
1'
0*
b1000 +
#238500000000
0!
0'
#238510000000
1!
b1001 %
1'
b1001 +
#238520000000
0!
0'
#238530000000
1!
b0 %
1'
b0 +
#238540000000
0!
0'
#238550000000
1!
1$
b1 %
1'
1*
b1 +
#238560000000
0!
0'
#238570000000
1!
b10 %
1'
b10 +
#238580000000
0!
0'
#238590000000
1!
b11 %
1'
b11 +
#238600000000
0!
0'
#238610000000
1!
b100 %
1'
b100 +
#238620000000
0!
0'
#238630000000
1!
b101 %
1'
b101 +
#238640000000
0!
0'
#238650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#238660000000
0!
0'
#238670000000
1!
b111 %
1'
b111 +
#238680000000
0!
0'
#238690000000
1!
b1000 %
1'
b1000 +
#238700000000
0!
0'
#238710000000
1!
b1001 %
1'
b1001 +
#238720000000
0!
0'
#238730000000
1!
b0 %
1'
b0 +
#238740000000
0!
0'
#238750000000
1!
1$
b1 %
1'
1*
b1 +
#238760000000
0!
0'
#238770000000
1!
b10 %
1'
b10 +
#238780000000
0!
0'
#238790000000
1!
b11 %
1'
b11 +
#238800000000
0!
0'
#238810000000
1!
b100 %
1'
b100 +
#238820000000
0!
0'
#238830000000
1!
b101 %
1'
b101 +
#238840000000
0!
0'
#238850000000
1!
0$
b110 %
1'
0*
b110 +
#238860000000
1"
1(
#238870000000
0!
0"
b100 &
0'
0(
b100 ,
#238880000000
1!
1$
b111 %
1'
1*
b111 +
#238890000000
0!
0'
#238900000000
1!
0$
b1000 %
1'
0*
b1000 +
#238910000000
0!
0'
#238920000000
1!
b1001 %
1'
b1001 +
#238930000000
0!
0'
#238940000000
1!
b0 %
1'
b0 +
#238950000000
0!
0'
#238960000000
1!
1$
b1 %
1'
1*
b1 +
#238970000000
0!
0'
#238980000000
1!
b10 %
1'
b10 +
#238990000000
0!
0'
#239000000000
1!
b11 %
1'
b11 +
#239010000000
0!
0'
#239020000000
1!
b100 %
1'
b100 +
#239030000000
0!
0'
#239040000000
1!
b101 %
1'
b101 +
#239050000000
0!
0'
#239060000000
1!
b110 %
1'
b110 +
#239070000000
0!
0'
#239080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#239090000000
0!
0'
#239100000000
1!
b1000 %
1'
b1000 +
#239110000000
0!
0'
#239120000000
1!
b1001 %
1'
b1001 +
#239130000000
0!
0'
#239140000000
1!
b0 %
1'
b0 +
#239150000000
0!
0'
#239160000000
1!
1$
b1 %
1'
1*
b1 +
#239170000000
0!
0'
#239180000000
1!
b10 %
1'
b10 +
#239190000000
0!
0'
#239200000000
1!
b11 %
1'
b11 +
#239210000000
0!
0'
#239220000000
1!
b100 %
1'
b100 +
#239230000000
0!
0'
#239240000000
1!
b101 %
1'
b101 +
#239250000000
0!
0'
#239260000000
1!
0$
b110 %
1'
0*
b110 +
#239270000000
0!
0'
#239280000000
1!
b111 %
1'
b111 +
#239290000000
1"
1(
#239300000000
0!
0"
b100 &
0'
0(
b100 ,
#239310000000
1!
b1000 %
1'
b1000 +
#239320000000
0!
0'
#239330000000
1!
b1001 %
1'
b1001 +
#239340000000
0!
0'
#239350000000
1!
b0 %
1'
b0 +
#239360000000
0!
0'
#239370000000
1!
1$
b1 %
1'
1*
b1 +
#239380000000
0!
0'
#239390000000
1!
b10 %
1'
b10 +
#239400000000
0!
0'
#239410000000
1!
b11 %
1'
b11 +
#239420000000
0!
0'
#239430000000
1!
b100 %
1'
b100 +
#239440000000
0!
0'
#239450000000
1!
b101 %
1'
b101 +
#239460000000
0!
0'
#239470000000
1!
b110 %
1'
b110 +
#239480000000
0!
0'
#239490000000
1!
b111 %
1'
b111 +
#239500000000
0!
0'
#239510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#239520000000
0!
0'
#239530000000
1!
b1001 %
1'
b1001 +
#239540000000
0!
0'
#239550000000
1!
b0 %
1'
b0 +
#239560000000
0!
0'
#239570000000
1!
1$
b1 %
1'
1*
b1 +
#239580000000
0!
0'
#239590000000
1!
b10 %
1'
b10 +
#239600000000
0!
0'
#239610000000
1!
b11 %
1'
b11 +
#239620000000
0!
0'
#239630000000
1!
b100 %
1'
b100 +
#239640000000
0!
0'
#239650000000
1!
b101 %
1'
b101 +
#239660000000
0!
0'
#239670000000
1!
0$
b110 %
1'
0*
b110 +
#239680000000
0!
0'
#239690000000
1!
b111 %
1'
b111 +
#239700000000
0!
0'
#239710000000
1!
b1000 %
1'
b1000 +
#239720000000
1"
1(
#239730000000
0!
0"
b100 &
0'
0(
b100 ,
#239740000000
1!
b1001 %
1'
b1001 +
#239750000000
0!
0'
#239760000000
1!
b0 %
1'
b0 +
#239770000000
0!
0'
#239780000000
1!
1$
b1 %
1'
1*
b1 +
#239790000000
0!
0'
#239800000000
1!
b10 %
1'
b10 +
#239810000000
0!
0'
#239820000000
1!
b11 %
1'
b11 +
#239830000000
0!
0'
#239840000000
1!
b100 %
1'
b100 +
#239850000000
0!
0'
#239860000000
1!
b101 %
1'
b101 +
#239870000000
0!
0'
#239880000000
1!
b110 %
1'
b110 +
#239890000000
0!
0'
#239900000000
1!
b111 %
1'
b111 +
#239910000000
0!
0'
#239920000000
1!
0$
b1000 %
1'
0*
b1000 +
#239930000000
0!
0'
#239940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#239950000000
0!
0'
#239960000000
1!
b0 %
1'
b0 +
#239970000000
0!
0'
#239980000000
1!
1$
b1 %
1'
1*
b1 +
#239990000000
0!
0'
#240000000000
1!
b10 %
1'
b10 +
#240010000000
0!
0'
#240020000000
1!
b11 %
1'
b11 +
#240030000000
0!
0'
#240040000000
1!
b100 %
1'
b100 +
#240050000000
0!
0'
#240060000000
1!
b101 %
1'
b101 +
#240070000000
0!
0'
#240080000000
1!
0$
b110 %
1'
0*
b110 +
#240090000000
0!
0'
#240100000000
1!
b111 %
1'
b111 +
#240110000000
0!
0'
#240120000000
1!
b1000 %
1'
b1000 +
#240130000000
0!
0'
#240140000000
1!
b1001 %
1'
b1001 +
#240150000000
1"
1(
#240160000000
0!
0"
b100 &
0'
0(
b100 ,
#240170000000
1!
b0 %
1'
b0 +
#240180000000
0!
0'
#240190000000
1!
1$
b1 %
1'
1*
b1 +
#240200000000
0!
0'
#240210000000
1!
b10 %
1'
b10 +
#240220000000
0!
0'
#240230000000
1!
b11 %
1'
b11 +
#240240000000
0!
0'
#240250000000
1!
b100 %
1'
b100 +
#240260000000
0!
0'
#240270000000
1!
b101 %
1'
b101 +
#240280000000
0!
0'
#240290000000
1!
b110 %
1'
b110 +
#240300000000
0!
0'
#240310000000
1!
b111 %
1'
b111 +
#240320000000
0!
0'
#240330000000
1!
0$
b1000 %
1'
0*
b1000 +
#240340000000
0!
0'
#240350000000
1!
b1001 %
1'
b1001 +
#240360000000
0!
0'
#240370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#240380000000
0!
0'
#240390000000
1!
1$
b1 %
1'
1*
b1 +
#240400000000
0!
0'
#240410000000
1!
b10 %
1'
b10 +
#240420000000
0!
0'
#240430000000
1!
b11 %
1'
b11 +
#240440000000
0!
0'
#240450000000
1!
b100 %
1'
b100 +
#240460000000
0!
0'
#240470000000
1!
b101 %
1'
b101 +
#240480000000
0!
0'
#240490000000
1!
0$
b110 %
1'
0*
b110 +
#240500000000
0!
0'
#240510000000
1!
b111 %
1'
b111 +
#240520000000
0!
0'
#240530000000
1!
b1000 %
1'
b1000 +
#240540000000
0!
0'
#240550000000
1!
b1001 %
1'
b1001 +
#240560000000
0!
0'
#240570000000
1!
b0 %
1'
b0 +
#240580000000
1"
1(
#240590000000
0!
0"
b100 &
0'
0(
b100 ,
#240600000000
1!
1$
b1 %
1'
1*
b1 +
#240610000000
0!
0'
#240620000000
1!
b10 %
1'
b10 +
#240630000000
0!
0'
#240640000000
1!
b11 %
1'
b11 +
#240650000000
0!
0'
#240660000000
1!
b100 %
1'
b100 +
#240670000000
0!
0'
#240680000000
1!
b101 %
1'
b101 +
#240690000000
0!
0'
#240700000000
1!
b110 %
1'
b110 +
#240710000000
0!
0'
#240720000000
1!
b111 %
1'
b111 +
#240730000000
0!
0'
#240740000000
1!
0$
b1000 %
1'
0*
b1000 +
#240750000000
0!
0'
#240760000000
1!
b1001 %
1'
b1001 +
#240770000000
0!
0'
#240780000000
1!
b0 %
1'
b0 +
#240790000000
0!
0'
#240800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#240810000000
0!
0'
#240820000000
1!
b10 %
1'
b10 +
#240830000000
0!
0'
#240840000000
1!
b11 %
1'
b11 +
#240850000000
0!
0'
#240860000000
1!
b100 %
1'
b100 +
#240870000000
0!
0'
#240880000000
1!
b101 %
1'
b101 +
#240890000000
0!
0'
#240900000000
1!
0$
b110 %
1'
0*
b110 +
#240910000000
0!
0'
#240920000000
1!
b111 %
1'
b111 +
#240930000000
0!
0'
#240940000000
1!
b1000 %
1'
b1000 +
#240950000000
0!
0'
#240960000000
1!
b1001 %
1'
b1001 +
#240970000000
0!
0'
#240980000000
1!
b0 %
1'
b0 +
#240990000000
0!
0'
#241000000000
1!
1$
b1 %
1'
1*
b1 +
#241010000000
1"
1(
#241020000000
0!
0"
b100 &
0'
0(
b100 ,
#241030000000
1!
b10 %
1'
b10 +
#241040000000
0!
0'
#241050000000
1!
b11 %
1'
b11 +
#241060000000
0!
0'
#241070000000
1!
b100 %
1'
b100 +
#241080000000
0!
0'
#241090000000
1!
b101 %
1'
b101 +
#241100000000
0!
0'
#241110000000
1!
b110 %
1'
b110 +
#241120000000
0!
0'
#241130000000
1!
b111 %
1'
b111 +
#241140000000
0!
0'
#241150000000
1!
0$
b1000 %
1'
0*
b1000 +
#241160000000
0!
0'
#241170000000
1!
b1001 %
1'
b1001 +
#241180000000
0!
0'
#241190000000
1!
b0 %
1'
b0 +
#241200000000
0!
0'
#241210000000
1!
1$
b1 %
1'
1*
b1 +
#241220000000
0!
0'
#241230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#241240000000
0!
0'
#241250000000
1!
b11 %
1'
b11 +
#241260000000
0!
0'
#241270000000
1!
b100 %
1'
b100 +
#241280000000
0!
0'
#241290000000
1!
b101 %
1'
b101 +
#241300000000
0!
0'
#241310000000
1!
0$
b110 %
1'
0*
b110 +
#241320000000
0!
0'
#241330000000
1!
b111 %
1'
b111 +
#241340000000
0!
0'
#241350000000
1!
b1000 %
1'
b1000 +
#241360000000
0!
0'
#241370000000
1!
b1001 %
1'
b1001 +
#241380000000
0!
0'
#241390000000
1!
b0 %
1'
b0 +
#241400000000
0!
0'
#241410000000
1!
1$
b1 %
1'
1*
b1 +
#241420000000
0!
0'
#241430000000
1!
b10 %
1'
b10 +
#241440000000
1"
1(
#241450000000
0!
0"
b100 &
0'
0(
b100 ,
#241460000000
1!
b11 %
1'
b11 +
#241470000000
0!
0'
#241480000000
1!
b100 %
1'
b100 +
#241490000000
0!
0'
#241500000000
1!
b101 %
1'
b101 +
#241510000000
0!
0'
#241520000000
1!
b110 %
1'
b110 +
#241530000000
0!
0'
#241540000000
1!
b111 %
1'
b111 +
#241550000000
0!
0'
#241560000000
1!
0$
b1000 %
1'
0*
b1000 +
#241570000000
0!
0'
#241580000000
1!
b1001 %
1'
b1001 +
#241590000000
0!
0'
#241600000000
1!
b0 %
1'
b0 +
#241610000000
0!
0'
#241620000000
1!
1$
b1 %
1'
1*
b1 +
#241630000000
0!
0'
#241640000000
1!
b10 %
1'
b10 +
#241650000000
0!
0'
#241660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#241670000000
0!
0'
#241680000000
1!
b100 %
1'
b100 +
#241690000000
0!
0'
#241700000000
1!
b101 %
1'
b101 +
#241710000000
0!
0'
#241720000000
1!
0$
b110 %
1'
0*
b110 +
#241730000000
0!
0'
#241740000000
1!
b111 %
1'
b111 +
#241750000000
0!
0'
#241760000000
1!
b1000 %
1'
b1000 +
#241770000000
0!
0'
#241780000000
1!
b1001 %
1'
b1001 +
#241790000000
0!
0'
#241800000000
1!
b0 %
1'
b0 +
#241810000000
0!
0'
#241820000000
1!
1$
b1 %
1'
1*
b1 +
#241830000000
0!
0'
#241840000000
1!
b10 %
1'
b10 +
#241850000000
0!
0'
#241860000000
1!
b11 %
1'
b11 +
#241870000000
1"
1(
#241880000000
0!
0"
b100 &
0'
0(
b100 ,
#241890000000
1!
b100 %
1'
b100 +
#241900000000
0!
0'
#241910000000
1!
b101 %
1'
b101 +
#241920000000
0!
0'
#241930000000
1!
b110 %
1'
b110 +
#241940000000
0!
0'
#241950000000
1!
b111 %
1'
b111 +
#241960000000
0!
0'
#241970000000
1!
0$
b1000 %
1'
0*
b1000 +
#241980000000
0!
0'
#241990000000
1!
b1001 %
1'
b1001 +
#242000000000
0!
0'
#242010000000
1!
b0 %
1'
b0 +
#242020000000
0!
0'
#242030000000
1!
1$
b1 %
1'
1*
b1 +
#242040000000
0!
0'
#242050000000
1!
b10 %
1'
b10 +
#242060000000
0!
0'
#242070000000
1!
b11 %
1'
b11 +
#242080000000
0!
0'
#242090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#242100000000
0!
0'
#242110000000
1!
b101 %
1'
b101 +
#242120000000
0!
0'
#242130000000
1!
0$
b110 %
1'
0*
b110 +
#242140000000
0!
0'
#242150000000
1!
b111 %
1'
b111 +
#242160000000
0!
0'
#242170000000
1!
b1000 %
1'
b1000 +
#242180000000
0!
0'
#242190000000
1!
b1001 %
1'
b1001 +
#242200000000
0!
0'
#242210000000
1!
b0 %
1'
b0 +
#242220000000
0!
0'
#242230000000
1!
1$
b1 %
1'
1*
b1 +
#242240000000
0!
0'
#242250000000
1!
b10 %
1'
b10 +
#242260000000
0!
0'
#242270000000
1!
b11 %
1'
b11 +
#242280000000
0!
0'
#242290000000
1!
b100 %
1'
b100 +
#242300000000
1"
1(
#242310000000
0!
0"
b100 &
0'
0(
b100 ,
#242320000000
1!
b101 %
1'
b101 +
#242330000000
0!
0'
#242340000000
1!
b110 %
1'
b110 +
#242350000000
0!
0'
#242360000000
1!
b111 %
1'
b111 +
#242370000000
0!
0'
#242380000000
1!
0$
b1000 %
1'
0*
b1000 +
#242390000000
0!
0'
#242400000000
1!
b1001 %
1'
b1001 +
#242410000000
0!
0'
#242420000000
1!
b0 %
1'
b0 +
#242430000000
0!
0'
#242440000000
1!
1$
b1 %
1'
1*
b1 +
#242450000000
0!
0'
#242460000000
1!
b10 %
1'
b10 +
#242470000000
0!
0'
#242480000000
1!
b11 %
1'
b11 +
#242490000000
0!
0'
#242500000000
1!
b100 %
1'
b100 +
#242510000000
0!
0'
#242520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#242530000000
0!
0'
#242540000000
1!
0$
b110 %
1'
0*
b110 +
#242550000000
0!
0'
#242560000000
1!
b111 %
1'
b111 +
#242570000000
0!
0'
#242580000000
1!
b1000 %
1'
b1000 +
#242590000000
0!
0'
#242600000000
1!
b1001 %
1'
b1001 +
#242610000000
0!
0'
#242620000000
1!
b0 %
1'
b0 +
#242630000000
0!
0'
#242640000000
1!
1$
b1 %
1'
1*
b1 +
#242650000000
0!
0'
#242660000000
1!
b10 %
1'
b10 +
#242670000000
0!
0'
#242680000000
1!
b11 %
1'
b11 +
#242690000000
0!
0'
#242700000000
1!
b100 %
1'
b100 +
#242710000000
0!
0'
#242720000000
1!
b101 %
1'
b101 +
#242730000000
1"
1(
#242740000000
0!
0"
b100 &
0'
0(
b100 ,
#242750000000
1!
b110 %
1'
b110 +
#242760000000
0!
0'
#242770000000
1!
b111 %
1'
b111 +
#242780000000
0!
0'
#242790000000
1!
0$
b1000 %
1'
0*
b1000 +
#242800000000
0!
0'
#242810000000
1!
b1001 %
1'
b1001 +
#242820000000
0!
0'
#242830000000
1!
b0 %
1'
b0 +
#242840000000
0!
0'
#242850000000
1!
1$
b1 %
1'
1*
b1 +
#242860000000
0!
0'
#242870000000
1!
b10 %
1'
b10 +
#242880000000
0!
0'
#242890000000
1!
b11 %
1'
b11 +
#242900000000
0!
0'
#242910000000
1!
b100 %
1'
b100 +
#242920000000
0!
0'
#242930000000
1!
b101 %
1'
b101 +
#242940000000
0!
0'
#242950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#242960000000
0!
0'
#242970000000
1!
b111 %
1'
b111 +
#242980000000
0!
0'
#242990000000
1!
b1000 %
1'
b1000 +
#243000000000
0!
0'
#243010000000
1!
b1001 %
1'
b1001 +
#243020000000
0!
0'
#243030000000
1!
b0 %
1'
b0 +
#243040000000
0!
0'
#243050000000
1!
1$
b1 %
1'
1*
b1 +
#243060000000
0!
0'
#243070000000
1!
b10 %
1'
b10 +
#243080000000
0!
0'
#243090000000
1!
b11 %
1'
b11 +
#243100000000
0!
0'
#243110000000
1!
b100 %
1'
b100 +
#243120000000
0!
0'
#243130000000
1!
b101 %
1'
b101 +
#243140000000
0!
0'
#243150000000
1!
0$
b110 %
1'
0*
b110 +
#243160000000
1"
1(
#243170000000
0!
0"
b100 &
0'
0(
b100 ,
#243180000000
1!
1$
b111 %
1'
1*
b111 +
#243190000000
0!
0'
#243200000000
1!
0$
b1000 %
1'
0*
b1000 +
#243210000000
0!
0'
#243220000000
1!
b1001 %
1'
b1001 +
#243230000000
0!
0'
#243240000000
1!
b0 %
1'
b0 +
#243250000000
0!
0'
#243260000000
1!
1$
b1 %
1'
1*
b1 +
#243270000000
0!
0'
#243280000000
1!
b10 %
1'
b10 +
#243290000000
0!
0'
#243300000000
1!
b11 %
1'
b11 +
#243310000000
0!
0'
#243320000000
1!
b100 %
1'
b100 +
#243330000000
0!
0'
#243340000000
1!
b101 %
1'
b101 +
#243350000000
0!
0'
#243360000000
1!
b110 %
1'
b110 +
#243370000000
0!
0'
#243380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#243390000000
0!
0'
#243400000000
1!
b1000 %
1'
b1000 +
#243410000000
0!
0'
#243420000000
1!
b1001 %
1'
b1001 +
#243430000000
0!
0'
#243440000000
1!
b0 %
1'
b0 +
#243450000000
0!
0'
#243460000000
1!
1$
b1 %
1'
1*
b1 +
#243470000000
0!
0'
#243480000000
1!
b10 %
1'
b10 +
#243490000000
0!
0'
#243500000000
1!
b11 %
1'
b11 +
#243510000000
0!
0'
#243520000000
1!
b100 %
1'
b100 +
#243530000000
0!
0'
#243540000000
1!
b101 %
1'
b101 +
#243550000000
0!
0'
#243560000000
1!
0$
b110 %
1'
0*
b110 +
#243570000000
0!
0'
#243580000000
1!
b111 %
1'
b111 +
#243590000000
1"
1(
#243600000000
0!
0"
b100 &
0'
0(
b100 ,
#243610000000
1!
b1000 %
1'
b1000 +
#243620000000
0!
0'
#243630000000
1!
b1001 %
1'
b1001 +
#243640000000
0!
0'
#243650000000
1!
b0 %
1'
b0 +
#243660000000
0!
0'
#243670000000
1!
1$
b1 %
1'
1*
b1 +
#243680000000
0!
0'
#243690000000
1!
b10 %
1'
b10 +
#243700000000
0!
0'
#243710000000
1!
b11 %
1'
b11 +
#243720000000
0!
0'
#243730000000
1!
b100 %
1'
b100 +
#243740000000
0!
0'
#243750000000
1!
b101 %
1'
b101 +
#243760000000
0!
0'
#243770000000
1!
b110 %
1'
b110 +
#243780000000
0!
0'
#243790000000
1!
b111 %
1'
b111 +
#243800000000
0!
0'
#243810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#243820000000
0!
0'
#243830000000
1!
b1001 %
1'
b1001 +
#243840000000
0!
0'
#243850000000
1!
b0 %
1'
b0 +
#243860000000
0!
0'
#243870000000
1!
1$
b1 %
1'
1*
b1 +
#243880000000
0!
0'
#243890000000
1!
b10 %
1'
b10 +
#243900000000
0!
0'
#243910000000
1!
b11 %
1'
b11 +
#243920000000
0!
0'
#243930000000
1!
b100 %
1'
b100 +
#243940000000
0!
0'
#243950000000
1!
b101 %
1'
b101 +
#243960000000
0!
0'
#243970000000
1!
0$
b110 %
1'
0*
b110 +
#243980000000
0!
0'
#243990000000
1!
b111 %
1'
b111 +
#244000000000
0!
0'
#244010000000
1!
b1000 %
1'
b1000 +
#244020000000
1"
1(
#244030000000
0!
0"
b100 &
0'
0(
b100 ,
#244040000000
1!
b1001 %
1'
b1001 +
#244050000000
0!
0'
#244060000000
1!
b0 %
1'
b0 +
#244070000000
0!
0'
#244080000000
1!
1$
b1 %
1'
1*
b1 +
#244090000000
0!
0'
#244100000000
1!
b10 %
1'
b10 +
#244110000000
0!
0'
#244120000000
1!
b11 %
1'
b11 +
#244130000000
0!
0'
#244140000000
1!
b100 %
1'
b100 +
#244150000000
0!
0'
#244160000000
1!
b101 %
1'
b101 +
#244170000000
0!
0'
#244180000000
1!
b110 %
1'
b110 +
#244190000000
0!
0'
#244200000000
1!
b111 %
1'
b111 +
#244210000000
0!
0'
#244220000000
1!
0$
b1000 %
1'
0*
b1000 +
#244230000000
0!
0'
#244240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#244250000000
0!
0'
#244260000000
1!
b0 %
1'
b0 +
#244270000000
0!
0'
#244280000000
1!
1$
b1 %
1'
1*
b1 +
#244290000000
0!
0'
#244300000000
1!
b10 %
1'
b10 +
#244310000000
0!
0'
#244320000000
1!
b11 %
1'
b11 +
#244330000000
0!
0'
#244340000000
1!
b100 %
1'
b100 +
#244350000000
0!
0'
#244360000000
1!
b101 %
1'
b101 +
#244370000000
0!
0'
#244380000000
1!
0$
b110 %
1'
0*
b110 +
#244390000000
0!
0'
#244400000000
1!
b111 %
1'
b111 +
#244410000000
0!
0'
#244420000000
1!
b1000 %
1'
b1000 +
#244430000000
0!
0'
#244440000000
1!
b1001 %
1'
b1001 +
#244450000000
1"
1(
#244460000000
0!
0"
b100 &
0'
0(
b100 ,
#244470000000
1!
b0 %
1'
b0 +
#244480000000
0!
0'
#244490000000
1!
1$
b1 %
1'
1*
b1 +
#244500000000
0!
0'
#244510000000
1!
b10 %
1'
b10 +
#244520000000
0!
0'
#244530000000
1!
b11 %
1'
b11 +
#244540000000
0!
0'
#244550000000
1!
b100 %
1'
b100 +
#244560000000
0!
0'
#244570000000
1!
b101 %
1'
b101 +
#244580000000
0!
0'
#244590000000
1!
b110 %
1'
b110 +
#244600000000
0!
0'
#244610000000
1!
b111 %
1'
b111 +
#244620000000
0!
0'
#244630000000
1!
0$
b1000 %
1'
0*
b1000 +
#244640000000
0!
0'
#244650000000
1!
b1001 %
1'
b1001 +
#244660000000
0!
0'
#244670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#244680000000
0!
0'
#244690000000
1!
1$
b1 %
1'
1*
b1 +
#244700000000
0!
0'
#244710000000
1!
b10 %
1'
b10 +
#244720000000
0!
0'
#244730000000
1!
b11 %
1'
b11 +
#244740000000
0!
0'
#244750000000
1!
b100 %
1'
b100 +
#244760000000
0!
0'
#244770000000
1!
b101 %
1'
b101 +
#244780000000
0!
0'
#244790000000
1!
0$
b110 %
1'
0*
b110 +
#244800000000
0!
0'
#244810000000
1!
b111 %
1'
b111 +
#244820000000
0!
0'
#244830000000
1!
b1000 %
1'
b1000 +
#244840000000
0!
0'
#244850000000
1!
b1001 %
1'
b1001 +
#244860000000
0!
0'
#244870000000
1!
b0 %
1'
b0 +
#244880000000
1"
1(
#244890000000
0!
0"
b100 &
0'
0(
b100 ,
#244900000000
1!
1$
b1 %
1'
1*
b1 +
#244910000000
0!
0'
#244920000000
1!
b10 %
1'
b10 +
#244930000000
0!
0'
#244940000000
1!
b11 %
1'
b11 +
#244950000000
0!
0'
#244960000000
1!
b100 %
1'
b100 +
#244970000000
0!
0'
#244980000000
1!
b101 %
1'
b101 +
#244990000000
0!
0'
#245000000000
1!
b110 %
1'
b110 +
#245010000000
0!
0'
#245020000000
1!
b111 %
1'
b111 +
#245030000000
0!
0'
#245040000000
1!
0$
b1000 %
1'
0*
b1000 +
#245050000000
0!
0'
#245060000000
1!
b1001 %
1'
b1001 +
#245070000000
0!
0'
#245080000000
1!
b0 %
1'
b0 +
#245090000000
0!
0'
#245100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#245110000000
0!
0'
#245120000000
1!
b10 %
1'
b10 +
#245130000000
0!
0'
#245140000000
1!
b11 %
1'
b11 +
#245150000000
0!
0'
#245160000000
1!
b100 %
1'
b100 +
#245170000000
0!
0'
#245180000000
1!
b101 %
1'
b101 +
#245190000000
0!
0'
#245200000000
1!
0$
b110 %
1'
0*
b110 +
#245210000000
0!
0'
#245220000000
1!
b111 %
1'
b111 +
#245230000000
0!
0'
#245240000000
1!
b1000 %
1'
b1000 +
#245250000000
0!
0'
#245260000000
1!
b1001 %
1'
b1001 +
#245270000000
0!
0'
#245280000000
1!
b0 %
1'
b0 +
#245290000000
0!
0'
#245300000000
1!
1$
b1 %
1'
1*
b1 +
#245310000000
1"
1(
#245320000000
0!
0"
b100 &
0'
0(
b100 ,
#245330000000
1!
b10 %
1'
b10 +
#245340000000
0!
0'
#245350000000
1!
b11 %
1'
b11 +
#245360000000
0!
0'
#245370000000
1!
b100 %
1'
b100 +
#245380000000
0!
0'
#245390000000
1!
b101 %
1'
b101 +
#245400000000
0!
0'
#245410000000
1!
b110 %
1'
b110 +
#245420000000
0!
0'
#245430000000
1!
b111 %
1'
b111 +
#245440000000
0!
0'
#245450000000
1!
0$
b1000 %
1'
0*
b1000 +
#245460000000
0!
0'
#245470000000
1!
b1001 %
1'
b1001 +
#245480000000
0!
0'
#245490000000
1!
b0 %
1'
b0 +
#245500000000
0!
0'
#245510000000
1!
1$
b1 %
1'
1*
b1 +
#245520000000
0!
0'
#245530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#245540000000
0!
0'
#245550000000
1!
b11 %
1'
b11 +
#245560000000
0!
0'
#245570000000
1!
b100 %
1'
b100 +
#245580000000
0!
0'
#245590000000
1!
b101 %
1'
b101 +
#245600000000
0!
0'
#245610000000
1!
0$
b110 %
1'
0*
b110 +
#245620000000
0!
0'
#245630000000
1!
b111 %
1'
b111 +
#245640000000
0!
0'
#245650000000
1!
b1000 %
1'
b1000 +
#245660000000
0!
0'
#245670000000
1!
b1001 %
1'
b1001 +
#245680000000
0!
0'
#245690000000
1!
b0 %
1'
b0 +
#245700000000
0!
0'
#245710000000
1!
1$
b1 %
1'
1*
b1 +
#245720000000
0!
0'
#245730000000
1!
b10 %
1'
b10 +
#245740000000
1"
1(
#245750000000
0!
0"
b100 &
0'
0(
b100 ,
#245760000000
1!
b11 %
1'
b11 +
#245770000000
0!
0'
#245780000000
1!
b100 %
1'
b100 +
#245790000000
0!
0'
#245800000000
1!
b101 %
1'
b101 +
#245810000000
0!
0'
#245820000000
1!
b110 %
1'
b110 +
#245830000000
0!
0'
#245840000000
1!
b111 %
1'
b111 +
#245850000000
0!
0'
#245860000000
1!
0$
b1000 %
1'
0*
b1000 +
#245870000000
0!
0'
#245880000000
1!
b1001 %
1'
b1001 +
#245890000000
0!
0'
#245900000000
1!
b0 %
1'
b0 +
#245910000000
0!
0'
#245920000000
1!
1$
b1 %
1'
1*
b1 +
#245930000000
0!
0'
#245940000000
1!
b10 %
1'
b10 +
#245950000000
0!
0'
#245960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#245970000000
0!
0'
#245980000000
1!
b100 %
1'
b100 +
#245990000000
0!
0'
#246000000000
1!
b101 %
1'
b101 +
#246010000000
0!
0'
#246020000000
1!
0$
b110 %
1'
0*
b110 +
#246030000000
0!
0'
#246040000000
1!
b111 %
1'
b111 +
#246050000000
0!
0'
#246060000000
1!
b1000 %
1'
b1000 +
#246070000000
0!
0'
#246080000000
1!
b1001 %
1'
b1001 +
#246090000000
0!
0'
#246100000000
1!
b0 %
1'
b0 +
#246110000000
0!
0'
#246120000000
1!
1$
b1 %
1'
1*
b1 +
#246130000000
0!
0'
#246140000000
1!
b10 %
1'
b10 +
#246150000000
0!
0'
#246160000000
1!
b11 %
1'
b11 +
#246170000000
1"
1(
#246180000000
0!
0"
b100 &
0'
0(
b100 ,
#246190000000
1!
b100 %
1'
b100 +
#246200000000
0!
0'
#246210000000
1!
b101 %
1'
b101 +
#246220000000
0!
0'
#246230000000
1!
b110 %
1'
b110 +
#246240000000
0!
0'
#246250000000
1!
b111 %
1'
b111 +
#246260000000
0!
0'
#246270000000
1!
0$
b1000 %
1'
0*
b1000 +
#246280000000
0!
0'
#246290000000
1!
b1001 %
1'
b1001 +
#246300000000
0!
0'
#246310000000
1!
b0 %
1'
b0 +
#246320000000
0!
0'
#246330000000
1!
1$
b1 %
1'
1*
b1 +
#246340000000
0!
0'
#246350000000
1!
b10 %
1'
b10 +
#246360000000
0!
0'
#246370000000
1!
b11 %
1'
b11 +
#246380000000
0!
0'
#246390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#246400000000
0!
0'
#246410000000
1!
b101 %
1'
b101 +
#246420000000
0!
0'
#246430000000
1!
0$
b110 %
1'
0*
b110 +
#246440000000
0!
0'
#246450000000
1!
b111 %
1'
b111 +
#246460000000
0!
0'
#246470000000
1!
b1000 %
1'
b1000 +
#246480000000
0!
0'
#246490000000
1!
b1001 %
1'
b1001 +
#246500000000
0!
0'
#246510000000
1!
b0 %
1'
b0 +
#246520000000
0!
0'
#246530000000
1!
1$
b1 %
1'
1*
b1 +
#246540000000
0!
0'
#246550000000
1!
b10 %
1'
b10 +
#246560000000
0!
0'
#246570000000
1!
b11 %
1'
b11 +
#246580000000
0!
0'
#246590000000
1!
b100 %
1'
b100 +
#246600000000
1"
1(
#246610000000
0!
0"
b100 &
0'
0(
b100 ,
#246620000000
1!
b101 %
1'
b101 +
#246630000000
0!
0'
#246640000000
1!
b110 %
1'
b110 +
#246650000000
0!
0'
#246660000000
1!
b111 %
1'
b111 +
#246670000000
0!
0'
#246680000000
1!
0$
b1000 %
1'
0*
b1000 +
#246690000000
0!
0'
#246700000000
1!
b1001 %
1'
b1001 +
#246710000000
0!
0'
#246720000000
1!
b0 %
1'
b0 +
#246730000000
0!
0'
#246740000000
1!
1$
b1 %
1'
1*
b1 +
#246750000000
0!
0'
#246760000000
1!
b10 %
1'
b10 +
#246770000000
0!
0'
#246780000000
1!
b11 %
1'
b11 +
#246790000000
0!
0'
#246800000000
1!
b100 %
1'
b100 +
#246810000000
0!
0'
#246820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#246830000000
0!
0'
#246840000000
1!
0$
b110 %
1'
0*
b110 +
#246850000000
0!
0'
#246860000000
1!
b111 %
1'
b111 +
#246870000000
0!
0'
#246880000000
1!
b1000 %
1'
b1000 +
#246890000000
0!
0'
#246900000000
1!
b1001 %
1'
b1001 +
#246910000000
0!
0'
#246920000000
1!
b0 %
1'
b0 +
#246930000000
0!
0'
#246940000000
1!
1$
b1 %
1'
1*
b1 +
#246950000000
0!
0'
#246960000000
1!
b10 %
1'
b10 +
#246970000000
0!
0'
#246980000000
1!
b11 %
1'
b11 +
#246990000000
0!
0'
#247000000000
1!
b100 %
1'
b100 +
#247010000000
0!
0'
#247020000000
1!
b101 %
1'
b101 +
#247030000000
1"
1(
#247040000000
0!
0"
b100 &
0'
0(
b100 ,
#247050000000
1!
b110 %
1'
b110 +
#247060000000
0!
0'
#247070000000
1!
b111 %
1'
b111 +
#247080000000
0!
0'
#247090000000
1!
0$
b1000 %
1'
0*
b1000 +
#247100000000
0!
0'
#247110000000
1!
b1001 %
1'
b1001 +
#247120000000
0!
0'
#247130000000
1!
b0 %
1'
b0 +
#247140000000
0!
0'
#247150000000
1!
1$
b1 %
1'
1*
b1 +
#247160000000
0!
0'
#247170000000
1!
b10 %
1'
b10 +
#247180000000
0!
0'
#247190000000
1!
b11 %
1'
b11 +
#247200000000
0!
0'
#247210000000
1!
b100 %
1'
b100 +
#247220000000
0!
0'
#247230000000
1!
b101 %
1'
b101 +
#247240000000
0!
0'
#247250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#247260000000
0!
0'
#247270000000
1!
b111 %
1'
b111 +
#247280000000
0!
0'
#247290000000
1!
b1000 %
1'
b1000 +
#247300000000
0!
0'
#247310000000
1!
b1001 %
1'
b1001 +
#247320000000
0!
0'
#247330000000
1!
b0 %
1'
b0 +
#247340000000
0!
0'
#247350000000
1!
1$
b1 %
1'
1*
b1 +
#247360000000
0!
0'
#247370000000
1!
b10 %
1'
b10 +
#247380000000
0!
0'
#247390000000
1!
b11 %
1'
b11 +
#247400000000
0!
0'
#247410000000
1!
b100 %
1'
b100 +
#247420000000
0!
0'
#247430000000
1!
b101 %
1'
b101 +
#247440000000
0!
0'
#247450000000
1!
0$
b110 %
1'
0*
b110 +
#247460000000
1"
1(
#247470000000
0!
0"
b100 &
0'
0(
b100 ,
#247480000000
1!
1$
b111 %
1'
1*
b111 +
#247490000000
0!
0'
#247500000000
1!
0$
b1000 %
1'
0*
b1000 +
#247510000000
0!
0'
#247520000000
1!
b1001 %
1'
b1001 +
#247530000000
0!
0'
#247540000000
1!
b0 %
1'
b0 +
#247550000000
0!
0'
#247560000000
1!
1$
b1 %
1'
1*
b1 +
#247570000000
0!
0'
#247580000000
1!
b10 %
1'
b10 +
#247590000000
0!
0'
#247600000000
1!
b11 %
1'
b11 +
#247610000000
0!
0'
#247620000000
1!
b100 %
1'
b100 +
#247630000000
0!
0'
#247640000000
1!
b101 %
1'
b101 +
#247650000000
0!
0'
#247660000000
1!
b110 %
1'
b110 +
#247670000000
0!
0'
#247680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#247690000000
0!
0'
#247700000000
1!
b1000 %
1'
b1000 +
#247710000000
0!
0'
#247720000000
1!
b1001 %
1'
b1001 +
#247730000000
0!
0'
#247740000000
1!
b0 %
1'
b0 +
#247750000000
0!
0'
#247760000000
1!
1$
b1 %
1'
1*
b1 +
#247770000000
0!
0'
#247780000000
1!
b10 %
1'
b10 +
#247790000000
0!
0'
#247800000000
1!
b11 %
1'
b11 +
#247810000000
0!
0'
#247820000000
1!
b100 %
1'
b100 +
#247830000000
0!
0'
#247840000000
1!
b101 %
1'
b101 +
#247850000000
0!
0'
#247860000000
1!
0$
b110 %
1'
0*
b110 +
#247870000000
0!
0'
#247880000000
1!
b111 %
1'
b111 +
#247890000000
1"
1(
#247900000000
0!
0"
b100 &
0'
0(
b100 ,
#247910000000
1!
b1000 %
1'
b1000 +
#247920000000
0!
0'
#247930000000
1!
b1001 %
1'
b1001 +
#247940000000
0!
0'
#247950000000
1!
b0 %
1'
b0 +
#247960000000
0!
0'
#247970000000
1!
1$
b1 %
1'
1*
b1 +
#247980000000
0!
0'
#247990000000
1!
b10 %
1'
b10 +
#248000000000
0!
0'
#248010000000
1!
b11 %
1'
b11 +
#248020000000
0!
0'
#248030000000
1!
b100 %
1'
b100 +
#248040000000
0!
0'
#248050000000
1!
b101 %
1'
b101 +
#248060000000
0!
0'
#248070000000
1!
b110 %
1'
b110 +
#248080000000
0!
0'
#248090000000
1!
b111 %
1'
b111 +
#248100000000
0!
0'
#248110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#248120000000
0!
0'
#248130000000
1!
b1001 %
1'
b1001 +
#248140000000
0!
0'
#248150000000
1!
b0 %
1'
b0 +
#248160000000
0!
0'
#248170000000
1!
1$
b1 %
1'
1*
b1 +
#248180000000
0!
0'
#248190000000
1!
b10 %
1'
b10 +
#248200000000
0!
0'
#248210000000
1!
b11 %
1'
b11 +
#248220000000
0!
0'
#248230000000
1!
b100 %
1'
b100 +
#248240000000
0!
0'
#248250000000
1!
b101 %
1'
b101 +
#248260000000
0!
0'
#248270000000
1!
0$
b110 %
1'
0*
b110 +
#248280000000
0!
0'
#248290000000
1!
b111 %
1'
b111 +
#248300000000
0!
0'
#248310000000
1!
b1000 %
1'
b1000 +
#248320000000
1"
1(
#248330000000
0!
0"
b100 &
0'
0(
b100 ,
#248340000000
1!
b1001 %
1'
b1001 +
#248350000000
0!
0'
#248360000000
1!
b0 %
1'
b0 +
#248370000000
0!
0'
#248380000000
1!
1$
b1 %
1'
1*
b1 +
#248390000000
0!
0'
#248400000000
1!
b10 %
1'
b10 +
#248410000000
0!
0'
#248420000000
1!
b11 %
1'
b11 +
#248430000000
0!
0'
#248440000000
1!
b100 %
1'
b100 +
#248450000000
0!
0'
#248460000000
1!
b101 %
1'
b101 +
#248470000000
0!
0'
#248480000000
1!
b110 %
1'
b110 +
#248490000000
0!
0'
#248500000000
1!
b111 %
1'
b111 +
#248510000000
0!
0'
#248520000000
1!
0$
b1000 %
1'
0*
b1000 +
#248530000000
0!
0'
#248540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#248550000000
0!
0'
#248560000000
1!
b0 %
1'
b0 +
#248570000000
0!
0'
#248580000000
1!
1$
b1 %
1'
1*
b1 +
#248590000000
0!
0'
#248600000000
1!
b10 %
1'
b10 +
#248610000000
0!
0'
#248620000000
1!
b11 %
1'
b11 +
#248630000000
0!
0'
#248640000000
1!
b100 %
1'
b100 +
#248650000000
0!
0'
#248660000000
1!
b101 %
1'
b101 +
#248670000000
0!
0'
#248680000000
1!
0$
b110 %
1'
0*
b110 +
#248690000000
0!
0'
#248700000000
1!
b111 %
1'
b111 +
#248710000000
0!
0'
#248720000000
1!
b1000 %
1'
b1000 +
#248730000000
0!
0'
#248740000000
1!
b1001 %
1'
b1001 +
#248750000000
1"
1(
#248760000000
0!
0"
b100 &
0'
0(
b100 ,
#248770000000
1!
b0 %
1'
b0 +
#248780000000
0!
0'
#248790000000
1!
1$
b1 %
1'
1*
b1 +
#248800000000
0!
0'
#248810000000
1!
b10 %
1'
b10 +
#248820000000
0!
0'
#248830000000
1!
b11 %
1'
b11 +
#248840000000
0!
0'
#248850000000
1!
b100 %
1'
b100 +
#248860000000
0!
0'
#248870000000
1!
b101 %
1'
b101 +
#248880000000
0!
0'
#248890000000
1!
b110 %
1'
b110 +
#248900000000
0!
0'
#248910000000
1!
b111 %
1'
b111 +
#248920000000
0!
0'
#248930000000
1!
0$
b1000 %
1'
0*
b1000 +
#248940000000
0!
0'
#248950000000
1!
b1001 %
1'
b1001 +
#248960000000
0!
0'
#248970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#248980000000
0!
0'
#248990000000
1!
1$
b1 %
1'
1*
b1 +
#249000000000
0!
0'
#249010000000
1!
b10 %
1'
b10 +
#249020000000
0!
0'
#249030000000
1!
b11 %
1'
b11 +
#249040000000
0!
0'
#249050000000
1!
b100 %
1'
b100 +
#249060000000
0!
0'
#249070000000
1!
b101 %
1'
b101 +
#249080000000
0!
0'
#249090000000
1!
0$
b110 %
1'
0*
b110 +
#249100000000
0!
0'
#249110000000
1!
b111 %
1'
b111 +
#249120000000
0!
0'
#249130000000
1!
b1000 %
1'
b1000 +
#249140000000
0!
0'
#249150000000
1!
b1001 %
1'
b1001 +
#249160000000
0!
0'
#249170000000
1!
b0 %
1'
b0 +
#249180000000
1"
1(
#249190000000
0!
0"
b100 &
0'
0(
b100 ,
#249200000000
1!
1$
b1 %
1'
1*
b1 +
#249210000000
0!
0'
#249220000000
1!
b10 %
1'
b10 +
#249230000000
0!
0'
#249240000000
1!
b11 %
1'
b11 +
#249250000000
0!
0'
#249260000000
1!
b100 %
1'
b100 +
#249270000000
0!
0'
#249280000000
1!
b101 %
1'
b101 +
#249290000000
0!
0'
#249300000000
1!
b110 %
1'
b110 +
#249310000000
0!
0'
#249320000000
1!
b111 %
1'
b111 +
#249330000000
0!
0'
#249340000000
1!
0$
b1000 %
1'
0*
b1000 +
#249350000000
0!
0'
#249360000000
1!
b1001 %
1'
b1001 +
#249370000000
0!
0'
#249380000000
1!
b0 %
1'
b0 +
#249390000000
0!
0'
#249400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#249410000000
0!
0'
#249420000000
1!
b10 %
1'
b10 +
#249430000000
0!
0'
#249440000000
1!
b11 %
1'
b11 +
#249450000000
0!
0'
#249460000000
1!
b100 %
1'
b100 +
#249470000000
0!
0'
#249480000000
1!
b101 %
1'
b101 +
#249490000000
0!
0'
#249500000000
1!
0$
b110 %
1'
0*
b110 +
#249510000000
0!
0'
#249520000000
1!
b111 %
1'
b111 +
#249530000000
0!
0'
#249540000000
1!
b1000 %
1'
b1000 +
#249550000000
0!
0'
#249560000000
1!
b1001 %
1'
b1001 +
#249570000000
0!
0'
#249580000000
1!
b0 %
1'
b0 +
#249590000000
0!
0'
#249600000000
1!
1$
b1 %
1'
1*
b1 +
#249610000000
1"
1(
#249620000000
0!
0"
b100 &
0'
0(
b100 ,
#249630000000
1!
b10 %
1'
b10 +
#249640000000
0!
0'
#249650000000
1!
b11 %
1'
b11 +
#249660000000
0!
0'
#249670000000
1!
b100 %
1'
b100 +
#249680000000
0!
0'
#249690000000
1!
b101 %
1'
b101 +
#249700000000
0!
0'
#249710000000
1!
b110 %
1'
b110 +
#249720000000
0!
0'
#249730000000
1!
b111 %
1'
b111 +
#249740000000
0!
0'
#249750000000
1!
0$
b1000 %
1'
0*
b1000 +
#249760000000
0!
0'
#249770000000
1!
b1001 %
1'
b1001 +
#249780000000
0!
0'
#249790000000
1!
b0 %
1'
b0 +
#249800000000
0!
0'
#249810000000
1!
1$
b1 %
1'
1*
b1 +
#249820000000
0!
0'
#249830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#249840000000
0!
0'
#249850000000
1!
b11 %
1'
b11 +
#249860000000
0!
0'
#249870000000
1!
b100 %
1'
b100 +
#249880000000
0!
0'
#249890000000
1!
b101 %
1'
b101 +
#249900000000
0!
0'
#249910000000
1!
0$
b110 %
1'
0*
b110 +
#249920000000
0!
0'
#249930000000
1!
b111 %
1'
b111 +
#249940000000
0!
0'
#249950000000
1!
b1000 %
1'
b1000 +
#249960000000
0!
0'
#249970000000
1!
b1001 %
1'
b1001 +
#249980000000
0!
0'
#249990000000
1!
b0 %
1'
b0 +
#250000000000
0!
0'
#250010000000
1!
1$
b1 %
1'
1*
b1 +
#250020000000
0!
0'
#250030000000
1!
b10 %
1'
b10 +
#250040000000
1"
1(
#250050000000
0!
0"
b100 &
0'
0(
b100 ,
#250060000000
1!
b11 %
1'
b11 +
#250070000000
0!
0'
#250080000000
1!
b100 %
1'
b100 +
#250090000000
0!
0'
#250100000000
1!
b101 %
1'
b101 +
#250110000000
0!
0'
#250120000000
1!
b110 %
1'
b110 +
#250130000000
0!
0'
#250140000000
1!
b111 %
1'
b111 +
#250150000000
0!
0'
#250160000000
1!
0$
b1000 %
1'
0*
b1000 +
#250170000000
0!
0'
#250180000000
1!
b1001 %
1'
b1001 +
#250190000000
0!
0'
#250200000000
1!
b0 %
1'
b0 +
#250210000000
0!
0'
#250220000000
1!
1$
b1 %
1'
1*
b1 +
#250230000000
0!
0'
#250240000000
1!
b10 %
1'
b10 +
#250250000000
0!
0'
#250260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#250270000000
0!
0'
#250280000000
1!
b100 %
1'
b100 +
#250290000000
0!
0'
#250300000000
1!
b101 %
1'
b101 +
#250310000000
0!
0'
#250320000000
1!
0$
b110 %
1'
0*
b110 +
#250330000000
0!
0'
#250340000000
1!
b111 %
1'
b111 +
#250350000000
0!
0'
#250360000000
1!
b1000 %
1'
b1000 +
#250370000000
0!
0'
#250380000000
1!
b1001 %
1'
b1001 +
#250390000000
0!
0'
#250400000000
1!
b0 %
1'
b0 +
#250410000000
0!
0'
#250420000000
1!
1$
b1 %
1'
1*
b1 +
#250430000000
0!
0'
#250440000000
1!
b10 %
1'
b10 +
#250450000000
0!
0'
#250460000000
1!
b11 %
1'
b11 +
#250470000000
1"
1(
#250480000000
0!
0"
b100 &
0'
0(
b100 ,
#250490000000
1!
b100 %
1'
b100 +
#250500000000
0!
0'
#250510000000
1!
b101 %
1'
b101 +
#250520000000
0!
0'
#250530000000
1!
b110 %
1'
b110 +
#250540000000
0!
0'
#250550000000
1!
b111 %
1'
b111 +
#250560000000
0!
0'
#250570000000
1!
0$
b1000 %
1'
0*
b1000 +
#250580000000
0!
0'
#250590000000
1!
b1001 %
1'
b1001 +
#250600000000
0!
0'
#250610000000
1!
b0 %
1'
b0 +
#250620000000
0!
0'
#250630000000
1!
1$
b1 %
1'
1*
b1 +
#250640000000
0!
0'
#250650000000
1!
b10 %
1'
b10 +
#250660000000
0!
0'
#250670000000
1!
b11 %
1'
b11 +
#250680000000
0!
0'
#250690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#250700000000
0!
0'
#250710000000
1!
b101 %
1'
b101 +
#250720000000
0!
0'
#250730000000
1!
0$
b110 %
1'
0*
b110 +
#250740000000
0!
0'
#250750000000
1!
b111 %
1'
b111 +
#250760000000
0!
0'
#250770000000
1!
b1000 %
1'
b1000 +
#250780000000
0!
0'
#250790000000
1!
b1001 %
1'
b1001 +
#250800000000
0!
0'
#250810000000
1!
b0 %
1'
b0 +
#250820000000
0!
0'
#250830000000
1!
1$
b1 %
1'
1*
b1 +
#250840000000
0!
0'
#250850000000
1!
b10 %
1'
b10 +
#250860000000
0!
0'
#250870000000
1!
b11 %
1'
b11 +
#250880000000
0!
0'
#250890000000
1!
b100 %
1'
b100 +
#250900000000
1"
1(
#250910000000
0!
0"
b100 &
0'
0(
b100 ,
#250920000000
1!
b101 %
1'
b101 +
#250930000000
0!
0'
#250940000000
1!
b110 %
1'
b110 +
#250950000000
0!
0'
#250960000000
1!
b111 %
1'
b111 +
#250970000000
0!
0'
#250980000000
1!
0$
b1000 %
1'
0*
b1000 +
#250990000000
0!
0'
#251000000000
1!
b1001 %
1'
b1001 +
#251010000000
0!
0'
#251020000000
1!
b0 %
1'
b0 +
#251030000000
0!
0'
#251040000000
1!
1$
b1 %
1'
1*
b1 +
#251050000000
0!
0'
#251060000000
1!
b10 %
1'
b10 +
#251070000000
0!
0'
#251080000000
1!
b11 %
1'
b11 +
#251090000000
0!
0'
#251100000000
1!
b100 %
1'
b100 +
#251110000000
0!
0'
#251120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#251130000000
0!
0'
#251140000000
1!
0$
b110 %
1'
0*
b110 +
#251150000000
0!
0'
#251160000000
1!
b111 %
1'
b111 +
#251170000000
0!
0'
#251180000000
1!
b1000 %
1'
b1000 +
#251190000000
0!
0'
#251200000000
1!
b1001 %
1'
b1001 +
#251210000000
0!
0'
#251220000000
1!
b0 %
1'
b0 +
#251230000000
0!
0'
#251240000000
1!
1$
b1 %
1'
1*
b1 +
#251250000000
0!
0'
#251260000000
1!
b10 %
1'
b10 +
#251270000000
0!
0'
#251280000000
1!
b11 %
1'
b11 +
#251290000000
0!
0'
#251300000000
1!
b100 %
1'
b100 +
#251310000000
0!
0'
#251320000000
1!
b101 %
1'
b101 +
#251330000000
1"
1(
#251340000000
0!
0"
b100 &
0'
0(
b100 ,
#251350000000
1!
b110 %
1'
b110 +
#251360000000
0!
0'
#251370000000
1!
b111 %
1'
b111 +
#251380000000
0!
0'
#251390000000
1!
0$
b1000 %
1'
0*
b1000 +
#251400000000
0!
0'
#251410000000
1!
b1001 %
1'
b1001 +
#251420000000
0!
0'
#251430000000
1!
b0 %
1'
b0 +
#251440000000
0!
0'
#251450000000
1!
1$
b1 %
1'
1*
b1 +
#251460000000
0!
0'
#251470000000
1!
b10 %
1'
b10 +
#251480000000
0!
0'
#251490000000
1!
b11 %
1'
b11 +
#251500000000
0!
0'
#251510000000
1!
b100 %
1'
b100 +
#251520000000
0!
0'
#251530000000
1!
b101 %
1'
b101 +
#251540000000
0!
0'
#251550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#251560000000
0!
0'
#251570000000
1!
b111 %
1'
b111 +
#251580000000
0!
0'
#251590000000
1!
b1000 %
1'
b1000 +
#251600000000
0!
0'
#251610000000
1!
b1001 %
1'
b1001 +
#251620000000
0!
0'
#251630000000
1!
b0 %
1'
b0 +
#251640000000
0!
0'
#251650000000
1!
1$
b1 %
1'
1*
b1 +
#251660000000
0!
0'
#251670000000
1!
b10 %
1'
b10 +
#251680000000
0!
0'
#251690000000
1!
b11 %
1'
b11 +
#251700000000
0!
0'
#251710000000
1!
b100 %
1'
b100 +
#251720000000
0!
0'
#251730000000
1!
b101 %
1'
b101 +
#251740000000
0!
0'
#251750000000
1!
0$
b110 %
1'
0*
b110 +
#251760000000
1"
1(
#251770000000
0!
0"
b100 &
0'
0(
b100 ,
#251780000000
1!
1$
b111 %
1'
1*
b111 +
#251790000000
0!
0'
#251800000000
1!
0$
b1000 %
1'
0*
b1000 +
#251810000000
0!
0'
#251820000000
1!
b1001 %
1'
b1001 +
#251830000000
0!
0'
#251840000000
1!
b0 %
1'
b0 +
#251850000000
0!
0'
#251860000000
1!
1$
b1 %
1'
1*
b1 +
#251870000000
0!
0'
#251880000000
1!
b10 %
1'
b10 +
#251890000000
0!
0'
#251900000000
1!
b11 %
1'
b11 +
#251910000000
0!
0'
#251920000000
1!
b100 %
1'
b100 +
#251930000000
0!
0'
#251940000000
1!
b101 %
1'
b101 +
#251950000000
0!
0'
#251960000000
1!
b110 %
1'
b110 +
#251970000000
0!
0'
#251980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#251990000000
0!
0'
#252000000000
1!
b1000 %
1'
b1000 +
#252010000000
0!
0'
#252020000000
1!
b1001 %
1'
b1001 +
#252030000000
0!
0'
#252040000000
1!
b0 %
1'
b0 +
#252050000000
0!
0'
#252060000000
1!
1$
b1 %
1'
1*
b1 +
#252070000000
0!
0'
#252080000000
1!
b10 %
1'
b10 +
#252090000000
0!
0'
#252100000000
1!
b11 %
1'
b11 +
#252110000000
0!
0'
#252120000000
1!
b100 %
1'
b100 +
#252130000000
0!
0'
#252140000000
1!
b101 %
1'
b101 +
#252150000000
0!
0'
#252160000000
1!
0$
b110 %
1'
0*
b110 +
#252170000000
0!
0'
#252180000000
1!
b111 %
1'
b111 +
#252190000000
1"
1(
#252200000000
0!
0"
b100 &
0'
0(
b100 ,
#252210000000
1!
b1000 %
1'
b1000 +
#252220000000
0!
0'
#252230000000
1!
b1001 %
1'
b1001 +
#252240000000
0!
0'
#252250000000
1!
b0 %
1'
b0 +
#252260000000
0!
0'
#252270000000
1!
1$
b1 %
1'
1*
b1 +
#252280000000
0!
0'
#252290000000
1!
b10 %
1'
b10 +
#252300000000
0!
0'
#252310000000
1!
b11 %
1'
b11 +
#252320000000
0!
0'
#252330000000
1!
b100 %
1'
b100 +
#252340000000
0!
0'
#252350000000
1!
b101 %
1'
b101 +
#252360000000
0!
0'
#252370000000
1!
b110 %
1'
b110 +
#252380000000
0!
0'
#252390000000
1!
b111 %
1'
b111 +
#252400000000
0!
0'
#252410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#252420000000
0!
0'
#252430000000
1!
b1001 %
1'
b1001 +
#252440000000
0!
0'
#252450000000
1!
b0 %
1'
b0 +
#252460000000
0!
0'
#252470000000
1!
1$
b1 %
1'
1*
b1 +
#252480000000
0!
0'
#252490000000
1!
b10 %
1'
b10 +
#252500000000
0!
0'
#252510000000
1!
b11 %
1'
b11 +
#252520000000
0!
0'
#252530000000
1!
b100 %
1'
b100 +
#252540000000
0!
0'
#252550000000
1!
b101 %
1'
b101 +
#252560000000
0!
0'
#252570000000
1!
0$
b110 %
1'
0*
b110 +
#252580000000
0!
0'
#252590000000
1!
b111 %
1'
b111 +
#252600000000
0!
0'
#252610000000
1!
b1000 %
1'
b1000 +
#252620000000
1"
1(
#252630000000
0!
0"
b100 &
0'
0(
b100 ,
#252640000000
1!
b1001 %
1'
b1001 +
#252650000000
0!
0'
#252660000000
1!
b0 %
1'
b0 +
#252670000000
0!
0'
#252680000000
1!
1$
b1 %
1'
1*
b1 +
#252690000000
0!
0'
#252700000000
1!
b10 %
1'
b10 +
#252710000000
0!
0'
#252720000000
1!
b11 %
1'
b11 +
#252730000000
0!
0'
#252740000000
1!
b100 %
1'
b100 +
#252750000000
0!
0'
#252760000000
1!
b101 %
1'
b101 +
#252770000000
0!
0'
#252780000000
1!
b110 %
1'
b110 +
#252790000000
0!
0'
#252800000000
1!
b111 %
1'
b111 +
#252810000000
0!
0'
#252820000000
1!
0$
b1000 %
1'
0*
b1000 +
#252830000000
0!
0'
#252840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#252850000000
0!
0'
#252860000000
1!
b0 %
1'
b0 +
#252870000000
0!
0'
#252880000000
1!
1$
b1 %
1'
1*
b1 +
#252890000000
0!
0'
#252900000000
1!
b10 %
1'
b10 +
#252910000000
0!
0'
#252920000000
1!
b11 %
1'
b11 +
#252930000000
0!
0'
#252940000000
1!
b100 %
1'
b100 +
#252950000000
0!
0'
#252960000000
1!
b101 %
1'
b101 +
#252970000000
0!
0'
#252980000000
1!
0$
b110 %
1'
0*
b110 +
#252990000000
0!
0'
#253000000000
1!
b111 %
1'
b111 +
#253010000000
0!
0'
#253020000000
1!
b1000 %
1'
b1000 +
#253030000000
0!
0'
#253040000000
1!
b1001 %
1'
b1001 +
#253050000000
1"
1(
#253060000000
0!
0"
b100 &
0'
0(
b100 ,
#253070000000
1!
b0 %
1'
b0 +
#253080000000
0!
0'
#253090000000
1!
1$
b1 %
1'
1*
b1 +
#253100000000
0!
0'
#253110000000
1!
b10 %
1'
b10 +
#253120000000
0!
0'
#253130000000
1!
b11 %
1'
b11 +
#253140000000
0!
0'
#253150000000
1!
b100 %
1'
b100 +
#253160000000
0!
0'
#253170000000
1!
b101 %
1'
b101 +
#253180000000
0!
0'
#253190000000
1!
b110 %
1'
b110 +
#253200000000
0!
0'
#253210000000
1!
b111 %
1'
b111 +
#253220000000
0!
0'
#253230000000
1!
0$
b1000 %
1'
0*
b1000 +
#253240000000
0!
0'
#253250000000
1!
b1001 %
1'
b1001 +
#253260000000
0!
0'
#253270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#253280000000
0!
0'
#253290000000
1!
1$
b1 %
1'
1*
b1 +
#253300000000
0!
0'
#253310000000
1!
b10 %
1'
b10 +
#253320000000
0!
0'
#253330000000
1!
b11 %
1'
b11 +
#253340000000
0!
0'
#253350000000
1!
b100 %
1'
b100 +
#253360000000
0!
0'
#253370000000
1!
b101 %
1'
b101 +
#253380000000
0!
0'
#253390000000
1!
0$
b110 %
1'
0*
b110 +
#253400000000
0!
0'
#253410000000
1!
b111 %
1'
b111 +
#253420000000
0!
0'
#253430000000
1!
b1000 %
1'
b1000 +
#253440000000
0!
0'
#253450000000
1!
b1001 %
1'
b1001 +
#253460000000
0!
0'
#253470000000
1!
b0 %
1'
b0 +
#253480000000
1"
1(
#253490000000
0!
0"
b100 &
0'
0(
b100 ,
#253500000000
1!
1$
b1 %
1'
1*
b1 +
#253510000000
0!
0'
#253520000000
1!
b10 %
1'
b10 +
#253530000000
0!
0'
#253540000000
1!
b11 %
1'
b11 +
#253550000000
0!
0'
#253560000000
1!
b100 %
1'
b100 +
#253570000000
0!
0'
#253580000000
1!
b101 %
1'
b101 +
#253590000000
0!
0'
#253600000000
1!
b110 %
1'
b110 +
#253610000000
0!
0'
#253620000000
1!
b111 %
1'
b111 +
#253630000000
0!
0'
#253640000000
1!
0$
b1000 %
1'
0*
b1000 +
#253650000000
0!
0'
#253660000000
1!
b1001 %
1'
b1001 +
#253670000000
0!
0'
#253680000000
1!
b0 %
1'
b0 +
#253690000000
0!
0'
#253700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#253710000000
0!
0'
#253720000000
1!
b10 %
1'
b10 +
#253730000000
0!
0'
#253740000000
1!
b11 %
1'
b11 +
#253750000000
0!
0'
#253760000000
1!
b100 %
1'
b100 +
#253770000000
0!
0'
#253780000000
1!
b101 %
1'
b101 +
#253790000000
0!
0'
#253800000000
1!
0$
b110 %
1'
0*
b110 +
#253810000000
0!
0'
#253820000000
1!
b111 %
1'
b111 +
#253830000000
0!
0'
#253840000000
1!
b1000 %
1'
b1000 +
#253850000000
0!
0'
#253860000000
1!
b1001 %
1'
b1001 +
#253870000000
0!
0'
#253880000000
1!
b0 %
1'
b0 +
#253890000000
0!
0'
#253900000000
1!
1$
b1 %
1'
1*
b1 +
#253910000000
1"
1(
#253920000000
0!
0"
b100 &
0'
0(
b100 ,
#253930000000
1!
b10 %
1'
b10 +
#253940000000
0!
0'
#253950000000
1!
b11 %
1'
b11 +
#253960000000
0!
0'
#253970000000
1!
b100 %
1'
b100 +
#253980000000
0!
0'
#253990000000
1!
b101 %
1'
b101 +
#254000000000
0!
0'
#254010000000
1!
b110 %
1'
b110 +
#254020000000
0!
0'
#254030000000
1!
b111 %
1'
b111 +
#254040000000
0!
0'
#254050000000
1!
0$
b1000 %
1'
0*
b1000 +
#254060000000
0!
0'
#254070000000
1!
b1001 %
1'
b1001 +
#254080000000
0!
0'
#254090000000
1!
b0 %
1'
b0 +
#254100000000
0!
0'
#254110000000
1!
1$
b1 %
1'
1*
b1 +
#254120000000
0!
0'
#254130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#254140000000
0!
0'
#254150000000
1!
b11 %
1'
b11 +
#254160000000
0!
0'
#254170000000
1!
b100 %
1'
b100 +
#254180000000
0!
0'
#254190000000
1!
b101 %
1'
b101 +
#254200000000
0!
0'
#254210000000
1!
0$
b110 %
1'
0*
b110 +
#254220000000
0!
0'
#254230000000
1!
b111 %
1'
b111 +
#254240000000
0!
0'
#254250000000
1!
b1000 %
1'
b1000 +
#254260000000
0!
0'
#254270000000
1!
b1001 %
1'
b1001 +
#254280000000
0!
0'
#254290000000
1!
b0 %
1'
b0 +
#254300000000
0!
0'
#254310000000
1!
1$
b1 %
1'
1*
b1 +
#254320000000
0!
0'
#254330000000
1!
b10 %
1'
b10 +
#254340000000
1"
1(
#254350000000
0!
0"
b100 &
0'
0(
b100 ,
#254360000000
1!
b11 %
1'
b11 +
#254370000000
0!
0'
#254380000000
1!
b100 %
1'
b100 +
#254390000000
0!
0'
#254400000000
1!
b101 %
1'
b101 +
#254410000000
0!
0'
#254420000000
1!
b110 %
1'
b110 +
#254430000000
0!
0'
#254440000000
1!
b111 %
1'
b111 +
#254450000000
0!
0'
#254460000000
1!
0$
b1000 %
1'
0*
b1000 +
#254470000000
0!
0'
#254480000000
1!
b1001 %
1'
b1001 +
#254490000000
0!
0'
#254500000000
1!
b0 %
1'
b0 +
#254510000000
0!
0'
#254520000000
1!
1$
b1 %
1'
1*
b1 +
#254530000000
0!
0'
#254540000000
1!
b10 %
1'
b10 +
#254550000000
0!
0'
#254560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#254570000000
0!
0'
#254580000000
1!
b100 %
1'
b100 +
#254590000000
0!
0'
#254600000000
1!
b101 %
1'
b101 +
#254610000000
0!
0'
#254620000000
1!
0$
b110 %
1'
0*
b110 +
#254630000000
0!
0'
#254640000000
1!
b111 %
1'
b111 +
#254650000000
0!
0'
#254660000000
1!
b1000 %
1'
b1000 +
#254670000000
0!
0'
#254680000000
1!
b1001 %
1'
b1001 +
#254690000000
0!
0'
#254700000000
1!
b0 %
1'
b0 +
#254710000000
0!
0'
#254720000000
1!
1$
b1 %
1'
1*
b1 +
#254730000000
0!
0'
#254740000000
1!
b10 %
1'
b10 +
#254750000000
0!
0'
#254760000000
1!
b11 %
1'
b11 +
#254770000000
1"
1(
#254780000000
0!
0"
b100 &
0'
0(
b100 ,
#254790000000
1!
b100 %
1'
b100 +
#254800000000
0!
0'
#254810000000
1!
b101 %
1'
b101 +
#254820000000
0!
0'
#254830000000
1!
b110 %
1'
b110 +
#254840000000
0!
0'
#254850000000
1!
b111 %
1'
b111 +
#254860000000
0!
0'
#254870000000
1!
0$
b1000 %
1'
0*
b1000 +
#254880000000
0!
0'
#254890000000
1!
b1001 %
1'
b1001 +
#254900000000
0!
0'
#254910000000
1!
b0 %
1'
b0 +
#254920000000
0!
0'
#254930000000
1!
1$
b1 %
1'
1*
b1 +
#254940000000
0!
0'
#254950000000
1!
b10 %
1'
b10 +
#254960000000
0!
0'
#254970000000
1!
b11 %
1'
b11 +
#254980000000
0!
0'
#254990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#255000000000
0!
0'
#255010000000
1!
b101 %
1'
b101 +
#255020000000
0!
0'
#255030000000
1!
0$
b110 %
1'
0*
b110 +
#255040000000
0!
0'
#255050000000
1!
b111 %
1'
b111 +
#255060000000
0!
0'
#255070000000
1!
b1000 %
1'
b1000 +
#255080000000
0!
0'
#255090000000
1!
b1001 %
1'
b1001 +
#255100000000
0!
0'
#255110000000
1!
b0 %
1'
b0 +
#255120000000
0!
0'
#255130000000
1!
1$
b1 %
1'
1*
b1 +
#255140000000
0!
0'
#255150000000
1!
b10 %
1'
b10 +
#255160000000
0!
0'
#255170000000
1!
b11 %
1'
b11 +
#255180000000
0!
0'
#255190000000
1!
b100 %
1'
b100 +
#255200000000
1"
1(
#255210000000
0!
0"
b100 &
0'
0(
b100 ,
#255220000000
1!
b101 %
1'
b101 +
#255230000000
0!
0'
#255240000000
1!
b110 %
1'
b110 +
#255250000000
0!
0'
#255260000000
1!
b111 %
1'
b111 +
#255270000000
0!
0'
#255280000000
1!
0$
b1000 %
1'
0*
b1000 +
#255290000000
0!
0'
#255300000000
1!
b1001 %
1'
b1001 +
#255310000000
0!
0'
#255320000000
1!
b0 %
1'
b0 +
#255330000000
0!
0'
#255340000000
1!
1$
b1 %
1'
1*
b1 +
#255350000000
0!
0'
#255360000000
1!
b10 %
1'
b10 +
#255370000000
0!
0'
#255380000000
1!
b11 %
1'
b11 +
#255390000000
0!
0'
#255400000000
1!
b100 %
1'
b100 +
#255410000000
0!
0'
#255420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#255430000000
0!
0'
#255440000000
1!
0$
b110 %
1'
0*
b110 +
#255450000000
0!
0'
#255460000000
1!
b111 %
1'
b111 +
#255470000000
0!
0'
#255480000000
1!
b1000 %
1'
b1000 +
#255490000000
0!
0'
#255500000000
1!
b1001 %
1'
b1001 +
#255510000000
0!
0'
#255520000000
1!
b0 %
1'
b0 +
#255530000000
0!
0'
#255540000000
1!
1$
b1 %
1'
1*
b1 +
#255550000000
0!
0'
#255560000000
1!
b10 %
1'
b10 +
#255570000000
0!
0'
#255580000000
1!
b11 %
1'
b11 +
#255590000000
0!
0'
#255600000000
1!
b100 %
1'
b100 +
#255610000000
0!
0'
#255620000000
1!
b101 %
1'
b101 +
#255630000000
1"
1(
#255640000000
0!
0"
b100 &
0'
0(
b100 ,
#255650000000
1!
b110 %
1'
b110 +
#255660000000
0!
0'
#255670000000
1!
b111 %
1'
b111 +
#255680000000
0!
0'
#255690000000
1!
0$
b1000 %
1'
0*
b1000 +
#255700000000
0!
0'
#255710000000
1!
b1001 %
1'
b1001 +
#255720000000
0!
0'
#255730000000
1!
b0 %
1'
b0 +
#255740000000
0!
0'
#255750000000
1!
1$
b1 %
1'
1*
b1 +
#255760000000
0!
0'
#255770000000
1!
b10 %
1'
b10 +
#255780000000
0!
0'
#255790000000
1!
b11 %
1'
b11 +
#255800000000
0!
0'
#255810000000
1!
b100 %
1'
b100 +
#255820000000
0!
0'
#255830000000
1!
b101 %
1'
b101 +
#255840000000
0!
0'
#255850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#255860000000
0!
0'
#255870000000
1!
b111 %
1'
b111 +
#255880000000
0!
0'
#255890000000
1!
b1000 %
1'
b1000 +
#255900000000
0!
0'
#255910000000
1!
b1001 %
1'
b1001 +
#255920000000
0!
0'
#255930000000
1!
b0 %
1'
b0 +
#255940000000
0!
0'
#255950000000
1!
1$
b1 %
1'
1*
b1 +
#255960000000
0!
0'
#255970000000
1!
b10 %
1'
b10 +
#255980000000
0!
0'
#255990000000
1!
b11 %
1'
b11 +
#256000000000
0!
0'
#256010000000
1!
b100 %
1'
b100 +
#256020000000
0!
0'
#256030000000
1!
b101 %
1'
b101 +
#256040000000
0!
0'
#256050000000
1!
0$
b110 %
1'
0*
b110 +
#256060000000
1"
1(
#256070000000
0!
0"
b100 &
0'
0(
b100 ,
#256080000000
1!
1$
b111 %
1'
1*
b111 +
#256090000000
0!
0'
#256100000000
1!
0$
b1000 %
1'
0*
b1000 +
#256110000000
0!
0'
#256120000000
1!
b1001 %
1'
b1001 +
#256130000000
0!
0'
#256140000000
1!
b0 %
1'
b0 +
#256150000000
0!
0'
#256160000000
1!
1$
b1 %
1'
1*
b1 +
#256170000000
0!
0'
#256180000000
1!
b10 %
1'
b10 +
#256190000000
0!
0'
#256200000000
1!
b11 %
1'
b11 +
#256210000000
0!
0'
#256220000000
1!
b100 %
1'
b100 +
#256230000000
0!
0'
#256240000000
1!
b101 %
1'
b101 +
#256250000000
0!
0'
#256260000000
1!
b110 %
1'
b110 +
#256270000000
0!
0'
#256280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#256290000000
0!
0'
#256300000000
1!
b1000 %
1'
b1000 +
#256310000000
0!
0'
#256320000000
1!
b1001 %
1'
b1001 +
#256330000000
0!
0'
#256340000000
1!
b0 %
1'
b0 +
#256350000000
0!
0'
#256360000000
1!
1$
b1 %
1'
1*
b1 +
#256370000000
0!
0'
#256380000000
1!
b10 %
1'
b10 +
#256390000000
0!
0'
#256400000000
1!
b11 %
1'
b11 +
#256410000000
0!
0'
#256420000000
1!
b100 %
1'
b100 +
#256430000000
0!
0'
#256440000000
1!
b101 %
1'
b101 +
#256450000000
0!
0'
#256460000000
1!
0$
b110 %
1'
0*
b110 +
#256470000000
0!
0'
#256480000000
1!
b111 %
1'
b111 +
#256490000000
1"
1(
#256500000000
0!
0"
b100 &
0'
0(
b100 ,
#256510000000
1!
b1000 %
1'
b1000 +
#256520000000
0!
0'
#256530000000
1!
b1001 %
1'
b1001 +
#256540000000
0!
0'
#256550000000
1!
b0 %
1'
b0 +
#256560000000
0!
0'
#256570000000
1!
1$
b1 %
1'
1*
b1 +
#256580000000
0!
0'
#256590000000
1!
b10 %
1'
b10 +
#256600000000
0!
0'
#256610000000
1!
b11 %
1'
b11 +
#256620000000
0!
0'
#256630000000
1!
b100 %
1'
b100 +
#256640000000
0!
0'
#256650000000
1!
b101 %
1'
b101 +
#256660000000
0!
0'
#256670000000
1!
b110 %
1'
b110 +
#256680000000
0!
0'
#256690000000
1!
b111 %
1'
b111 +
#256700000000
0!
0'
#256710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#256720000000
0!
0'
#256730000000
1!
b1001 %
1'
b1001 +
#256740000000
0!
0'
#256750000000
1!
b0 %
1'
b0 +
#256760000000
0!
0'
#256770000000
1!
1$
b1 %
1'
1*
b1 +
#256780000000
0!
0'
#256790000000
1!
b10 %
1'
b10 +
#256800000000
0!
0'
#256810000000
1!
b11 %
1'
b11 +
#256820000000
0!
0'
#256830000000
1!
b100 %
1'
b100 +
#256840000000
0!
0'
#256850000000
1!
b101 %
1'
b101 +
#256860000000
0!
0'
#256870000000
1!
0$
b110 %
1'
0*
b110 +
#256880000000
0!
0'
#256890000000
1!
b111 %
1'
b111 +
#256900000000
0!
0'
#256910000000
1!
b1000 %
1'
b1000 +
#256920000000
1"
1(
#256930000000
0!
0"
b100 &
0'
0(
b100 ,
#256940000000
1!
b1001 %
1'
b1001 +
#256950000000
0!
0'
#256960000000
1!
b0 %
1'
b0 +
#256970000000
0!
0'
#256980000000
1!
1$
b1 %
1'
1*
b1 +
#256990000000
0!
0'
#257000000000
1!
b10 %
1'
b10 +
#257010000000
0!
0'
#257020000000
1!
b11 %
1'
b11 +
#257030000000
0!
0'
#257040000000
1!
b100 %
1'
b100 +
#257050000000
0!
0'
#257060000000
1!
b101 %
1'
b101 +
#257070000000
0!
0'
#257080000000
1!
b110 %
1'
b110 +
#257090000000
0!
0'
#257100000000
1!
b111 %
1'
b111 +
#257110000000
0!
0'
#257120000000
1!
0$
b1000 %
1'
0*
b1000 +
#257130000000
0!
0'
#257140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#257150000000
0!
0'
#257160000000
1!
b0 %
1'
b0 +
#257170000000
0!
0'
#257180000000
1!
1$
b1 %
1'
1*
b1 +
#257190000000
0!
0'
#257200000000
1!
b10 %
1'
b10 +
#257210000000
0!
0'
#257220000000
1!
b11 %
1'
b11 +
#257230000000
0!
0'
#257240000000
1!
b100 %
1'
b100 +
#257250000000
0!
0'
#257260000000
1!
b101 %
1'
b101 +
#257270000000
0!
0'
#257280000000
1!
0$
b110 %
1'
0*
b110 +
#257290000000
0!
0'
#257300000000
1!
b111 %
1'
b111 +
#257310000000
0!
0'
#257320000000
1!
b1000 %
1'
b1000 +
#257330000000
0!
0'
#257340000000
1!
b1001 %
1'
b1001 +
#257350000000
1"
1(
#257360000000
0!
0"
b100 &
0'
0(
b100 ,
#257370000000
1!
b0 %
1'
b0 +
#257380000000
0!
0'
#257390000000
1!
1$
b1 %
1'
1*
b1 +
#257400000000
0!
0'
#257410000000
1!
b10 %
1'
b10 +
#257420000000
0!
0'
#257430000000
1!
b11 %
1'
b11 +
#257440000000
0!
0'
#257450000000
1!
b100 %
1'
b100 +
#257460000000
0!
0'
#257470000000
1!
b101 %
1'
b101 +
#257480000000
0!
0'
#257490000000
1!
b110 %
1'
b110 +
#257500000000
0!
0'
#257510000000
1!
b111 %
1'
b111 +
#257520000000
0!
0'
#257530000000
1!
0$
b1000 %
1'
0*
b1000 +
#257540000000
0!
0'
#257550000000
1!
b1001 %
1'
b1001 +
#257560000000
0!
0'
#257570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#257580000000
0!
0'
#257590000000
1!
1$
b1 %
1'
1*
b1 +
#257600000000
0!
0'
#257610000000
1!
b10 %
1'
b10 +
#257620000000
0!
0'
#257630000000
1!
b11 %
1'
b11 +
#257640000000
0!
0'
#257650000000
1!
b100 %
1'
b100 +
#257660000000
0!
0'
#257670000000
1!
b101 %
1'
b101 +
#257680000000
0!
0'
#257690000000
1!
0$
b110 %
1'
0*
b110 +
#257700000000
0!
0'
#257710000000
1!
b111 %
1'
b111 +
#257720000000
0!
0'
#257730000000
1!
b1000 %
1'
b1000 +
#257740000000
0!
0'
#257750000000
1!
b1001 %
1'
b1001 +
#257760000000
0!
0'
#257770000000
1!
b0 %
1'
b0 +
#257780000000
1"
1(
#257790000000
0!
0"
b100 &
0'
0(
b100 ,
#257800000000
1!
1$
b1 %
1'
1*
b1 +
#257810000000
0!
0'
#257820000000
1!
b10 %
1'
b10 +
#257830000000
0!
0'
#257840000000
1!
b11 %
1'
b11 +
#257850000000
0!
0'
#257860000000
1!
b100 %
1'
b100 +
#257870000000
0!
0'
#257880000000
1!
b101 %
1'
b101 +
#257890000000
0!
0'
#257900000000
1!
b110 %
1'
b110 +
#257910000000
0!
0'
#257920000000
1!
b111 %
1'
b111 +
#257930000000
0!
0'
#257940000000
1!
0$
b1000 %
1'
0*
b1000 +
#257950000000
0!
0'
#257960000000
1!
b1001 %
1'
b1001 +
#257970000000
0!
0'
#257980000000
1!
b0 %
1'
b0 +
#257990000000
0!
0'
#258000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#258010000000
0!
0'
#258020000000
1!
b10 %
1'
b10 +
#258030000000
0!
0'
#258040000000
1!
b11 %
1'
b11 +
#258050000000
0!
0'
#258060000000
1!
b100 %
1'
b100 +
#258070000000
0!
0'
#258080000000
1!
b101 %
1'
b101 +
#258090000000
0!
0'
#258100000000
1!
0$
b110 %
1'
0*
b110 +
#258110000000
0!
0'
#258120000000
1!
b111 %
1'
b111 +
#258130000000
0!
0'
#258140000000
1!
b1000 %
1'
b1000 +
#258150000000
0!
0'
#258160000000
1!
b1001 %
1'
b1001 +
#258170000000
0!
0'
#258180000000
1!
b0 %
1'
b0 +
#258190000000
0!
0'
#258200000000
1!
1$
b1 %
1'
1*
b1 +
#258210000000
1"
1(
#258220000000
0!
0"
b100 &
0'
0(
b100 ,
#258230000000
1!
b10 %
1'
b10 +
#258240000000
0!
0'
#258250000000
1!
b11 %
1'
b11 +
#258260000000
0!
0'
#258270000000
1!
b100 %
1'
b100 +
#258280000000
0!
0'
#258290000000
1!
b101 %
1'
b101 +
#258300000000
0!
0'
#258310000000
1!
b110 %
1'
b110 +
#258320000000
0!
0'
#258330000000
1!
b111 %
1'
b111 +
#258340000000
0!
0'
#258350000000
1!
0$
b1000 %
1'
0*
b1000 +
#258360000000
0!
0'
#258370000000
1!
b1001 %
1'
b1001 +
#258380000000
0!
0'
#258390000000
1!
b0 %
1'
b0 +
#258400000000
0!
0'
#258410000000
1!
1$
b1 %
1'
1*
b1 +
#258420000000
0!
0'
#258430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#258440000000
0!
0'
#258450000000
1!
b11 %
1'
b11 +
#258460000000
0!
0'
#258470000000
1!
b100 %
1'
b100 +
#258480000000
0!
0'
#258490000000
1!
b101 %
1'
b101 +
#258500000000
0!
0'
#258510000000
1!
0$
b110 %
1'
0*
b110 +
#258520000000
0!
0'
#258530000000
1!
b111 %
1'
b111 +
#258540000000
0!
0'
#258550000000
1!
b1000 %
1'
b1000 +
#258560000000
0!
0'
#258570000000
1!
b1001 %
1'
b1001 +
#258580000000
0!
0'
#258590000000
1!
b0 %
1'
b0 +
#258600000000
0!
0'
#258610000000
1!
1$
b1 %
1'
1*
b1 +
#258620000000
0!
0'
#258630000000
1!
b10 %
1'
b10 +
#258640000000
1"
1(
#258650000000
0!
0"
b100 &
0'
0(
b100 ,
#258660000000
1!
b11 %
1'
b11 +
#258670000000
0!
0'
#258680000000
1!
b100 %
1'
b100 +
#258690000000
0!
0'
#258700000000
1!
b101 %
1'
b101 +
#258710000000
0!
0'
#258720000000
1!
b110 %
1'
b110 +
#258730000000
0!
0'
#258740000000
1!
b111 %
1'
b111 +
#258750000000
0!
0'
#258760000000
1!
0$
b1000 %
1'
0*
b1000 +
#258770000000
0!
0'
#258780000000
1!
b1001 %
1'
b1001 +
#258790000000
0!
0'
#258800000000
1!
b0 %
1'
b0 +
#258810000000
0!
0'
#258820000000
1!
1$
b1 %
1'
1*
b1 +
#258830000000
0!
0'
#258840000000
1!
b10 %
1'
b10 +
#258850000000
0!
0'
#258860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#258870000000
0!
0'
#258880000000
1!
b100 %
1'
b100 +
#258890000000
0!
0'
#258900000000
1!
b101 %
1'
b101 +
#258910000000
0!
0'
#258920000000
1!
0$
b110 %
1'
0*
b110 +
#258930000000
0!
0'
#258940000000
1!
b111 %
1'
b111 +
#258950000000
0!
0'
#258960000000
1!
b1000 %
1'
b1000 +
#258970000000
0!
0'
#258980000000
1!
b1001 %
1'
b1001 +
#258990000000
0!
0'
#259000000000
1!
b0 %
1'
b0 +
#259010000000
0!
0'
#259020000000
1!
1$
b1 %
1'
1*
b1 +
#259030000000
0!
0'
#259040000000
1!
b10 %
1'
b10 +
#259050000000
0!
0'
#259060000000
1!
b11 %
1'
b11 +
#259070000000
1"
1(
#259080000000
0!
0"
b100 &
0'
0(
b100 ,
#259090000000
1!
b100 %
1'
b100 +
#259100000000
0!
0'
#259110000000
1!
b101 %
1'
b101 +
#259120000000
0!
0'
#259130000000
1!
b110 %
1'
b110 +
#259140000000
0!
0'
#259150000000
1!
b111 %
1'
b111 +
#259160000000
0!
0'
#259170000000
1!
0$
b1000 %
1'
0*
b1000 +
#259180000000
0!
0'
#259190000000
1!
b1001 %
1'
b1001 +
#259200000000
0!
0'
#259210000000
1!
b0 %
1'
b0 +
#259220000000
0!
0'
#259230000000
1!
1$
b1 %
1'
1*
b1 +
#259240000000
0!
0'
#259250000000
1!
b10 %
1'
b10 +
#259260000000
0!
0'
#259270000000
1!
b11 %
1'
b11 +
#259280000000
0!
0'
#259290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#259300000000
0!
0'
#259310000000
1!
b101 %
1'
b101 +
#259320000000
0!
0'
#259330000000
1!
0$
b110 %
1'
0*
b110 +
#259340000000
0!
0'
#259350000000
1!
b111 %
1'
b111 +
#259360000000
0!
0'
#259370000000
1!
b1000 %
1'
b1000 +
#259380000000
0!
0'
#259390000000
1!
b1001 %
1'
b1001 +
#259400000000
0!
0'
#259410000000
1!
b0 %
1'
b0 +
#259420000000
0!
0'
#259430000000
1!
1$
b1 %
1'
1*
b1 +
#259440000000
0!
0'
#259450000000
1!
b10 %
1'
b10 +
#259460000000
0!
0'
#259470000000
1!
b11 %
1'
b11 +
#259480000000
0!
0'
#259490000000
1!
b100 %
1'
b100 +
#259500000000
1"
1(
#259510000000
0!
0"
b100 &
0'
0(
b100 ,
#259520000000
1!
b101 %
1'
b101 +
#259530000000
0!
0'
#259540000000
1!
b110 %
1'
b110 +
#259550000000
0!
0'
#259560000000
1!
b111 %
1'
b111 +
#259570000000
0!
0'
#259580000000
1!
0$
b1000 %
1'
0*
b1000 +
#259590000000
0!
0'
#259600000000
1!
b1001 %
1'
b1001 +
#259610000000
0!
0'
#259620000000
1!
b0 %
1'
b0 +
#259630000000
0!
0'
#259640000000
1!
1$
b1 %
1'
1*
b1 +
#259650000000
0!
0'
#259660000000
1!
b10 %
1'
b10 +
#259670000000
0!
0'
#259680000000
1!
b11 %
1'
b11 +
#259690000000
0!
0'
#259700000000
1!
b100 %
1'
b100 +
#259710000000
0!
0'
#259720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#259730000000
0!
0'
#259740000000
1!
0$
b110 %
1'
0*
b110 +
#259750000000
0!
0'
#259760000000
1!
b111 %
1'
b111 +
#259770000000
0!
0'
#259780000000
1!
b1000 %
1'
b1000 +
#259790000000
0!
0'
#259800000000
1!
b1001 %
1'
b1001 +
#259810000000
0!
0'
#259820000000
1!
b0 %
1'
b0 +
#259830000000
0!
0'
#259840000000
1!
1$
b1 %
1'
1*
b1 +
#259850000000
0!
0'
#259860000000
1!
b10 %
1'
b10 +
#259870000000
0!
0'
#259880000000
1!
b11 %
1'
b11 +
#259890000000
0!
0'
#259900000000
1!
b100 %
1'
b100 +
#259910000000
0!
0'
#259920000000
1!
b101 %
1'
b101 +
#259930000000
1"
1(
#259940000000
0!
0"
b100 &
0'
0(
b100 ,
#259950000000
1!
b110 %
1'
b110 +
#259960000000
0!
0'
#259970000000
1!
b111 %
1'
b111 +
#259980000000
0!
0'
#259990000000
1!
0$
b1000 %
1'
0*
b1000 +
#260000000000
0!
0'
#260010000000
1!
b1001 %
1'
b1001 +
#260020000000
0!
0'
#260030000000
1!
b0 %
1'
b0 +
#260040000000
0!
0'
#260050000000
1!
1$
b1 %
1'
1*
b1 +
#260060000000
0!
0'
#260070000000
1!
b10 %
1'
b10 +
#260080000000
0!
0'
#260090000000
1!
b11 %
1'
b11 +
#260100000000
0!
0'
#260110000000
1!
b100 %
1'
b100 +
#260120000000
0!
0'
#260130000000
1!
b101 %
1'
b101 +
#260140000000
0!
0'
#260150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#260160000000
0!
0'
#260170000000
1!
b111 %
1'
b111 +
#260180000000
0!
0'
#260190000000
1!
b1000 %
1'
b1000 +
#260200000000
0!
0'
#260210000000
1!
b1001 %
1'
b1001 +
#260220000000
0!
0'
#260230000000
1!
b0 %
1'
b0 +
#260240000000
0!
0'
#260250000000
1!
1$
b1 %
1'
1*
b1 +
#260260000000
0!
0'
#260270000000
1!
b10 %
1'
b10 +
#260280000000
0!
0'
#260290000000
1!
b11 %
1'
b11 +
#260300000000
0!
0'
#260310000000
1!
b100 %
1'
b100 +
#260320000000
0!
0'
#260330000000
1!
b101 %
1'
b101 +
#260340000000
0!
0'
#260350000000
1!
0$
b110 %
1'
0*
b110 +
#260360000000
1"
1(
#260370000000
0!
0"
b100 &
0'
0(
b100 ,
#260380000000
1!
1$
b111 %
1'
1*
b111 +
#260390000000
0!
0'
#260400000000
1!
0$
b1000 %
1'
0*
b1000 +
#260410000000
0!
0'
#260420000000
1!
b1001 %
1'
b1001 +
#260430000000
0!
0'
#260440000000
1!
b0 %
1'
b0 +
#260450000000
0!
0'
#260460000000
1!
1$
b1 %
1'
1*
b1 +
#260470000000
0!
0'
#260480000000
1!
b10 %
1'
b10 +
#260490000000
0!
0'
#260500000000
1!
b11 %
1'
b11 +
#260510000000
0!
0'
#260520000000
1!
b100 %
1'
b100 +
#260530000000
0!
0'
#260540000000
1!
b101 %
1'
b101 +
#260550000000
0!
0'
#260560000000
1!
b110 %
1'
b110 +
#260570000000
0!
0'
#260580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#260590000000
0!
0'
#260600000000
1!
b1000 %
1'
b1000 +
#260610000000
0!
0'
#260620000000
1!
b1001 %
1'
b1001 +
#260630000000
0!
0'
#260640000000
1!
b0 %
1'
b0 +
#260650000000
0!
0'
#260660000000
1!
1$
b1 %
1'
1*
b1 +
#260670000000
0!
0'
#260680000000
1!
b10 %
1'
b10 +
#260690000000
0!
0'
#260700000000
1!
b11 %
1'
b11 +
#260710000000
0!
0'
#260720000000
1!
b100 %
1'
b100 +
#260730000000
0!
0'
#260740000000
1!
b101 %
1'
b101 +
#260750000000
0!
0'
#260760000000
1!
0$
b110 %
1'
0*
b110 +
#260770000000
0!
0'
#260780000000
1!
b111 %
1'
b111 +
#260790000000
1"
1(
#260800000000
0!
0"
b100 &
0'
0(
b100 ,
#260810000000
1!
b1000 %
1'
b1000 +
#260820000000
0!
0'
#260830000000
1!
b1001 %
1'
b1001 +
#260840000000
0!
0'
#260850000000
1!
b0 %
1'
b0 +
#260860000000
0!
0'
#260870000000
1!
1$
b1 %
1'
1*
b1 +
#260880000000
0!
0'
#260890000000
1!
b10 %
1'
b10 +
#260900000000
0!
0'
#260910000000
1!
b11 %
1'
b11 +
#260920000000
0!
0'
#260930000000
1!
b100 %
1'
b100 +
#260940000000
0!
0'
#260950000000
1!
b101 %
1'
b101 +
#260960000000
0!
0'
#260970000000
1!
b110 %
1'
b110 +
#260980000000
0!
0'
#260990000000
1!
b111 %
1'
b111 +
#261000000000
0!
0'
#261010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#261020000000
0!
0'
#261030000000
1!
b1001 %
1'
b1001 +
#261040000000
0!
0'
#261050000000
1!
b0 %
1'
b0 +
#261060000000
0!
0'
#261070000000
1!
1$
b1 %
1'
1*
b1 +
#261080000000
0!
0'
#261090000000
1!
b10 %
1'
b10 +
#261100000000
0!
0'
#261110000000
1!
b11 %
1'
b11 +
#261120000000
0!
0'
#261130000000
1!
b100 %
1'
b100 +
#261140000000
0!
0'
#261150000000
1!
b101 %
1'
b101 +
#261160000000
0!
0'
#261170000000
1!
0$
b110 %
1'
0*
b110 +
#261180000000
0!
0'
#261190000000
1!
b111 %
1'
b111 +
#261200000000
0!
0'
#261210000000
1!
b1000 %
1'
b1000 +
#261220000000
1"
1(
#261230000000
0!
0"
b100 &
0'
0(
b100 ,
#261240000000
1!
b1001 %
1'
b1001 +
#261250000000
0!
0'
#261260000000
1!
b0 %
1'
b0 +
#261270000000
0!
0'
#261280000000
1!
1$
b1 %
1'
1*
b1 +
#261290000000
0!
0'
#261300000000
1!
b10 %
1'
b10 +
#261310000000
0!
0'
#261320000000
1!
b11 %
1'
b11 +
#261330000000
0!
0'
#261340000000
1!
b100 %
1'
b100 +
#261350000000
0!
0'
#261360000000
1!
b101 %
1'
b101 +
#261370000000
0!
0'
#261380000000
1!
b110 %
1'
b110 +
#261390000000
0!
0'
#261400000000
1!
b111 %
1'
b111 +
#261410000000
0!
0'
#261420000000
1!
0$
b1000 %
1'
0*
b1000 +
#261430000000
0!
0'
#261440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#261450000000
0!
0'
#261460000000
1!
b0 %
1'
b0 +
#261470000000
0!
0'
#261480000000
1!
1$
b1 %
1'
1*
b1 +
#261490000000
0!
0'
#261500000000
1!
b10 %
1'
b10 +
#261510000000
0!
0'
#261520000000
1!
b11 %
1'
b11 +
#261530000000
0!
0'
#261540000000
1!
b100 %
1'
b100 +
#261550000000
0!
0'
#261560000000
1!
b101 %
1'
b101 +
#261570000000
0!
0'
#261580000000
1!
0$
b110 %
1'
0*
b110 +
#261590000000
0!
0'
#261600000000
1!
b111 %
1'
b111 +
#261610000000
0!
0'
#261620000000
1!
b1000 %
1'
b1000 +
#261630000000
0!
0'
#261640000000
1!
b1001 %
1'
b1001 +
#261650000000
1"
1(
#261660000000
0!
0"
b100 &
0'
0(
b100 ,
#261670000000
1!
b0 %
1'
b0 +
#261680000000
0!
0'
#261690000000
1!
1$
b1 %
1'
1*
b1 +
#261700000000
0!
0'
#261710000000
1!
b10 %
1'
b10 +
#261720000000
0!
0'
#261730000000
1!
b11 %
1'
b11 +
#261740000000
0!
0'
#261750000000
1!
b100 %
1'
b100 +
#261760000000
0!
0'
#261770000000
1!
b101 %
1'
b101 +
#261780000000
0!
0'
#261790000000
1!
b110 %
1'
b110 +
#261800000000
0!
0'
#261810000000
1!
b111 %
1'
b111 +
#261820000000
0!
0'
#261830000000
1!
0$
b1000 %
1'
0*
b1000 +
#261840000000
0!
0'
#261850000000
1!
b1001 %
1'
b1001 +
#261860000000
0!
0'
#261870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#261880000000
0!
0'
#261890000000
1!
1$
b1 %
1'
1*
b1 +
#261900000000
0!
0'
#261910000000
1!
b10 %
1'
b10 +
#261920000000
0!
0'
#261930000000
1!
b11 %
1'
b11 +
#261940000000
0!
0'
#261950000000
1!
b100 %
1'
b100 +
#261960000000
0!
0'
#261970000000
1!
b101 %
1'
b101 +
#261980000000
0!
0'
#261990000000
1!
0$
b110 %
1'
0*
b110 +
#262000000000
0!
0'
#262010000000
1!
b111 %
1'
b111 +
#262020000000
0!
0'
#262030000000
1!
b1000 %
1'
b1000 +
#262040000000
0!
0'
#262050000000
1!
b1001 %
1'
b1001 +
#262060000000
0!
0'
#262070000000
1!
b0 %
1'
b0 +
#262080000000
1"
1(
#262090000000
0!
0"
b100 &
0'
0(
b100 ,
#262100000000
1!
1$
b1 %
1'
1*
b1 +
#262110000000
0!
0'
#262120000000
1!
b10 %
1'
b10 +
#262130000000
0!
0'
#262140000000
1!
b11 %
1'
b11 +
#262150000000
0!
0'
#262160000000
1!
b100 %
1'
b100 +
#262170000000
0!
0'
#262180000000
1!
b101 %
1'
b101 +
#262190000000
0!
0'
#262200000000
1!
b110 %
1'
b110 +
#262210000000
0!
0'
#262220000000
1!
b111 %
1'
b111 +
#262230000000
0!
0'
#262240000000
1!
0$
b1000 %
1'
0*
b1000 +
#262250000000
0!
0'
#262260000000
1!
b1001 %
1'
b1001 +
#262270000000
0!
0'
#262280000000
1!
b0 %
1'
b0 +
#262290000000
0!
0'
#262300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#262310000000
0!
0'
#262320000000
1!
b10 %
1'
b10 +
#262330000000
0!
0'
#262340000000
1!
b11 %
1'
b11 +
#262350000000
0!
0'
#262360000000
1!
b100 %
1'
b100 +
#262370000000
0!
0'
#262380000000
1!
b101 %
1'
b101 +
#262390000000
0!
0'
#262400000000
1!
0$
b110 %
1'
0*
b110 +
#262410000000
0!
0'
#262420000000
1!
b111 %
1'
b111 +
#262430000000
0!
0'
#262440000000
1!
b1000 %
1'
b1000 +
#262450000000
0!
0'
#262460000000
1!
b1001 %
1'
b1001 +
#262470000000
0!
0'
#262480000000
1!
b0 %
1'
b0 +
#262490000000
0!
0'
#262500000000
1!
1$
b1 %
1'
1*
b1 +
#262510000000
1"
1(
#262520000000
0!
0"
b100 &
0'
0(
b100 ,
#262530000000
1!
b10 %
1'
b10 +
#262540000000
0!
0'
#262550000000
1!
b11 %
1'
b11 +
#262560000000
0!
0'
#262570000000
1!
b100 %
1'
b100 +
#262580000000
0!
0'
#262590000000
1!
b101 %
1'
b101 +
#262600000000
0!
0'
#262610000000
1!
b110 %
1'
b110 +
#262620000000
0!
0'
#262630000000
1!
b111 %
1'
b111 +
#262640000000
0!
0'
#262650000000
1!
0$
b1000 %
1'
0*
b1000 +
#262660000000
0!
0'
#262670000000
1!
b1001 %
1'
b1001 +
#262680000000
0!
0'
#262690000000
1!
b0 %
1'
b0 +
#262700000000
0!
0'
#262710000000
1!
1$
b1 %
1'
1*
b1 +
#262720000000
0!
0'
#262730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#262740000000
0!
0'
#262750000000
1!
b11 %
1'
b11 +
#262760000000
0!
0'
#262770000000
1!
b100 %
1'
b100 +
#262780000000
0!
0'
#262790000000
1!
b101 %
1'
b101 +
#262800000000
0!
0'
#262810000000
1!
0$
b110 %
1'
0*
b110 +
#262820000000
0!
0'
#262830000000
1!
b111 %
1'
b111 +
#262840000000
0!
0'
#262850000000
1!
b1000 %
1'
b1000 +
#262860000000
0!
0'
#262870000000
1!
b1001 %
1'
b1001 +
#262880000000
0!
0'
#262890000000
1!
b0 %
1'
b0 +
#262900000000
0!
0'
#262910000000
1!
1$
b1 %
1'
1*
b1 +
#262920000000
0!
0'
#262930000000
1!
b10 %
1'
b10 +
#262940000000
1"
1(
#262950000000
0!
0"
b100 &
0'
0(
b100 ,
#262960000000
1!
b11 %
1'
b11 +
#262970000000
0!
0'
#262980000000
1!
b100 %
1'
b100 +
#262990000000
0!
0'
#263000000000
1!
b101 %
1'
b101 +
#263010000000
0!
0'
#263020000000
1!
b110 %
1'
b110 +
#263030000000
0!
0'
#263040000000
1!
b111 %
1'
b111 +
#263050000000
0!
0'
#263060000000
1!
0$
b1000 %
1'
0*
b1000 +
#263070000000
0!
0'
#263080000000
1!
b1001 %
1'
b1001 +
#263090000000
0!
0'
#263100000000
1!
b0 %
1'
b0 +
#263110000000
0!
0'
#263120000000
1!
1$
b1 %
1'
1*
b1 +
#263130000000
0!
0'
#263140000000
1!
b10 %
1'
b10 +
#263150000000
0!
0'
#263160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#263170000000
0!
0'
#263180000000
1!
b100 %
1'
b100 +
#263190000000
0!
0'
#263200000000
1!
b101 %
1'
b101 +
#263210000000
0!
0'
#263220000000
1!
0$
b110 %
1'
0*
b110 +
#263230000000
0!
0'
#263240000000
1!
b111 %
1'
b111 +
#263250000000
0!
0'
#263260000000
1!
b1000 %
1'
b1000 +
#263270000000
0!
0'
#263280000000
1!
b1001 %
1'
b1001 +
#263290000000
0!
0'
#263300000000
1!
b0 %
1'
b0 +
#263310000000
0!
0'
#263320000000
1!
1$
b1 %
1'
1*
b1 +
#263330000000
0!
0'
#263340000000
1!
b10 %
1'
b10 +
#263350000000
0!
0'
#263360000000
1!
b11 %
1'
b11 +
#263370000000
1"
1(
#263380000000
0!
0"
b100 &
0'
0(
b100 ,
#263390000000
1!
b100 %
1'
b100 +
#263400000000
0!
0'
#263410000000
1!
b101 %
1'
b101 +
#263420000000
0!
0'
#263430000000
1!
b110 %
1'
b110 +
#263440000000
0!
0'
#263450000000
1!
b111 %
1'
b111 +
#263460000000
0!
0'
#263470000000
1!
0$
b1000 %
1'
0*
b1000 +
#263480000000
0!
0'
#263490000000
1!
b1001 %
1'
b1001 +
#263500000000
0!
0'
#263510000000
1!
b0 %
1'
b0 +
#263520000000
0!
0'
#263530000000
1!
1$
b1 %
1'
1*
b1 +
#263540000000
0!
0'
#263550000000
1!
b10 %
1'
b10 +
#263560000000
0!
0'
#263570000000
1!
b11 %
1'
b11 +
#263580000000
0!
0'
#263590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#263600000000
0!
0'
#263610000000
1!
b101 %
1'
b101 +
#263620000000
0!
0'
#263630000000
1!
0$
b110 %
1'
0*
b110 +
#263640000000
0!
0'
#263650000000
1!
b111 %
1'
b111 +
#263660000000
0!
0'
#263670000000
1!
b1000 %
1'
b1000 +
#263680000000
0!
0'
#263690000000
1!
b1001 %
1'
b1001 +
#263700000000
0!
0'
#263710000000
1!
b0 %
1'
b0 +
#263720000000
0!
0'
#263730000000
1!
1$
b1 %
1'
1*
b1 +
#263740000000
0!
0'
#263750000000
1!
b10 %
1'
b10 +
#263760000000
0!
0'
#263770000000
1!
b11 %
1'
b11 +
#263780000000
0!
0'
#263790000000
1!
b100 %
1'
b100 +
#263800000000
1"
1(
#263810000000
0!
0"
b100 &
0'
0(
b100 ,
#263820000000
1!
b101 %
1'
b101 +
#263830000000
0!
0'
#263840000000
1!
b110 %
1'
b110 +
#263850000000
0!
0'
#263860000000
1!
b111 %
1'
b111 +
#263870000000
0!
0'
#263880000000
1!
0$
b1000 %
1'
0*
b1000 +
#263890000000
0!
0'
#263900000000
1!
b1001 %
1'
b1001 +
#263910000000
0!
0'
#263920000000
1!
b0 %
1'
b0 +
#263930000000
0!
0'
#263940000000
1!
1$
b1 %
1'
1*
b1 +
#263950000000
0!
0'
#263960000000
1!
b10 %
1'
b10 +
#263970000000
0!
0'
#263980000000
1!
b11 %
1'
b11 +
#263990000000
0!
0'
#264000000000
1!
b100 %
1'
b100 +
#264010000000
0!
0'
#264020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#264030000000
0!
0'
#264040000000
1!
0$
b110 %
1'
0*
b110 +
#264050000000
0!
0'
#264060000000
1!
b111 %
1'
b111 +
#264070000000
0!
0'
#264080000000
1!
b1000 %
1'
b1000 +
#264090000000
0!
0'
#264100000000
1!
b1001 %
1'
b1001 +
#264110000000
0!
0'
#264120000000
1!
b0 %
1'
b0 +
#264130000000
0!
0'
#264140000000
1!
1$
b1 %
1'
1*
b1 +
#264150000000
0!
0'
#264160000000
1!
b10 %
1'
b10 +
#264170000000
0!
0'
#264180000000
1!
b11 %
1'
b11 +
#264190000000
0!
0'
#264200000000
1!
b100 %
1'
b100 +
#264210000000
0!
0'
#264220000000
1!
b101 %
1'
b101 +
#264230000000
1"
1(
#264240000000
0!
0"
b100 &
0'
0(
b100 ,
#264250000000
1!
b110 %
1'
b110 +
#264260000000
0!
0'
#264270000000
1!
b111 %
1'
b111 +
#264280000000
0!
0'
#264290000000
1!
0$
b1000 %
1'
0*
b1000 +
#264300000000
0!
0'
#264310000000
1!
b1001 %
1'
b1001 +
#264320000000
0!
0'
#264330000000
1!
b0 %
1'
b0 +
#264340000000
0!
0'
#264350000000
1!
1$
b1 %
1'
1*
b1 +
#264360000000
0!
0'
#264370000000
1!
b10 %
1'
b10 +
#264380000000
0!
0'
#264390000000
1!
b11 %
1'
b11 +
#264400000000
0!
0'
#264410000000
1!
b100 %
1'
b100 +
#264420000000
0!
0'
#264430000000
1!
b101 %
1'
b101 +
#264440000000
0!
0'
#264450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#264460000000
0!
0'
#264470000000
1!
b111 %
1'
b111 +
#264480000000
0!
0'
#264490000000
1!
b1000 %
1'
b1000 +
#264500000000
0!
0'
#264510000000
1!
b1001 %
1'
b1001 +
#264520000000
0!
0'
#264530000000
1!
b0 %
1'
b0 +
#264540000000
0!
0'
#264550000000
1!
1$
b1 %
1'
1*
b1 +
#264560000000
0!
0'
#264570000000
1!
b10 %
1'
b10 +
#264580000000
0!
0'
#264590000000
1!
b11 %
1'
b11 +
#264600000000
0!
0'
#264610000000
1!
b100 %
1'
b100 +
#264620000000
0!
0'
#264630000000
1!
b101 %
1'
b101 +
#264640000000
0!
0'
#264650000000
1!
0$
b110 %
1'
0*
b110 +
#264660000000
1"
1(
#264670000000
0!
0"
b100 &
0'
0(
b100 ,
#264680000000
1!
1$
b111 %
1'
1*
b111 +
#264690000000
0!
0'
#264700000000
1!
0$
b1000 %
1'
0*
b1000 +
#264710000000
0!
0'
#264720000000
1!
b1001 %
1'
b1001 +
#264730000000
0!
0'
#264740000000
1!
b0 %
1'
b0 +
#264750000000
0!
0'
#264760000000
1!
1$
b1 %
1'
1*
b1 +
#264770000000
0!
0'
#264780000000
1!
b10 %
1'
b10 +
#264790000000
0!
0'
#264800000000
1!
b11 %
1'
b11 +
#264810000000
0!
0'
#264820000000
1!
b100 %
1'
b100 +
#264830000000
0!
0'
#264840000000
1!
b101 %
1'
b101 +
#264850000000
0!
0'
#264860000000
1!
b110 %
1'
b110 +
#264870000000
0!
0'
#264880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#264890000000
0!
0'
#264900000000
1!
b1000 %
1'
b1000 +
#264910000000
0!
0'
#264920000000
1!
b1001 %
1'
b1001 +
#264930000000
0!
0'
#264940000000
1!
b0 %
1'
b0 +
#264950000000
0!
0'
#264960000000
1!
1$
b1 %
1'
1*
b1 +
#264970000000
0!
0'
#264980000000
1!
b10 %
1'
b10 +
#264990000000
0!
0'
#265000000000
1!
b11 %
1'
b11 +
#265010000000
0!
0'
#265020000000
1!
b100 %
1'
b100 +
#265030000000
0!
0'
#265040000000
1!
b101 %
1'
b101 +
#265050000000
0!
0'
#265060000000
1!
0$
b110 %
1'
0*
b110 +
#265070000000
0!
0'
#265080000000
1!
b111 %
1'
b111 +
#265090000000
1"
1(
#265100000000
0!
0"
b100 &
0'
0(
b100 ,
#265110000000
1!
b1000 %
1'
b1000 +
#265120000000
0!
0'
#265130000000
1!
b1001 %
1'
b1001 +
#265140000000
0!
0'
#265150000000
1!
b0 %
1'
b0 +
#265160000000
0!
0'
#265170000000
1!
1$
b1 %
1'
1*
b1 +
#265180000000
0!
0'
#265190000000
1!
b10 %
1'
b10 +
#265200000000
0!
0'
#265210000000
1!
b11 %
1'
b11 +
#265220000000
0!
0'
#265230000000
1!
b100 %
1'
b100 +
#265240000000
0!
0'
#265250000000
1!
b101 %
1'
b101 +
#265260000000
0!
0'
#265270000000
1!
b110 %
1'
b110 +
#265280000000
0!
0'
#265290000000
1!
b111 %
1'
b111 +
#265300000000
0!
0'
#265310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#265320000000
0!
0'
#265330000000
1!
b1001 %
1'
b1001 +
#265340000000
0!
0'
#265350000000
1!
b0 %
1'
b0 +
#265360000000
0!
0'
#265370000000
1!
1$
b1 %
1'
1*
b1 +
#265380000000
0!
0'
#265390000000
1!
b10 %
1'
b10 +
#265400000000
0!
0'
#265410000000
1!
b11 %
1'
b11 +
#265420000000
0!
0'
#265430000000
1!
b100 %
1'
b100 +
#265440000000
0!
0'
#265450000000
1!
b101 %
1'
b101 +
#265460000000
0!
0'
#265470000000
1!
0$
b110 %
1'
0*
b110 +
#265480000000
0!
0'
#265490000000
1!
b111 %
1'
b111 +
#265500000000
0!
0'
#265510000000
1!
b1000 %
1'
b1000 +
#265520000000
1"
1(
#265530000000
0!
0"
b100 &
0'
0(
b100 ,
#265540000000
1!
b1001 %
1'
b1001 +
#265550000000
0!
0'
#265560000000
1!
b0 %
1'
b0 +
#265570000000
0!
0'
#265580000000
1!
1$
b1 %
1'
1*
b1 +
#265590000000
0!
0'
#265600000000
1!
b10 %
1'
b10 +
#265610000000
0!
0'
#265620000000
1!
b11 %
1'
b11 +
#265630000000
0!
0'
#265640000000
1!
b100 %
1'
b100 +
#265650000000
0!
0'
#265660000000
1!
b101 %
1'
b101 +
#265670000000
0!
0'
#265680000000
1!
b110 %
1'
b110 +
#265690000000
0!
0'
#265700000000
1!
b111 %
1'
b111 +
#265710000000
0!
0'
#265720000000
1!
0$
b1000 %
1'
0*
b1000 +
#265730000000
0!
0'
#265740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#265750000000
0!
0'
#265760000000
1!
b0 %
1'
b0 +
#265770000000
0!
0'
#265780000000
1!
1$
b1 %
1'
1*
b1 +
#265790000000
0!
0'
#265800000000
1!
b10 %
1'
b10 +
#265810000000
0!
0'
#265820000000
1!
b11 %
1'
b11 +
#265830000000
0!
0'
#265840000000
1!
b100 %
1'
b100 +
#265850000000
0!
0'
#265860000000
1!
b101 %
1'
b101 +
#265870000000
0!
0'
#265880000000
1!
0$
b110 %
1'
0*
b110 +
#265890000000
0!
0'
#265900000000
1!
b111 %
1'
b111 +
#265910000000
0!
0'
#265920000000
1!
b1000 %
1'
b1000 +
#265930000000
0!
0'
#265940000000
1!
b1001 %
1'
b1001 +
#265950000000
1"
1(
#265960000000
0!
0"
b100 &
0'
0(
b100 ,
#265970000000
1!
b0 %
1'
b0 +
#265980000000
0!
0'
#265990000000
1!
1$
b1 %
1'
1*
b1 +
#266000000000
0!
0'
#266010000000
1!
b10 %
1'
b10 +
#266020000000
0!
0'
#266030000000
1!
b11 %
1'
b11 +
#266040000000
0!
0'
#266050000000
1!
b100 %
1'
b100 +
#266060000000
0!
0'
#266070000000
1!
b101 %
1'
b101 +
#266080000000
0!
0'
#266090000000
1!
b110 %
1'
b110 +
#266100000000
0!
0'
#266110000000
1!
b111 %
1'
b111 +
#266120000000
0!
0'
#266130000000
1!
0$
b1000 %
1'
0*
b1000 +
#266140000000
0!
0'
#266150000000
1!
b1001 %
1'
b1001 +
#266160000000
0!
0'
#266170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#266180000000
0!
0'
#266190000000
1!
1$
b1 %
1'
1*
b1 +
#266200000000
0!
0'
#266210000000
1!
b10 %
1'
b10 +
#266220000000
0!
0'
#266230000000
1!
b11 %
1'
b11 +
#266240000000
0!
0'
#266250000000
1!
b100 %
1'
b100 +
#266260000000
0!
0'
#266270000000
1!
b101 %
1'
b101 +
#266280000000
0!
0'
#266290000000
1!
0$
b110 %
1'
0*
b110 +
#266300000000
0!
0'
#266310000000
1!
b111 %
1'
b111 +
#266320000000
0!
0'
#266330000000
1!
b1000 %
1'
b1000 +
#266340000000
0!
0'
#266350000000
1!
b1001 %
1'
b1001 +
#266360000000
0!
0'
#266370000000
1!
b0 %
1'
b0 +
#266380000000
1"
1(
#266390000000
0!
0"
b100 &
0'
0(
b100 ,
#266400000000
1!
1$
b1 %
1'
1*
b1 +
#266410000000
0!
0'
#266420000000
1!
b10 %
1'
b10 +
#266430000000
0!
0'
#266440000000
1!
b11 %
1'
b11 +
#266450000000
0!
0'
#266460000000
1!
b100 %
1'
b100 +
#266470000000
0!
0'
#266480000000
1!
b101 %
1'
b101 +
#266490000000
0!
0'
#266500000000
1!
b110 %
1'
b110 +
#266510000000
0!
0'
#266520000000
1!
b111 %
1'
b111 +
#266530000000
0!
0'
#266540000000
1!
0$
b1000 %
1'
0*
b1000 +
#266550000000
0!
0'
#266560000000
1!
b1001 %
1'
b1001 +
#266570000000
0!
0'
#266580000000
1!
b0 %
1'
b0 +
#266590000000
0!
0'
#266600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#266610000000
0!
0'
#266620000000
1!
b10 %
1'
b10 +
#266630000000
0!
0'
#266640000000
1!
b11 %
1'
b11 +
#266650000000
0!
0'
#266660000000
1!
b100 %
1'
b100 +
#266670000000
0!
0'
#266680000000
1!
b101 %
1'
b101 +
#266690000000
0!
0'
#266700000000
1!
0$
b110 %
1'
0*
b110 +
#266710000000
0!
0'
#266720000000
1!
b111 %
1'
b111 +
#266730000000
0!
0'
#266740000000
1!
b1000 %
1'
b1000 +
#266750000000
0!
0'
#266760000000
1!
b1001 %
1'
b1001 +
#266770000000
0!
0'
#266780000000
1!
b0 %
1'
b0 +
#266790000000
0!
0'
#266800000000
1!
1$
b1 %
1'
1*
b1 +
#266810000000
1"
1(
#266820000000
0!
0"
b100 &
0'
0(
b100 ,
#266830000000
1!
b10 %
1'
b10 +
#266840000000
0!
0'
#266850000000
1!
b11 %
1'
b11 +
#266860000000
0!
0'
#266870000000
1!
b100 %
1'
b100 +
#266880000000
0!
0'
#266890000000
1!
b101 %
1'
b101 +
#266900000000
0!
0'
#266910000000
1!
b110 %
1'
b110 +
#266920000000
0!
0'
#266930000000
1!
b111 %
1'
b111 +
#266940000000
0!
0'
#266950000000
1!
0$
b1000 %
1'
0*
b1000 +
#266960000000
0!
0'
#266970000000
1!
b1001 %
1'
b1001 +
#266980000000
0!
0'
#266990000000
1!
b0 %
1'
b0 +
#267000000000
0!
0'
#267010000000
1!
1$
b1 %
1'
1*
b1 +
#267020000000
0!
0'
#267030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#267040000000
0!
0'
#267050000000
1!
b11 %
1'
b11 +
#267060000000
0!
0'
#267070000000
1!
b100 %
1'
b100 +
#267080000000
0!
0'
#267090000000
1!
b101 %
1'
b101 +
#267100000000
0!
0'
#267110000000
1!
0$
b110 %
1'
0*
b110 +
#267120000000
0!
0'
#267130000000
1!
b111 %
1'
b111 +
#267140000000
0!
0'
#267150000000
1!
b1000 %
1'
b1000 +
#267160000000
0!
0'
#267170000000
1!
b1001 %
1'
b1001 +
#267180000000
0!
0'
#267190000000
1!
b0 %
1'
b0 +
#267200000000
0!
0'
#267210000000
1!
1$
b1 %
1'
1*
b1 +
#267220000000
0!
0'
#267230000000
1!
b10 %
1'
b10 +
#267240000000
1"
1(
#267250000000
0!
0"
b100 &
0'
0(
b100 ,
#267260000000
1!
b11 %
1'
b11 +
#267270000000
0!
0'
#267280000000
1!
b100 %
1'
b100 +
#267290000000
0!
0'
#267300000000
1!
b101 %
1'
b101 +
#267310000000
0!
0'
#267320000000
1!
b110 %
1'
b110 +
#267330000000
0!
0'
#267340000000
1!
b111 %
1'
b111 +
#267350000000
0!
0'
#267360000000
1!
0$
b1000 %
1'
0*
b1000 +
#267370000000
0!
0'
#267380000000
1!
b1001 %
1'
b1001 +
#267390000000
0!
0'
#267400000000
1!
b0 %
1'
b0 +
#267410000000
0!
0'
#267420000000
1!
1$
b1 %
1'
1*
b1 +
#267430000000
0!
0'
#267440000000
1!
b10 %
1'
b10 +
#267450000000
0!
0'
#267460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#267470000000
0!
0'
#267480000000
1!
b100 %
1'
b100 +
#267490000000
0!
0'
#267500000000
1!
b101 %
1'
b101 +
#267510000000
0!
0'
#267520000000
1!
0$
b110 %
1'
0*
b110 +
#267530000000
0!
0'
#267540000000
1!
b111 %
1'
b111 +
#267550000000
0!
0'
#267560000000
1!
b1000 %
1'
b1000 +
#267570000000
0!
0'
#267580000000
1!
b1001 %
1'
b1001 +
#267590000000
0!
0'
#267600000000
1!
b0 %
1'
b0 +
#267610000000
0!
0'
#267620000000
1!
1$
b1 %
1'
1*
b1 +
#267630000000
0!
0'
#267640000000
1!
b10 %
1'
b10 +
#267650000000
0!
0'
#267660000000
1!
b11 %
1'
b11 +
#267670000000
1"
1(
#267680000000
0!
0"
b100 &
0'
0(
b100 ,
#267690000000
1!
b100 %
1'
b100 +
#267700000000
0!
0'
#267710000000
1!
b101 %
1'
b101 +
#267720000000
0!
0'
#267730000000
1!
b110 %
1'
b110 +
#267740000000
0!
0'
#267750000000
1!
b111 %
1'
b111 +
#267760000000
0!
0'
#267770000000
1!
0$
b1000 %
1'
0*
b1000 +
#267780000000
0!
0'
#267790000000
1!
b1001 %
1'
b1001 +
#267800000000
0!
0'
#267810000000
1!
b0 %
1'
b0 +
#267820000000
0!
0'
#267830000000
1!
1$
b1 %
1'
1*
b1 +
#267840000000
0!
0'
#267850000000
1!
b10 %
1'
b10 +
#267860000000
0!
0'
#267870000000
1!
b11 %
1'
b11 +
#267880000000
0!
0'
#267890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#267900000000
0!
0'
#267910000000
1!
b101 %
1'
b101 +
#267920000000
0!
0'
#267930000000
1!
0$
b110 %
1'
0*
b110 +
#267940000000
0!
0'
#267950000000
1!
b111 %
1'
b111 +
#267960000000
0!
0'
#267970000000
1!
b1000 %
1'
b1000 +
#267980000000
0!
0'
#267990000000
1!
b1001 %
1'
b1001 +
#268000000000
0!
0'
#268010000000
1!
b0 %
1'
b0 +
#268020000000
0!
0'
#268030000000
1!
1$
b1 %
1'
1*
b1 +
#268040000000
0!
0'
#268050000000
1!
b10 %
1'
b10 +
#268060000000
0!
0'
#268070000000
1!
b11 %
1'
b11 +
#268080000000
0!
0'
#268090000000
1!
b100 %
1'
b100 +
#268100000000
1"
1(
#268110000000
0!
0"
b100 &
0'
0(
b100 ,
#268120000000
1!
b101 %
1'
b101 +
#268130000000
0!
0'
#268140000000
1!
b110 %
1'
b110 +
#268150000000
0!
0'
#268160000000
1!
b111 %
1'
b111 +
#268170000000
0!
0'
#268180000000
1!
0$
b1000 %
1'
0*
b1000 +
#268190000000
0!
0'
#268200000000
1!
b1001 %
1'
b1001 +
#268210000000
0!
0'
#268220000000
1!
b0 %
1'
b0 +
#268230000000
0!
0'
#268240000000
1!
1$
b1 %
1'
1*
b1 +
#268250000000
0!
0'
#268260000000
1!
b10 %
1'
b10 +
#268270000000
0!
0'
#268280000000
1!
b11 %
1'
b11 +
#268290000000
0!
0'
#268300000000
1!
b100 %
1'
b100 +
#268310000000
0!
0'
#268320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#268330000000
0!
0'
#268340000000
1!
0$
b110 %
1'
0*
b110 +
#268350000000
0!
0'
#268360000000
1!
b111 %
1'
b111 +
#268370000000
0!
0'
#268380000000
1!
b1000 %
1'
b1000 +
#268390000000
0!
0'
#268400000000
1!
b1001 %
1'
b1001 +
#268410000000
0!
0'
#268420000000
1!
b0 %
1'
b0 +
#268430000000
0!
0'
#268440000000
1!
1$
b1 %
1'
1*
b1 +
#268450000000
0!
0'
#268460000000
1!
b10 %
1'
b10 +
#268470000000
0!
0'
#268480000000
1!
b11 %
1'
b11 +
#268490000000
0!
0'
#268500000000
1!
b100 %
1'
b100 +
#268510000000
0!
0'
#268520000000
1!
b101 %
1'
b101 +
#268530000000
1"
1(
#268540000000
0!
0"
b100 &
0'
0(
b100 ,
#268550000000
1!
b110 %
1'
b110 +
#268560000000
0!
0'
#268570000000
1!
b111 %
1'
b111 +
#268580000000
0!
0'
#268590000000
1!
0$
b1000 %
1'
0*
b1000 +
#268600000000
0!
0'
#268610000000
1!
b1001 %
1'
b1001 +
#268620000000
0!
0'
#268630000000
1!
b0 %
1'
b0 +
#268640000000
0!
0'
#268650000000
1!
1$
b1 %
1'
1*
b1 +
#268660000000
0!
0'
#268670000000
1!
b10 %
1'
b10 +
#268680000000
0!
0'
#268690000000
1!
b11 %
1'
b11 +
#268700000000
0!
0'
#268710000000
1!
b100 %
1'
b100 +
#268720000000
0!
0'
#268730000000
1!
b101 %
1'
b101 +
#268740000000
0!
0'
#268750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#268760000000
0!
0'
#268770000000
1!
b111 %
1'
b111 +
#268780000000
0!
0'
#268790000000
1!
b1000 %
1'
b1000 +
#268800000000
0!
0'
#268810000000
1!
b1001 %
1'
b1001 +
#268820000000
0!
0'
#268830000000
1!
b0 %
1'
b0 +
#268840000000
0!
0'
#268850000000
1!
1$
b1 %
1'
1*
b1 +
#268860000000
0!
0'
#268870000000
1!
b10 %
1'
b10 +
#268880000000
0!
0'
#268890000000
1!
b11 %
1'
b11 +
#268900000000
0!
0'
#268910000000
1!
b100 %
1'
b100 +
#268920000000
0!
0'
#268930000000
1!
b101 %
1'
b101 +
#268940000000
0!
0'
#268950000000
1!
0$
b110 %
1'
0*
b110 +
#268960000000
1"
1(
#268970000000
0!
0"
b100 &
0'
0(
b100 ,
#268980000000
1!
1$
b111 %
1'
1*
b111 +
#268990000000
0!
0'
#269000000000
1!
0$
b1000 %
1'
0*
b1000 +
#269010000000
0!
0'
#269020000000
1!
b1001 %
1'
b1001 +
#269030000000
0!
0'
#269040000000
1!
b0 %
1'
b0 +
#269050000000
0!
0'
#269060000000
1!
1$
b1 %
1'
1*
b1 +
#269070000000
0!
0'
#269080000000
1!
b10 %
1'
b10 +
#269090000000
0!
0'
#269100000000
1!
b11 %
1'
b11 +
#269110000000
0!
0'
#269120000000
1!
b100 %
1'
b100 +
#269130000000
0!
0'
#269140000000
1!
b101 %
1'
b101 +
#269150000000
0!
0'
#269160000000
1!
b110 %
1'
b110 +
#269170000000
0!
0'
#269180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#269190000000
0!
0'
#269200000000
1!
b1000 %
1'
b1000 +
#269210000000
0!
0'
#269220000000
1!
b1001 %
1'
b1001 +
#269230000000
0!
0'
#269240000000
1!
b0 %
1'
b0 +
#269250000000
0!
0'
#269260000000
1!
1$
b1 %
1'
1*
b1 +
#269270000000
0!
0'
#269280000000
1!
b10 %
1'
b10 +
#269290000000
0!
0'
#269300000000
1!
b11 %
1'
b11 +
#269310000000
0!
0'
#269320000000
1!
b100 %
1'
b100 +
#269330000000
0!
0'
#269340000000
1!
b101 %
1'
b101 +
#269350000000
0!
0'
#269360000000
1!
0$
b110 %
1'
0*
b110 +
#269370000000
0!
0'
#269380000000
1!
b111 %
1'
b111 +
#269390000000
1"
1(
#269400000000
0!
0"
b100 &
0'
0(
b100 ,
#269410000000
1!
b1000 %
1'
b1000 +
#269420000000
0!
0'
#269430000000
1!
b1001 %
1'
b1001 +
#269440000000
0!
0'
#269450000000
1!
b0 %
1'
b0 +
#269460000000
0!
0'
#269470000000
1!
1$
b1 %
1'
1*
b1 +
#269480000000
0!
0'
#269490000000
1!
b10 %
1'
b10 +
#269500000000
0!
0'
#269510000000
1!
b11 %
1'
b11 +
#269520000000
0!
0'
#269530000000
1!
b100 %
1'
b100 +
#269540000000
0!
0'
#269550000000
1!
b101 %
1'
b101 +
#269560000000
0!
0'
#269570000000
1!
b110 %
1'
b110 +
#269580000000
0!
0'
#269590000000
1!
b111 %
1'
b111 +
#269600000000
0!
0'
#269610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#269620000000
0!
0'
#269630000000
1!
b1001 %
1'
b1001 +
#269640000000
0!
0'
#269650000000
1!
b0 %
1'
b0 +
#269660000000
0!
0'
#269670000000
1!
1$
b1 %
1'
1*
b1 +
#269680000000
0!
0'
#269690000000
1!
b10 %
1'
b10 +
#269700000000
0!
0'
#269710000000
1!
b11 %
1'
b11 +
#269720000000
0!
0'
#269730000000
1!
b100 %
1'
b100 +
#269740000000
0!
0'
#269750000000
1!
b101 %
1'
b101 +
#269760000000
0!
0'
#269770000000
1!
0$
b110 %
1'
0*
b110 +
#269780000000
0!
0'
#269790000000
1!
b111 %
1'
b111 +
#269800000000
0!
0'
#269810000000
1!
b1000 %
1'
b1000 +
#269820000000
1"
1(
#269830000000
0!
0"
b100 &
0'
0(
b100 ,
#269840000000
1!
b1001 %
1'
b1001 +
#269850000000
0!
0'
#269860000000
1!
b0 %
1'
b0 +
#269870000000
0!
0'
#269880000000
1!
1$
b1 %
1'
1*
b1 +
#269890000000
0!
0'
#269900000000
1!
b10 %
1'
b10 +
#269910000000
0!
0'
#269920000000
1!
b11 %
1'
b11 +
#269930000000
0!
0'
#269940000000
1!
b100 %
1'
b100 +
#269950000000
0!
0'
#269960000000
1!
b101 %
1'
b101 +
#269970000000
0!
0'
#269980000000
1!
b110 %
1'
b110 +
#269990000000
0!
0'
#270000000000
1!
b111 %
1'
b111 +
#270010000000
0!
0'
#270020000000
1!
0$
b1000 %
1'
0*
b1000 +
#270030000000
0!
0'
#270040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#270050000000
0!
0'
#270060000000
1!
b0 %
1'
b0 +
#270070000000
0!
0'
#270080000000
1!
1$
b1 %
1'
1*
b1 +
#270090000000
0!
0'
#270100000000
1!
b10 %
1'
b10 +
#270110000000
0!
0'
#270120000000
1!
b11 %
1'
b11 +
#270130000000
0!
0'
#270140000000
1!
b100 %
1'
b100 +
#270150000000
0!
0'
#270160000000
1!
b101 %
1'
b101 +
#270170000000
0!
0'
#270180000000
1!
0$
b110 %
1'
0*
b110 +
#270190000000
0!
0'
#270200000000
1!
b111 %
1'
b111 +
#270210000000
0!
0'
#270220000000
1!
b1000 %
1'
b1000 +
#270230000000
0!
0'
#270240000000
1!
b1001 %
1'
b1001 +
#270250000000
1"
1(
#270260000000
0!
0"
b100 &
0'
0(
b100 ,
#270270000000
1!
b0 %
1'
b0 +
#270280000000
0!
0'
#270290000000
1!
1$
b1 %
1'
1*
b1 +
#270300000000
0!
0'
#270310000000
1!
b10 %
1'
b10 +
#270320000000
0!
0'
#270330000000
1!
b11 %
1'
b11 +
#270340000000
0!
0'
#270350000000
1!
b100 %
1'
b100 +
#270360000000
0!
0'
#270370000000
1!
b101 %
1'
b101 +
#270380000000
0!
0'
#270390000000
1!
b110 %
1'
b110 +
#270400000000
0!
0'
#270410000000
1!
b111 %
1'
b111 +
#270420000000
0!
0'
#270430000000
1!
0$
b1000 %
1'
0*
b1000 +
#270440000000
0!
0'
#270450000000
1!
b1001 %
1'
b1001 +
#270460000000
0!
0'
#270470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#270480000000
0!
0'
#270490000000
1!
1$
b1 %
1'
1*
b1 +
#270500000000
0!
0'
#270510000000
1!
b10 %
1'
b10 +
#270520000000
0!
0'
#270530000000
1!
b11 %
1'
b11 +
#270540000000
0!
0'
#270550000000
1!
b100 %
1'
b100 +
#270560000000
0!
0'
#270570000000
1!
b101 %
1'
b101 +
#270580000000
0!
0'
#270590000000
1!
0$
b110 %
1'
0*
b110 +
#270600000000
0!
0'
#270610000000
1!
b111 %
1'
b111 +
#270620000000
0!
0'
#270630000000
1!
b1000 %
1'
b1000 +
#270640000000
0!
0'
#270650000000
1!
b1001 %
1'
b1001 +
#270660000000
0!
0'
#270670000000
1!
b0 %
1'
b0 +
#270680000000
1"
1(
#270690000000
0!
0"
b100 &
0'
0(
b100 ,
#270700000000
1!
1$
b1 %
1'
1*
b1 +
#270710000000
0!
0'
#270720000000
1!
b10 %
1'
b10 +
#270730000000
0!
0'
#270740000000
1!
b11 %
1'
b11 +
#270750000000
0!
0'
#270760000000
1!
b100 %
1'
b100 +
#270770000000
0!
0'
#270780000000
1!
b101 %
1'
b101 +
#270790000000
0!
0'
#270800000000
1!
b110 %
1'
b110 +
#270810000000
0!
0'
#270820000000
1!
b111 %
1'
b111 +
#270830000000
0!
0'
#270840000000
1!
0$
b1000 %
1'
0*
b1000 +
#270850000000
0!
0'
#270860000000
1!
b1001 %
1'
b1001 +
#270870000000
0!
0'
#270880000000
1!
b0 %
1'
b0 +
#270890000000
0!
0'
#270900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#270910000000
0!
0'
#270920000000
1!
b10 %
1'
b10 +
#270930000000
0!
0'
#270940000000
1!
b11 %
1'
b11 +
#270950000000
0!
0'
#270960000000
1!
b100 %
1'
b100 +
#270970000000
0!
0'
#270980000000
1!
b101 %
1'
b101 +
#270990000000
0!
0'
#271000000000
1!
0$
b110 %
1'
0*
b110 +
#271010000000
0!
0'
#271020000000
1!
b111 %
1'
b111 +
#271030000000
0!
0'
#271040000000
1!
b1000 %
1'
b1000 +
#271050000000
0!
0'
#271060000000
1!
b1001 %
1'
b1001 +
#271070000000
0!
0'
#271080000000
1!
b0 %
1'
b0 +
#271090000000
0!
0'
#271100000000
1!
1$
b1 %
1'
1*
b1 +
#271110000000
1"
1(
#271120000000
0!
0"
b100 &
0'
0(
b100 ,
#271130000000
1!
b10 %
1'
b10 +
#271140000000
0!
0'
#271150000000
1!
b11 %
1'
b11 +
#271160000000
0!
0'
#271170000000
1!
b100 %
1'
b100 +
#271180000000
0!
0'
#271190000000
1!
b101 %
1'
b101 +
#271200000000
0!
0'
#271210000000
1!
b110 %
1'
b110 +
#271220000000
0!
0'
#271230000000
1!
b111 %
1'
b111 +
#271240000000
0!
0'
#271250000000
1!
0$
b1000 %
1'
0*
b1000 +
#271260000000
0!
0'
#271270000000
1!
b1001 %
1'
b1001 +
#271280000000
0!
0'
#271290000000
1!
b0 %
1'
b0 +
#271300000000
0!
0'
#271310000000
1!
1$
b1 %
1'
1*
b1 +
#271320000000
0!
0'
#271330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#271340000000
0!
0'
#271350000000
1!
b11 %
1'
b11 +
#271360000000
0!
0'
#271370000000
1!
b100 %
1'
b100 +
#271380000000
0!
0'
#271390000000
1!
b101 %
1'
b101 +
#271400000000
0!
0'
#271410000000
1!
0$
b110 %
1'
0*
b110 +
#271420000000
0!
0'
#271430000000
1!
b111 %
1'
b111 +
#271440000000
0!
0'
#271450000000
1!
b1000 %
1'
b1000 +
#271460000000
0!
0'
#271470000000
1!
b1001 %
1'
b1001 +
#271480000000
0!
0'
#271490000000
1!
b0 %
1'
b0 +
#271500000000
0!
0'
#271510000000
1!
1$
b1 %
1'
1*
b1 +
#271520000000
0!
0'
#271530000000
1!
b10 %
1'
b10 +
#271540000000
1"
1(
#271550000000
0!
0"
b100 &
0'
0(
b100 ,
#271560000000
1!
b11 %
1'
b11 +
#271570000000
0!
0'
#271580000000
1!
b100 %
1'
b100 +
#271590000000
0!
0'
#271600000000
1!
b101 %
1'
b101 +
#271610000000
0!
0'
#271620000000
1!
b110 %
1'
b110 +
#271630000000
0!
0'
#271640000000
1!
b111 %
1'
b111 +
#271650000000
0!
0'
#271660000000
1!
0$
b1000 %
1'
0*
b1000 +
#271670000000
0!
0'
#271680000000
1!
b1001 %
1'
b1001 +
#271690000000
0!
0'
#271700000000
1!
b0 %
1'
b0 +
#271710000000
0!
0'
#271720000000
1!
1$
b1 %
1'
1*
b1 +
#271730000000
0!
0'
#271740000000
1!
b10 %
1'
b10 +
#271750000000
0!
0'
#271760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#271770000000
0!
0'
#271780000000
1!
b100 %
1'
b100 +
#271790000000
0!
0'
#271800000000
1!
b101 %
1'
b101 +
#271810000000
0!
0'
#271820000000
1!
0$
b110 %
1'
0*
b110 +
#271830000000
0!
0'
#271840000000
1!
b111 %
1'
b111 +
#271850000000
0!
0'
#271860000000
1!
b1000 %
1'
b1000 +
#271870000000
0!
0'
#271880000000
1!
b1001 %
1'
b1001 +
#271890000000
0!
0'
#271900000000
1!
b0 %
1'
b0 +
#271910000000
0!
0'
#271920000000
1!
1$
b1 %
1'
1*
b1 +
#271930000000
0!
0'
#271940000000
1!
b10 %
1'
b10 +
#271950000000
0!
0'
#271960000000
1!
b11 %
1'
b11 +
#271970000000
1"
1(
#271980000000
0!
0"
b100 &
0'
0(
b100 ,
#271990000000
1!
b100 %
1'
b100 +
#272000000000
0!
0'
#272010000000
1!
b101 %
1'
b101 +
#272020000000
0!
0'
#272030000000
1!
b110 %
1'
b110 +
#272040000000
0!
0'
#272050000000
1!
b111 %
1'
b111 +
#272060000000
0!
0'
#272070000000
1!
0$
b1000 %
1'
0*
b1000 +
#272080000000
0!
0'
#272090000000
1!
b1001 %
1'
b1001 +
#272100000000
0!
0'
#272110000000
1!
b0 %
1'
b0 +
#272120000000
0!
0'
#272130000000
1!
1$
b1 %
1'
1*
b1 +
#272140000000
0!
0'
#272150000000
1!
b10 %
1'
b10 +
#272160000000
0!
0'
#272170000000
1!
b11 %
1'
b11 +
#272180000000
0!
0'
#272190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#272200000000
0!
0'
#272210000000
1!
b101 %
1'
b101 +
#272220000000
0!
0'
#272230000000
1!
0$
b110 %
1'
0*
b110 +
#272240000000
0!
0'
#272250000000
1!
b111 %
1'
b111 +
#272260000000
0!
0'
#272270000000
1!
b1000 %
1'
b1000 +
#272280000000
0!
0'
#272290000000
1!
b1001 %
1'
b1001 +
#272300000000
0!
0'
#272310000000
1!
b0 %
1'
b0 +
#272320000000
0!
0'
#272330000000
1!
1$
b1 %
1'
1*
b1 +
#272340000000
0!
0'
#272350000000
1!
b10 %
1'
b10 +
#272360000000
0!
0'
#272370000000
1!
b11 %
1'
b11 +
#272380000000
0!
0'
#272390000000
1!
b100 %
1'
b100 +
#272400000000
1"
1(
#272410000000
0!
0"
b100 &
0'
0(
b100 ,
#272420000000
1!
b101 %
1'
b101 +
#272430000000
0!
0'
#272440000000
1!
b110 %
1'
b110 +
#272450000000
0!
0'
#272460000000
1!
b111 %
1'
b111 +
#272470000000
0!
0'
#272480000000
1!
0$
b1000 %
1'
0*
b1000 +
#272490000000
0!
0'
#272500000000
1!
b1001 %
1'
b1001 +
#272510000000
0!
0'
#272520000000
1!
b0 %
1'
b0 +
#272530000000
0!
0'
#272540000000
1!
1$
b1 %
1'
1*
b1 +
#272550000000
0!
0'
#272560000000
1!
b10 %
1'
b10 +
#272570000000
0!
0'
#272580000000
1!
b11 %
1'
b11 +
#272590000000
0!
0'
#272600000000
1!
b100 %
1'
b100 +
#272610000000
0!
0'
#272620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#272630000000
0!
0'
#272640000000
1!
0$
b110 %
1'
0*
b110 +
#272650000000
0!
0'
#272660000000
1!
b111 %
1'
b111 +
#272670000000
0!
0'
#272680000000
1!
b1000 %
1'
b1000 +
#272690000000
0!
0'
#272700000000
1!
b1001 %
1'
b1001 +
#272710000000
0!
0'
#272720000000
1!
b0 %
1'
b0 +
#272730000000
0!
0'
#272740000000
1!
1$
b1 %
1'
1*
b1 +
#272750000000
0!
0'
#272760000000
1!
b10 %
1'
b10 +
#272770000000
0!
0'
#272780000000
1!
b11 %
1'
b11 +
#272790000000
0!
0'
#272800000000
1!
b100 %
1'
b100 +
#272810000000
0!
0'
#272820000000
1!
b101 %
1'
b101 +
#272830000000
1"
1(
#272840000000
0!
0"
b100 &
0'
0(
b100 ,
#272850000000
1!
b110 %
1'
b110 +
#272860000000
0!
0'
#272870000000
1!
b111 %
1'
b111 +
#272880000000
0!
0'
#272890000000
1!
0$
b1000 %
1'
0*
b1000 +
#272900000000
0!
0'
#272910000000
1!
b1001 %
1'
b1001 +
#272920000000
0!
0'
#272930000000
1!
b0 %
1'
b0 +
#272940000000
0!
0'
#272950000000
1!
1$
b1 %
1'
1*
b1 +
#272960000000
0!
0'
#272970000000
1!
b10 %
1'
b10 +
#272980000000
0!
0'
#272990000000
1!
b11 %
1'
b11 +
#273000000000
0!
0'
#273010000000
1!
b100 %
1'
b100 +
#273020000000
0!
0'
#273030000000
1!
b101 %
1'
b101 +
#273040000000
0!
0'
#273050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#273060000000
0!
0'
#273070000000
1!
b111 %
1'
b111 +
#273080000000
0!
0'
#273090000000
1!
b1000 %
1'
b1000 +
#273100000000
0!
0'
#273110000000
1!
b1001 %
1'
b1001 +
#273120000000
0!
0'
#273130000000
1!
b0 %
1'
b0 +
#273140000000
0!
0'
#273150000000
1!
1$
b1 %
1'
1*
b1 +
#273160000000
0!
0'
#273170000000
1!
b10 %
1'
b10 +
#273180000000
0!
0'
#273190000000
1!
b11 %
1'
b11 +
#273200000000
0!
0'
#273210000000
1!
b100 %
1'
b100 +
#273220000000
0!
0'
#273230000000
1!
b101 %
1'
b101 +
#273240000000
0!
0'
#273250000000
1!
0$
b110 %
1'
0*
b110 +
#273260000000
1"
1(
#273270000000
0!
0"
b100 &
0'
0(
b100 ,
#273280000000
1!
1$
b111 %
1'
1*
b111 +
#273290000000
0!
0'
#273300000000
1!
0$
b1000 %
1'
0*
b1000 +
#273310000000
0!
0'
#273320000000
1!
b1001 %
1'
b1001 +
#273330000000
0!
0'
#273340000000
1!
b0 %
1'
b0 +
#273350000000
0!
0'
#273360000000
1!
1$
b1 %
1'
1*
b1 +
#273370000000
0!
0'
#273380000000
1!
b10 %
1'
b10 +
#273390000000
0!
0'
#273400000000
1!
b11 %
1'
b11 +
#273410000000
0!
0'
#273420000000
1!
b100 %
1'
b100 +
#273430000000
0!
0'
#273440000000
1!
b101 %
1'
b101 +
#273450000000
0!
0'
#273460000000
1!
b110 %
1'
b110 +
#273470000000
0!
0'
#273480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#273490000000
0!
0'
#273500000000
1!
b1000 %
1'
b1000 +
#273510000000
0!
0'
#273520000000
1!
b1001 %
1'
b1001 +
#273530000000
0!
0'
#273540000000
1!
b0 %
1'
b0 +
#273550000000
0!
0'
#273560000000
1!
1$
b1 %
1'
1*
b1 +
#273570000000
0!
0'
#273580000000
1!
b10 %
1'
b10 +
#273590000000
0!
0'
#273600000000
1!
b11 %
1'
b11 +
#273610000000
0!
0'
#273620000000
1!
b100 %
1'
b100 +
#273630000000
0!
0'
#273640000000
1!
b101 %
1'
b101 +
#273650000000
0!
0'
#273660000000
1!
0$
b110 %
1'
0*
b110 +
#273670000000
0!
0'
#273680000000
1!
b111 %
1'
b111 +
#273690000000
1"
1(
#273700000000
0!
0"
b100 &
0'
0(
b100 ,
#273710000000
1!
b1000 %
1'
b1000 +
#273720000000
0!
0'
#273730000000
1!
b1001 %
1'
b1001 +
#273740000000
0!
0'
#273750000000
1!
b0 %
1'
b0 +
#273760000000
0!
0'
#273770000000
1!
1$
b1 %
1'
1*
b1 +
#273780000000
0!
0'
#273790000000
1!
b10 %
1'
b10 +
#273800000000
0!
0'
#273810000000
1!
b11 %
1'
b11 +
#273820000000
0!
0'
#273830000000
1!
b100 %
1'
b100 +
#273840000000
0!
0'
#273850000000
1!
b101 %
1'
b101 +
#273860000000
0!
0'
#273870000000
1!
b110 %
1'
b110 +
#273880000000
0!
0'
#273890000000
1!
b111 %
1'
b111 +
#273900000000
0!
0'
#273910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#273920000000
0!
0'
#273930000000
1!
b1001 %
1'
b1001 +
#273940000000
0!
0'
#273950000000
1!
b0 %
1'
b0 +
#273960000000
0!
0'
#273970000000
1!
1$
b1 %
1'
1*
b1 +
#273980000000
0!
0'
#273990000000
1!
b10 %
1'
b10 +
#274000000000
0!
0'
#274010000000
1!
b11 %
1'
b11 +
#274020000000
0!
0'
#274030000000
1!
b100 %
1'
b100 +
#274040000000
0!
0'
#274050000000
1!
b101 %
1'
b101 +
#274060000000
0!
0'
#274070000000
1!
0$
b110 %
1'
0*
b110 +
#274080000000
0!
0'
#274090000000
1!
b111 %
1'
b111 +
#274100000000
0!
0'
#274110000000
1!
b1000 %
1'
b1000 +
#274120000000
1"
1(
#274130000000
0!
0"
b100 &
0'
0(
b100 ,
#274140000000
1!
b1001 %
1'
b1001 +
#274150000000
0!
0'
#274160000000
1!
b0 %
1'
b0 +
#274170000000
0!
0'
#274180000000
1!
1$
b1 %
1'
1*
b1 +
#274190000000
0!
0'
#274200000000
1!
b10 %
1'
b10 +
#274210000000
0!
0'
#274220000000
1!
b11 %
1'
b11 +
#274230000000
0!
0'
#274240000000
1!
b100 %
1'
b100 +
#274250000000
0!
0'
#274260000000
1!
b101 %
1'
b101 +
#274270000000
0!
0'
#274280000000
1!
b110 %
1'
b110 +
#274290000000
0!
0'
#274300000000
1!
b111 %
1'
b111 +
#274310000000
0!
0'
#274320000000
1!
0$
b1000 %
1'
0*
b1000 +
#274330000000
0!
0'
#274340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#274350000000
0!
0'
#274360000000
1!
b0 %
1'
b0 +
#274370000000
0!
0'
#274380000000
1!
1$
b1 %
1'
1*
b1 +
#274390000000
0!
0'
#274400000000
1!
b10 %
1'
b10 +
#274410000000
0!
0'
#274420000000
1!
b11 %
1'
b11 +
#274430000000
0!
0'
#274440000000
1!
b100 %
1'
b100 +
#274450000000
0!
0'
#274460000000
1!
b101 %
1'
b101 +
#274470000000
0!
0'
#274480000000
1!
0$
b110 %
1'
0*
b110 +
#274490000000
0!
0'
#274500000000
1!
b111 %
1'
b111 +
#274510000000
0!
0'
#274520000000
1!
b1000 %
1'
b1000 +
#274530000000
0!
0'
#274540000000
1!
b1001 %
1'
b1001 +
#274550000000
1"
1(
#274560000000
0!
0"
b100 &
0'
0(
b100 ,
#274570000000
1!
b0 %
1'
b0 +
#274580000000
0!
0'
#274590000000
1!
1$
b1 %
1'
1*
b1 +
#274600000000
0!
0'
#274610000000
1!
b10 %
1'
b10 +
#274620000000
0!
0'
#274630000000
1!
b11 %
1'
b11 +
#274640000000
0!
0'
#274650000000
1!
b100 %
1'
b100 +
#274660000000
0!
0'
#274670000000
1!
b101 %
1'
b101 +
#274680000000
0!
0'
#274690000000
1!
b110 %
1'
b110 +
#274700000000
0!
0'
#274710000000
1!
b111 %
1'
b111 +
#274720000000
0!
0'
#274730000000
1!
0$
b1000 %
1'
0*
b1000 +
#274740000000
0!
0'
#274750000000
1!
b1001 %
1'
b1001 +
#274760000000
0!
0'
#274770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#274780000000
0!
0'
#274790000000
1!
1$
b1 %
1'
1*
b1 +
#274800000000
0!
0'
#274810000000
1!
b10 %
1'
b10 +
#274820000000
0!
0'
#274830000000
1!
b11 %
1'
b11 +
#274840000000
0!
0'
#274850000000
1!
b100 %
1'
b100 +
#274860000000
0!
0'
#274870000000
1!
b101 %
1'
b101 +
#274880000000
0!
0'
#274890000000
1!
0$
b110 %
1'
0*
b110 +
#274900000000
0!
0'
#274910000000
1!
b111 %
1'
b111 +
#274920000000
0!
0'
#274930000000
1!
b1000 %
1'
b1000 +
#274940000000
0!
0'
#274950000000
1!
b1001 %
1'
b1001 +
#274960000000
0!
0'
#274970000000
1!
b0 %
1'
b0 +
#274980000000
1"
1(
#274990000000
0!
0"
b100 &
0'
0(
b100 ,
#275000000000
1!
1$
b1 %
1'
1*
b1 +
#275010000000
0!
0'
#275020000000
1!
b10 %
1'
b10 +
#275030000000
0!
0'
#275040000000
1!
b11 %
1'
b11 +
#275050000000
0!
0'
#275060000000
1!
b100 %
1'
b100 +
#275070000000
0!
0'
#275080000000
1!
b101 %
1'
b101 +
#275090000000
0!
0'
#275100000000
1!
b110 %
1'
b110 +
#275110000000
0!
0'
#275120000000
1!
b111 %
1'
b111 +
#275130000000
0!
0'
#275140000000
1!
0$
b1000 %
1'
0*
b1000 +
#275150000000
0!
0'
#275160000000
1!
b1001 %
1'
b1001 +
#275170000000
0!
0'
#275180000000
1!
b0 %
1'
b0 +
#275190000000
0!
0'
#275200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#275210000000
0!
0'
#275220000000
1!
b10 %
1'
b10 +
#275230000000
0!
0'
#275240000000
1!
b11 %
1'
b11 +
#275250000000
0!
0'
#275260000000
1!
b100 %
1'
b100 +
#275270000000
0!
0'
#275280000000
1!
b101 %
1'
b101 +
#275290000000
0!
0'
#275300000000
1!
0$
b110 %
1'
0*
b110 +
#275310000000
0!
0'
#275320000000
1!
b111 %
1'
b111 +
#275330000000
0!
0'
#275340000000
1!
b1000 %
1'
b1000 +
#275350000000
0!
0'
#275360000000
1!
b1001 %
1'
b1001 +
#275370000000
0!
0'
#275380000000
1!
b0 %
1'
b0 +
#275390000000
0!
0'
#275400000000
1!
1$
b1 %
1'
1*
b1 +
#275410000000
1"
1(
#275420000000
0!
0"
b100 &
0'
0(
b100 ,
#275430000000
1!
b10 %
1'
b10 +
#275440000000
0!
0'
#275450000000
1!
b11 %
1'
b11 +
#275460000000
0!
0'
#275470000000
1!
b100 %
1'
b100 +
#275480000000
0!
0'
#275490000000
1!
b101 %
1'
b101 +
#275500000000
0!
0'
#275510000000
1!
b110 %
1'
b110 +
#275520000000
0!
0'
#275530000000
1!
b111 %
1'
b111 +
#275540000000
0!
0'
#275550000000
1!
0$
b1000 %
1'
0*
b1000 +
#275560000000
0!
0'
#275570000000
1!
b1001 %
1'
b1001 +
#275580000000
0!
0'
#275590000000
1!
b0 %
1'
b0 +
#275600000000
0!
0'
#275610000000
1!
1$
b1 %
1'
1*
b1 +
#275620000000
0!
0'
#275630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#275640000000
0!
0'
#275650000000
1!
b11 %
1'
b11 +
#275660000000
0!
0'
#275670000000
1!
b100 %
1'
b100 +
#275680000000
0!
0'
#275690000000
1!
b101 %
1'
b101 +
#275700000000
0!
0'
#275710000000
1!
0$
b110 %
1'
0*
b110 +
#275720000000
0!
0'
#275730000000
1!
b111 %
1'
b111 +
#275740000000
0!
0'
#275750000000
1!
b1000 %
1'
b1000 +
#275760000000
0!
0'
#275770000000
1!
b1001 %
1'
b1001 +
#275780000000
0!
0'
#275790000000
1!
b0 %
1'
b0 +
#275800000000
0!
0'
#275810000000
1!
1$
b1 %
1'
1*
b1 +
#275820000000
0!
0'
#275830000000
1!
b10 %
1'
b10 +
#275840000000
1"
1(
#275850000000
0!
0"
b100 &
0'
0(
b100 ,
#275860000000
1!
b11 %
1'
b11 +
#275870000000
0!
0'
#275880000000
1!
b100 %
1'
b100 +
#275890000000
0!
0'
#275900000000
1!
b101 %
1'
b101 +
#275910000000
0!
0'
#275920000000
1!
b110 %
1'
b110 +
#275930000000
0!
0'
#275940000000
1!
b111 %
1'
b111 +
#275950000000
0!
0'
#275960000000
1!
0$
b1000 %
1'
0*
b1000 +
#275970000000
0!
0'
#275980000000
1!
b1001 %
1'
b1001 +
#275990000000
0!
0'
#276000000000
1!
b0 %
1'
b0 +
#276010000000
0!
0'
#276020000000
1!
1$
b1 %
1'
1*
b1 +
#276030000000
0!
0'
#276040000000
1!
b10 %
1'
b10 +
#276050000000
0!
0'
#276060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#276070000000
0!
0'
#276080000000
1!
b100 %
1'
b100 +
#276090000000
0!
0'
#276100000000
1!
b101 %
1'
b101 +
#276110000000
0!
0'
#276120000000
1!
0$
b110 %
1'
0*
b110 +
#276130000000
0!
0'
#276140000000
1!
b111 %
1'
b111 +
#276150000000
0!
0'
#276160000000
1!
b1000 %
1'
b1000 +
#276170000000
0!
0'
#276180000000
1!
b1001 %
1'
b1001 +
#276190000000
0!
0'
#276200000000
1!
b0 %
1'
b0 +
#276210000000
0!
0'
#276220000000
1!
1$
b1 %
1'
1*
b1 +
#276230000000
0!
0'
#276240000000
1!
b10 %
1'
b10 +
#276250000000
0!
0'
#276260000000
1!
b11 %
1'
b11 +
#276270000000
1"
1(
#276280000000
0!
0"
b100 &
0'
0(
b100 ,
#276290000000
1!
b100 %
1'
b100 +
#276300000000
0!
0'
#276310000000
1!
b101 %
1'
b101 +
#276320000000
0!
0'
#276330000000
1!
b110 %
1'
b110 +
#276340000000
0!
0'
#276350000000
1!
b111 %
1'
b111 +
#276360000000
0!
0'
#276370000000
1!
0$
b1000 %
1'
0*
b1000 +
#276380000000
0!
0'
#276390000000
1!
b1001 %
1'
b1001 +
#276400000000
0!
0'
#276410000000
1!
b0 %
1'
b0 +
#276420000000
0!
0'
#276430000000
1!
1$
b1 %
1'
1*
b1 +
#276440000000
0!
0'
#276450000000
1!
b10 %
1'
b10 +
#276460000000
0!
0'
#276470000000
1!
b11 %
1'
b11 +
#276480000000
0!
0'
#276490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#276500000000
0!
0'
#276510000000
1!
b101 %
1'
b101 +
#276520000000
0!
0'
#276530000000
1!
0$
b110 %
1'
0*
b110 +
#276540000000
0!
0'
#276550000000
1!
b111 %
1'
b111 +
#276560000000
0!
0'
#276570000000
1!
b1000 %
1'
b1000 +
#276580000000
0!
0'
#276590000000
1!
b1001 %
1'
b1001 +
#276600000000
0!
0'
#276610000000
1!
b0 %
1'
b0 +
#276620000000
0!
0'
#276630000000
1!
1$
b1 %
1'
1*
b1 +
#276640000000
0!
0'
#276650000000
1!
b10 %
1'
b10 +
#276660000000
0!
0'
#276670000000
1!
b11 %
1'
b11 +
#276680000000
0!
0'
#276690000000
1!
b100 %
1'
b100 +
#276700000000
1"
1(
#276710000000
0!
0"
b100 &
0'
0(
b100 ,
#276720000000
1!
b101 %
1'
b101 +
#276730000000
0!
0'
#276740000000
1!
b110 %
1'
b110 +
#276750000000
0!
0'
#276760000000
1!
b111 %
1'
b111 +
#276770000000
0!
0'
#276780000000
1!
0$
b1000 %
1'
0*
b1000 +
#276790000000
0!
0'
#276800000000
1!
b1001 %
1'
b1001 +
#276810000000
0!
0'
#276820000000
1!
b0 %
1'
b0 +
#276830000000
0!
0'
#276840000000
1!
1$
b1 %
1'
1*
b1 +
#276850000000
0!
0'
#276860000000
1!
b10 %
1'
b10 +
#276870000000
0!
0'
#276880000000
1!
b11 %
1'
b11 +
#276890000000
0!
0'
#276900000000
1!
b100 %
1'
b100 +
#276910000000
0!
0'
#276920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#276930000000
0!
0'
#276940000000
1!
0$
b110 %
1'
0*
b110 +
#276950000000
0!
0'
#276960000000
1!
b111 %
1'
b111 +
#276970000000
0!
0'
#276980000000
1!
b1000 %
1'
b1000 +
#276990000000
0!
0'
#277000000000
1!
b1001 %
1'
b1001 +
#277010000000
0!
0'
#277020000000
1!
b0 %
1'
b0 +
#277030000000
0!
0'
#277040000000
1!
1$
b1 %
1'
1*
b1 +
#277050000000
0!
0'
#277060000000
1!
b10 %
1'
b10 +
#277070000000
0!
0'
#277080000000
1!
b11 %
1'
b11 +
#277090000000
0!
0'
#277100000000
1!
b100 %
1'
b100 +
#277110000000
0!
0'
#277120000000
1!
b101 %
1'
b101 +
#277130000000
1"
1(
#277140000000
0!
0"
b100 &
0'
0(
b100 ,
#277150000000
1!
b110 %
1'
b110 +
#277160000000
0!
0'
#277170000000
1!
b111 %
1'
b111 +
#277180000000
0!
0'
#277190000000
1!
0$
b1000 %
1'
0*
b1000 +
#277200000000
0!
0'
#277210000000
1!
b1001 %
1'
b1001 +
#277220000000
0!
0'
#277230000000
1!
b0 %
1'
b0 +
#277240000000
0!
0'
#277250000000
1!
1$
b1 %
1'
1*
b1 +
#277260000000
0!
0'
#277270000000
1!
b10 %
1'
b10 +
#277280000000
0!
0'
#277290000000
1!
b11 %
1'
b11 +
#277300000000
0!
0'
#277310000000
1!
b100 %
1'
b100 +
#277320000000
0!
0'
#277330000000
1!
b101 %
1'
b101 +
#277340000000
0!
0'
#277350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#277360000000
0!
0'
#277370000000
1!
b111 %
1'
b111 +
#277380000000
0!
0'
#277390000000
1!
b1000 %
1'
b1000 +
#277400000000
0!
0'
#277410000000
1!
b1001 %
1'
b1001 +
#277420000000
0!
0'
#277430000000
1!
b0 %
1'
b0 +
#277440000000
0!
0'
#277450000000
1!
1$
b1 %
1'
1*
b1 +
#277460000000
0!
0'
#277470000000
1!
b10 %
1'
b10 +
#277480000000
0!
0'
#277490000000
1!
b11 %
1'
b11 +
#277500000000
0!
0'
#277510000000
1!
b100 %
1'
b100 +
#277520000000
0!
0'
#277530000000
1!
b101 %
1'
b101 +
#277540000000
0!
0'
#277550000000
1!
0$
b110 %
1'
0*
b110 +
#277560000000
1"
1(
#277570000000
0!
0"
b100 &
0'
0(
b100 ,
#277580000000
1!
1$
b111 %
1'
1*
b111 +
#277590000000
0!
0'
#277600000000
1!
0$
b1000 %
1'
0*
b1000 +
#277610000000
0!
0'
#277620000000
1!
b1001 %
1'
b1001 +
#277630000000
0!
0'
#277640000000
1!
b0 %
1'
b0 +
#277650000000
0!
0'
#277660000000
1!
1$
b1 %
1'
1*
b1 +
#277670000000
0!
0'
#277680000000
1!
b10 %
1'
b10 +
#277690000000
0!
0'
#277700000000
1!
b11 %
1'
b11 +
#277710000000
0!
0'
#277720000000
1!
b100 %
1'
b100 +
#277730000000
0!
0'
#277740000000
1!
b101 %
1'
b101 +
#277750000000
0!
0'
#277760000000
1!
b110 %
1'
b110 +
#277770000000
0!
0'
#277780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#277790000000
0!
0'
#277800000000
1!
b1000 %
1'
b1000 +
#277810000000
0!
0'
#277820000000
1!
b1001 %
1'
b1001 +
#277830000000
0!
0'
#277840000000
1!
b0 %
1'
b0 +
#277850000000
0!
0'
#277860000000
1!
1$
b1 %
1'
1*
b1 +
#277870000000
0!
0'
#277880000000
1!
b10 %
1'
b10 +
#277890000000
0!
0'
#277900000000
1!
b11 %
1'
b11 +
#277910000000
0!
0'
#277920000000
1!
b100 %
1'
b100 +
#277930000000
0!
0'
#277940000000
1!
b101 %
1'
b101 +
#277950000000
0!
0'
#277960000000
1!
0$
b110 %
1'
0*
b110 +
#277970000000
0!
0'
#277980000000
1!
b111 %
1'
b111 +
#277990000000
1"
1(
#278000000000
0!
0"
b100 &
0'
0(
b100 ,
#278010000000
1!
b1000 %
1'
b1000 +
#278020000000
0!
0'
#278030000000
1!
b1001 %
1'
b1001 +
#278040000000
0!
0'
#278050000000
1!
b0 %
1'
b0 +
#278060000000
0!
0'
#278070000000
1!
1$
b1 %
1'
1*
b1 +
#278080000000
0!
0'
#278090000000
1!
b10 %
1'
b10 +
#278100000000
0!
0'
#278110000000
1!
b11 %
1'
b11 +
#278120000000
0!
0'
#278130000000
1!
b100 %
1'
b100 +
#278140000000
0!
0'
#278150000000
1!
b101 %
1'
b101 +
#278160000000
0!
0'
#278170000000
1!
b110 %
1'
b110 +
#278180000000
0!
0'
#278190000000
1!
b111 %
1'
b111 +
#278200000000
0!
0'
#278210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#278220000000
0!
0'
#278230000000
1!
b1001 %
1'
b1001 +
#278240000000
0!
0'
#278250000000
1!
b0 %
1'
b0 +
#278260000000
0!
0'
#278270000000
1!
1$
b1 %
1'
1*
b1 +
#278280000000
0!
0'
#278290000000
1!
b10 %
1'
b10 +
#278300000000
0!
0'
#278310000000
1!
b11 %
1'
b11 +
#278320000000
0!
0'
#278330000000
1!
b100 %
1'
b100 +
#278340000000
0!
0'
#278350000000
1!
b101 %
1'
b101 +
#278360000000
0!
0'
#278370000000
1!
0$
b110 %
1'
0*
b110 +
#278380000000
0!
0'
#278390000000
1!
b111 %
1'
b111 +
#278400000000
0!
0'
#278410000000
1!
b1000 %
1'
b1000 +
#278420000000
1"
1(
#278430000000
0!
0"
b100 &
0'
0(
b100 ,
#278440000000
1!
b1001 %
1'
b1001 +
#278450000000
0!
0'
#278460000000
1!
b0 %
1'
b0 +
#278470000000
0!
0'
#278480000000
1!
1$
b1 %
1'
1*
b1 +
#278490000000
0!
0'
#278500000000
1!
b10 %
1'
b10 +
#278510000000
0!
0'
#278520000000
1!
b11 %
1'
b11 +
#278530000000
0!
0'
#278540000000
1!
b100 %
1'
b100 +
#278550000000
0!
0'
#278560000000
1!
b101 %
1'
b101 +
#278570000000
0!
0'
#278580000000
1!
b110 %
1'
b110 +
#278590000000
0!
0'
#278600000000
1!
b111 %
1'
b111 +
#278610000000
0!
0'
#278620000000
1!
0$
b1000 %
1'
0*
b1000 +
#278630000000
0!
0'
#278640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#278650000000
0!
0'
#278660000000
1!
b0 %
1'
b0 +
#278670000000
0!
0'
#278680000000
1!
1$
b1 %
1'
1*
b1 +
#278690000000
0!
0'
#278700000000
1!
b10 %
1'
b10 +
#278710000000
0!
0'
#278720000000
1!
b11 %
1'
b11 +
#278730000000
0!
0'
#278740000000
1!
b100 %
1'
b100 +
#278750000000
0!
0'
#278760000000
1!
b101 %
1'
b101 +
#278770000000
0!
0'
#278780000000
1!
0$
b110 %
1'
0*
b110 +
#278790000000
0!
0'
#278800000000
1!
b111 %
1'
b111 +
#278810000000
0!
0'
#278820000000
1!
b1000 %
1'
b1000 +
#278830000000
0!
0'
#278840000000
1!
b1001 %
1'
b1001 +
#278850000000
1"
1(
#278860000000
0!
0"
b100 &
0'
0(
b100 ,
#278870000000
1!
b0 %
1'
b0 +
#278880000000
0!
0'
#278890000000
1!
1$
b1 %
1'
1*
b1 +
#278900000000
0!
0'
#278910000000
1!
b10 %
1'
b10 +
#278920000000
0!
0'
#278930000000
1!
b11 %
1'
b11 +
#278940000000
0!
0'
#278950000000
1!
b100 %
1'
b100 +
#278960000000
0!
0'
#278970000000
1!
b101 %
1'
b101 +
#278980000000
0!
0'
#278990000000
1!
b110 %
1'
b110 +
#279000000000
0!
0'
#279010000000
1!
b111 %
1'
b111 +
#279020000000
0!
0'
#279030000000
1!
0$
b1000 %
1'
0*
b1000 +
#279040000000
0!
0'
#279050000000
1!
b1001 %
1'
b1001 +
#279060000000
0!
0'
#279070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#279080000000
0!
0'
#279090000000
1!
1$
b1 %
1'
1*
b1 +
#279100000000
0!
0'
#279110000000
1!
b10 %
1'
b10 +
#279120000000
0!
0'
#279130000000
1!
b11 %
1'
b11 +
#279140000000
0!
0'
#279150000000
1!
b100 %
1'
b100 +
#279160000000
0!
0'
#279170000000
1!
b101 %
1'
b101 +
#279180000000
0!
0'
#279190000000
1!
0$
b110 %
1'
0*
b110 +
#279200000000
0!
0'
#279210000000
1!
b111 %
1'
b111 +
#279220000000
0!
0'
#279230000000
1!
b1000 %
1'
b1000 +
#279240000000
0!
0'
#279250000000
1!
b1001 %
1'
b1001 +
#279260000000
0!
0'
#279270000000
1!
b0 %
1'
b0 +
#279280000000
1"
1(
#279290000000
0!
0"
b100 &
0'
0(
b100 ,
#279300000000
1!
1$
b1 %
1'
1*
b1 +
#279310000000
0!
0'
#279320000000
1!
b10 %
1'
b10 +
#279330000000
0!
0'
#279340000000
1!
b11 %
1'
b11 +
#279350000000
0!
0'
#279360000000
1!
b100 %
1'
b100 +
#279370000000
0!
0'
#279380000000
1!
b101 %
1'
b101 +
#279390000000
0!
0'
#279400000000
1!
b110 %
1'
b110 +
#279410000000
0!
0'
#279420000000
1!
b111 %
1'
b111 +
#279430000000
0!
0'
#279440000000
1!
0$
b1000 %
1'
0*
b1000 +
#279450000000
0!
0'
#279460000000
1!
b1001 %
1'
b1001 +
#279470000000
0!
0'
#279480000000
1!
b0 %
1'
b0 +
#279490000000
0!
0'
#279500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#279510000000
0!
0'
#279520000000
1!
b10 %
1'
b10 +
#279530000000
0!
0'
#279540000000
1!
b11 %
1'
b11 +
#279550000000
0!
0'
#279560000000
1!
b100 %
1'
b100 +
#279570000000
0!
0'
#279580000000
1!
b101 %
1'
b101 +
#279590000000
0!
0'
#279600000000
1!
0$
b110 %
1'
0*
b110 +
#279610000000
0!
0'
#279620000000
1!
b111 %
1'
b111 +
#279630000000
0!
0'
#279640000000
1!
b1000 %
1'
b1000 +
#279650000000
0!
0'
#279660000000
1!
b1001 %
1'
b1001 +
#279670000000
0!
0'
#279680000000
1!
b0 %
1'
b0 +
#279690000000
0!
0'
#279700000000
1!
1$
b1 %
1'
1*
b1 +
#279710000000
1"
1(
#279720000000
0!
0"
b100 &
0'
0(
b100 ,
#279730000000
1!
b10 %
1'
b10 +
#279740000000
0!
0'
#279750000000
1!
b11 %
1'
b11 +
#279760000000
0!
0'
#279770000000
1!
b100 %
1'
b100 +
#279780000000
0!
0'
#279790000000
1!
b101 %
1'
b101 +
#279800000000
0!
0'
#279810000000
1!
b110 %
1'
b110 +
#279820000000
0!
0'
#279830000000
1!
b111 %
1'
b111 +
#279840000000
0!
0'
#279850000000
1!
0$
b1000 %
1'
0*
b1000 +
#279860000000
0!
0'
#279870000000
1!
b1001 %
1'
b1001 +
#279880000000
0!
0'
#279890000000
1!
b0 %
1'
b0 +
#279900000000
0!
0'
#279910000000
1!
1$
b1 %
1'
1*
b1 +
#279920000000
0!
0'
#279930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#279940000000
0!
0'
#279950000000
1!
b11 %
1'
b11 +
#279960000000
0!
0'
#279970000000
1!
b100 %
1'
b100 +
#279980000000
0!
0'
#279990000000
1!
b101 %
1'
b101 +
#280000000000
0!
0'
#280010000000
1!
0$
b110 %
1'
0*
b110 +
#280020000000
0!
0'
#280030000000
1!
b111 %
1'
b111 +
#280040000000
0!
0'
#280050000000
1!
b1000 %
1'
b1000 +
#280060000000
0!
0'
#280070000000
1!
b1001 %
1'
b1001 +
#280080000000
0!
0'
#280090000000
1!
b0 %
1'
b0 +
#280100000000
0!
0'
#280110000000
1!
1$
b1 %
1'
1*
b1 +
#280120000000
0!
0'
#280130000000
1!
b10 %
1'
b10 +
#280140000000
1"
1(
#280150000000
0!
0"
b100 &
0'
0(
b100 ,
#280160000000
1!
b11 %
1'
b11 +
#280170000000
0!
0'
#280180000000
1!
b100 %
1'
b100 +
#280190000000
0!
0'
#280200000000
1!
b101 %
1'
b101 +
#280210000000
0!
0'
#280220000000
1!
b110 %
1'
b110 +
#280230000000
0!
0'
#280240000000
1!
b111 %
1'
b111 +
#280250000000
0!
0'
#280260000000
1!
0$
b1000 %
1'
0*
b1000 +
#280270000000
0!
0'
#280280000000
1!
b1001 %
1'
b1001 +
#280290000000
0!
0'
#280300000000
1!
b0 %
1'
b0 +
#280310000000
0!
0'
#280320000000
1!
1$
b1 %
1'
1*
b1 +
#280330000000
0!
0'
#280340000000
1!
b10 %
1'
b10 +
#280350000000
0!
0'
#280360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#280370000000
0!
0'
#280380000000
1!
b100 %
1'
b100 +
#280390000000
0!
0'
#280400000000
1!
b101 %
1'
b101 +
#280410000000
0!
0'
#280420000000
1!
0$
b110 %
1'
0*
b110 +
#280430000000
0!
0'
#280440000000
1!
b111 %
1'
b111 +
#280450000000
0!
0'
#280460000000
1!
b1000 %
1'
b1000 +
#280470000000
0!
0'
#280480000000
1!
b1001 %
1'
b1001 +
#280490000000
0!
0'
#280500000000
1!
b0 %
1'
b0 +
#280510000000
0!
0'
#280520000000
1!
1$
b1 %
1'
1*
b1 +
#280530000000
0!
0'
#280540000000
1!
b10 %
1'
b10 +
#280550000000
0!
0'
#280560000000
1!
b11 %
1'
b11 +
#280570000000
1"
1(
#280580000000
0!
0"
b100 &
0'
0(
b100 ,
#280590000000
1!
b100 %
1'
b100 +
#280600000000
0!
0'
#280610000000
1!
b101 %
1'
b101 +
#280620000000
0!
0'
#280630000000
1!
b110 %
1'
b110 +
#280640000000
0!
0'
#280650000000
1!
b111 %
1'
b111 +
#280660000000
0!
0'
#280670000000
1!
0$
b1000 %
1'
0*
b1000 +
#280680000000
0!
0'
#280690000000
1!
b1001 %
1'
b1001 +
#280700000000
0!
0'
#280710000000
1!
b0 %
1'
b0 +
#280720000000
0!
0'
#280730000000
1!
1$
b1 %
1'
1*
b1 +
#280740000000
0!
0'
#280750000000
1!
b10 %
1'
b10 +
#280760000000
0!
0'
#280770000000
1!
b11 %
1'
b11 +
#280780000000
0!
0'
#280790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#280800000000
0!
0'
#280810000000
1!
b101 %
1'
b101 +
#280820000000
0!
0'
#280830000000
1!
0$
b110 %
1'
0*
b110 +
#280840000000
0!
0'
#280850000000
1!
b111 %
1'
b111 +
#280860000000
0!
0'
#280870000000
1!
b1000 %
1'
b1000 +
#280880000000
0!
0'
#280890000000
1!
b1001 %
1'
b1001 +
#280900000000
0!
0'
#280910000000
1!
b0 %
1'
b0 +
#280920000000
0!
0'
#280930000000
1!
1$
b1 %
1'
1*
b1 +
#280940000000
0!
0'
#280950000000
1!
b10 %
1'
b10 +
#280960000000
0!
0'
#280970000000
1!
b11 %
1'
b11 +
#280980000000
0!
0'
#280990000000
1!
b100 %
1'
b100 +
#281000000000
1"
1(
#281010000000
0!
0"
b100 &
0'
0(
b100 ,
#281020000000
1!
b101 %
1'
b101 +
#281030000000
0!
0'
#281040000000
1!
b110 %
1'
b110 +
#281050000000
0!
0'
#281060000000
1!
b111 %
1'
b111 +
#281070000000
0!
0'
#281080000000
1!
0$
b1000 %
1'
0*
b1000 +
#281090000000
0!
0'
#281100000000
1!
b1001 %
1'
b1001 +
#281110000000
0!
0'
#281120000000
1!
b0 %
1'
b0 +
#281130000000
0!
0'
#281140000000
1!
1$
b1 %
1'
1*
b1 +
#281150000000
0!
0'
#281160000000
1!
b10 %
1'
b10 +
#281170000000
0!
0'
#281180000000
1!
b11 %
1'
b11 +
#281190000000
0!
0'
#281200000000
1!
b100 %
1'
b100 +
#281210000000
0!
0'
#281220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#281230000000
0!
0'
#281240000000
1!
0$
b110 %
1'
0*
b110 +
#281250000000
0!
0'
#281260000000
1!
b111 %
1'
b111 +
#281270000000
0!
0'
#281280000000
1!
b1000 %
1'
b1000 +
#281290000000
0!
0'
#281300000000
1!
b1001 %
1'
b1001 +
#281310000000
0!
0'
#281320000000
1!
b0 %
1'
b0 +
#281330000000
0!
0'
#281340000000
1!
1$
b1 %
1'
1*
b1 +
#281350000000
0!
0'
#281360000000
1!
b10 %
1'
b10 +
#281370000000
0!
0'
#281380000000
1!
b11 %
1'
b11 +
#281390000000
0!
0'
#281400000000
1!
b100 %
1'
b100 +
#281410000000
0!
0'
#281420000000
1!
b101 %
1'
b101 +
#281430000000
1"
1(
#281440000000
0!
0"
b100 &
0'
0(
b100 ,
#281450000000
1!
b110 %
1'
b110 +
#281460000000
0!
0'
#281470000000
1!
b111 %
1'
b111 +
#281480000000
0!
0'
#281490000000
1!
0$
b1000 %
1'
0*
b1000 +
#281500000000
0!
0'
#281510000000
1!
b1001 %
1'
b1001 +
#281520000000
0!
0'
#281530000000
1!
b0 %
1'
b0 +
#281540000000
0!
0'
#281550000000
1!
1$
b1 %
1'
1*
b1 +
#281560000000
0!
0'
#281570000000
1!
b10 %
1'
b10 +
#281580000000
0!
0'
#281590000000
1!
b11 %
1'
b11 +
#281600000000
0!
0'
#281610000000
1!
b100 %
1'
b100 +
#281620000000
0!
0'
#281630000000
1!
b101 %
1'
b101 +
#281640000000
0!
0'
#281650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#281660000000
0!
0'
#281670000000
1!
b111 %
1'
b111 +
#281680000000
0!
0'
#281690000000
1!
b1000 %
1'
b1000 +
#281700000000
0!
0'
#281710000000
1!
b1001 %
1'
b1001 +
#281720000000
0!
0'
#281730000000
1!
b0 %
1'
b0 +
#281740000000
0!
0'
#281750000000
1!
1$
b1 %
1'
1*
b1 +
#281760000000
0!
0'
#281770000000
1!
b10 %
1'
b10 +
#281780000000
0!
0'
#281790000000
1!
b11 %
1'
b11 +
#281800000000
0!
0'
#281810000000
1!
b100 %
1'
b100 +
#281820000000
0!
0'
#281830000000
1!
b101 %
1'
b101 +
#281840000000
0!
0'
#281850000000
1!
0$
b110 %
1'
0*
b110 +
#281860000000
1"
1(
#281870000000
0!
0"
b100 &
0'
0(
b100 ,
#281880000000
1!
1$
b111 %
1'
1*
b111 +
#281890000000
0!
0'
#281900000000
1!
0$
b1000 %
1'
0*
b1000 +
#281910000000
0!
0'
#281920000000
1!
b1001 %
1'
b1001 +
#281930000000
0!
0'
#281940000000
1!
b0 %
1'
b0 +
#281950000000
0!
0'
#281960000000
1!
1$
b1 %
1'
1*
b1 +
#281970000000
0!
0'
#281980000000
1!
b10 %
1'
b10 +
#281990000000
0!
0'
#282000000000
1!
b11 %
1'
b11 +
#282010000000
0!
0'
#282020000000
1!
b100 %
1'
b100 +
#282030000000
0!
0'
#282040000000
1!
b101 %
1'
b101 +
#282050000000
0!
0'
#282060000000
1!
b110 %
1'
b110 +
#282070000000
0!
0'
#282080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#282090000000
0!
0'
#282100000000
1!
b1000 %
1'
b1000 +
#282110000000
0!
0'
#282120000000
1!
b1001 %
1'
b1001 +
#282130000000
0!
0'
#282140000000
1!
b0 %
1'
b0 +
#282150000000
0!
0'
#282160000000
1!
1$
b1 %
1'
1*
b1 +
#282170000000
0!
0'
#282180000000
1!
b10 %
1'
b10 +
#282190000000
0!
0'
#282200000000
1!
b11 %
1'
b11 +
#282210000000
0!
0'
#282220000000
1!
b100 %
1'
b100 +
#282230000000
0!
0'
#282240000000
1!
b101 %
1'
b101 +
#282250000000
0!
0'
#282260000000
1!
0$
b110 %
1'
0*
b110 +
#282270000000
0!
0'
#282280000000
1!
b111 %
1'
b111 +
#282290000000
1"
1(
#282300000000
0!
0"
b100 &
0'
0(
b100 ,
#282310000000
1!
b1000 %
1'
b1000 +
#282320000000
0!
0'
#282330000000
1!
b1001 %
1'
b1001 +
#282340000000
0!
0'
#282350000000
1!
b0 %
1'
b0 +
#282360000000
0!
0'
#282370000000
1!
1$
b1 %
1'
1*
b1 +
#282380000000
0!
0'
#282390000000
1!
b10 %
1'
b10 +
#282400000000
0!
0'
#282410000000
1!
b11 %
1'
b11 +
#282420000000
0!
0'
#282430000000
1!
b100 %
1'
b100 +
#282440000000
0!
0'
#282450000000
1!
b101 %
1'
b101 +
#282460000000
0!
0'
#282470000000
1!
b110 %
1'
b110 +
#282480000000
0!
0'
#282490000000
1!
b111 %
1'
b111 +
#282500000000
0!
0'
#282510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#282520000000
0!
0'
#282530000000
1!
b1001 %
1'
b1001 +
#282540000000
0!
0'
#282550000000
1!
b0 %
1'
b0 +
#282560000000
0!
0'
#282570000000
1!
1$
b1 %
1'
1*
b1 +
#282580000000
0!
0'
#282590000000
1!
b10 %
1'
b10 +
#282600000000
0!
0'
#282610000000
1!
b11 %
1'
b11 +
#282620000000
0!
0'
#282630000000
1!
b100 %
1'
b100 +
#282640000000
0!
0'
#282650000000
1!
b101 %
1'
b101 +
#282660000000
0!
0'
#282670000000
1!
0$
b110 %
1'
0*
b110 +
#282680000000
0!
0'
#282690000000
1!
b111 %
1'
b111 +
#282700000000
0!
0'
#282710000000
1!
b1000 %
1'
b1000 +
#282720000000
1"
1(
#282730000000
0!
0"
b100 &
0'
0(
b100 ,
#282740000000
1!
b1001 %
1'
b1001 +
#282750000000
0!
0'
#282760000000
1!
b0 %
1'
b0 +
#282770000000
0!
0'
#282780000000
1!
1$
b1 %
1'
1*
b1 +
#282790000000
0!
0'
#282800000000
1!
b10 %
1'
b10 +
#282810000000
0!
0'
#282820000000
1!
b11 %
1'
b11 +
#282830000000
0!
0'
#282840000000
1!
b100 %
1'
b100 +
#282850000000
0!
0'
#282860000000
1!
b101 %
1'
b101 +
#282870000000
0!
0'
#282880000000
1!
b110 %
1'
b110 +
#282890000000
0!
0'
#282900000000
1!
b111 %
1'
b111 +
#282910000000
0!
0'
#282920000000
1!
0$
b1000 %
1'
0*
b1000 +
#282930000000
0!
0'
#282940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#282950000000
0!
0'
#282960000000
1!
b0 %
1'
b0 +
#282970000000
0!
0'
#282980000000
1!
1$
b1 %
1'
1*
b1 +
#282990000000
0!
0'
#283000000000
1!
b10 %
1'
b10 +
#283010000000
0!
0'
#283020000000
1!
b11 %
1'
b11 +
#283030000000
0!
0'
#283040000000
1!
b100 %
1'
b100 +
#283050000000
0!
0'
#283060000000
1!
b101 %
1'
b101 +
#283070000000
0!
0'
#283080000000
1!
0$
b110 %
1'
0*
b110 +
#283090000000
0!
0'
#283100000000
1!
b111 %
1'
b111 +
#283110000000
0!
0'
#283120000000
1!
b1000 %
1'
b1000 +
#283130000000
0!
0'
#283140000000
1!
b1001 %
1'
b1001 +
#283150000000
1"
1(
#283160000000
0!
0"
b100 &
0'
0(
b100 ,
#283170000000
1!
b0 %
1'
b0 +
#283180000000
0!
0'
#283190000000
1!
1$
b1 %
1'
1*
b1 +
#283200000000
0!
0'
#283210000000
1!
b10 %
1'
b10 +
#283220000000
0!
0'
#283230000000
1!
b11 %
1'
b11 +
#283240000000
0!
0'
#283250000000
1!
b100 %
1'
b100 +
#283260000000
0!
0'
#283270000000
1!
b101 %
1'
b101 +
#283280000000
0!
0'
#283290000000
1!
b110 %
1'
b110 +
#283300000000
0!
0'
#283310000000
1!
b111 %
1'
b111 +
#283320000000
0!
0'
#283330000000
1!
0$
b1000 %
1'
0*
b1000 +
#283340000000
0!
0'
#283350000000
1!
b1001 %
1'
b1001 +
#283360000000
0!
0'
#283370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#283380000000
0!
0'
#283390000000
1!
1$
b1 %
1'
1*
b1 +
#283400000000
0!
0'
#283410000000
1!
b10 %
1'
b10 +
#283420000000
0!
0'
#283430000000
1!
b11 %
1'
b11 +
#283440000000
0!
0'
#283450000000
1!
b100 %
1'
b100 +
#283460000000
0!
0'
#283470000000
1!
b101 %
1'
b101 +
#283480000000
0!
0'
#283490000000
1!
0$
b110 %
1'
0*
b110 +
#283500000000
0!
0'
#283510000000
1!
b111 %
1'
b111 +
#283520000000
0!
0'
#283530000000
1!
b1000 %
1'
b1000 +
#283540000000
0!
0'
#283550000000
1!
b1001 %
1'
b1001 +
#283560000000
0!
0'
#283570000000
1!
b0 %
1'
b0 +
#283580000000
1"
1(
#283590000000
0!
0"
b100 &
0'
0(
b100 ,
#283600000000
1!
1$
b1 %
1'
1*
b1 +
#283610000000
0!
0'
#283620000000
1!
b10 %
1'
b10 +
#283630000000
0!
0'
#283640000000
1!
b11 %
1'
b11 +
#283650000000
0!
0'
#283660000000
1!
b100 %
1'
b100 +
#283670000000
0!
0'
#283680000000
1!
b101 %
1'
b101 +
#283690000000
0!
0'
#283700000000
1!
b110 %
1'
b110 +
#283710000000
0!
0'
#283720000000
1!
b111 %
1'
b111 +
#283730000000
0!
0'
#283740000000
1!
0$
b1000 %
1'
0*
b1000 +
#283750000000
0!
0'
#283760000000
1!
b1001 %
1'
b1001 +
#283770000000
0!
0'
#283780000000
1!
b0 %
1'
b0 +
#283790000000
0!
0'
#283800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#283810000000
0!
0'
#283820000000
1!
b10 %
1'
b10 +
#283830000000
0!
0'
#283840000000
1!
b11 %
1'
b11 +
#283850000000
0!
0'
#283860000000
1!
b100 %
1'
b100 +
#283870000000
0!
0'
#283880000000
1!
b101 %
1'
b101 +
#283890000000
0!
0'
#283900000000
1!
0$
b110 %
1'
0*
b110 +
#283910000000
0!
0'
#283920000000
1!
b111 %
1'
b111 +
#283930000000
0!
0'
#283940000000
1!
b1000 %
1'
b1000 +
#283950000000
0!
0'
#283960000000
1!
b1001 %
1'
b1001 +
#283970000000
0!
0'
#283980000000
1!
b0 %
1'
b0 +
#283990000000
0!
0'
#284000000000
1!
1$
b1 %
1'
1*
b1 +
#284010000000
1"
1(
#284020000000
0!
0"
b100 &
0'
0(
b100 ,
#284030000000
1!
b10 %
1'
b10 +
#284040000000
0!
0'
#284050000000
1!
b11 %
1'
b11 +
#284060000000
0!
0'
#284070000000
1!
b100 %
1'
b100 +
#284080000000
0!
0'
#284090000000
1!
b101 %
1'
b101 +
#284100000000
0!
0'
#284110000000
1!
b110 %
1'
b110 +
#284120000000
0!
0'
#284130000000
1!
b111 %
1'
b111 +
#284140000000
0!
0'
#284150000000
1!
0$
b1000 %
1'
0*
b1000 +
#284160000000
0!
0'
#284170000000
1!
b1001 %
1'
b1001 +
#284180000000
0!
0'
#284190000000
1!
b0 %
1'
b0 +
#284200000000
0!
0'
#284210000000
1!
1$
b1 %
1'
1*
b1 +
#284220000000
0!
0'
#284230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#284240000000
0!
0'
#284250000000
1!
b11 %
1'
b11 +
#284260000000
0!
0'
#284270000000
1!
b100 %
1'
b100 +
#284280000000
0!
0'
#284290000000
1!
b101 %
1'
b101 +
#284300000000
0!
0'
#284310000000
1!
0$
b110 %
1'
0*
b110 +
#284320000000
0!
0'
#284330000000
1!
b111 %
1'
b111 +
#284340000000
0!
0'
#284350000000
1!
b1000 %
1'
b1000 +
#284360000000
0!
0'
#284370000000
1!
b1001 %
1'
b1001 +
#284380000000
0!
0'
#284390000000
1!
b0 %
1'
b0 +
#284400000000
0!
0'
#284410000000
1!
1$
b1 %
1'
1*
b1 +
#284420000000
0!
0'
#284430000000
1!
b10 %
1'
b10 +
#284440000000
1"
1(
#284450000000
0!
0"
b100 &
0'
0(
b100 ,
#284460000000
1!
b11 %
1'
b11 +
#284470000000
0!
0'
#284480000000
1!
b100 %
1'
b100 +
#284490000000
0!
0'
#284500000000
1!
b101 %
1'
b101 +
#284510000000
0!
0'
#284520000000
1!
b110 %
1'
b110 +
#284530000000
0!
0'
#284540000000
1!
b111 %
1'
b111 +
#284550000000
0!
0'
#284560000000
1!
0$
b1000 %
1'
0*
b1000 +
#284570000000
0!
0'
#284580000000
1!
b1001 %
1'
b1001 +
#284590000000
0!
0'
#284600000000
1!
b0 %
1'
b0 +
#284610000000
0!
0'
#284620000000
1!
1$
b1 %
1'
1*
b1 +
#284630000000
0!
0'
#284640000000
1!
b10 %
1'
b10 +
#284650000000
0!
0'
#284660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#284670000000
0!
0'
#284680000000
1!
b100 %
1'
b100 +
#284690000000
0!
0'
#284700000000
1!
b101 %
1'
b101 +
#284710000000
0!
0'
#284720000000
1!
0$
b110 %
1'
0*
b110 +
#284730000000
0!
0'
#284740000000
1!
b111 %
1'
b111 +
#284750000000
0!
0'
#284760000000
1!
b1000 %
1'
b1000 +
#284770000000
0!
0'
#284780000000
1!
b1001 %
1'
b1001 +
#284790000000
0!
0'
#284800000000
1!
b0 %
1'
b0 +
#284810000000
0!
0'
#284820000000
1!
1$
b1 %
1'
1*
b1 +
#284830000000
0!
0'
#284840000000
1!
b10 %
1'
b10 +
#284850000000
0!
0'
#284860000000
1!
b11 %
1'
b11 +
#284870000000
1"
1(
#284880000000
0!
0"
b100 &
0'
0(
b100 ,
#284890000000
1!
b100 %
1'
b100 +
#284900000000
0!
0'
#284910000000
1!
b101 %
1'
b101 +
#284920000000
0!
0'
#284930000000
1!
b110 %
1'
b110 +
#284940000000
0!
0'
#284950000000
1!
b111 %
1'
b111 +
#284960000000
0!
0'
#284970000000
1!
0$
b1000 %
1'
0*
b1000 +
#284980000000
0!
0'
#284990000000
1!
b1001 %
1'
b1001 +
#285000000000
0!
0'
#285010000000
1!
b0 %
1'
b0 +
#285020000000
0!
0'
#285030000000
1!
1$
b1 %
1'
1*
b1 +
#285040000000
0!
0'
#285050000000
1!
b10 %
1'
b10 +
#285060000000
0!
0'
#285070000000
1!
b11 %
1'
b11 +
#285080000000
0!
0'
#285090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#285100000000
0!
0'
#285110000000
1!
b101 %
1'
b101 +
#285120000000
0!
0'
#285130000000
1!
0$
b110 %
1'
0*
b110 +
#285140000000
0!
0'
#285150000000
1!
b111 %
1'
b111 +
#285160000000
0!
0'
#285170000000
1!
b1000 %
1'
b1000 +
#285180000000
0!
0'
#285190000000
1!
b1001 %
1'
b1001 +
#285200000000
0!
0'
#285210000000
1!
b0 %
1'
b0 +
#285220000000
0!
0'
#285230000000
1!
1$
b1 %
1'
1*
b1 +
#285240000000
0!
0'
#285250000000
1!
b10 %
1'
b10 +
#285260000000
0!
0'
#285270000000
1!
b11 %
1'
b11 +
#285280000000
0!
0'
#285290000000
1!
b100 %
1'
b100 +
#285300000000
1"
1(
#285310000000
0!
0"
b100 &
0'
0(
b100 ,
#285320000000
1!
b101 %
1'
b101 +
#285330000000
0!
0'
#285340000000
1!
b110 %
1'
b110 +
#285350000000
0!
0'
#285360000000
1!
b111 %
1'
b111 +
#285370000000
0!
0'
#285380000000
1!
0$
b1000 %
1'
0*
b1000 +
#285390000000
0!
0'
#285400000000
1!
b1001 %
1'
b1001 +
#285410000000
0!
0'
#285420000000
1!
b0 %
1'
b0 +
#285430000000
0!
0'
#285440000000
1!
1$
b1 %
1'
1*
b1 +
#285450000000
0!
0'
#285460000000
1!
b10 %
1'
b10 +
#285470000000
0!
0'
#285480000000
1!
b11 %
1'
b11 +
#285490000000
0!
0'
#285500000000
1!
b100 %
1'
b100 +
#285510000000
0!
0'
#285520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#285530000000
0!
0'
#285540000000
1!
0$
b110 %
1'
0*
b110 +
#285550000000
0!
0'
#285560000000
1!
b111 %
1'
b111 +
#285570000000
0!
0'
#285580000000
1!
b1000 %
1'
b1000 +
#285590000000
0!
0'
#285600000000
1!
b1001 %
1'
b1001 +
#285610000000
0!
0'
#285620000000
1!
b0 %
1'
b0 +
#285630000000
0!
0'
#285640000000
1!
1$
b1 %
1'
1*
b1 +
#285650000000
0!
0'
#285660000000
1!
b10 %
1'
b10 +
#285670000000
0!
0'
#285680000000
1!
b11 %
1'
b11 +
#285690000000
0!
0'
#285700000000
1!
b100 %
1'
b100 +
#285710000000
0!
0'
#285720000000
1!
b101 %
1'
b101 +
#285730000000
1"
1(
#285740000000
0!
0"
b100 &
0'
0(
b100 ,
#285750000000
1!
b110 %
1'
b110 +
#285760000000
0!
0'
#285770000000
1!
b111 %
1'
b111 +
#285780000000
0!
0'
#285790000000
1!
0$
b1000 %
1'
0*
b1000 +
#285800000000
0!
0'
#285810000000
1!
b1001 %
1'
b1001 +
#285820000000
0!
0'
#285830000000
1!
b0 %
1'
b0 +
#285840000000
0!
0'
#285850000000
1!
1$
b1 %
1'
1*
b1 +
#285860000000
0!
0'
#285870000000
1!
b10 %
1'
b10 +
#285880000000
0!
0'
#285890000000
1!
b11 %
1'
b11 +
#285900000000
0!
0'
#285910000000
1!
b100 %
1'
b100 +
#285920000000
0!
0'
#285930000000
1!
b101 %
1'
b101 +
#285940000000
0!
0'
#285950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#285960000000
0!
0'
#285970000000
1!
b111 %
1'
b111 +
#285980000000
0!
0'
#285990000000
1!
b1000 %
1'
b1000 +
#286000000000
0!
0'
#286010000000
1!
b1001 %
1'
b1001 +
#286020000000
0!
0'
#286030000000
1!
b0 %
1'
b0 +
#286040000000
0!
0'
#286050000000
1!
1$
b1 %
1'
1*
b1 +
#286060000000
0!
0'
#286070000000
1!
b10 %
1'
b10 +
#286080000000
0!
0'
#286090000000
1!
b11 %
1'
b11 +
#286100000000
0!
0'
#286110000000
1!
b100 %
1'
b100 +
#286120000000
0!
0'
#286130000000
1!
b101 %
1'
b101 +
#286140000000
0!
0'
#286150000000
1!
0$
b110 %
1'
0*
b110 +
#286160000000
1"
1(
#286170000000
0!
0"
b100 &
0'
0(
b100 ,
#286180000000
1!
1$
b111 %
1'
1*
b111 +
#286190000000
0!
0'
#286200000000
1!
0$
b1000 %
1'
0*
b1000 +
#286210000000
0!
0'
#286220000000
1!
b1001 %
1'
b1001 +
#286230000000
0!
0'
#286240000000
1!
b0 %
1'
b0 +
#286250000000
0!
0'
#286260000000
1!
1$
b1 %
1'
1*
b1 +
#286270000000
0!
0'
#286280000000
1!
b10 %
1'
b10 +
#286290000000
0!
0'
#286300000000
1!
b11 %
1'
b11 +
#286310000000
0!
0'
#286320000000
1!
b100 %
1'
b100 +
#286330000000
0!
0'
#286340000000
1!
b101 %
1'
b101 +
#286350000000
0!
0'
#286360000000
1!
b110 %
1'
b110 +
#286370000000
0!
0'
#286380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#286390000000
0!
0'
#286400000000
1!
b1000 %
1'
b1000 +
#286410000000
0!
0'
#286420000000
1!
b1001 %
1'
b1001 +
#286430000000
0!
0'
#286440000000
1!
b0 %
1'
b0 +
#286450000000
0!
0'
#286460000000
1!
1$
b1 %
1'
1*
b1 +
#286470000000
0!
0'
#286480000000
1!
b10 %
1'
b10 +
#286490000000
0!
0'
#286500000000
1!
b11 %
1'
b11 +
#286510000000
0!
0'
#286520000000
1!
b100 %
1'
b100 +
#286530000000
0!
0'
#286540000000
1!
b101 %
1'
b101 +
#286550000000
0!
0'
#286560000000
1!
0$
b110 %
1'
0*
b110 +
#286570000000
0!
0'
#286580000000
1!
b111 %
1'
b111 +
#286590000000
1"
1(
#286600000000
0!
0"
b100 &
0'
0(
b100 ,
#286610000000
1!
b1000 %
1'
b1000 +
#286620000000
0!
0'
#286630000000
1!
b1001 %
1'
b1001 +
#286640000000
0!
0'
#286650000000
1!
b0 %
1'
b0 +
#286660000000
0!
0'
#286670000000
1!
1$
b1 %
1'
1*
b1 +
#286680000000
0!
0'
#286690000000
1!
b10 %
1'
b10 +
#286700000000
0!
0'
#286710000000
1!
b11 %
1'
b11 +
#286720000000
0!
0'
#286730000000
1!
b100 %
1'
b100 +
#286740000000
0!
0'
#286750000000
1!
b101 %
1'
b101 +
#286760000000
0!
0'
#286770000000
1!
b110 %
1'
b110 +
#286780000000
0!
0'
#286790000000
1!
b111 %
1'
b111 +
#286800000000
0!
0'
#286810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#286820000000
0!
0'
#286830000000
1!
b1001 %
1'
b1001 +
#286840000000
0!
0'
#286850000000
1!
b0 %
1'
b0 +
#286860000000
0!
0'
#286870000000
1!
1$
b1 %
1'
1*
b1 +
#286880000000
0!
0'
#286890000000
1!
b10 %
1'
b10 +
#286900000000
0!
0'
#286910000000
1!
b11 %
1'
b11 +
#286920000000
0!
0'
#286930000000
1!
b100 %
1'
b100 +
#286940000000
0!
0'
#286950000000
1!
b101 %
1'
b101 +
#286960000000
0!
0'
#286970000000
1!
0$
b110 %
1'
0*
b110 +
#286980000000
0!
0'
#286990000000
1!
b111 %
1'
b111 +
#287000000000
0!
0'
#287010000000
1!
b1000 %
1'
b1000 +
#287020000000
1"
1(
#287030000000
0!
0"
b100 &
0'
0(
b100 ,
#287040000000
1!
b1001 %
1'
b1001 +
#287050000000
0!
0'
#287060000000
1!
b0 %
1'
b0 +
#287070000000
0!
0'
#287080000000
1!
1$
b1 %
1'
1*
b1 +
#287090000000
0!
0'
#287100000000
1!
b10 %
1'
b10 +
#287110000000
0!
0'
#287120000000
1!
b11 %
1'
b11 +
#287130000000
0!
0'
#287140000000
1!
b100 %
1'
b100 +
#287150000000
0!
0'
#287160000000
1!
b101 %
1'
b101 +
#287170000000
0!
0'
#287180000000
1!
b110 %
1'
b110 +
#287190000000
0!
0'
#287200000000
1!
b111 %
1'
b111 +
#287210000000
0!
0'
#287220000000
1!
0$
b1000 %
1'
0*
b1000 +
#287230000000
0!
0'
#287240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#287250000000
0!
0'
#287260000000
1!
b0 %
1'
b0 +
#287270000000
0!
0'
#287280000000
1!
1$
b1 %
1'
1*
b1 +
#287290000000
0!
0'
#287300000000
1!
b10 %
1'
b10 +
#287310000000
0!
0'
#287320000000
1!
b11 %
1'
b11 +
#287330000000
0!
0'
#287340000000
1!
b100 %
1'
b100 +
#287350000000
0!
0'
#287360000000
1!
b101 %
1'
b101 +
#287370000000
0!
0'
#287380000000
1!
0$
b110 %
1'
0*
b110 +
#287390000000
0!
0'
#287400000000
1!
b111 %
1'
b111 +
#287410000000
0!
0'
#287420000000
1!
b1000 %
1'
b1000 +
#287430000000
0!
0'
#287440000000
1!
b1001 %
1'
b1001 +
#287450000000
1"
1(
#287460000000
0!
0"
b100 &
0'
0(
b100 ,
#287470000000
1!
b0 %
1'
b0 +
#287480000000
0!
0'
#287490000000
1!
1$
b1 %
1'
1*
b1 +
#287500000000
0!
0'
#287510000000
1!
b10 %
1'
b10 +
#287520000000
0!
0'
#287530000000
1!
b11 %
1'
b11 +
#287540000000
0!
0'
#287550000000
1!
b100 %
1'
b100 +
#287560000000
0!
0'
#287570000000
1!
b101 %
1'
b101 +
#287580000000
0!
0'
#287590000000
1!
b110 %
1'
b110 +
#287600000000
0!
0'
#287610000000
1!
b111 %
1'
b111 +
#287620000000
0!
0'
#287630000000
1!
0$
b1000 %
1'
0*
b1000 +
#287640000000
0!
0'
#287650000000
1!
b1001 %
1'
b1001 +
#287660000000
0!
0'
#287670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#287680000000
0!
0'
#287690000000
1!
1$
b1 %
1'
1*
b1 +
#287700000000
0!
0'
#287710000000
1!
b10 %
1'
b10 +
#287720000000
0!
0'
#287730000000
1!
b11 %
1'
b11 +
#287740000000
0!
0'
#287750000000
1!
b100 %
1'
b100 +
#287760000000
0!
0'
#287770000000
1!
b101 %
1'
b101 +
#287780000000
0!
0'
#287790000000
1!
0$
b110 %
1'
0*
b110 +
#287800000000
0!
0'
#287810000000
1!
b111 %
1'
b111 +
#287820000000
0!
0'
#287830000000
1!
b1000 %
1'
b1000 +
#287840000000
0!
0'
#287850000000
1!
b1001 %
1'
b1001 +
#287860000000
0!
0'
#287870000000
1!
b0 %
1'
b0 +
#287880000000
1"
1(
#287890000000
0!
0"
b100 &
0'
0(
b100 ,
#287900000000
1!
1$
b1 %
1'
1*
b1 +
#287910000000
0!
0'
#287920000000
1!
b10 %
1'
b10 +
#287930000000
0!
0'
#287940000000
1!
b11 %
1'
b11 +
#287950000000
0!
0'
#287960000000
1!
b100 %
1'
b100 +
#287970000000
0!
0'
#287980000000
1!
b101 %
1'
b101 +
#287990000000
0!
0'
#288000000000
1!
b110 %
1'
b110 +
#288010000000
0!
0'
#288020000000
1!
b111 %
1'
b111 +
#288030000000
0!
0'
#288040000000
1!
0$
b1000 %
1'
0*
b1000 +
#288050000000
0!
0'
#288060000000
1!
b1001 %
1'
b1001 +
#288070000000
0!
0'
#288080000000
1!
b0 %
1'
b0 +
#288090000000
0!
0'
#288100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#288110000000
0!
0'
#288120000000
1!
b10 %
1'
b10 +
#288130000000
0!
0'
#288140000000
1!
b11 %
1'
b11 +
#288150000000
0!
0'
#288160000000
1!
b100 %
1'
b100 +
#288170000000
0!
0'
#288180000000
1!
b101 %
1'
b101 +
#288190000000
0!
0'
#288200000000
1!
0$
b110 %
1'
0*
b110 +
#288210000000
0!
0'
#288220000000
1!
b111 %
1'
b111 +
#288230000000
0!
0'
#288240000000
1!
b1000 %
1'
b1000 +
#288250000000
0!
0'
#288260000000
1!
b1001 %
1'
b1001 +
#288270000000
0!
0'
#288280000000
1!
b0 %
1'
b0 +
#288290000000
0!
0'
#288300000000
1!
1$
b1 %
1'
1*
b1 +
#288310000000
1"
1(
#288320000000
0!
0"
b100 &
0'
0(
b100 ,
#288330000000
1!
b10 %
1'
b10 +
#288340000000
0!
0'
#288350000000
1!
b11 %
1'
b11 +
#288360000000
0!
0'
#288370000000
1!
b100 %
1'
b100 +
#288380000000
0!
0'
#288390000000
1!
b101 %
1'
b101 +
#288400000000
0!
0'
#288410000000
1!
b110 %
1'
b110 +
#288420000000
0!
0'
#288430000000
1!
b111 %
1'
b111 +
#288440000000
0!
0'
#288450000000
1!
0$
b1000 %
1'
0*
b1000 +
#288460000000
0!
0'
#288470000000
1!
b1001 %
1'
b1001 +
#288480000000
0!
0'
#288490000000
1!
b0 %
1'
b0 +
#288500000000
0!
0'
#288510000000
1!
1$
b1 %
1'
1*
b1 +
#288520000000
0!
0'
#288530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#288540000000
0!
0'
#288550000000
1!
b11 %
1'
b11 +
#288560000000
0!
0'
#288570000000
1!
b100 %
1'
b100 +
#288580000000
0!
0'
#288590000000
1!
b101 %
1'
b101 +
#288600000000
0!
0'
#288610000000
1!
0$
b110 %
1'
0*
b110 +
#288620000000
0!
0'
#288630000000
1!
b111 %
1'
b111 +
#288640000000
0!
0'
#288650000000
1!
b1000 %
1'
b1000 +
#288660000000
0!
0'
#288670000000
1!
b1001 %
1'
b1001 +
#288680000000
0!
0'
#288690000000
1!
b0 %
1'
b0 +
#288700000000
0!
0'
#288710000000
1!
1$
b1 %
1'
1*
b1 +
#288720000000
0!
0'
#288730000000
1!
b10 %
1'
b10 +
#288740000000
1"
1(
#288750000000
0!
0"
b100 &
0'
0(
b100 ,
#288760000000
1!
b11 %
1'
b11 +
#288770000000
0!
0'
#288780000000
1!
b100 %
1'
b100 +
#288790000000
0!
0'
#288800000000
1!
b101 %
1'
b101 +
#288810000000
0!
0'
#288820000000
1!
b110 %
1'
b110 +
#288830000000
0!
0'
#288840000000
1!
b111 %
1'
b111 +
#288850000000
0!
0'
#288860000000
1!
0$
b1000 %
1'
0*
b1000 +
#288870000000
0!
0'
#288880000000
1!
b1001 %
1'
b1001 +
#288890000000
0!
0'
#288900000000
1!
b0 %
1'
b0 +
#288910000000
0!
0'
#288920000000
1!
1$
b1 %
1'
1*
b1 +
#288930000000
0!
0'
#288940000000
1!
b10 %
1'
b10 +
#288950000000
0!
0'
#288960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#288970000000
0!
0'
#288980000000
1!
b100 %
1'
b100 +
#288990000000
0!
0'
#289000000000
1!
b101 %
1'
b101 +
#289010000000
0!
0'
#289020000000
1!
0$
b110 %
1'
0*
b110 +
#289030000000
0!
0'
#289040000000
1!
b111 %
1'
b111 +
#289050000000
0!
0'
#289060000000
1!
b1000 %
1'
b1000 +
#289070000000
0!
0'
#289080000000
1!
b1001 %
1'
b1001 +
#289090000000
0!
0'
#289100000000
1!
b0 %
1'
b0 +
#289110000000
0!
0'
#289120000000
1!
1$
b1 %
1'
1*
b1 +
#289130000000
0!
0'
#289140000000
1!
b10 %
1'
b10 +
#289150000000
0!
0'
#289160000000
1!
b11 %
1'
b11 +
#289170000000
1"
1(
#289180000000
0!
0"
b100 &
0'
0(
b100 ,
#289190000000
1!
b100 %
1'
b100 +
#289200000000
0!
0'
#289210000000
1!
b101 %
1'
b101 +
#289220000000
0!
0'
#289230000000
1!
b110 %
1'
b110 +
#289240000000
0!
0'
#289250000000
1!
b111 %
1'
b111 +
#289260000000
0!
0'
#289270000000
1!
0$
b1000 %
1'
0*
b1000 +
#289280000000
0!
0'
#289290000000
1!
b1001 %
1'
b1001 +
#289300000000
0!
0'
#289310000000
1!
b0 %
1'
b0 +
#289320000000
0!
0'
#289330000000
1!
1$
b1 %
1'
1*
b1 +
#289340000000
0!
0'
#289350000000
1!
b10 %
1'
b10 +
#289360000000
0!
0'
#289370000000
1!
b11 %
1'
b11 +
#289380000000
0!
0'
#289390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#289400000000
0!
0'
#289410000000
1!
b101 %
1'
b101 +
#289420000000
0!
0'
#289430000000
1!
0$
b110 %
1'
0*
b110 +
#289440000000
0!
0'
#289450000000
1!
b111 %
1'
b111 +
#289460000000
0!
0'
#289470000000
1!
b1000 %
1'
b1000 +
#289480000000
0!
0'
#289490000000
1!
b1001 %
1'
b1001 +
#289500000000
0!
0'
#289510000000
1!
b0 %
1'
b0 +
#289520000000
0!
0'
#289530000000
1!
1$
b1 %
1'
1*
b1 +
#289540000000
0!
0'
#289550000000
1!
b10 %
1'
b10 +
#289560000000
0!
0'
#289570000000
1!
b11 %
1'
b11 +
#289580000000
0!
0'
#289590000000
1!
b100 %
1'
b100 +
#289600000000
1"
1(
#289610000000
0!
0"
b100 &
0'
0(
b100 ,
#289620000000
1!
b101 %
1'
b101 +
#289630000000
0!
0'
#289640000000
1!
b110 %
1'
b110 +
#289650000000
0!
0'
#289660000000
1!
b111 %
1'
b111 +
#289670000000
0!
0'
#289680000000
1!
0$
b1000 %
1'
0*
b1000 +
#289690000000
0!
0'
#289700000000
1!
b1001 %
1'
b1001 +
#289710000000
0!
0'
#289720000000
1!
b0 %
1'
b0 +
#289730000000
0!
0'
#289740000000
1!
1$
b1 %
1'
1*
b1 +
#289750000000
0!
0'
#289760000000
1!
b10 %
1'
b10 +
#289770000000
0!
0'
#289780000000
1!
b11 %
1'
b11 +
#289790000000
0!
0'
#289800000000
1!
b100 %
1'
b100 +
#289810000000
0!
0'
#289820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#289830000000
0!
0'
#289840000000
1!
0$
b110 %
1'
0*
b110 +
#289850000000
0!
0'
#289860000000
1!
b111 %
1'
b111 +
#289870000000
0!
0'
#289880000000
1!
b1000 %
1'
b1000 +
#289890000000
0!
0'
#289900000000
1!
b1001 %
1'
b1001 +
#289910000000
0!
0'
#289920000000
1!
b0 %
1'
b0 +
#289930000000
0!
0'
#289940000000
1!
1$
b1 %
1'
1*
b1 +
#289950000000
0!
0'
#289960000000
1!
b10 %
1'
b10 +
#289970000000
0!
0'
#289980000000
1!
b11 %
1'
b11 +
#289990000000
0!
0'
#290000000000
1!
b100 %
1'
b100 +
#290010000000
0!
0'
#290020000000
1!
b101 %
1'
b101 +
#290030000000
1"
1(
#290040000000
0!
0"
b100 &
0'
0(
b100 ,
#290050000000
1!
b110 %
1'
b110 +
#290060000000
0!
0'
#290070000000
1!
b111 %
1'
b111 +
#290080000000
0!
0'
#290090000000
1!
0$
b1000 %
1'
0*
b1000 +
#290100000000
0!
0'
#290110000000
1!
b1001 %
1'
b1001 +
#290120000000
0!
0'
#290130000000
1!
b0 %
1'
b0 +
#290140000000
0!
0'
#290150000000
1!
1$
b1 %
1'
1*
b1 +
#290160000000
0!
0'
#290170000000
1!
b10 %
1'
b10 +
#290180000000
0!
0'
#290190000000
1!
b11 %
1'
b11 +
#290200000000
0!
0'
#290210000000
1!
b100 %
1'
b100 +
#290220000000
0!
0'
#290230000000
1!
b101 %
1'
b101 +
#290240000000
0!
0'
#290250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#290260000000
0!
0'
#290270000000
1!
b111 %
1'
b111 +
#290280000000
0!
0'
#290290000000
1!
b1000 %
1'
b1000 +
#290300000000
0!
0'
#290310000000
1!
b1001 %
1'
b1001 +
#290320000000
0!
0'
#290330000000
1!
b0 %
1'
b0 +
#290340000000
0!
0'
#290350000000
1!
1$
b1 %
1'
1*
b1 +
#290360000000
0!
0'
#290370000000
1!
b10 %
1'
b10 +
#290380000000
0!
0'
#290390000000
1!
b11 %
1'
b11 +
#290400000000
0!
0'
#290410000000
1!
b100 %
1'
b100 +
#290420000000
0!
0'
#290430000000
1!
b101 %
1'
b101 +
#290440000000
0!
0'
#290450000000
1!
0$
b110 %
1'
0*
b110 +
#290460000000
1"
1(
#290470000000
0!
0"
b100 &
0'
0(
b100 ,
#290480000000
1!
1$
b111 %
1'
1*
b111 +
#290490000000
0!
0'
#290500000000
1!
0$
b1000 %
1'
0*
b1000 +
#290510000000
0!
0'
#290520000000
1!
b1001 %
1'
b1001 +
#290530000000
0!
0'
#290540000000
1!
b0 %
1'
b0 +
#290550000000
0!
0'
#290560000000
1!
1$
b1 %
1'
1*
b1 +
#290570000000
0!
0'
#290580000000
1!
b10 %
1'
b10 +
#290590000000
0!
0'
#290600000000
1!
b11 %
1'
b11 +
#290610000000
0!
0'
#290620000000
1!
b100 %
1'
b100 +
#290630000000
0!
0'
#290640000000
1!
b101 %
1'
b101 +
#290650000000
0!
0'
#290660000000
1!
b110 %
1'
b110 +
#290670000000
0!
0'
#290680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#290690000000
0!
0'
#290700000000
1!
b1000 %
1'
b1000 +
#290710000000
0!
0'
#290720000000
1!
b1001 %
1'
b1001 +
#290730000000
0!
0'
#290740000000
1!
b0 %
1'
b0 +
#290750000000
0!
0'
#290760000000
1!
1$
b1 %
1'
1*
b1 +
#290770000000
0!
0'
#290780000000
1!
b10 %
1'
b10 +
#290790000000
0!
0'
#290800000000
1!
b11 %
1'
b11 +
#290810000000
0!
0'
#290820000000
1!
b100 %
1'
b100 +
#290830000000
0!
0'
#290840000000
1!
b101 %
1'
b101 +
#290850000000
0!
0'
#290860000000
1!
0$
b110 %
1'
0*
b110 +
#290870000000
0!
0'
#290880000000
1!
b111 %
1'
b111 +
#290890000000
1"
1(
#290900000000
0!
0"
b100 &
0'
0(
b100 ,
#290910000000
1!
b1000 %
1'
b1000 +
#290920000000
0!
0'
#290930000000
1!
b1001 %
1'
b1001 +
#290940000000
0!
0'
#290950000000
1!
b0 %
1'
b0 +
#290960000000
0!
0'
#290970000000
1!
1$
b1 %
1'
1*
b1 +
#290980000000
0!
0'
#290990000000
1!
b10 %
1'
b10 +
#291000000000
0!
0'
#291010000000
1!
b11 %
1'
b11 +
#291020000000
0!
0'
#291030000000
1!
b100 %
1'
b100 +
#291040000000
0!
0'
#291050000000
1!
b101 %
1'
b101 +
#291060000000
0!
0'
#291070000000
1!
b110 %
1'
b110 +
#291080000000
0!
0'
#291090000000
1!
b111 %
1'
b111 +
#291100000000
0!
0'
#291110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#291120000000
0!
0'
#291130000000
1!
b1001 %
1'
b1001 +
#291140000000
0!
0'
#291150000000
1!
b0 %
1'
b0 +
#291160000000
0!
0'
#291170000000
1!
1$
b1 %
1'
1*
b1 +
#291180000000
0!
0'
#291190000000
1!
b10 %
1'
b10 +
#291200000000
0!
0'
#291210000000
1!
b11 %
1'
b11 +
#291220000000
0!
0'
#291230000000
1!
b100 %
1'
b100 +
#291240000000
0!
0'
#291250000000
1!
b101 %
1'
b101 +
#291260000000
0!
0'
#291270000000
1!
0$
b110 %
1'
0*
b110 +
#291280000000
0!
0'
#291290000000
1!
b111 %
1'
b111 +
#291300000000
0!
0'
#291310000000
1!
b1000 %
1'
b1000 +
#291320000000
1"
1(
#291330000000
0!
0"
b100 &
0'
0(
b100 ,
#291340000000
1!
b1001 %
1'
b1001 +
#291350000000
0!
0'
#291360000000
1!
b0 %
1'
b0 +
#291370000000
0!
0'
#291380000000
1!
1$
b1 %
1'
1*
b1 +
#291390000000
0!
0'
#291400000000
1!
b10 %
1'
b10 +
#291410000000
0!
0'
#291420000000
1!
b11 %
1'
b11 +
#291430000000
0!
0'
#291440000000
1!
b100 %
1'
b100 +
#291450000000
0!
0'
#291460000000
1!
b101 %
1'
b101 +
#291470000000
0!
0'
#291480000000
1!
b110 %
1'
b110 +
#291490000000
0!
0'
#291500000000
1!
b111 %
1'
b111 +
#291510000000
0!
0'
#291520000000
1!
0$
b1000 %
1'
0*
b1000 +
#291530000000
0!
0'
#291540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#291550000000
0!
0'
#291560000000
1!
b0 %
1'
b0 +
#291570000000
0!
0'
#291580000000
1!
1$
b1 %
1'
1*
b1 +
#291590000000
0!
0'
#291600000000
1!
b10 %
1'
b10 +
#291610000000
0!
0'
#291620000000
1!
b11 %
1'
b11 +
#291630000000
0!
0'
#291640000000
1!
b100 %
1'
b100 +
#291650000000
0!
0'
#291660000000
1!
b101 %
1'
b101 +
#291670000000
0!
0'
#291680000000
1!
0$
b110 %
1'
0*
b110 +
#291690000000
0!
0'
#291700000000
1!
b111 %
1'
b111 +
#291710000000
0!
0'
#291720000000
1!
b1000 %
1'
b1000 +
#291730000000
0!
0'
#291740000000
1!
b1001 %
1'
b1001 +
#291750000000
1"
1(
#291760000000
0!
0"
b100 &
0'
0(
b100 ,
#291770000000
1!
b0 %
1'
b0 +
#291780000000
0!
0'
#291790000000
1!
1$
b1 %
1'
1*
b1 +
#291800000000
0!
0'
#291810000000
1!
b10 %
1'
b10 +
#291820000000
0!
0'
#291830000000
1!
b11 %
1'
b11 +
#291840000000
0!
0'
#291850000000
1!
b100 %
1'
b100 +
#291860000000
0!
0'
#291870000000
1!
b101 %
1'
b101 +
#291880000000
0!
0'
#291890000000
1!
b110 %
1'
b110 +
#291900000000
0!
0'
#291910000000
1!
b111 %
1'
b111 +
#291920000000
0!
0'
#291930000000
1!
0$
b1000 %
1'
0*
b1000 +
#291940000000
0!
0'
#291950000000
1!
b1001 %
1'
b1001 +
#291960000000
0!
0'
#291970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#291980000000
0!
0'
#291990000000
1!
1$
b1 %
1'
1*
b1 +
#292000000000
0!
0'
#292010000000
1!
b10 %
1'
b10 +
#292020000000
0!
0'
#292030000000
1!
b11 %
1'
b11 +
#292040000000
0!
0'
#292050000000
1!
b100 %
1'
b100 +
#292060000000
0!
0'
#292070000000
1!
b101 %
1'
b101 +
#292080000000
0!
0'
#292090000000
1!
0$
b110 %
1'
0*
b110 +
#292100000000
0!
0'
#292110000000
1!
b111 %
1'
b111 +
#292120000000
0!
0'
#292130000000
1!
b1000 %
1'
b1000 +
#292140000000
0!
0'
#292150000000
1!
b1001 %
1'
b1001 +
#292160000000
0!
0'
#292170000000
1!
b0 %
1'
b0 +
#292180000000
1"
1(
#292190000000
0!
0"
b100 &
0'
0(
b100 ,
#292200000000
1!
1$
b1 %
1'
1*
b1 +
#292210000000
0!
0'
#292220000000
1!
b10 %
1'
b10 +
#292230000000
0!
0'
#292240000000
1!
b11 %
1'
b11 +
#292250000000
0!
0'
#292260000000
1!
b100 %
1'
b100 +
#292270000000
0!
0'
#292280000000
1!
b101 %
1'
b101 +
#292290000000
0!
0'
#292300000000
1!
b110 %
1'
b110 +
#292310000000
0!
0'
#292320000000
1!
b111 %
1'
b111 +
#292330000000
0!
0'
#292340000000
1!
0$
b1000 %
1'
0*
b1000 +
#292350000000
0!
0'
#292360000000
1!
b1001 %
1'
b1001 +
#292370000000
0!
0'
#292380000000
1!
b0 %
1'
b0 +
#292390000000
0!
0'
#292400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#292410000000
0!
0'
#292420000000
1!
b10 %
1'
b10 +
#292430000000
0!
0'
#292440000000
1!
b11 %
1'
b11 +
#292450000000
0!
0'
#292460000000
1!
b100 %
1'
b100 +
#292470000000
0!
0'
#292480000000
1!
b101 %
1'
b101 +
#292490000000
0!
0'
#292500000000
1!
0$
b110 %
1'
0*
b110 +
#292510000000
0!
0'
#292520000000
1!
b111 %
1'
b111 +
#292530000000
0!
0'
#292540000000
1!
b1000 %
1'
b1000 +
#292550000000
0!
0'
#292560000000
1!
b1001 %
1'
b1001 +
#292570000000
0!
0'
#292580000000
1!
b0 %
1'
b0 +
#292590000000
0!
0'
#292600000000
1!
1$
b1 %
1'
1*
b1 +
#292610000000
1"
1(
#292620000000
0!
0"
b100 &
0'
0(
b100 ,
#292630000000
1!
b10 %
1'
b10 +
#292640000000
0!
0'
#292650000000
1!
b11 %
1'
b11 +
#292660000000
0!
0'
#292670000000
1!
b100 %
1'
b100 +
#292680000000
0!
0'
#292690000000
1!
b101 %
1'
b101 +
#292700000000
0!
0'
#292710000000
1!
b110 %
1'
b110 +
#292720000000
0!
0'
#292730000000
1!
b111 %
1'
b111 +
#292740000000
0!
0'
#292750000000
1!
0$
b1000 %
1'
0*
b1000 +
#292760000000
0!
0'
#292770000000
1!
b1001 %
1'
b1001 +
#292780000000
0!
0'
#292790000000
1!
b0 %
1'
b0 +
#292800000000
0!
0'
#292810000000
1!
1$
b1 %
1'
1*
b1 +
#292820000000
0!
0'
#292830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#292840000000
0!
0'
#292850000000
1!
b11 %
1'
b11 +
#292860000000
0!
0'
#292870000000
1!
b100 %
1'
b100 +
#292880000000
0!
0'
#292890000000
1!
b101 %
1'
b101 +
#292900000000
0!
0'
#292910000000
1!
0$
b110 %
1'
0*
b110 +
#292920000000
0!
0'
#292930000000
1!
b111 %
1'
b111 +
#292940000000
0!
0'
#292950000000
1!
b1000 %
1'
b1000 +
#292960000000
0!
0'
#292970000000
1!
b1001 %
1'
b1001 +
#292980000000
0!
0'
#292990000000
1!
b0 %
1'
b0 +
#293000000000
0!
0'
#293010000000
1!
1$
b1 %
1'
1*
b1 +
#293020000000
0!
0'
#293030000000
1!
b10 %
1'
b10 +
#293040000000
1"
1(
#293050000000
0!
0"
b100 &
0'
0(
b100 ,
#293060000000
1!
b11 %
1'
b11 +
#293070000000
0!
0'
#293080000000
1!
b100 %
1'
b100 +
#293090000000
0!
0'
#293100000000
1!
b101 %
1'
b101 +
#293110000000
0!
0'
#293120000000
1!
b110 %
1'
b110 +
#293130000000
0!
0'
#293140000000
1!
b111 %
1'
b111 +
#293150000000
0!
0'
#293160000000
1!
0$
b1000 %
1'
0*
b1000 +
#293170000000
0!
0'
#293180000000
1!
b1001 %
1'
b1001 +
#293190000000
0!
0'
#293200000000
1!
b0 %
1'
b0 +
#293210000000
0!
0'
#293220000000
1!
1$
b1 %
1'
1*
b1 +
#293230000000
0!
0'
#293240000000
1!
b10 %
1'
b10 +
#293250000000
0!
0'
#293260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#293270000000
0!
0'
#293280000000
1!
b100 %
1'
b100 +
#293290000000
0!
0'
#293300000000
1!
b101 %
1'
b101 +
#293310000000
0!
0'
#293320000000
1!
0$
b110 %
1'
0*
b110 +
#293330000000
0!
0'
#293340000000
1!
b111 %
1'
b111 +
#293350000000
0!
0'
#293360000000
1!
b1000 %
1'
b1000 +
#293370000000
0!
0'
#293380000000
1!
b1001 %
1'
b1001 +
#293390000000
0!
0'
#293400000000
1!
b0 %
1'
b0 +
#293410000000
0!
0'
#293420000000
1!
1$
b1 %
1'
1*
b1 +
#293430000000
0!
0'
#293440000000
1!
b10 %
1'
b10 +
#293450000000
0!
0'
#293460000000
1!
b11 %
1'
b11 +
#293470000000
1"
1(
#293480000000
0!
0"
b100 &
0'
0(
b100 ,
#293490000000
1!
b100 %
1'
b100 +
#293500000000
0!
0'
#293510000000
1!
b101 %
1'
b101 +
#293520000000
0!
0'
#293530000000
1!
b110 %
1'
b110 +
#293540000000
0!
0'
#293550000000
1!
b111 %
1'
b111 +
#293560000000
0!
0'
#293570000000
1!
0$
b1000 %
1'
0*
b1000 +
#293580000000
0!
0'
#293590000000
1!
b1001 %
1'
b1001 +
#293600000000
0!
0'
#293610000000
1!
b0 %
1'
b0 +
#293620000000
0!
0'
#293630000000
1!
1$
b1 %
1'
1*
b1 +
#293640000000
0!
0'
#293650000000
1!
b10 %
1'
b10 +
#293660000000
0!
0'
#293670000000
1!
b11 %
1'
b11 +
#293680000000
0!
0'
#293690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#293700000000
0!
0'
#293710000000
1!
b101 %
1'
b101 +
#293720000000
0!
0'
#293730000000
1!
0$
b110 %
1'
0*
b110 +
#293740000000
0!
0'
#293750000000
1!
b111 %
1'
b111 +
#293760000000
0!
0'
#293770000000
1!
b1000 %
1'
b1000 +
#293780000000
0!
0'
#293790000000
1!
b1001 %
1'
b1001 +
#293800000000
0!
0'
#293810000000
1!
b0 %
1'
b0 +
#293820000000
0!
0'
#293830000000
1!
1$
b1 %
1'
1*
b1 +
#293840000000
0!
0'
#293850000000
1!
b10 %
1'
b10 +
#293860000000
0!
0'
#293870000000
1!
b11 %
1'
b11 +
#293880000000
0!
0'
#293890000000
1!
b100 %
1'
b100 +
#293900000000
1"
1(
#293910000000
0!
0"
b100 &
0'
0(
b100 ,
#293920000000
1!
b101 %
1'
b101 +
#293930000000
0!
0'
#293940000000
1!
b110 %
1'
b110 +
#293950000000
0!
0'
#293960000000
1!
b111 %
1'
b111 +
#293970000000
0!
0'
#293980000000
1!
0$
b1000 %
1'
0*
b1000 +
#293990000000
0!
0'
#294000000000
1!
b1001 %
1'
b1001 +
#294010000000
0!
0'
#294020000000
1!
b0 %
1'
b0 +
#294030000000
0!
0'
#294040000000
1!
1$
b1 %
1'
1*
b1 +
#294050000000
0!
0'
#294060000000
1!
b10 %
1'
b10 +
#294070000000
0!
0'
#294080000000
1!
b11 %
1'
b11 +
#294090000000
0!
0'
#294100000000
1!
b100 %
1'
b100 +
#294110000000
0!
0'
#294120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#294130000000
0!
0'
#294140000000
1!
0$
b110 %
1'
0*
b110 +
#294150000000
0!
0'
#294160000000
1!
b111 %
1'
b111 +
#294170000000
0!
0'
#294180000000
1!
b1000 %
1'
b1000 +
#294190000000
0!
0'
#294200000000
1!
b1001 %
1'
b1001 +
#294210000000
0!
0'
#294220000000
1!
b0 %
1'
b0 +
#294230000000
0!
0'
#294240000000
1!
1$
b1 %
1'
1*
b1 +
#294250000000
0!
0'
#294260000000
1!
b10 %
1'
b10 +
#294270000000
0!
0'
#294280000000
1!
b11 %
1'
b11 +
#294290000000
0!
0'
#294300000000
1!
b100 %
1'
b100 +
#294310000000
0!
0'
#294320000000
1!
b101 %
1'
b101 +
#294330000000
1"
1(
#294340000000
0!
0"
b100 &
0'
0(
b100 ,
#294350000000
1!
b110 %
1'
b110 +
#294360000000
0!
0'
#294370000000
1!
b111 %
1'
b111 +
#294380000000
0!
0'
#294390000000
1!
0$
b1000 %
1'
0*
b1000 +
#294400000000
0!
0'
#294410000000
1!
b1001 %
1'
b1001 +
#294420000000
0!
0'
#294430000000
1!
b0 %
1'
b0 +
#294440000000
0!
0'
#294450000000
1!
1$
b1 %
1'
1*
b1 +
#294460000000
0!
0'
#294470000000
1!
b10 %
1'
b10 +
#294480000000
0!
0'
#294490000000
1!
b11 %
1'
b11 +
#294500000000
0!
0'
#294510000000
1!
b100 %
1'
b100 +
#294520000000
0!
0'
#294530000000
1!
b101 %
1'
b101 +
#294540000000
0!
0'
#294550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#294560000000
0!
0'
#294570000000
1!
b111 %
1'
b111 +
#294580000000
0!
0'
#294590000000
1!
b1000 %
1'
b1000 +
#294600000000
0!
0'
#294610000000
1!
b1001 %
1'
b1001 +
#294620000000
0!
0'
#294630000000
1!
b0 %
1'
b0 +
#294640000000
0!
0'
#294650000000
1!
1$
b1 %
1'
1*
b1 +
#294660000000
0!
0'
#294670000000
1!
b10 %
1'
b10 +
#294680000000
0!
0'
#294690000000
1!
b11 %
1'
b11 +
#294700000000
0!
0'
#294710000000
1!
b100 %
1'
b100 +
#294720000000
0!
0'
#294730000000
1!
b101 %
1'
b101 +
#294740000000
0!
0'
#294750000000
1!
0$
b110 %
1'
0*
b110 +
#294760000000
1"
1(
#294770000000
0!
0"
b100 &
0'
0(
b100 ,
#294780000000
1!
1$
b111 %
1'
1*
b111 +
#294790000000
0!
0'
#294800000000
1!
0$
b1000 %
1'
0*
b1000 +
#294810000000
0!
0'
#294820000000
1!
b1001 %
1'
b1001 +
#294830000000
0!
0'
#294840000000
1!
b0 %
1'
b0 +
#294850000000
0!
0'
#294860000000
1!
1$
b1 %
1'
1*
b1 +
#294870000000
0!
0'
#294880000000
1!
b10 %
1'
b10 +
#294890000000
0!
0'
#294900000000
1!
b11 %
1'
b11 +
#294910000000
0!
0'
#294920000000
1!
b100 %
1'
b100 +
#294930000000
0!
0'
#294940000000
1!
b101 %
1'
b101 +
#294950000000
0!
0'
#294960000000
1!
b110 %
1'
b110 +
#294970000000
0!
0'
#294980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#294990000000
0!
0'
#295000000000
1!
b1000 %
1'
b1000 +
#295010000000
0!
0'
#295020000000
1!
b1001 %
1'
b1001 +
#295030000000
0!
0'
#295040000000
1!
b0 %
1'
b0 +
#295050000000
0!
0'
#295060000000
1!
1$
b1 %
1'
1*
b1 +
#295070000000
0!
0'
#295080000000
1!
b10 %
1'
b10 +
#295090000000
0!
0'
#295100000000
1!
b11 %
1'
b11 +
#295110000000
0!
0'
#295120000000
1!
b100 %
1'
b100 +
#295130000000
0!
0'
#295140000000
1!
b101 %
1'
b101 +
#295150000000
0!
0'
#295160000000
1!
0$
b110 %
1'
0*
b110 +
#295170000000
0!
0'
#295180000000
1!
b111 %
1'
b111 +
#295190000000
1"
1(
#295200000000
0!
0"
b100 &
0'
0(
b100 ,
#295210000000
1!
b1000 %
1'
b1000 +
#295220000000
0!
0'
#295230000000
1!
b1001 %
1'
b1001 +
#295240000000
0!
0'
#295250000000
1!
b0 %
1'
b0 +
#295260000000
0!
0'
#295270000000
1!
1$
b1 %
1'
1*
b1 +
#295280000000
0!
0'
#295290000000
1!
b10 %
1'
b10 +
#295300000000
0!
0'
#295310000000
1!
b11 %
1'
b11 +
#295320000000
0!
0'
#295330000000
1!
b100 %
1'
b100 +
#295340000000
0!
0'
#295350000000
1!
b101 %
1'
b101 +
#295360000000
0!
0'
#295370000000
1!
b110 %
1'
b110 +
#295380000000
0!
0'
#295390000000
1!
b111 %
1'
b111 +
#295400000000
0!
0'
#295410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#295420000000
0!
0'
#295430000000
1!
b1001 %
1'
b1001 +
#295440000000
0!
0'
#295450000000
1!
b0 %
1'
b0 +
#295460000000
0!
0'
#295470000000
1!
1$
b1 %
1'
1*
b1 +
#295480000000
0!
0'
#295490000000
1!
b10 %
1'
b10 +
#295500000000
0!
0'
#295510000000
1!
b11 %
1'
b11 +
#295520000000
0!
0'
#295530000000
1!
b100 %
1'
b100 +
#295540000000
0!
0'
#295550000000
1!
b101 %
1'
b101 +
#295560000000
0!
0'
#295570000000
1!
0$
b110 %
1'
0*
b110 +
#295580000000
0!
0'
#295590000000
1!
b111 %
1'
b111 +
#295600000000
0!
0'
#295610000000
1!
b1000 %
1'
b1000 +
#295620000000
1"
1(
#295630000000
0!
0"
b100 &
0'
0(
b100 ,
#295640000000
1!
b1001 %
1'
b1001 +
#295650000000
0!
0'
#295660000000
1!
b0 %
1'
b0 +
#295670000000
0!
0'
#295680000000
1!
1$
b1 %
1'
1*
b1 +
#295690000000
0!
0'
#295700000000
1!
b10 %
1'
b10 +
#295710000000
0!
0'
#295720000000
1!
b11 %
1'
b11 +
#295730000000
0!
0'
#295740000000
1!
b100 %
1'
b100 +
#295750000000
0!
0'
#295760000000
1!
b101 %
1'
b101 +
#295770000000
0!
0'
#295780000000
1!
b110 %
1'
b110 +
#295790000000
0!
0'
#295800000000
1!
b111 %
1'
b111 +
#295810000000
0!
0'
#295820000000
1!
0$
b1000 %
1'
0*
b1000 +
#295830000000
0!
0'
#295840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#295850000000
0!
0'
#295860000000
1!
b0 %
1'
b0 +
#295870000000
0!
0'
#295880000000
1!
1$
b1 %
1'
1*
b1 +
#295890000000
0!
0'
#295900000000
1!
b10 %
1'
b10 +
#295910000000
0!
0'
#295920000000
1!
b11 %
1'
b11 +
#295930000000
0!
0'
#295940000000
1!
b100 %
1'
b100 +
#295950000000
0!
0'
#295960000000
1!
b101 %
1'
b101 +
#295970000000
0!
0'
#295980000000
1!
0$
b110 %
1'
0*
b110 +
#295990000000
0!
0'
#296000000000
1!
b111 %
1'
b111 +
#296010000000
0!
0'
#296020000000
1!
b1000 %
1'
b1000 +
#296030000000
0!
0'
#296040000000
1!
b1001 %
1'
b1001 +
#296050000000
1"
1(
#296060000000
0!
0"
b100 &
0'
0(
b100 ,
#296070000000
1!
b0 %
1'
b0 +
#296080000000
0!
0'
#296090000000
1!
1$
b1 %
1'
1*
b1 +
#296100000000
0!
0'
#296110000000
1!
b10 %
1'
b10 +
#296120000000
0!
0'
#296130000000
1!
b11 %
1'
b11 +
#296140000000
0!
0'
#296150000000
1!
b100 %
1'
b100 +
#296160000000
0!
0'
#296170000000
1!
b101 %
1'
b101 +
#296180000000
0!
0'
#296190000000
1!
b110 %
1'
b110 +
#296200000000
0!
0'
#296210000000
1!
b111 %
1'
b111 +
#296220000000
0!
0'
#296230000000
1!
0$
b1000 %
1'
0*
b1000 +
#296240000000
0!
0'
#296250000000
1!
b1001 %
1'
b1001 +
#296260000000
0!
0'
#296270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#296280000000
0!
0'
#296290000000
1!
1$
b1 %
1'
1*
b1 +
#296300000000
0!
0'
#296310000000
1!
b10 %
1'
b10 +
#296320000000
0!
0'
#296330000000
1!
b11 %
1'
b11 +
#296340000000
0!
0'
#296350000000
1!
b100 %
1'
b100 +
#296360000000
0!
0'
#296370000000
1!
b101 %
1'
b101 +
#296380000000
0!
0'
#296390000000
1!
0$
b110 %
1'
0*
b110 +
#296400000000
0!
0'
#296410000000
1!
b111 %
1'
b111 +
#296420000000
0!
0'
#296430000000
1!
b1000 %
1'
b1000 +
#296440000000
0!
0'
#296450000000
1!
b1001 %
1'
b1001 +
#296460000000
0!
0'
#296470000000
1!
b0 %
1'
b0 +
#296480000000
1"
1(
#296490000000
0!
0"
b100 &
0'
0(
b100 ,
#296500000000
1!
1$
b1 %
1'
1*
b1 +
#296510000000
0!
0'
#296520000000
1!
b10 %
1'
b10 +
#296530000000
0!
0'
#296540000000
1!
b11 %
1'
b11 +
#296550000000
0!
0'
#296560000000
1!
b100 %
1'
b100 +
#296570000000
0!
0'
#296580000000
1!
b101 %
1'
b101 +
#296590000000
0!
0'
#296600000000
1!
b110 %
1'
b110 +
#296610000000
0!
0'
#296620000000
1!
b111 %
1'
b111 +
#296630000000
0!
0'
#296640000000
1!
0$
b1000 %
1'
0*
b1000 +
#296650000000
0!
0'
#296660000000
1!
b1001 %
1'
b1001 +
#296670000000
0!
0'
#296680000000
1!
b0 %
1'
b0 +
#296690000000
0!
0'
#296700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#296710000000
0!
0'
#296720000000
1!
b10 %
1'
b10 +
#296730000000
0!
0'
#296740000000
1!
b11 %
1'
b11 +
#296750000000
0!
0'
#296760000000
1!
b100 %
1'
b100 +
#296770000000
0!
0'
#296780000000
1!
b101 %
1'
b101 +
#296790000000
0!
0'
#296800000000
1!
0$
b110 %
1'
0*
b110 +
#296810000000
0!
0'
#296820000000
1!
b111 %
1'
b111 +
#296830000000
0!
0'
#296840000000
1!
b1000 %
1'
b1000 +
#296850000000
0!
0'
#296860000000
1!
b1001 %
1'
b1001 +
#296870000000
0!
0'
#296880000000
1!
b0 %
1'
b0 +
#296890000000
0!
0'
#296900000000
1!
1$
b1 %
1'
1*
b1 +
#296910000000
1"
1(
#296920000000
0!
0"
b100 &
0'
0(
b100 ,
#296930000000
1!
b10 %
1'
b10 +
#296940000000
0!
0'
#296950000000
1!
b11 %
1'
b11 +
#296960000000
0!
0'
#296970000000
1!
b100 %
1'
b100 +
#296980000000
0!
0'
#296990000000
1!
b101 %
1'
b101 +
#297000000000
0!
0'
#297010000000
1!
b110 %
1'
b110 +
#297020000000
0!
0'
#297030000000
1!
b111 %
1'
b111 +
#297040000000
0!
0'
#297050000000
1!
0$
b1000 %
1'
0*
b1000 +
#297060000000
0!
0'
#297070000000
1!
b1001 %
1'
b1001 +
#297080000000
0!
0'
#297090000000
1!
b0 %
1'
b0 +
#297100000000
0!
0'
#297110000000
1!
1$
b1 %
1'
1*
b1 +
#297120000000
0!
0'
#297130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#297140000000
0!
0'
#297150000000
1!
b11 %
1'
b11 +
#297160000000
0!
0'
#297170000000
1!
b100 %
1'
b100 +
#297180000000
0!
0'
#297190000000
1!
b101 %
1'
b101 +
#297200000000
0!
0'
#297210000000
1!
0$
b110 %
1'
0*
b110 +
#297220000000
0!
0'
#297230000000
1!
b111 %
1'
b111 +
#297240000000
0!
0'
#297250000000
1!
b1000 %
1'
b1000 +
#297260000000
0!
0'
#297270000000
1!
b1001 %
1'
b1001 +
#297280000000
0!
0'
#297290000000
1!
b0 %
1'
b0 +
#297300000000
0!
0'
#297310000000
1!
1$
b1 %
1'
1*
b1 +
#297320000000
0!
0'
#297330000000
1!
b10 %
1'
b10 +
#297340000000
1"
1(
#297350000000
0!
0"
b100 &
0'
0(
b100 ,
#297360000000
1!
b11 %
1'
b11 +
#297370000000
0!
0'
#297380000000
1!
b100 %
1'
b100 +
#297390000000
0!
0'
#297400000000
1!
b101 %
1'
b101 +
#297410000000
0!
0'
#297420000000
1!
b110 %
1'
b110 +
#297430000000
0!
0'
#297440000000
1!
b111 %
1'
b111 +
#297450000000
0!
0'
#297460000000
1!
0$
b1000 %
1'
0*
b1000 +
#297470000000
0!
0'
#297480000000
1!
b1001 %
1'
b1001 +
#297490000000
0!
0'
#297500000000
1!
b0 %
1'
b0 +
#297510000000
0!
0'
#297520000000
1!
1$
b1 %
1'
1*
b1 +
#297530000000
0!
0'
#297540000000
1!
b10 %
1'
b10 +
#297550000000
0!
0'
#297560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#297570000000
0!
0'
#297580000000
1!
b100 %
1'
b100 +
#297590000000
0!
0'
#297600000000
1!
b101 %
1'
b101 +
#297610000000
0!
0'
#297620000000
1!
0$
b110 %
1'
0*
b110 +
#297630000000
0!
0'
#297640000000
1!
b111 %
1'
b111 +
#297650000000
0!
0'
#297660000000
1!
b1000 %
1'
b1000 +
#297670000000
0!
0'
#297680000000
1!
b1001 %
1'
b1001 +
#297690000000
0!
0'
#297700000000
1!
b0 %
1'
b0 +
#297710000000
0!
0'
#297720000000
1!
1$
b1 %
1'
1*
b1 +
#297730000000
0!
0'
#297740000000
1!
b10 %
1'
b10 +
#297750000000
0!
0'
#297760000000
1!
b11 %
1'
b11 +
#297770000000
1"
1(
#297780000000
0!
0"
b100 &
0'
0(
b100 ,
#297790000000
1!
b100 %
1'
b100 +
#297800000000
0!
0'
#297810000000
1!
b101 %
1'
b101 +
#297820000000
0!
0'
#297830000000
1!
b110 %
1'
b110 +
#297840000000
0!
0'
#297850000000
1!
b111 %
1'
b111 +
#297860000000
0!
0'
#297870000000
1!
0$
b1000 %
1'
0*
b1000 +
#297880000000
0!
0'
#297890000000
1!
b1001 %
1'
b1001 +
#297900000000
0!
0'
#297910000000
1!
b0 %
1'
b0 +
#297920000000
0!
0'
#297930000000
1!
1$
b1 %
1'
1*
b1 +
#297940000000
0!
0'
#297950000000
1!
b10 %
1'
b10 +
#297960000000
0!
0'
#297970000000
1!
b11 %
1'
b11 +
#297980000000
0!
0'
#297990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#298000000000
0!
0'
#298010000000
1!
b101 %
1'
b101 +
#298020000000
0!
0'
#298030000000
1!
0$
b110 %
1'
0*
b110 +
#298040000000
0!
0'
#298050000000
1!
b111 %
1'
b111 +
#298060000000
0!
0'
#298070000000
1!
b1000 %
1'
b1000 +
#298080000000
0!
0'
#298090000000
1!
b1001 %
1'
b1001 +
#298100000000
0!
0'
#298110000000
1!
b0 %
1'
b0 +
#298120000000
0!
0'
#298130000000
1!
1$
b1 %
1'
1*
b1 +
#298140000000
0!
0'
#298150000000
1!
b10 %
1'
b10 +
#298160000000
0!
0'
#298170000000
1!
b11 %
1'
b11 +
#298180000000
0!
0'
#298190000000
1!
b100 %
1'
b100 +
#298200000000
1"
1(
#298210000000
0!
0"
b100 &
0'
0(
b100 ,
#298220000000
1!
b101 %
1'
b101 +
#298230000000
0!
0'
#298240000000
1!
b110 %
1'
b110 +
#298250000000
0!
0'
#298260000000
1!
b111 %
1'
b111 +
#298270000000
0!
0'
#298280000000
1!
0$
b1000 %
1'
0*
b1000 +
#298290000000
0!
0'
#298300000000
1!
b1001 %
1'
b1001 +
#298310000000
0!
0'
#298320000000
1!
b0 %
1'
b0 +
#298330000000
0!
0'
#298340000000
1!
1$
b1 %
1'
1*
b1 +
#298350000000
0!
0'
#298360000000
1!
b10 %
1'
b10 +
#298370000000
0!
0'
#298380000000
1!
b11 %
1'
b11 +
#298390000000
0!
0'
#298400000000
1!
b100 %
1'
b100 +
#298410000000
0!
0'
#298420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#298430000000
0!
0'
#298440000000
1!
0$
b110 %
1'
0*
b110 +
#298450000000
0!
0'
#298460000000
1!
b111 %
1'
b111 +
#298470000000
0!
0'
#298480000000
1!
b1000 %
1'
b1000 +
#298490000000
0!
0'
#298500000000
1!
b1001 %
1'
b1001 +
#298510000000
0!
0'
#298520000000
1!
b0 %
1'
b0 +
#298530000000
0!
0'
#298540000000
1!
1$
b1 %
1'
1*
b1 +
#298550000000
0!
0'
#298560000000
1!
b10 %
1'
b10 +
#298570000000
0!
0'
#298580000000
1!
b11 %
1'
b11 +
#298590000000
0!
0'
#298600000000
1!
b100 %
1'
b100 +
#298610000000
0!
0'
#298620000000
1!
b101 %
1'
b101 +
#298630000000
1"
1(
#298640000000
0!
0"
b100 &
0'
0(
b100 ,
#298650000000
1!
b110 %
1'
b110 +
#298660000000
0!
0'
#298670000000
1!
b111 %
1'
b111 +
#298680000000
0!
0'
#298690000000
1!
0$
b1000 %
1'
0*
b1000 +
#298700000000
0!
0'
#298710000000
1!
b1001 %
1'
b1001 +
#298720000000
0!
0'
#298730000000
1!
b0 %
1'
b0 +
#298740000000
0!
0'
#298750000000
1!
1$
b1 %
1'
1*
b1 +
#298760000000
0!
0'
#298770000000
1!
b10 %
1'
b10 +
#298780000000
0!
0'
#298790000000
1!
b11 %
1'
b11 +
#298800000000
0!
0'
#298810000000
1!
b100 %
1'
b100 +
#298820000000
0!
0'
#298830000000
1!
b101 %
1'
b101 +
#298840000000
0!
0'
#298850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#298860000000
0!
0'
#298870000000
1!
b111 %
1'
b111 +
#298880000000
0!
0'
#298890000000
1!
b1000 %
1'
b1000 +
#298900000000
0!
0'
#298910000000
1!
b1001 %
1'
b1001 +
#298920000000
0!
0'
#298930000000
1!
b0 %
1'
b0 +
#298940000000
0!
0'
#298950000000
1!
1$
b1 %
1'
1*
b1 +
#298960000000
0!
0'
#298970000000
1!
b10 %
1'
b10 +
#298980000000
0!
0'
#298990000000
1!
b11 %
1'
b11 +
#299000000000
0!
0'
#299010000000
1!
b100 %
1'
b100 +
#299020000000
0!
0'
#299030000000
1!
b101 %
1'
b101 +
#299040000000
0!
0'
#299050000000
1!
0$
b110 %
1'
0*
b110 +
#299060000000
1"
1(
#299070000000
0!
0"
b100 &
0'
0(
b100 ,
#299080000000
1!
1$
b111 %
1'
1*
b111 +
#299090000000
0!
0'
#299100000000
1!
0$
b1000 %
1'
0*
b1000 +
#299110000000
0!
0'
#299120000000
1!
b1001 %
1'
b1001 +
#299130000000
0!
0'
#299140000000
1!
b0 %
1'
b0 +
#299150000000
0!
0'
#299160000000
1!
1$
b1 %
1'
1*
b1 +
#299170000000
0!
0'
#299180000000
1!
b10 %
1'
b10 +
#299190000000
0!
0'
#299200000000
1!
b11 %
1'
b11 +
#299210000000
0!
0'
#299220000000
1!
b100 %
1'
b100 +
#299230000000
0!
0'
#299240000000
1!
b101 %
1'
b101 +
#299250000000
0!
0'
#299260000000
1!
b110 %
1'
b110 +
#299270000000
0!
0'
#299280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#299290000000
0!
0'
#299300000000
1!
b1000 %
1'
b1000 +
#299310000000
0!
0'
#299320000000
1!
b1001 %
1'
b1001 +
#299330000000
0!
0'
#299340000000
1!
b0 %
1'
b0 +
#299350000000
0!
0'
#299360000000
1!
1$
b1 %
1'
1*
b1 +
#299370000000
0!
0'
#299380000000
1!
b10 %
1'
b10 +
#299390000000
0!
0'
#299400000000
1!
b11 %
1'
b11 +
#299410000000
0!
0'
#299420000000
1!
b100 %
1'
b100 +
#299430000000
0!
0'
#299440000000
1!
b101 %
1'
b101 +
#299450000000
0!
0'
#299460000000
1!
0$
b110 %
1'
0*
b110 +
#299470000000
0!
0'
#299480000000
1!
b111 %
1'
b111 +
#299490000000
1"
1(
#299500000000
0!
0"
b100 &
0'
0(
b100 ,
#299510000000
1!
b1000 %
1'
b1000 +
#299520000000
0!
0'
#299530000000
1!
b1001 %
1'
b1001 +
#299540000000
0!
0'
#299550000000
1!
b0 %
1'
b0 +
#299560000000
0!
0'
#299570000000
1!
1$
b1 %
1'
1*
b1 +
#299580000000
0!
0'
#299590000000
1!
b10 %
1'
b10 +
#299600000000
0!
0'
#299610000000
1!
b11 %
1'
b11 +
#299620000000
0!
0'
#299630000000
1!
b100 %
1'
b100 +
#299640000000
0!
0'
#299650000000
1!
b101 %
1'
b101 +
#299660000000
0!
0'
#299670000000
1!
b110 %
1'
b110 +
#299680000000
0!
0'
#299690000000
1!
b111 %
1'
b111 +
#299700000000
0!
0'
#299710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#299720000000
0!
0'
#299730000000
1!
b1001 %
1'
b1001 +
#299740000000
0!
0'
#299750000000
1!
b0 %
1'
b0 +
#299760000000
0!
0'
#299770000000
1!
1$
b1 %
1'
1*
b1 +
#299780000000
0!
0'
#299790000000
1!
b10 %
1'
b10 +
#299800000000
0!
0'
#299810000000
1!
b11 %
1'
b11 +
#299820000000
0!
0'
#299830000000
1!
b100 %
1'
b100 +
#299840000000
0!
0'
#299850000000
1!
b101 %
1'
b101 +
#299860000000
0!
0'
#299870000000
1!
0$
b110 %
1'
0*
b110 +
#299880000000
0!
0'
#299890000000
1!
b111 %
1'
b111 +
#299900000000
0!
0'
#299910000000
1!
b1000 %
1'
b1000 +
#299920000000
1"
1(
#299930000000
0!
0"
b100 &
0'
0(
b100 ,
#299940000000
1!
b1001 %
1'
b1001 +
#299950000000
0!
0'
#299960000000
1!
b0 %
1'
b0 +
#299970000000
0!
0'
#299980000000
1!
1$
b1 %
1'
1*
b1 +
#299990000000
0!
0'
#300000000000
1!
b10 %
1'
b10 +
#300010000000
0!
0'
#300020000000
1!
b11 %
1'
b11 +
#300030000000
0!
0'
#300040000000
1!
b100 %
1'
b100 +
#300050000000
0!
0'
#300060000000
1!
b101 %
1'
b101 +
#300070000000
0!
0'
#300080000000
1!
b110 %
1'
b110 +
#300090000000
0!
0'
#300100000000
1!
b111 %
1'
b111 +
#300110000000
0!
0'
#300120000000
1!
0$
b1000 %
1'
0*
b1000 +
#300130000000
0!
0'
#300140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#300150000000
0!
0'
#300160000000
1!
b0 %
1'
b0 +
#300170000000
0!
0'
#300180000000
1!
1$
b1 %
1'
1*
b1 +
#300190000000
0!
0'
#300200000000
1!
b10 %
1'
b10 +
#300210000000
0!
0'
#300220000000
1!
b11 %
1'
b11 +
#300230000000
0!
0'
#300240000000
1!
b100 %
1'
b100 +
#300250000000
0!
0'
#300260000000
1!
b101 %
1'
b101 +
#300270000000
0!
0'
#300280000000
1!
0$
b110 %
1'
0*
b110 +
#300290000000
0!
0'
#300300000000
1!
b111 %
1'
b111 +
#300310000000
0!
0'
#300320000000
1!
b1000 %
1'
b1000 +
#300330000000
0!
0'
#300340000000
1!
b1001 %
1'
b1001 +
#300350000000
1"
1(
#300360000000
0!
0"
b100 &
0'
0(
b100 ,
#300370000000
1!
b0 %
1'
b0 +
#300380000000
0!
0'
#300390000000
1!
1$
b1 %
1'
1*
b1 +
#300400000000
0!
0'
#300410000000
1!
b10 %
1'
b10 +
#300420000000
0!
0'
#300430000000
1!
b11 %
1'
b11 +
#300440000000
0!
0'
#300450000000
1!
b100 %
1'
b100 +
#300460000000
0!
0'
#300470000000
1!
b101 %
1'
b101 +
#300480000000
0!
0'
#300490000000
1!
b110 %
1'
b110 +
#300500000000
0!
0'
#300510000000
1!
b111 %
1'
b111 +
#300520000000
0!
0'
#300530000000
1!
0$
b1000 %
1'
0*
b1000 +
#300540000000
0!
0'
#300550000000
1!
b1001 %
1'
b1001 +
#300560000000
0!
0'
#300570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#300580000000
0!
0'
#300590000000
1!
1$
b1 %
1'
1*
b1 +
#300600000000
0!
0'
#300610000000
1!
b10 %
1'
b10 +
#300620000000
0!
0'
#300630000000
1!
b11 %
1'
b11 +
#300640000000
0!
0'
#300650000000
1!
b100 %
1'
b100 +
#300660000000
0!
0'
#300670000000
1!
b101 %
1'
b101 +
#300680000000
0!
0'
#300690000000
1!
0$
b110 %
1'
0*
b110 +
#300700000000
0!
0'
#300710000000
1!
b111 %
1'
b111 +
#300720000000
0!
0'
#300730000000
1!
b1000 %
1'
b1000 +
#300740000000
0!
0'
#300750000000
1!
b1001 %
1'
b1001 +
#300760000000
0!
0'
#300770000000
1!
b0 %
1'
b0 +
#300780000000
1"
1(
#300790000000
0!
0"
b100 &
0'
0(
b100 ,
#300800000000
1!
1$
b1 %
1'
1*
b1 +
#300810000000
0!
0'
#300820000000
1!
b10 %
1'
b10 +
#300830000000
0!
0'
#300840000000
1!
b11 %
1'
b11 +
#300850000000
0!
0'
#300860000000
1!
b100 %
1'
b100 +
#300870000000
0!
0'
#300880000000
1!
b101 %
1'
b101 +
#300890000000
0!
0'
#300900000000
1!
b110 %
1'
b110 +
#300910000000
0!
0'
#300920000000
1!
b111 %
1'
b111 +
#300930000000
0!
0'
#300940000000
1!
0$
b1000 %
1'
0*
b1000 +
#300950000000
0!
0'
#300960000000
1!
b1001 %
1'
b1001 +
#300970000000
0!
0'
#300980000000
1!
b0 %
1'
b0 +
#300990000000
0!
0'
#301000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#301010000000
0!
0'
#301020000000
1!
b10 %
1'
b10 +
#301030000000
0!
0'
#301040000000
1!
b11 %
1'
b11 +
#301050000000
0!
0'
#301060000000
1!
b100 %
1'
b100 +
#301070000000
0!
0'
#301080000000
1!
b101 %
1'
b101 +
#301090000000
0!
0'
#301100000000
1!
0$
b110 %
1'
0*
b110 +
#301110000000
0!
0'
#301120000000
1!
b111 %
1'
b111 +
#301130000000
0!
0'
#301140000000
1!
b1000 %
1'
b1000 +
#301150000000
0!
0'
#301160000000
1!
b1001 %
1'
b1001 +
#301170000000
0!
0'
#301180000000
1!
b0 %
1'
b0 +
#301190000000
0!
0'
#301200000000
1!
1$
b1 %
1'
1*
b1 +
#301210000000
1"
1(
#301220000000
0!
0"
b100 &
0'
0(
b100 ,
#301230000000
1!
b10 %
1'
b10 +
#301240000000
0!
0'
#301250000000
1!
b11 %
1'
b11 +
#301260000000
0!
0'
#301270000000
1!
b100 %
1'
b100 +
#301280000000
0!
0'
#301290000000
1!
b101 %
1'
b101 +
#301300000000
0!
0'
#301310000000
1!
b110 %
1'
b110 +
#301320000000
0!
0'
#301330000000
1!
b111 %
1'
b111 +
#301340000000
0!
0'
#301350000000
1!
0$
b1000 %
1'
0*
b1000 +
#301360000000
0!
0'
#301370000000
1!
b1001 %
1'
b1001 +
#301380000000
0!
0'
#301390000000
1!
b0 %
1'
b0 +
#301400000000
0!
0'
#301410000000
1!
1$
b1 %
1'
1*
b1 +
#301420000000
0!
0'
#301430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#301440000000
0!
0'
#301450000000
1!
b11 %
1'
b11 +
#301460000000
0!
0'
#301470000000
1!
b100 %
1'
b100 +
#301480000000
0!
0'
#301490000000
1!
b101 %
1'
b101 +
#301500000000
0!
0'
#301510000000
1!
0$
b110 %
1'
0*
b110 +
#301520000000
0!
0'
#301530000000
1!
b111 %
1'
b111 +
#301540000000
0!
0'
#301550000000
1!
b1000 %
1'
b1000 +
#301560000000
0!
0'
#301570000000
1!
b1001 %
1'
b1001 +
#301580000000
0!
0'
#301590000000
1!
b0 %
1'
b0 +
#301600000000
0!
0'
#301610000000
1!
1$
b1 %
1'
1*
b1 +
#301620000000
0!
0'
#301630000000
1!
b10 %
1'
b10 +
#301640000000
1"
1(
#301650000000
0!
0"
b100 &
0'
0(
b100 ,
#301660000000
1!
b11 %
1'
b11 +
#301670000000
0!
0'
#301680000000
1!
b100 %
1'
b100 +
#301690000000
0!
0'
#301700000000
1!
b101 %
1'
b101 +
#301710000000
0!
0'
#301720000000
1!
b110 %
1'
b110 +
#301730000000
0!
0'
#301740000000
1!
b111 %
1'
b111 +
#301750000000
0!
0'
#301760000000
1!
0$
b1000 %
1'
0*
b1000 +
#301770000000
0!
0'
#301780000000
1!
b1001 %
1'
b1001 +
#301790000000
0!
0'
#301800000000
1!
b0 %
1'
b0 +
#301810000000
0!
0'
#301820000000
1!
1$
b1 %
1'
1*
b1 +
#301830000000
0!
0'
#301840000000
1!
b10 %
1'
b10 +
#301850000000
0!
0'
#301860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#301870000000
0!
0'
#301880000000
1!
b100 %
1'
b100 +
#301890000000
0!
0'
#301900000000
1!
b101 %
1'
b101 +
#301910000000
0!
0'
#301920000000
1!
0$
b110 %
1'
0*
b110 +
#301930000000
0!
0'
#301940000000
1!
b111 %
1'
b111 +
#301950000000
0!
0'
#301960000000
1!
b1000 %
1'
b1000 +
#301970000000
0!
0'
#301980000000
1!
b1001 %
1'
b1001 +
#301990000000
0!
0'
#302000000000
1!
b0 %
1'
b0 +
#302010000000
0!
0'
#302020000000
1!
1$
b1 %
1'
1*
b1 +
#302030000000
0!
0'
#302040000000
1!
b10 %
1'
b10 +
#302050000000
0!
0'
#302060000000
1!
b11 %
1'
b11 +
#302070000000
1"
1(
#302080000000
0!
0"
b100 &
0'
0(
b100 ,
#302090000000
1!
b100 %
1'
b100 +
#302100000000
0!
0'
#302110000000
1!
b101 %
1'
b101 +
#302120000000
0!
0'
#302130000000
1!
b110 %
1'
b110 +
#302140000000
0!
0'
#302150000000
1!
b111 %
1'
b111 +
#302160000000
0!
0'
#302170000000
1!
0$
b1000 %
1'
0*
b1000 +
#302180000000
0!
0'
#302190000000
1!
b1001 %
1'
b1001 +
#302200000000
0!
0'
#302210000000
1!
b0 %
1'
b0 +
#302220000000
0!
0'
#302230000000
1!
1$
b1 %
1'
1*
b1 +
#302240000000
0!
0'
#302250000000
1!
b10 %
1'
b10 +
#302260000000
0!
0'
#302270000000
1!
b11 %
1'
b11 +
#302280000000
0!
0'
#302290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#302300000000
0!
0'
#302310000000
1!
b101 %
1'
b101 +
#302320000000
0!
0'
#302330000000
1!
0$
b110 %
1'
0*
b110 +
#302340000000
0!
0'
#302350000000
1!
b111 %
1'
b111 +
#302360000000
0!
0'
#302370000000
1!
b1000 %
1'
b1000 +
#302380000000
0!
0'
#302390000000
1!
b1001 %
1'
b1001 +
#302400000000
0!
0'
#302410000000
1!
b0 %
1'
b0 +
#302420000000
0!
0'
#302430000000
1!
1$
b1 %
1'
1*
b1 +
#302440000000
0!
0'
#302450000000
1!
b10 %
1'
b10 +
#302460000000
0!
0'
#302470000000
1!
b11 %
1'
b11 +
#302480000000
0!
0'
#302490000000
1!
b100 %
1'
b100 +
#302500000000
1"
1(
#302510000000
0!
0"
b100 &
0'
0(
b100 ,
#302520000000
1!
b101 %
1'
b101 +
#302530000000
0!
0'
#302540000000
1!
b110 %
1'
b110 +
#302550000000
0!
0'
#302560000000
1!
b111 %
1'
b111 +
#302570000000
0!
0'
#302580000000
1!
0$
b1000 %
1'
0*
b1000 +
#302590000000
0!
0'
#302600000000
1!
b1001 %
1'
b1001 +
#302610000000
0!
0'
#302620000000
1!
b0 %
1'
b0 +
#302630000000
0!
0'
#302640000000
1!
1$
b1 %
1'
1*
b1 +
#302650000000
0!
0'
#302660000000
1!
b10 %
1'
b10 +
#302670000000
0!
0'
#302680000000
1!
b11 %
1'
b11 +
#302690000000
0!
0'
#302700000000
1!
b100 %
1'
b100 +
#302710000000
0!
0'
#302720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#302730000000
0!
0'
#302740000000
1!
0$
b110 %
1'
0*
b110 +
#302750000000
0!
0'
#302760000000
1!
b111 %
1'
b111 +
#302770000000
0!
0'
#302780000000
1!
b1000 %
1'
b1000 +
#302790000000
0!
0'
#302800000000
1!
b1001 %
1'
b1001 +
#302810000000
0!
0'
#302820000000
1!
b0 %
1'
b0 +
#302830000000
0!
0'
#302840000000
1!
1$
b1 %
1'
1*
b1 +
#302850000000
0!
0'
#302860000000
1!
b10 %
1'
b10 +
#302870000000
0!
0'
#302880000000
1!
b11 %
1'
b11 +
#302890000000
0!
0'
#302900000000
1!
b100 %
1'
b100 +
#302910000000
0!
0'
#302920000000
1!
b101 %
1'
b101 +
#302930000000
1"
1(
#302940000000
0!
0"
b100 &
0'
0(
b100 ,
#302950000000
1!
b110 %
1'
b110 +
#302960000000
0!
0'
#302970000000
1!
b111 %
1'
b111 +
#302980000000
0!
0'
#302990000000
1!
0$
b1000 %
1'
0*
b1000 +
#303000000000
0!
0'
#303010000000
1!
b1001 %
1'
b1001 +
#303020000000
0!
0'
#303030000000
1!
b0 %
1'
b0 +
#303040000000
0!
0'
#303050000000
1!
1$
b1 %
1'
1*
b1 +
#303060000000
0!
0'
#303070000000
1!
b10 %
1'
b10 +
#303080000000
0!
0'
#303090000000
1!
b11 %
1'
b11 +
#303100000000
0!
0'
#303110000000
1!
b100 %
1'
b100 +
#303120000000
0!
0'
#303130000000
1!
b101 %
1'
b101 +
#303140000000
0!
0'
#303150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#303160000000
0!
0'
#303170000000
1!
b111 %
1'
b111 +
#303180000000
0!
0'
#303190000000
1!
b1000 %
1'
b1000 +
#303200000000
0!
0'
#303210000000
1!
b1001 %
1'
b1001 +
#303220000000
0!
0'
#303230000000
1!
b0 %
1'
b0 +
#303240000000
0!
0'
#303250000000
1!
1$
b1 %
1'
1*
b1 +
#303260000000
0!
0'
#303270000000
1!
b10 %
1'
b10 +
#303280000000
0!
0'
#303290000000
1!
b11 %
1'
b11 +
#303300000000
0!
0'
#303310000000
1!
b100 %
1'
b100 +
#303320000000
0!
0'
#303330000000
1!
b101 %
1'
b101 +
#303340000000
0!
0'
#303350000000
1!
0$
b110 %
1'
0*
b110 +
#303360000000
1"
1(
#303370000000
0!
0"
b100 &
0'
0(
b100 ,
#303380000000
1!
1$
b111 %
1'
1*
b111 +
#303390000000
0!
0'
#303400000000
1!
0$
b1000 %
1'
0*
b1000 +
#303410000000
0!
0'
#303420000000
1!
b1001 %
1'
b1001 +
#303430000000
0!
0'
#303440000000
1!
b0 %
1'
b0 +
#303450000000
0!
0'
#303460000000
1!
1$
b1 %
1'
1*
b1 +
#303470000000
0!
0'
#303480000000
1!
b10 %
1'
b10 +
#303490000000
0!
0'
#303500000000
1!
b11 %
1'
b11 +
#303510000000
0!
0'
#303520000000
1!
b100 %
1'
b100 +
#303530000000
0!
0'
#303540000000
1!
b101 %
1'
b101 +
#303550000000
0!
0'
#303560000000
1!
b110 %
1'
b110 +
#303570000000
0!
0'
#303580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#303590000000
0!
0'
#303600000000
1!
b1000 %
1'
b1000 +
#303610000000
0!
0'
#303620000000
1!
b1001 %
1'
b1001 +
#303630000000
0!
0'
#303640000000
1!
b0 %
1'
b0 +
#303650000000
0!
0'
#303660000000
1!
1$
b1 %
1'
1*
b1 +
#303670000000
0!
0'
#303680000000
1!
b10 %
1'
b10 +
#303690000000
0!
0'
#303700000000
1!
b11 %
1'
b11 +
#303710000000
0!
0'
#303720000000
1!
b100 %
1'
b100 +
#303730000000
0!
0'
#303740000000
1!
b101 %
1'
b101 +
#303750000000
0!
0'
#303760000000
1!
0$
b110 %
1'
0*
b110 +
#303770000000
0!
0'
#303780000000
1!
b111 %
1'
b111 +
#303790000000
1"
1(
#303800000000
0!
0"
b100 &
0'
0(
b100 ,
#303810000000
1!
b1000 %
1'
b1000 +
#303820000000
0!
0'
#303830000000
1!
b1001 %
1'
b1001 +
#303840000000
0!
0'
#303850000000
1!
b0 %
1'
b0 +
#303860000000
0!
0'
#303870000000
1!
1$
b1 %
1'
1*
b1 +
#303880000000
0!
0'
#303890000000
1!
b10 %
1'
b10 +
#303900000000
0!
0'
#303910000000
1!
b11 %
1'
b11 +
#303920000000
0!
0'
#303930000000
1!
b100 %
1'
b100 +
#303940000000
0!
0'
#303950000000
1!
b101 %
1'
b101 +
#303960000000
0!
0'
#303970000000
1!
b110 %
1'
b110 +
#303980000000
0!
0'
#303990000000
1!
b111 %
1'
b111 +
#304000000000
0!
0'
#304010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#304020000000
0!
0'
#304030000000
1!
b1001 %
1'
b1001 +
#304040000000
0!
0'
#304050000000
1!
b0 %
1'
b0 +
#304060000000
0!
0'
#304070000000
1!
1$
b1 %
1'
1*
b1 +
#304080000000
0!
0'
#304090000000
1!
b10 %
1'
b10 +
#304100000000
0!
0'
#304110000000
1!
b11 %
1'
b11 +
#304120000000
0!
0'
#304130000000
1!
b100 %
1'
b100 +
#304140000000
0!
0'
#304150000000
1!
b101 %
1'
b101 +
#304160000000
0!
0'
#304170000000
1!
0$
b110 %
1'
0*
b110 +
#304180000000
0!
0'
#304190000000
1!
b111 %
1'
b111 +
#304200000000
0!
0'
#304210000000
1!
b1000 %
1'
b1000 +
#304220000000
1"
1(
#304230000000
0!
0"
b100 &
0'
0(
b100 ,
#304240000000
1!
b1001 %
1'
b1001 +
#304250000000
0!
0'
#304260000000
1!
b0 %
1'
b0 +
#304270000000
0!
0'
#304280000000
1!
1$
b1 %
1'
1*
b1 +
#304290000000
0!
0'
#304300000000
1!
b10 %
1'
b10 +
#304310000000
0!
0'
#304320000000
1!
b11 %
1'
b11 +
#304330000000
0!
0'
#304340000000
1!
b100 %
1'
b100 +
#304350000000
0!
0'
#304360000000
1!
b101 %
1'
b101 +
#304370000000
0!
0'
#304380000000
1!
b110 %
1'
b110 +
#304390000000
0!
0'
#304400000000
1!
b111 %
1'
b111 +
#304410000000
0!
0'
#304420000000
1!
0$
b1000 %
1'
0*
b1000 +
#304430000000
0!
0'
#304440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#304450000000
0!
0'
#304460000000
1!
b0 %
1'
b0 +
#304470000000
0!
0'
#304480000000
1!
1$
b1 %
1'
1*
b1 +
#304490000000
0!
0'
#304500000000
1!
b10 %
1'
b10 +
#304510000000
0!
0'
#304520000000
1!
b11 %
1'
b11 +
#304530000000
0!
0'
#304540000000
1!
b100 %
1'
b100 +
#304550000000
0!
0'
#304560000000
1!
b101 %
1'
b101 +
#304570000000
0!
0'
#304580000000
1!
0$
b110 %
1'
0*
b110 +
#304590000000
0!
0'
#304600000000
1!
b111 %
1'
b111 +
#304610000000
0!
0'
#304620000000
1!
b1000 %
1'
b1000 +
#304630000000
0!
0'
#304640000000
1!
b1001 %
1'
b1001 +
#304650000000
1"
1(
#304660000000
0!
0"
b100 &
0'
0(
b100 ,
#304670000000
1!
b0 %
1'
b0 +
#304680000000
0!
0'
#304690000000
1!
1$
b1 %
1'
1*
b1 +
#304700000000
0!
0'
#304710000000
1!
b10 %
1'
b10 +
#304720000000
0!
0'
#304730000000
1!
b11 %
1'
b11 +
#304740000000
0!
0'
#304750000000
1!
b100 %
1'
b100 +
#304760000000
0!
0'
#304770000000
1!
b101 %
1'
b101 +
#304780000000
0!
0'
#304790000000
1!
b110 %
1'
b110 +
#304800000000
0!
0'
#304810000000
1!
b111 %
1'
b111 +
#304820000000
0!
0'
#304830000000
1!
0$
b1000 %
1'
0*
b1000 +
#304840000000
0!
0'
#304850000000
1!
b1001 %
1'
b1001 +
#304860000000
0!
0'
#304870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#304880000000
0!
0'
#304890000000
1!
1$
b1 %
1'
1*
b1 +
#304900000000
0!
0'
#304910000000
1!
b10 %
1'
b10 +
#304920000000
0!
0'
#304930000000
1!
b11 %
1'
b11 +
#304940000000
0!
0'
#304950000000
1!
b100 %
1'
b100 +
#304960000000
0!
0'
#304970000000
1!
b101 %
1'
b101 +
#304980000000
0!
0'
#304990000000
1!
0$
b110 %
1'
0*
b110 +
#305000000000
0!
0'
#305010000000
1!
b111 %
1'
b111 +
#305020000000
0!
0'
#305030000000
1!
b1000 %
1'
b1000 +
#305040000000
0!
0'
#305050000000
1!
b1001 %
1'
b1001 +
#305060000000
0!
0'
#305070000000
1!
b0 %
1'
b0 +
#305080000000
1"
1(
#305090000000
0!
0"
b100 &
0'
0(
b100 ,
#305100000000
1!
1$
b1 %
1'
1*
b1 +
#305110000000
0!
0'
#305120000000
1!
b10 %
1'
b10 +
#305130000000
0!
0'
#305140000000
1!
b11 %
1'
b11 +
#305150000000
0!
0'
#305160000000
1!
b100 %
1'
b100 +
#305170000000
0!
0'
#305180000000
1!
b101 %
1'
b101 +
#305190000000
0!
0'
#305200000000
1!
b110 %
1'
b110 +
#305210000000
0!
0'
#305220000000
1!
b111 %
1'
b111 +
#305230000000
0!
0'
#305240000000
1!
0$
b1000 %
1'
0*
b1000 +
#305250000000
0!
0'
#305260000000
1!
b1001 %
1'
b1001 +
#305270000000
0!
0'
#305280000000
1!
b0 %
1'
b0 +
#305290000000
0!
0'
#305300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#305310000000
0!
0'
#305320000000
1!
b10 %
1'
b10 +
#305330000000
0!
0'
#305340000000
1!
b11 %
1'
b11 +
#305350000000
0!
0'
#305360000000
1!
b100 %
1'
b100 +
#305370000000
0!
0'
#305380000000
1!
b101 %
1'
b101 +
#305390000000
0!
0'
#305400000000
1!
0$
b110 %
1'
0*
b110 +
#305410000000
0!
0'
#305420000000
1!
b111 %
1'
b111 +
#305430000000
0!
0'
#305440000000
1!
b1000 %
1'
b1000 +
#305450000000
0!
0'
#305460000000
1!
b1001 %
1'
b1001 +
#305470000000
0!
0'
#305480000000
1!
b0 %
1'
b0 +
#305490000000
0!
0'
#305500000000
1!
1$
b1 %
1'
1*
b1 +
#305510000000
1"
1(
#305520000000
0!
0"
b100 &
0'
0(
b100 ,
#305530000000
1!
b10 %
1'
b10 +
#305540000000
0!
0'
#305550000000
1!
b11 %
1'
b11 +
#305560000000
0!
0'
#305570000000
1!
b100 %
1'
b100 +
#305580000000
0!
0'
#305590000000
1!
b101 %
1'
b101 +
#305600000000
0!
0'
#305610000000
1!
b110 %
1'
b110 +
#305620000000
0!
0'
#305630000000
1!
b111 %
1'
b111 +
#305640000000
0!
0'
#305650000000
1!
0$
b1000 %
1'
0*
b1000 +
#305660000000
0!
0'
#305670000000
1!
b1001 %
1'
b1001 +
#305680000000
0!
0'
#305690000000
1!
b0 %
1'
b0 +
#305700000000
0!
0'
#305710000000
1!
1$
b1 %
1'
1*
b1 +
#305720000000
0!
0'
#305730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#305740000000
0!
0'
#305750000000
1!
b11 %
1'
b11 +
#305760000000
0!
0'
#305770000000
1!
b100 %
1'
b100 +
#305780000000
0!
0'
#305790000000
1!
b101 %
1'
b101 +
#305800000000
0!
0'
#305810000000
1!
0$
b110 %
1'
0*
b110 +
#305820000000
0!
0'
#305830000000
1!
b111 %
1'
b111 +
#305840000000
0!
0'
#305850000000
1!
b1000 %
1'
b1000 +
#305860000000
0!
0'
#305870000000
1!
b1001 %
1'
b1001 +
#305880000000
0!
0'
#305890000000
1!
b0 %
1'
b0 +
#305900000000
0!
0'
#305910000000
1!
1$
b1 %
1'
1*
b1 +
#305920000000
0!
0'
#305930000000
1!
b10 %
1'
b10 +
#305940000000
1"
1(
#305950000000
0!
0"
b100 &
0'
0(
b100 ,
#305960000000
1!
b11 %
1'
b11 +
#305970000000
0!
0'
#305980000000
1!
b100 %
1'
b100 +
#305990000000
0!
0'
#306000000000
1!
b101 %
1'
b101 +
#306010000000
0!
0'
#306020000000
1!
b110 %
1'
b110 +
#306030000000
0!
0'
#306040000000
1!
b111 %
1'
b111 +
#306050000000
0!
0'
#306060000000
1!
0$
b1000 %
1'
0*
b1000 +
#306070000000
0!
0'
#306080000000
1!
b1001 %
1'
b1001 +
#306090000000
0!
0'
#306100000000
1!
b0 %
1'
b0 +
#306110000000
0!
0'
#306120000000
1!
1$
b1 %
1'
1*
b1 +
#306130000000
0!
0'
#306140000000
1!
b10 %
1'
b10 +
#306150000000
0!
0'
#306160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#306170000000
0!
0'
#306180000000
1!
b100 %
1'
b100 +
#306190000000
0!
0'
#306200000000
1!
b101 %
1'
b101 +
#306210000000
0!
0'
#306220000000
1!
0$
b110 %
1'
0*
b110 +
#306230000000
0!
0'
#306240000000
1!
b111 %
1'
b111 +
#306250000000
0!
0'
#306260000000
1!
b1000 %
1'
b1000 +
#306270000000
0!
0'
#306280000000
1!
b1001 %
1'
b1001 +
#306290000000
0!
0'
#306300000000
1!
b0 %
1'
b0 +
#306310000000
0!
0'
#306320000000
1!
1$
b1 %
1'
1*
b1 +
#306330000000
0!
0'
#306340000000
1!
b10 %
1'
b10 +
#306350000000
0!
0'
#306360000000
1!
b11 %
1'
b11 +
#306370000000
1"
1(
#306380000000
0!
0"
b100 &
0'
0(
b100 ,
#306390000000
1!
b100 %
1'
b100 +
#306400000000
0!
0'
#306410000000
1!
b101 %
1'
b101 +
#306420000000
0!
0'
#306430000000
1!
b110 %
1'
b110 +
#306440000000
0!
0'
#306450000000
1!
b111 %
1'
b111 +
#306460000000
0!
0'
#306470000000
1!
0$
b1000 %
1'
0*
b1000 +
#306480000000
0!
0'
#306490000000
1!
b1001 %
1'
b1001 +
#306500000000
0!
0'
#306510000000
1!
b0 %
1'
b0 +
#306520000000
0!
0'
#306530000000
1!
1$
b1 %
1'
1*
b1 +
#306540000000
0!
0'
#306550000000
1!
b10 %
1'
b10 +
#306560000000
0!
0'
#306570000000
1!
b11 %
1'
b11 +
#306580000000
0!
0'
#306590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#306600000000
0!
0'
#306610000000
1!
b101 %
1'
b101 +
#306620000000
0!
0'
#306630000000
1!
0$
b110 %
1'
0*
b110 +
#306640000000
0!
0'
#306650000000
1!
b111 %
1'
b111 +
#306660000000
0!
0'
#306670000000
1!
b1000 %
1'
b1000 +
#306680000000
0!
0'
#306690000000
1!
b1001 %
1'
b1001 +
#306700000000
0!
0'
#306710000000
1!
b0 %
1'
b0 +
#306720000000
0!
0'
#306730000000
1!
1$
b1 %
1'
1*
b1 +
#306740000000
0!
0'
#306750000000
1!
b10 %
1'
b10 +
#306760000000
0!
0'
#306770000000
1!
b11 %
1'
b11 +
#306780000000
0!
0'
#306790000000
1!
b100 %
1'
b100 +
#306800000000
1"
1(
#306810000000
0!
0"
b100 &
0'
0(
b100 ,
#306820000000
1!
b101 %
1'
b101 +
#306830000000
0!
0'
#306840000000
1!
b110 %
1'
b110 +
#306850000000
0!
0'
#306860000000
1!
b111 %
1'
b111 +
#306870000000
0!
0'
#306880000000
1!
0$
b1000 %
1'
0*
b1000 +
#306890000000
0!
0'
#306900000000
1!
b1001 %
1'
b1001 +
#306910000000
0!
0'
#306920000000
1!
b0 %
1'
b0 +
#306930000000
0!
0'
#306940000000
1!
1$
b1 %
1'
1*
b1 +
#306950000000
0!
0'
#306960000000
1!
b10 %
1'
b10 +
#306970000000
0!
0'
#306980000000
1!
b11 %
1'
b11 +
#306990000000
0!
0'
#307000000000
1!
b100 %
1'
b100 +
#307010000000
0!
0'
#307020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#307030000000
0!
0'
#307040000000
1!
0$
b110 %
1'
0*
b110 +
#307050000000
0!
0'
#307060000000
1!
b111 %
1'
b111 +
#307070000000
0!
0'
#307080000000
1!
b1000 %
1'
b1000 +
#307090000000
0!
0'
#307100000000
1!
b1001 %
1'
b1001 +
#307110000000
0!
0'
#307120000000
1!
b0 %
1'
b0 +
#307130000000
0!
0'
#307140000000
1!
1$
b1 %
1'
1*
b1 +
#307150000000
0!
0'
#307160000000
1!
b10 %
1'
b10 +
#307170000000
0!
0'
#307180000000
1!
b11 %
1'
b11 +
#307190000000
0!
0'
#307200000000
1!
b100 %
1'
b100 +
#307210000000
0!
0'
#307220000000
1!
b101 %
1'
b101 +
#307230000000
1"
1(
#307240000000
0!
0"
b100 &
0'
0(
b100 ,
#307250000000
1!
b110 %
1'
b110 +
#307260000000
0!
0'
#307270000000
1!
b111 %
1'
b111 +
#307280000000
0!
0'
#307290000000
1!
0$
b1000 %
1'
0*
b1000 +
#307300000000
0!
0'
#307310000000
1!
b1001 %
1'
b1001 +
#307320000000
0!
0'
#307330000000
1!
b0 %
1'
b0 +
#307340000000
0!
0'
#307350000000
1!
1$
b1 %
1'
1*
b1 +
#307360000000
0!
0'
#307370000000
1!
b10 %
1'
b10 +
#307380000000
0!
0'
#307390000000
1!
b11 %
1'
b11 +
#307400000000
0!
0'
#307410000000
1!
b100 %
1'
b100 +
#307420000000
0!
0'
#307430000000
1!
b101 %
1'
b101 +
#307440000000
0!
0'
#307450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#307460000000
0!
0'
#307470000000
1!
b111 %
1'
b111 +
#307480000000
0!
0'
#307490000000
1!
b1000 %
1'
b1000 +
#307500000000
0!
0'
#307510000000
1!
b1001 %
1'
b1001 +
#307520000000
0!
0'
#307530000000
1!
b0 %
1'
b0 +
#307540000000
0!
0'
#307550000000
1!
1$
b1 %
1'
1*
b1 +
#307560000000
0!
0'
#307570000000
1!
b10 %
1'
b10 +
#307580000000
0!
0'
#307590000000
1!
b11 %
1'
b11 +
#307600000000
0!
0'
#307610000000
1!
b100 %
1'
b100 +
#307620000000
0!
0'
#307630000000
1!
b101 %
1'
b101 +
#307640000000
0!
0'
#307650000000
1!
0$
b110 %
1'
0*
b110 +
#307660000000
1"
1(
#307670000000
0!
0"
b100 &
0'
0(
b100 ,
#307680000000
1!
1$
b111 %
1'
1*
b111 +
#307690000000
0!
0'
#307700000000
1!
0$
b1000 %
1'
0*
b1000 +
#307710000000
0!
0'
#307720000000
1!
b1001 %
1'
b1001 +
#307730000000
0!
0'
#307740000000
1!
b0 %
1'
b0 +
#307750000000
0!
0'
#307760000000
1!
1$
b1 %
1'
1*
b1 +
#307770000000
0!
0'
#307780000000
1!
b10 %
1'
b10 +
#307790000000
0!
0'
#307800000000
1!
b11 %
1'
b11 +
#307810000000
0!
0'
#307820000000
1!
b100 %
1'
b100 +
#307830000000
0!
0'
#307840000000
1!
b101 %
1'
b101 +
#307850000000
0!
0'
#307860000000
1!
b110 %
1'
b110 +
#307870000000
0!
0'
#307880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#307890000000
0!
0'
#307900000000
1!
b1000 %
1'
b1000 +
#307910000000
0!
0'
#307920000000
1!
b1001 %
1'
b1001 +
#307930000000
0!
0'
#307940000000
1!
b0 %
1'
b0 +
#307950000000
0!
0'
#307960000000
1!
1$
b1 %
1'
1*
b1 +
#307970000000
0!
0'
#307980000000
1!
b10 %
1'
b10 +
#307990000000
0!
0'
#308000000000
1!
b11 %
1'
b11 +
#308010000000
0!
0'
#308020000000
1!
b100 %
1'
b100 +
#308030000000
0!
0'
#308040000000
1!
b101 %
1'
b101 +
#308050000000
0!
0'
#308060000000
1!
0$
b110 %
1'
0*
b110 +
#308070000000
0!
0'
#308080000000
1!
b111 %
1'
b111 +
#308090000000
1"
1(
#308100000000
0!
0"
b100 &
0'
0(
b100 ,
#308110000000
1!
b1000 %
1'
b1000 +
#308120000000
0!
0'
#308130000000
1!
b1001 %
1'
b1001 +
#308140000000
0!
0'
#308150000000
1!
b0 %
1'
b0 +
#308160000000
0!
0'
#308170000000
1!
1$
b1 %
1'
1*
b1 +
#308180000000
0!
0'
#308190000000
1!
b10 %
1'
b10 +
#308200000000
0!
0'
#308210000000
1!
b11 %
1'
b11 +
#308220000000
0!
0'
#308230000000
1!
b100 %
1'
b100 +
#308240000000
0!
0'
#308250000000
1!
b101 %
1'
b101 +
#308260000000
0!
0'
#308270000000
1!
b110 %
1'
b110 +
#308280000000
0!
0'
#308290000000
1!
b111 %
1'
b111 +
#308300000000
0!
0'
#308310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#308320000000
0!
0'
#308330000000
1!
b1001 %
1'
b1001 +
#308340000000
0!
0'
#308350000000
1!
b0 %
1'
b0 +
#308360000000
0!
0'
#308370000000
1!
1$
b1 %
1'
1*
b1 +
#308380000000
0!
0'
#308390000000
1!
b10 %
1'
b10 +
#308400000000
0!
0'
#308410000000
1!
b11 %
1'
b11 +
#308420000000
0!
0'
#308430000000
1!
b100 %
1'
b100 +
#308440000000
0!
0'
#308450000000
1!
b101 %
1'
b101 +
#308460000000
0!
0'
#308470000000
1!
0$
b110 %
1'
0*
b110 +
#308480000000
0!
0'
#308490000000
1!
b111 %
1'
b111 +
#308500000000
0!
0'
#308510000000
1!
b1000 %
1'
b1000 +
#308520000000
1"
1(
#308530000000
0!
0"
b100 &
0'
0(
b100 ,
#308540000000
1!
b1001 %
1'
b1001 +
#308550000000
0!
0'
#308560000000
1!
b0 %
1'
b0 +
#308570000000
0!
0'
#308580000000
1!
1$
b1 %
1'
1*
b1 +
#308590000000
0!
0'
#308600000000
1!
b10 %
1'
b10 +
#308610000000
0!
0'
#308620000000
1!
b11 %
1'
b11 +
#308630000000
0!
0'
#308640000000
1!
b100 %
1'
b100 +
#308650000000
0!
0'
#308660000000
1!
b101 %
1'
b101 +
#308670000000
0!
0'
#308680000000
1!
b110 %
1'
b110 +
#308690000000
0!
0'
#308700000000
1!
b111 %
1'
b111 +
#308710000000
0!
0'
#308720000000
1!
0$
b1000 %
1'
0*
b1000 +
#308730000000
0!
0'
#308740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#308750000000
0!
0'
#308760000000
1!
b0 %
1'
b0 +
#308770000000
0!
0'
#308780000000
1!
1$
b1 %
1'
1*
b1 +
#308790000000
0!
0'
#308800000000
1!
b10 %
1'
b10 +
#308810000000
0!
0'
#308820000000
1!
b11 %
1'
b11 +
#308830000000
0!
0'
#308840000000
1!
b100 %
1'
b100 +
#308850000000
0!
0'
#308860000000
1!
b101 %
1'
b101 +
#308870000000
0!
0'
#308880000000
1!
0$
b110 %
1'
0*
b110 +
#308890000000
0!
0'
#308900000000
1!
b111 %
1'
b111 +
#308910000000
0!
0'
#308920000000
1!
b1000 %
1'
b1000 +
#308930000000
0!
0'
#308940000000
1!
b1001 %
1'
b1001 +
#308950000000
1"
1(
#308960000000
0!
0"
b100 &
0'
0(
b100 ,
#308970000000
1!
b0 %
1'
b0 +
#308980000000
0!
0'
#308990000000
1!
1$
b1 %
1'
1*
b1 +
#309000000000
0!
0'
#309010000000
1!
b10 %
1'
b10 +
#309020000000
0!
0'
#309030000000
1!
b11 %
1'
b11 +
#309040000000
0!
0'
#309050000000
1!
b100 %
1'
b100 +
#309060000000
0!
0'
#309070000000
1!
b101 %
1'
b101 +
#309080000000
0!
0'
#309090000000
1!
b110 %
1'
b110 +
#309100000000
0!
0'
#309110000000
1!
b111 %
1'
b111 +
#309120000000
0!
0'
#309130000000
1!
0$
b1000 %
1'
0*
b1000 +
#309140000000
0!
0'
#309150000000
1!
b1001 %
1'
b1001 +
#309160000000
0!
0'
#309170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#309180000000
0!
0'
#309190000000
1!
1$
b1 %
1'
1*
b1 +
#309200000000
0!
0'
#309210000000
1!
b10 %
1'
b10 +
#309220000000
0!
0'
#309230000000
1!
b11 %
1'
b11 +
#309240000000
0!
0'
#309250000000
1!
b100 %
1'
b100 +
#309260000000
0!
0'
#309270000000
1!
b101 %
1'
b101 +
#309280000000
0!
0'
#309290000000
1!
0$
b110 %
1'
0*
b110 +
#309300000000
0!
0'
#309310000000
1!
b111 %
1'
b111 +
#309320000000
0!
0'
#309330000000
1!
b1000 %
1'
b1000 +
#309340000000
0!
0'
#309350000000
1!
b1001 %
1'
b1001 +
#309360000000
0!
0'
#309370000000
1!
b0 %
1'
b0 +
#309380000000
1"
1(
#309390000000
0!
0"
b100 &
0'
0(
b100 ,
#309400000000
1!
1$
b1 %
1'
1*
b1 +
#309410000000
0!
0'
#309420000000
1!
b10 %
1'
b10 +
#309430000000
0!
0'
#309440000000
1!
b11 %
1'
b11 +
#309450000000
0!
0'
#309460000000
1!
b100 %
1'
b100 +
#309470000000
0!
0'
#309480000000
1!
b101 %
1'
b101 +
#309490000000
0!
0'
#309500000000
1!
b110 %
1'
b110 +
#309510000000
0!
0'
#309520000000
1!
b111 %
1'
b111 +
#309530000000
0!
0'
#309540000000
1!
0$
b1000 %
1'
0*
b1000 +
#309550000000
0!
0'
#309560000000
1!
b1001 %
1'
b1001 +
#309570000000
0!
0'
#309580000000
1!
b0 %
1'
b0 +
#309590000000
0!
0'
#309600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#309610000000
0!
0'
#309620000000
1!
b10 %
1'
b10 +
#309630000000
0!
0'
#309640000000
1!
b11 %
1'
b11 +
#309650000000
0!
0'
#309660000000
1!
b100 %
1'
b100 +
#309670000000
0!
0'
#309680000000
1!
b101 %
1'
b101 +
#309690000000
0!
0'
#309700000000
1!
0$
b110 %
1'
0*
b110 +
#309710000000
0!
0'
#309720000000
1!
b111 %
1'
b111 +
#309730000000
0!
0'
#309740000000
1!
b1000 %
1'
b1000 +
#309750000000
0!
0'
#309760000000
1!
b1001 %
1'
b1001 +
#309770000000
0!
0'
#309780000000
1!
b0 %
1'
b0 +
#309790000000
0!
0'
#309800000000
1!
1$
b1 %
1'
1*
b1 +
#309810000000
1"
1(
#309820000000
0!
0"
b100 &
0'
0(
b100 ,
#309830000000
1!
b10 %
1'
b10 +
#309840000000
0!
0'
#309850000000
1!
b11 %
1'
b11 +
#309860000000
0!
0'
#309870000000
1!
b100 %
1'
b100 +
#309880000000
0!
0'
#309890000000
1!
b101 %
1'
b101 +
#309900000000
0!
0'
#309910000000
1!
b110 %
1'
b110 +
#309920000000
0!
0'
#309930000000
1!
b111 %
1'
b111 +
#309940000000
0!
0'
#309950000000
1!
0$
b1000 %
1'
0*
b1000 +
#309960000000
0!
0'
#309970000000
1!
b1001 %
1'
b1001 +
#309980000000
0!
0'
#309990000000
1!
b0 %
1'
b0 +
#310000000000
0!
0'
#310010000000
1!
1$
b1 %
1'
1*
b1 +
#310020000000
0!
0'
#310030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#310040000000
0!
0'
#310050000000
1!
b11 %
1'
b11 +
#310060000000
0!
0'
#310070000000
1!
b100 %
1'
b100 +
#310080000000
0!
0'
#310090000000
1!
b101 %
1'
b101 +
#310100000000
0!
0'
#310110000000
1!
0$
b110 %
1'
0*
b110 +
#310120000000
0!
0'
#310130000000
1!
b111 %
1'
b111 +
#310140000000
0!
0'
#310150000000
1!
b1000 %
1'
b1000 +
#310160000000
0!
0'
#310170000000
1!
b1001 %
1'
b1001 +
#310180000000
0!
0'
#310190000000
1!
b0 %
1'
b0 +
#310200000000
0!
0'
#310210000000
1!
1$
b1 %
1'
1*
b1 +
#310220000000
0!
0'
#310230000000
1!
b10 %
1'
b10 +
#310240000000
1"
1(
#310250000000
0!
0"
b100 &
0'
0(
b100 ,
#310260000000
1!
b11 %
1'
b11 +
#310270000000
0!
0'
#310280000000
1!
b100 %
1'
b100 +
#310290000000
0!
0'
#310300000000
1!
b101 %
1'
b101 +
#310310000000
0!
0'
#310320000000
1!
b110 %
1'
b110 +
#310330000000
0!
0'
#310340000000
1!
b111 %
1'
b111 +
#310350000000
0!
0'
#310360000000
1!
0$
b1000 %
1'
0*
b1000 +
#310370000000
0!
0'
#310380000000
1!
b1001 %
1'
b1001 +
#310390000000
0!
0'
#310400000000
1!
b0 %
1'
b0 +
#310410000000
0!
0'
#310420000000
1!
1$
b1 %
1'
1*
b1 +
#310430000000
0!
0'
#310440000000
1!
b10 %
1'
b10 +
#310450000000
0!
0'
#310460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#310470000000
0!
0'
#310480000000
1!
b100 %
1'
b100 +
#310490000000
0!
0'
#310500000000
1!
b101 %
1'
b101 +
#310510000000
0!
0'
#310520000000
1!
0$
b110 %
1'
0*
b110 +
#310530000000
0!
0'
#310540000000
1!
b111 %
1'
b111 +
#310550000000
0!
0'
#310560000000
1!
b1000 %
1'
b1000 +
#310570000000
0!
0'
#310580000000
1!
b1001 %
1'
b1001 +
#310590000000
0!
0'
#310600000000
1!
b0 %
1'
b0 +
#310610000000
0!
0'
#310620000000
1!
1$
b1 %
1'
1*
b1 +
#310630000000
0!
0'
#310640000000
1!
b10 %
1'
b10 +
#310650000000
0!
0'
#310660000000
1!
b11 %
1'
b11 +
#310670000000
1"
1(
#310680000000
0!
0"
b100 &
0'
0(
b100 ,
#310690000000
1!
b100 %
1'
b100 +
#310700000000
0!
0'
#310710000000
1!
b101 %
1'
b101 +
#310720000000
0!
0'
#310730000000
1!
b110 %
1'
b110 +
#310740000000
0!
0'
#310750000000
1!
b111 %
1'
b111 +
#310760000000
0!
0'
#310770000000
1!
0$
b1000 %
1'
0*
b1000 +
#310780000000
0!
0'
#310790000000
1!
b1001 %
1'
b1001 +
#310800000000
0!
0'
#310810000000
1!
b0 %
1'
b0 +
#310820000000
0!
0'
#310830000000
1!
1$
b1 %
1'
1*
b1 +
#310840000000
0!
0'
#310850000000
1!
b10 %
1'
b10 +
#310860000000
0!
0'
#310870000000
1!
b11 %
1'
b11 +
#310880000000
0!
0'
#310890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#310900000000
0!
0'
#310910000000
1!
b101 %
1'
b101 +
#310920000000
0!
0'
#310930000000
1!
0$
b110 %
1'
0*
b110 +
#310940000000
0!
0'
#310950000000
1!
b111 %
1'
b111 +
#310960000000
0!
0'
#310970000000
1!
b1000 %
1'
b1000 +
#310980000000
0!
0'
#310990000000
1!
b1001 %
1'
b1001 +
#311000000000
0!
0'
#311010000000
1!
b0 %
1'
b0 +
#311020000000
0!
0'
#311030000000
1!
1$
b1 %
1'
1*
b1 +
#311040000000
0!
0'
#311050000000
1!
b10 %
1'
b10 +
#311060000000
0!
0'
#311070000000
1!
b11 %
1'
b11 +
#311080000000
0!
0'
#311090000000
1!
b100 %
1'
b100 +
#311100000000
1"
1(
#311110000000
0!
0"
b100 &
0'
0(
b100 ,
#311120000000
1!
b101 %
1'
b101 +
#311130000000
0!
0'
#311140000000
1!
b110 %
1'
b110 +
#311150000000
0!
0'
#311160000000
1!
b111 %
1'
b111 +
#311170000000
0!
0'
#311180000000
1!
0$
b1000 %
1'
0*
b1000 +
#311190000000
0!
0'
#311200000000
1!
b1001 %
1'
b1001 +
#311210000000
0!
0'
#311220000000
1!
b0 %
1'
b0 +
#311230000000
0!
0'
#311240000000
1!
1$
b1 %
1'
1*
b1 +
#311250000000
0!
0'
#311260000000
1!
b10 %
1'
b10 +
#311270000000
0!
0'
#311280000000
1!
b11 %
1'
b11 +
#311290000000
0!
0'
#311300000000
1!
b100 %
1'
b100 +
#311310000000
0!
0'
#311320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#311330000000
0!
0'
#311340000000
1!
0$
b110 %
1'
0*
b110 +
#311350000000
0!
0'
#311360000000
1!
b111 %
1'
b111 +
#311370000000
0!
0'
#311380000000
1!
b1000 %
1'
b1000 +
#311390000000
0!
0'
#311400000000
1!
b1001 %
1'
b1001 +
#311410000000
0!
0'
#311420000000
1!
b0 %
1'
b0 +
#311430000000
0!
0'
#311440000000
1!
1$
b1 %
1'
1*
b1 +
#311450000000
0!
0'
#311460000000
1!
b10 %
1'
b10 +
#311470000000
0!
0'
#311480000000
1!
b11 %
1'
b11 +
#311490000000
0!
0'
#311500000000
1!
b100 %
1'
b100 +
#311510000000
0!
0'
#311520000000
1!
b101 %
1'
b101 +
#311530000000
1"
1(
#311540000000
0!
0"
b100 &
0'
0(
b100 ,
#311550000000
1!
b110 %
1'
b110 +
#311560000000
0!
0'
#311570000000
1!
b111 %
1'
b111 +
#311580000000
0!
0'
#311590000000
1!
0$
b1000 %
1'
0*
b1000 +
#311600000000
0!
0'
#311610000000
1!
b1001 %
1'
b1001 +
#311620000000
0!
0'
#311630000000
1!
b0 %
1'
b0 +
#311640000000
0!
0'
#311650000000
1!
1$
b1 %
1'
1*
b1 +
#311660000000
0!
0'
#311670000000
1!
b10 %
1'
b10 +
#311680000000
0!
0'
#311690000000
1!
b11 %
1'
b11 +
#311700000000
0!
0'
#311710000000
1!
b100 %
1'
b100 +
#311720000000
0!
0'
#311730000000
1!
b101 %
1'
b101 +
#311740000000
0!
0'
#311750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#311760000000
0!
0'
#311770000000
1!
b111 %
1'
b111 +
#311780000000
0!
0'
#311790000000
1!
b1000 %
1'
b1000 +
#311800000000
0!
0'
#311810000000
1!
b1001 %
1'
b1001 +
#311820000000
0!
0'
#311830000000
1!
b0 %
1'
b0 +
#311840000000
0!
0'
#311850000000
1!
1$
b1 %
1'
1*
b1 +
#311860000000
0!
0'
#311870000000
1!
b10 %
1'
b10 +
#311880000000
0!
0'
#311890000000
1!
b11 %
1'
b11 +
#311900000000
0!
0'
#311910000000
1!
b100 %
1'
b100 +
#311920000000
0!
0'
#311930000000
1!
b101 %
1'
b101 +
#311940000000
0!
0'
#311950000000
1!
0$
b110 %
1'
0*
b110 +
#311960000000
1"
1(
#311970000000
0!
0"
b100 &
0'
0(
b100 ,
#311980000000
1!
1$
b111 %
1'
1*
b111 +
#311990000000
0!
0'
#312000000000
1!
0$
b1000 %
1'
0*
b1000 +
#312010000000
0!
0'
#312020000000
1!
b1001 %
1'
b1001 +
#312030000000
0!
0'
#312040000000
1!
b0 %
1'
b0 +
#312050000000
0!
0'
#312060000000
1!
1$
b1 %
1'
1*
b1 +
#312070000000
0!
0'
#312080000000
1!
b10 %
1'
b10 +
#312090000000
0!
0'
#312100000000
1!
b11 %
1'
b11 +
#312110000000
0!
0'
#312120000000
1!
b100 %
1'
b100 +
#312130000000
0!
0'
#312140000000
1!
b101 %
1'
b101 +
#312150000000
0!
0'
#312160000000
1!
b110 %
1'
b110 +
#312170000000
0!
0'
#312180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#312190000000
0!
0'
#312200000000
1!
b1000 %
1'
b1000 +
#312210000000
0!
0'
#312220000000
1!
b1001 %
1'
b1001 +
#312230000000
0!
0'
#312240000000
1!
b0 %
1'
b0 +
#312250000000
0!
0'
#312260000000
1!
1$
b1 %
1'
1*
b1 +
#312270000000
0!
0'
#312280000000
1!
b10 %
1'
b10 +
#312290000000
0!
0'
#312300000000
1!
b11 %
1'
b11 +
#312310000000
0!
0'
#312320000000
1!
b100 %
1'
b100 +
#312330000000
0!
0'
#312340000000
1!
b101 %
1'
b101 +
#312350000000
0!
0'
#312360000000
1!
0$
b110 %
1'
0*
b110 +
#312370000000
0!
0'
#312380000000
1!
b111 %
1'
b111 +
#312390000000
1"
1(
#312400000000
0!
0"
b100 &
0'
0(
b100 ,
#312410000000
1!
b1000 %
1'
b1000 +
#312420000000
0!
0'
#312430000000
1!
b1001 %
1'
b1001 +
#312440000000
0!
0'
#312450000000
1!
b0 %
1'
b0 +
#312460000000
0!
0'
#312470000000
1!
1$
b1 %
1'
1*
b1 +
#312480000000
0!
0'
#312490000000
1!
b10 %
1'
b10 +
#312500000000
0!
0'
#312510000000
1!
b11 %
1'
b11 +
#312520000000
0!
0'
#312530000000
1!
b100 %
1'
b100 +
#312540000000
0!
0'
#312550000000
1!
b101 %
1'
b101 +
#312560000000
0!
0'
#312570000000
1!
b110 %
1'
b110 +
#312580000000
0!
0'
#312590000000
1!
b111 %
1'
b111 +
#312600000000
0!
0'
#312610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#312620000000
0!
0'
#312630000000
1!
b1001 %
1'
b1001 +
#312640000000
0!
0'
#312650000000
1!
b0 %
1'
b0 +
#312660000000
0!
0'
#312670000000
1!
1$
b1 %
1'
1*
b1 +
#312680000000
0!
0'
#312690000000
1!
b10 %
1'
b10 +
#312700000000
0!
0'
#312710000000
1!
b11 %
1'
b11 +
#312720000000
0!
0'
#312730000000
1!
b100 %
1'
b100 +
#312740000000
0!
0'
#312750000000
1!
b101 %
1'
b101 +
#312760000000
0!
0'
#312770000000
1!
0$
b110 %
1'
0*
b110 +
#312780000000
0!
0'
#312790000000
1!
b111 %
1'
b111 +
#312800000000
0!
0'
#312810000000
1!
b1000 %
1'
b1000 +
#312820000000
1"
1(
#312830000000
0!
0"
b100 &
0'
0(
b100 ,
#312840000000
1!
b1001 %
1'
b1001 +
#312850000000
0!
0'
#312860000000
1!
b0 %
1'
b0 +
#312870000000
0!
0'
#312880000000
1!
1$
b1 %
1'
1*
b1 +
#312890000000
0!
0'
#312900000000
1!
b10 %
1'
b10 +
#312910000000
0!
0'
#312920000000
1!
b11 %
1'
b11 +
#312930000000
0!
0'
#312940000000
1!
b100 %
1'
b100 +
#312950000000
0!
0'
#312960000000
1!
b101 %
1'
b101 +
#312970000000
0!
0'
#312980000000
1!
b110 %
1'
b110 +
#312990000000
0!
0'
#313000000000
1!
b111 %
1'
b111 +
#313010000000
0!
0'
#313020000000
1!
0$
b1000 %
1'
0*
b1000 +
#313030000000
0!
0'
#313040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#313050000000
0!
0'
#313060000000
1!
b0 %
1'
b0 +
#313070000000
0!
0'
#313080000000
1!
1$
b1 %
1'
1*
b1 +
#313090000000
0!
0'
#313100000000
1!
b10 %
1'
b10 +
#313110000000
0!
0'
#313120000000
1!
b11 %
1'
b11 +
#313130000000
0!
0'
#313140000000
1!
b100 %
1'
b100 +
#313150000000
0!
0'
#313160000000
1!
b101 %
1'
b101 +
#313170000000
0!
0'
#313180000000
1!
0$
b110 %
1'
0*
b110 +
#313190000000
0!
0'
#313200000000
1!
b111 %
1'
b111 +
#313210000000
0!
0'
#313220000000
1!
b1000 %
1'
b1000 +
#313230000000
0!
0'
#313240000000
1!
b1001 %
1'
b1001 +
#313250000000
1"
1(
#313260000000
0!
0"
b100 &
0'
0(
b100 ,
#313270000000
1!
b0 %
1'
b0 +
#313280000000
0!
0'
#313290000000
1!
1$
b1 %
1'
1*
b1 +
#313300000000
0!
0'
#313310000000
1!
b10 %
1'
b10 +
#313320000000
0!
0'
#313330000000
1!
b11 %
1'
b11 +
#313340000000
0!
0'
#313350000000
1!
b100 %
1'
b100 +
#313360000000
0!
0'
#313370000000
1!
b101 %
1'
b101 +
#313380000000
0!
0'
#313390000000
1!
b110 %
1'
b110 +
#313400000000
0!
0'
#313410000000
1!
b111 %
1'
b111 +
#313420000000
0!
0'
#313430000000
1!
0$
b1000 %
1'
0*
b1000 +
#313440000000
0!
0'
#313450000000
1!
b1001 %
1'
b1001 +
#313460000000
0!
0'
#313470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#313480000000
0!
0'
#313490000000
1!
1$
b1 %
1'
1*
b1 +
#313500000000
0!
0'
#313510000000
1!
b10 %
1'
b10 +
#313520000000
0!
0'
#313530000000
1!
b11 %
1'
b11 +
#313540000000
0!
0'
#313550000000
1!
b100 %
1'
b100 +
#313560000000
0!
0'
#313570000000
1!
b101 %
1'
b101 +
#313580000000
0!
0'
#313590000000
1!
0$
b110 %
1'
0*
b110 +
#313600000000
0!
0'
#313610000000
1!
b111 %
1'
b111 +
#313620000000
0!
0'
#313630000000
1!
b1000 %
1'
b1000 +
#313640000000
0!
0'
#313650000000
1!
b1001 %
1'
b1001 +
#313660000000
0!
0'
#313670000000
1!
b0 %
1'
b0 +
#313680000000
1"
1(
#313690000000
0!
0"
b100 &
0'
0(
b100 ,
#313700000000
1!
1$
b1 %
1'
1*
b1 +
#313710000000
0!
0'
#313720000000
1!
b10 %
1'
b10 +
#313730000000
0!
0'
#313740000000
1!
b11 %
1'
b11 +
#313750000000
0!
0'
#313760000000
1!
b100 %
1'
b100 +
#313770000000
0!
0'
#313780000000
1!
b101 %
1'
b101 +
#313790000000
0!
0'
#313800000000
1!
b110 %
1'
b110 +
#313810000000
0!
0'
#313820000000
1!
b111 %
1'
b111 +
#313830000000
0!
0'
#313840000000
1!
0$
b1000 %
1'
0*
b1000 +
#313850000000
0!
0'
#313860000000
1!
b1001 %
1'
b1001 +
#313870000000
0!
0'
#313880000000
1!
b0 %
1'
b0 +
#313890000000
0!
0'
#313900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#313910000000
0!
0'
#313920000000
1!
b10 %
1'
b10 +
#313930000000
0!
0'
#313940000000
1!
b11 %
1'
b11 +
#313950000000
0!
0'
#313960000000
1!
b100 %
1'
b100 +
#313970000000
0!
0'
#313980000000
1!
b101 %
1'
b101 +
#313990000000
0!
0'
#314000000000
1!
0$
b110 %
1'
0*
b110 +
#314010000000
0!
0'
#314020000000
1!
b111 %
1'
b111 +
#314030000000
0!
0'
#314040000000
1!
b1000 %
1'
b1000 +
#314050000000
0!
0'
#314060000000
1!
b1001 %
1'
b1001 +
#314070000000
0!
0'
#314080000000
1!
b0 %
1'
b0 +
#314090000000
0!
0'
#314100000000
1!
1$
b1 %
1'
1*
b1 +
#314110000000
1"
1(
#314120000000
0!
0"
b100 &
0'
0(
b100 ,
#314130000000
1!
b10 %
1'
b10 +
#314140000000
0!
0'
#314150000000
1!
b11 %
1'
b11 +
#314160000000
0!
0'
#314170000000
1!
b100 %
1'
b100 +
#314180000000
0!
0'
#314190000000
1!
b101 %
1'
b101 +
#314200000000
0!
0'
#314210000000
1!
b110 %
1'
b110 +
#314220000000
0!
0'
#314230000000
1!
b111 %
1'
b111 +
#314240000000
0!
0'
#314250000000
1!
0$
b1000 %
1'
0*
b1000 +
#314260000000
0!
0'
#314270000000
1!
b1001 %
1'
b1001 +
#314280000000
0!
0'
#314290000000
1!
b0 %
1'
b0 +
#314300000000
0!
0'
#314310000000
1!
1$
b1 %
1'
1*
b1 +
#314320000000
0!
0'
#314330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#314340000000
0!
0'
#314350000000
1!
b11 %
1'
b11 +
#314360000000
0!
0'
#314370000000
1!
b100 %
1'
b100 +
#314380000000
0!
0'
#314390000000
1!
b101 %
1'
b101 +
#314400000000
0!
0'
#314410000000
1!
0$
b110 %
1'
0*
b110 +
#314420000000
0!
0'
#314430000000
1!
b111 %
1'
b111 +
#314440000000
0!
0'
#314450000000
1!
b1000 %
1'
b1000 +
#314460000000
0!
0'
#314470000000
1!
b1001 %
1'
b1001 +
#314480000000
0!
0'
#314490000000
1!
b0 %
1'
b0 +
#314500000000
0!
0'
#314510000000
1!
1$
b1 %
1'
1*
b1 +
#314520000000
0!
0'
#314530000000
1!
b10 %
1'
b10 +
#314540000000
1"
1(
#314550000000
0!
0"
b100 &
0'
0(
b100 ,
#314560000000
1!
b11 %
1'
b11 +
#314570000000
0!
0'
#314580000000
1!
b100 %
1'
b100 +
#314590000000
0!
0'
#314600000000
1!
b101 %
1'
b101 +
#314610000000
0!
0'
#314620000000
1!
b110 %
1'
b110 +
#314630000000
0!
0'
#314640000000
1!
b111 %
1'
b111 +
#314650000000
0!
0'
#314660000000
1!
0$
b1000 %
1'
0*
b1000 +
#314670000000
0!
0'
#314680000000
1!
b1001 %
1'
b1001 +
#314690000000
0!
0'
#314700000000
1!
b0 %
1'
b0 +
#314710000000
0!
0'
#314720000000
1!
1$
b1 %
1'
1*
b1 +
#314730000000
0!
0'
#314740000000
1!
b10 %
1'
b10 +
#314750000000
0!
0'
#314760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#314770000000
0!
0'
#314780000000
1!
b100 %
1'
b100 +
#314790000000
0!
0'
#314800000000
1!
b101 %
1'
b101 +
#314810000000
0!
0'
#314820000000
1!
0$
b110 %
1'
0*
b110 +
#314830000000
0!
0'
#314840000000
1!
b111 %
1'
b111 +
#314850000000
0!
0'
#314860000000
1!
b1000 %
1'
b1000 +
#314870000000
0!
0'
#314880000000
1!
b1001 %
1'
b1001 +
#314890000000
0!
0'
#314900000000
1!
b0 %
1'
b0 +
#314910000000
0!
0'
#314920000000
1!
1$
b1 %
1'
1*
b1 +
#314930000000
0!
0'
#314940000000
1!
b10 %
1'
b10 +
#314950000000
0!
0'
#314960000000
1!
b11 %
1'
b11 +
#314970000000
1"
1(
#314980000000
0!
0"
b100 &
0'
0(
b100 ,
#314990000000
1!
b100 %
1'
b100 +
#315000000000
0!
0'
#315010000000
1!
b101 %
1'
b101 +
#315020000000
0!
0'
#315030000000
1!
b110 %
1'
b110 +
#315040000000
0!
0'
#315050000000
1!
b111 %
1'
b111 +
#315060000000
0!
0'
#315070000000
1!
0$
b1000 %
1'
0*
b1000 +
#315080000000
0!
0'
#315090000000
1!
b1001 %
1'
b1001 +
#315100000000
0!
0'
#315110000000
1!
b0 %
1'
b0 +
#315120000000
0!
0'
#315130000000
1!
1$
b1 %
1'
1*
b1 +
#315140000000
0!
0'
#315150000000
1!
b10 %
1'
b10 +
#315160000000
0!
0'
#315170000000
1!
b11 %
1'
b11 +
#315180000000
0!
0'
#315190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#315200000000
0!
0'
#315210000000
1!
b101 %
1'
b101 +
#315220000000
0!
0'
#315230000000
1!
0$
b110 %
1'
0*
b110 +
#315240000000
0!
0'
#315250000000
1!
b111 %
1'
b111 +
#315260000000
0!
0'
#315270000000
1!
b1000 %
1'
b1000 +
#315280000000
0!
0'
#315290000000
1!
b1001 %
1'
b1001 +
#315300000000
0!
0'
#315310000000
1!
b0 %
1'
b0 +
#315320000000
0!
0'
#315330000000
1!
1$
b1 %
1'
1*
b1 +
#315340000000
0!
0'
#315350000000
1!
b10 %
1'
b10 +
#315360000000
0!
0'
#315370000000
1!
b11 %
1'
b11 +
#315380000000
0!
0'
#315390000000
1!
b100 %
1'
b100 +
#315400000000
1"
1(
#315410000000
0!
0"
b100 &
0'
0(
b100 ,
#315420000000
1!
b101 %
1'
b101 +
#315430000000
0!
0'
#315440000000
1!
b110 %
1'
b110 +
#315450000000
0!
0'
#315460000000
1!
b111 %
1'
b111 +
#315470000000
0!
0'
#315480000000
1!
0$
b1000 %
1'
0*
b1000 +
#315490000000
0!
0'
#315500000000
1!
b1001 %
1'
b1001 +
#315510000000
0!
0'
#315520000000
1!
b0 %
1'
b0 +
#315530000000
0!
0'
#315540000000
1!
1$
b1 %
1'
1*
b1 +
#315550000000
0!
0'
#315560000000
1!
b10 %
1'
b10 +
#315570000000
0!
0'
#315580000000
1!
b11 %
1'
b11 +
#315590000000
0!
0'
#315600000000
1!
b100 %
1'
b100 +
#315610000000
0!
0'
#315620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#315630000000
0!
0'
#315640000000
1!
0$
b110 %
1'
0*
b110 +
#315650000000
0!
0'
#315660000000
1!
b111 %
1'
b111 +
#315670000000
0!
0'
#315680000000
1!
b1000 %
1'
b1000 +
#315690000000
0!
0'
#315700000000
1!
b1001 %
1'
b1001 +
#315710000000
0!
0'
#315720000000
1!
b0 %
1'
b0 +
#315730000000
0!
0'
#315740000000
1!
1$
b1 %
1'
1*
b1 +
#315750000000
0!
0'
#315760000000
1!
b10 %
1'
b10 +
#315770000000
0!
0'
#315780000000
1!
b11 %
1'
b11 +
#315790000000
0!
0'
#315800000000
1!
b100 %
1'
b100 +
#315810000000
0!
0'
#315820000000
1!
b101 %
1'
b101 +
#315830000000
1"
1(
#315840000000
0!
0"
b100 &
0'
0(
b100 ,
#315850000000
1!
b110 %
1'
b110 +
#315860000000
0!
0'
#315870000000
1!
b111 %
1'
b111 +
#315880000000
0!
0'
#315890000000
1!
0$
b1000 %
1'
0*
b1000 +
#315900000000
0!
0'
#315910000000
1!
b1001 %
1'
b1001 +
#315920000000
0!
0'
#315930000000
1!
b0 %
1'
b0 +
#315940000000
0!
0'
#315950000000
1!
1$
b1 %
1'
1*
b1 +
#315960000000
0!
0'
#315970000000
1!
b10 %
1'
b10 +
#315980000000
0!
0'
#315990000000
1!
b11 %
1'
b11 +
#316000000000
0!
0'
#316010000000
1!
b100 %
1'
b100 +
#316020000000
0!
0'
#316030000000
1!
b101 %
1'
b101 +
#316040000000
0!
0'
#316050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#316060000000
0!
0'
#316070000000
1!
b111 %
1'
b111 +
#316080000000
0!
0'
#316090000000
1!
b1000 %
1'
b1000 +
#316100000000
0!
0'
#316110000000
1!
b1001 %
1'
b1001 +
#316120000000
0!
0'
#316130000000
1!
b0 %
1'
b0 +
#316140000000
0!
0'
#316150000000
1!
1$
b1 %
1'
1*
b1 +
#316160000000
0!
0'
#316170000000
1!
b10 %
1'
b10 +
#316180000000
0!
0'
#316190000000
1!
b11 %
1'
b11 +
#316200000000
0!
0'
#316210000000
1!
b100 %
1'
b100 +
#316220000000
0!
0'
#316230000000
1!
b101 %
1'
b101 +
#316240000000
0!
0'
#316250000000
1!
0$
b110 %
1'
0*
b110 +
#316260000000
1"
1(
#316270000000
0!
0"
b100 &
0'
0(
b100 ,
#316280000000
1!
1$
b111 %
1'
1*
b111 +
#316290000000
0!
0'
#316300000000
1!
0$
b1000 %
1'
0*
b1000 +
#316310000000
0!
0'
#316320000000
1!
b1001 %
1'
b1001 +
#316330000000
0!
0'
#316340000000
1!
b0 %
1'
b0 +
#316350000000
0!
0'
#316360000000
1!
1$
b1 %
1'
1*
b1 +
#316370000000
0!
0'
#316380000000
1!
b10 %
1'
b10 +
#316390000000
0!
0'
#316400000000
1!
b11 %
1'
b11 +
#316410000000
0!
0'
#316420000000
1!
b100 %
1'
b100 +
#316430000000
0!
0'
#316440000000
1!
b101 %
1'
b101 +
#316450000000
0!
0'
#316460000000
1!
b110 %
1'
b110 +
#316470000000
0!
0'
#316480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#316490000000
0!
0'
#316500000000
1!
b1000 %
1'
b1000 +
#316510000000
0!
0'
#316520000000
1!
b1001 %
1'
b1001 +
#316530000000
0!
0'
#316540000000
1!
b0 %
1'
b0 +
#316550000000
0!
0'
#316560000000
1!
1$
b1 %
1'
1*
b1 +
#316570000000
0!
0'
#316580000000
1!
b10 %
1'
b10 +
#316590000000
0!
0'
#316600000000
1!
b11 %
1'
b11 +
#316610000000
0!
0'
#316620000000
1!
b100 %
1'
b100 +
#316630000000
0!
0'
#316640000000
1!
b101 %
1'
b101 +
#316650000000
0!
0'
#316660000000
1!
0$
b110 %
1'
0*
b110 +
#316670000000
0!
0'
#316680000000
1!
b111 %
1'
b111 +
#316690000000
1"
1(
#316700000000
0!
0"
b100 &
0'
0(
b100 ,
#316710000000
1!
b1000 %
1'
b1000 +
#316720000000
0!
0'
#316730000000
1!
b1001 %
1'
b1001 +
#316740000000
0!
0'
#316750000000
1!
b0 %
1'
b0 +
#316760000000
0!
0'
#316770000000
1!
1$
b1 %
1'
1*
b1 +
#316780000000
0!
0'
#316790000000
1!
b10 %
1'
b10 +
#316800000000
0!
0'
#316810000000
1!
b11 %
1'
b11 +
#316820000000
0!
0'
#316830000000
1!
b100 %
1'
b100 +
#316840000000
0!
0'
#316850000000
1!
b101 %
1'
b101 +
#316860000000
0!
0'
#316870000000
1!
b110 %
1'
b110 +
#316880000000
0!
0'
#316890000000
1!
b111 %
1'
b111 +
#316900000000
0!
0'
#316910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#316920000000
0!
0'
#316930000000
1!
b1001 %
1'
b1001 +
#316940000000
0!
0'
#316950000000
1!
b0 %
1'
b0 +
#316960000000
0!
0'
#316970000000
1!
1$
b1 %
1'
1*
b1 +
#316980000000
0!
0'
#316990000000
1!
b10 %
1'
b10 +
#317000000000
0!
0'
#317010000000
1!
b11 %
1'
b11 +
#317020000000
0!
0'
#317030000000
1!
b100 %
1'
b100 +
#317040000000
0!
0'
#317050000000
1!
b101 %
1'
b101 +
#317060000000
0!
0'
#317070000000
1!
0$
b110 %
1'
0*
b110 +
#317080000000
0!
0'
#317090000000
1!
b111 %
1'
b111 +
#317100000000
0!
0'
#317110000000
1!
b1000 %
1'
b1000 +
#317120000000
1"
1(
#317130000000
0!
0"
b100 &
0'
0(
b100 ,
#317140000000
1!
b1001 %
1'
b1001 +
#317150000000
0!
0'
#317160000000
1!
b0 %
1'
b0 +
#317170000000
0!
0'
#317180000000
1!
1$
b1 %
1'
1*
b1 +
#317190000000
0!
0'
#317200000000
1!
b10 %
1'
b10 +
#317210000000
0!
0'
#317220000000
1!
b11 %
1'
b11 +
#317230000000
0!
0'
#317240000000
1!
b100 %
1'
b100 +
#317250000000
0!
0'
#317260000000
1!
b101 %
1'
b101 +
#317270000000
0!
0'
#317280000000
1!
b110 %
1'
b110 +
#317290000000
0!
0'
#317300000000
1!
b111 %
1'
b111 +
#317310000000
0!
0'
#317320000000
1!
0$
b1000 %
1'
0*
b1000 +
#317330000000
0!
0'
#317340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#317350000000
0!
0'
#317360000000
1!
b0 %
1'
b0 +
#317370000000
0!
0'
#317380000000
1!
1$
b1 %
1'
1*
b1 +
#317390000000
0!
0'
#317400000000
1!
b10 %
1'
b10 +
#317410000000
0!
0'
#317420000000
1!
b11 %
1'
b11 +
#317430000000
0!
0'
#317440000000
1!
b100 %
1'
b100 +
#317450000000
0!
0'
#317460000000
1!
b101 %
1'
b101 +
#317470000000
0!
0'
#317480000000
1!
0$
b110 %
1'
0*
b110 +
#317490000000
0!
0'
#317500000000
1!
b111 %
1'
b111 +
#317510000000
0!
0'
#317520000000
1!
b1000 %
1'
b1000 +
#317530000000
0!
0'
#317540000000
1!
b1001 %
1'
b1001 +
#317550000000
1"
1(
#317560000000
0!
0"
b100 &
0'
0(
b100 ,
#317570000000
1!
b0 %
1'
b0 +
#317580000000
0!
0'
#317590000000
1!
1$
b1 %
1'
1*
b1 +
#317600000000
0!
0'
#317610000000
1!
b10 %
1'
b10 +
#317620000000
0!
0'
#317630000000
1!
b11 %
1'
b11 +
#317640000000
0!
0'
#317650000000
1!
b100 %
1'
b100 +
#317660000000
0!
0'
#317670000000
1!
b101 %
1'
b101 +
#317680000000
0!
0'
#317690000000
1!
b110 %
1'
b110 +
#317700000000
0!
0'
#317710000000
1!
b111 %
1'
b111 +
#317720000000
0!
0'
#317730000000
1!
0$
b1000 %
1'
0*
b1000 +
#317740000000
0!
0'
#317750000000
1!
b1001 %
1'
b1001 +
#317760000000
0!
0'
#317770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#317780000000
0!
0'
#317790000000
1!
1$
b1 %
1'
1*
b1 +
#317800000000
0!
0'
#317810000000
1!
b10 %
1'
b10 +
#317820000000
0!
0'
#317830000000
1!
b11 %
1'
b11 +
#317840000000
0!
0'
#317850000000
1!
b100 %
1'
b100 +
#317860000000
0!
0'
#317870000000
1!
b101 %
1'
b101 +
#317880000000
0!
0'
#317890000000
1!
0$
b110 %
1'
0*
b110 +
#317900000000
0!
0'
#317910000000
1!
b111 %
1'
b111 +
#317920000000
0!
0'
#317930000000
1!
b1000 %
1'
b1000 +
#317940000000
0!
0'
#317950000000
1!
b1001 %
1'
b1001 +
#317960000000
0!
0'
#317970000000
1!
b0 %
1'
b0 +
#317980000000
1"
1(
#317990000000
0!
0"
b100 &
0'
0(
b100 ,
#318000000000
1!
1$
b1 %
1'
1*
b1 +
#318010000000
0!
0'
#318020000000
1!
b10 %
1'
b10 +
#318030000000
0!
0'
#318040000000
1!
b11 %
1'
b11 +
#318050000000
0!
0'
#318060000000
1!
b100 %
1'
b100 +
#318070000000
0!
0'
#318080000000
1!
b101 %
1'
b101 +
#318090000000
0!
0'
#318100000000
1!
b110 %
1'
b110 +
#318110000000
0!
0'
#318120000000
1!
b111 %
1'
b111 +
#318130000000
0!
0'
#318140000000
1!
0$
b1000 %
1'
0*
b1000 +
#318150000000
0!
0'
#318160000000
1!
b1001 %
1'
b1001 +
#318170000000
0!
0'
#318180000000
1!
b0 %
1'
b0 +
#318190000000
0!
0'
#318200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#318210000000
0!
0'
#318220000000
1!
b10 %
1'
b10 +
#318230000000
0!
0'
#318240000000
1!
b11 %
1'
b11 +
#318250000000
0!
0'
#318260000000
1!
b100 %
1'
b100 +
#318270000000
0!
0'
#318280000000
1!
b101 %
1'
b101 +
#318290000000
0!
0'
#318300000000
1!
0$
b110 %
1'
0*
b110 +
#318310000000
0!
0'
#318320000000
1!
b111 %
1'
b111 +
#318330000000
0!
0'
#318340000000
1!
b1000 %
1'
b1000 +
#318350000000
0!
0'
#318360000000
1!
b1001 %
1'
b1001 +
#318370000000
0!
0'
#318380000000
1!
b0 %
1'
b0 +
#318390000000
0!
0'
#318400000000
1!
1$
b1 %
1'
1*
b1 +
#318410000000
1"
1(
#318420000000
0!
0"
b100 &
0'
0(
b100 ,
#318430000000
1!
b10 %
1'
b10 +
#318440000000
0!
0'
#318450000000
1!
b11 %
1'
b11 +
#318460000000
0!
0'
#318470000000
1!
b100 %
1'
b100 +
#318480000000
0!
0'
#318490000000
1!
b101 %
1'
b101 +
#318500000000
0!
0'
#318510000000
1!
b110 %
1'
b110 +
#318520000000
0!
0'
#318530000000
1!
b111 %
1'
b111 +
#318540000000
0!
0'
#318550000000
1!
0$
b1000 %
1'
0*
b1000 +
#318560000000
0!
0'
#318570000000
1!
b1001 %
1'
b1001 +
#318580000000
0!
0'
#318590000000
1!
b0 %
1'
b0 +
#318600000000
0!
0'
#318610000000
1!
1$
b1 %
1'
1*
b1 +
#318620000000
0!
0'
#318630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#318640000000
0!
0'
#318650000000
1!
b11 %
1'
b11 +
#318660000000
0!
0'
#318670000000
1!
b100 %
1'
b100 +
#318680000000
0!
0'
#318690000000
1!
b101 %
1'
b101 +
#318700000000
0!
0'
#318710000000
1!
0$
b110 %
1'
0*
b110 +
#318720000000
0!
0'
#318730000000
1!
b111 %
1'
b111 +
#318740000000
0!
0'
#318750000000
1!
b1000 %
1'
b1000 +
#318760000000
0!
0'
#318770000000
1!
b1001 %
1'
b1001 +
#318780000000
0!
0'
#318790000000
1!
b0 %
1'
b0 +
#318800000000
0!
0'
#318810000000
1!
1$
b1 %
1'
1*
b1 +
#318820000000
0!
0'
#318830000000
1!
b10 %
1'
b10 +
#318840000000
1"
1(
#318850000000
0!
0"
b100 &
0'
0(
b100 ,
#318860000000
1!
b11 %
1'
b11 +
#318870000000
0!
0'
#318880000000
1!
b100 %
1'
b100 +
#318890000000
0!
0'
#318900000000
1!
b101 %
1'
b101 +
#318910000000
0!
0'
#318920000000
1!
b110 %
1'
b110 +
#318930000000
0!
0'
#318940000000
1!
b111 %
1'
b111 +
#318950000000
0!
0'
#318960000000
1!
0$
b1000 %
1'
0*
b1000 +
#318970000000
0!
0'
#318980000000
1!
b1001 %
1'
b1001 +
#318990000000
0!
0'
#319000000000
1!
b0 %
1'
b0 +
#319010000000
0!
0'
#319020000000
1!
1$
b1 %
1'
1*
b1 +
#319030000000
0!
0'
#319040000000
1!
b10 %
1'
b10 +
#319050000000
0!
0'
#319060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#319070000000
0!
0'
#319080000000
1!
b100 %
1'
b100 +
#319090000000
0!
0'
#319100000000
1!
b101 %
1'
b101 +
#319110000000
0!
0'
#319120000000
1!
0$
b110 %
1'
0*
b110 +
#319130000000
0!
0'
#319140000000
1!
b111 %
1'
b111 +
#319150000000
0!
0'
#319160000000
1!
b1000 %
1'
b1000 +
#319170000000
0!
0'
#319180000000
1!
b1001 %
1'
b1001 +
#319190000000
0!
0'
#319200000000
1!
b0 %
1'
b0 +
#319210000000
0!
0'
#319220000000
1!
1$
b1 %
1'
1*
b1 +
#319230000000
0!
0'
#319240000000
1!
b10 %
1'
b10 +
#319250000000
0!
0'
#319260000000
1!
b11 %
1'
b11 +
#319270000000
1"
1(
#319280000000
0!
0"
b100 &
0'
0(
b100 ,
#319290000000
1!
b100 %
1'
b100 +
#319300000000
0!
0'
#319310000000
1!
b101 %
1'
b101 +
#319320000000
0!
0'
#319330000000
1!
b110 %
1'
b110 +
#319340000000
0!
0'
#319350000000
1!
b111 %
1'
b111 +
#319360000000
0!
0'
#319370000000
1!
0$
b1000 %
1'
0*
b1000 +
#319380000000
0!
0'
#319390000000
1!
b1001 %
1'
b1001 +
#319400000000
0!
0'
#319410000000
1!
b0 %
1'
b0 +
#319420000000
0!
0'
#319430000000
1!
1$
b1 %
1'
1*
b1 +
#319440000000
0!
0'
#319450000000
1!
b10 %
1'
b10 +
#319460000000
0!
0'
#319470000000
1!
b11 %
1'
b11 +
#319480000000
0!
0'
#319490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#319500000000
0!
0'
#319510000000
1!
b101 %
1'
b101 +
#319520000000
0!
0'
#319530000000
1!
0$
b110 %
1'
0*
b110 +
#319540000000
0!
0'
#319550000000
1!
b111 %
1'
b111 +
#319560000000
0!
0'
#319570000000
1!
b1000 %
1'
b1000 +
#319580000000
0!
0'
#319590000000
1!
b1001 %
1'
b1001 +
#319600000000
0!
0'
#319610000000
1!
b0 %
1'
b0 +
#319620000000
0!
0'
#319630000000
1!
1$
b1 %
1'
1*
b1 +
#319640000000
0!
0'
#319650000000
1!
b10 %
1'
b10 +
#319660000000
0!
0'
#319670000000
1!
b11 %
1'
b11 +
#319680000000
0!
0'
#319690000000
1!
b100 %
1'
b100 +
#319700000000
1"
1(
#319710000000
0!
0"
b100 &
0'
0(
b100 ,
#319720000000
1!
b101 %
1'
b101 +
#319730000000
0!
0'
#319740000000
1!
b110 %
1'
b110 +
#319750000000
0!
0'
#319760000000
1!
b111 %
1'
b111 +
#319770000000
0!
0'
#319780000000
1!
0$
b1000 %
1'
0*
b1000 +
#319790000000
0!
0'
#319800000000
1!
b1001 %
1'
b1001 +
#319810000000
0!
0'
#319820000000
1!
b0 %
1'
b0 +
#319830000000
0!
0'
#319840000000
1!
1$
b1 %
1'
1*
b1 +
#319850000000
0!
0'
#319860000000
1!
b10 %
1'
b10 +
#319870000000
0!
0'
#319880000000
1!
b11 %
1'
b11 +
#319890000000
0!
0'
#319900000000
1!
b100 %
1'
b100 +
#319910000000
0!
0'
#319920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#319930000000
0!
0'
#319940000000
1!
0$
b110 %
1'
0*
b110 +
#319950000000
0!
0'
#319960000000
1!
b111 %
1'
b111 +
#319970000000
0!
0'
#319980000000
1!
b1000 %
1'
b1000 +
#319990000000
0!
0'
#320000000000
1!
b1001 %
1'
b1001 +
#320010000000
0!
0'
#320020000000
1!
b0 %
1'
b0 +
#320030000000
0!
0'
#320040000000
1!
1$
b1 %
1'
1*
b1 +
#320050000000
0!
0'
#320060000000
1!
b10 %
1'
b10 +
#320070000000
0!
0'
#320080000000
1!
b11 %
1'
b11 +
#320090000000
0!
0'
#320100000000
1!
b100 %
1'
b100 +
#320110000000
0!
0'
#320120000000
1!
b101 %
1'
b101 +
#320130000000
1"
1(
#320140000000
0!
0"
b100 &
0'
0(
b100 ,
#320150000000
1!
b110 %
1'
b110 +
#320160000000
0!
0'
#320170000000
1!
b111 %
1'
b111 +
#320180000000
0!
0'
#320190000000
1!
0$
b1000 %
1'
0*
b1000 +
#320200000000
0!
0'
#320210000000
1!
b1001 %
1'
b1001 +
#320220000000
0!
0'
#320230000000
1!
b0 %
1'
b0 +
#320240000000
0!
0'
#320250000000
1!
1$
b1 %
1'
1*
b1 +
#320260000000
0!
0'
#320270000000
1!
b10 %
1'
b10 +
#320280000000
0!
0'
#320290000000
1!
b11 %
1'
b11 +
#320300000000
0!
0'
#320310000000
1!
b100 %
1'
b100 +
#320320000000
0!
0'
#320330000000
1!
b101 %
1'
b101 +
#320340000000
0!
0'
#320350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#320360000000
0!
0'
#320370000000
1!
b111 %
1'
b111 +
#320380000000
0!
0'
#320390000000
1!
b1000 %
1'
b1000 +
#320400000000
0!
0'
#320410000000
1!
b1001 %
1'
b1001 +
#320420000000
0!
0'
#320430000000
1!
b0 %
1'
b0 +
#320440000000
0!
0'
#320450000000
1!
1$
b1 %
1'
1*
b1 +
#320460000000
0!
0'
#320470000000
1!
b10 %
1'
b10 +
#320480000000
0!
0'
#320490000000
1!
b11 %
1'
b11 +
#320500000000
0!
0'
#320510000000
1!
b100 %
1'
b100 +
#320520000000
0!
0'
#320530000000
1!
b101 %
1'
b101 +
#320540000000
0!
0'
#320550000000
1!
0$
b110 %
1'
0*
b110 +
#320560000000
1"
1(
#320570000000
0!
0"
b100 &
0'
0(
b100 ,
#320580000000
1!
1$
b111 %
1'
1*
b111 +
#320590000000
0!
0'
#320600000000
1!
0$
b1000 %
1'
0*
b1000 +
#320610000000
0!
0'
#320620000000
1!
b1001 %
1'
b1001 +
#320630000000
0!
0'
#320640000000
1!
b0 %
1'
b0 +
#320650000000
0!
0'
#320660000000
1!
1$
b1 %
1'
1*
b1 +
#320670000000
0!
0'
#320680000000
1!
b10 %
1'
b10 +
#320690000000
0!
0'
#320700000000
1!
b11 %
1'
b11 +
#320710000000
0!
0'
#320720000000
1!
b100 %
1'
b100 +
#320730000000
0!
0'
#320740000000
1!
b101 %
1'
b101 +
#320750000000
0!
0'
#320760000000
1!
b110 %
1'
b110 +
#320770000000
0!
0'
#320780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#320790000000
0!
0'
#320800000000
1!
b1000 %
1'
b1000 +
#320810000000
0!
0'
#320820000000
1!
b1001 %
1'
b1001 +
#320830000000
0!
0'
#320840000000
1!
b0 %
1'
b0 +
#320850000000
0!
0'
#320860000000
1!
1$
b1 %
1'
1*
b1 +
#320870000000
0!
0'
#320880000000
1!
b10 %
1'
b10 +
#320890000000
0!
0'
#320900000000
1!
b11 %
1'
b11 +
#320910000000
0!
0'
#320920000000
1!
b100 %
1'
b100 +
#320930000000
0!
0'
#320940000000
1!
b101 %
1'
b101 +
#320950000000
0!
0'
#320960000000
1!
0$
b110 %
1'
0*
b110 +
#320970000000
0!
0'
#320980000000
1!
b111 %
1'
b111 +
#320990000000
1"
1(
#321000000000
0!
0"
b100 &
0'
0(
b100 ,
#321010000000
1!
b1000 %
1'
b1000 +
#321020000000
0!
0'
#321030000000
1!
b1001 %
1'
b1001 +
#321040000000
0!
0'
#321050000000
1!
b0 %
1'
b0 +
#321060000000
0!
0'
#321070000000
1!
1$
b1 %
1'
1*
b1 +
#321080000000
0!
0'
#321090000000
1!
b10 %
1'
b10 +
#321100000000
0!
0'
#321110000000
1!
b11 %
1'
b11 +
#321120000000
0!
0'
#321130000000
1!
b100 %
1'
b100 +
#321140000000
0!
0'
#321150000000
1!
b101 %
1'
b101 +
#321160000000
0!
0'
#321170000000
1!
b110 %
1'
b110 +
#321180000000
0!
0'
#321190000000
1!
b111 %
1'
b111 +
#321200000000
0!
0'
#321210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#321220000000
0!
0'
#321230000000
1!
b1001 %
1'
b1001 +
#321240000000
0!
0'
#321250000000
1!
b0 %
1'
b0 +
#321260000000
0!
0'
#321270000000
1!
1$
b1 %
1'
1*
b1 +
#321280000000
0!
0'
#321290000000
1!
b10 %
1'
b10 +
#321300000000
0!
0'
#321310000000
1!
b11 %
1'
b11 +
#321320000000
0!
0'
#321330000000
1!
b100 %
1'
b100 +
#321340000000
0!
0'
#321350000000
1!
b101 %
1'
b101 +
#321360000000
0!
0'
#321370000000
1!
0$
b110 %
1'
0*
b110 +
#321380000000
0!
0'
#321390000000
1!
b111 %
1'
b111 +
#321400000000
0!
0'
#321410000000
1!
b1000 %
1'
b1000 +
#321420000000
1"
1(
#321430000000
0!
0"
b100 &
0'
0(
b100 ,
#321440000000
1!
b1001 %
1'
b1001 +
#321450000000
0!
0'
#321460000000
1!
b0 %
1'
b0 +
#321470000000
0!
0'
#321480000000
1!
1$
b1 %
1'
1*
b1 +
#321490000000
0!
0'
#321500000000
1!
b10 %
1'
b10 +
#321510000000
0!
0'
#321520000000
1!
b11 %
1'
b11 +
#321530000000
0!
0'
#321540000000
1!
b100 %
1'
b100 +
#321550000000
0!
0'
#321560000000
1!
b101 %
1'
b101 +
#321570000000
0!
0'
#321580000000
1!
b110 %
1'
b110 +
#321590000000
0!
0'
#321600000000
1!
b111 %
1'
b111 +
#321610000000
0!
0'
#321620000000
1!
0$
b1000 %
1'
0*
b1000 +
#321630000000
0!
0'
#321640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#321650000000
0!
0'
#321660000000
1!
b0 %
1'
b0 +
#321670000000
0!
0'
#321680000000
1!
1$
b1 %
1'
1*
b1 +
#321690000000
0!
0'
#321700000000
1!
b10 %
1'
b10 +
#321710000000
0!
0'
#321720000000
1!
b11 %
1'
b11 +
#321730000000
0!
0'
#321740000000
1!
b100 %
1'
b100 +
#321750000000
0!
0'
#321760000000
1!
b101 %
1'
b101 +
#321770000000
0!
0'
#321780000000
1!
0$
b110 %
1'
0*
b110 +
#321790000000
0!
0'
#321800000000
1!
b111 %
1'
b111 +
#321810000000
0!
0'
#321820000000
1!
b1000 %
1'
b1000 +
#321830000000
0!
0'
#321840000000
1!
b1001 %
1'
b1001 +
#321850000000
1"
1(
#321860000000
0!
0"
b100 &
0'
0(
b100 ,
#321870000000
1!
b0 %
1'
b0 +
#321880000000
0!
0'
#321890000000
1!
1$
b1 %
1'
1*
b1 +
#321900000000
0!
0'
#321910000000
1!
b10 %
1'
b10 +
#321920000000
0!
0'
#321930000000
1!
b11 %
1'
b11 +
#321940000000
0!
0'
#321950000000
1!
b100 %
1'
b100 +
#321960000000
0!
0'
#321970000000
1!
b101 %
1'
b101 +
#321980000000
0!
0'
#321990000000
1!
b110 %
1'
b110 +
#322000000000
0!
0'
#322010000000
1!
b111 %
1'
b111 +
#322020000000
0!
0'
#322030000000
1!
0$
b1000 %
1'
0*
b1000 +
#322040000000
0!
0'
#322050000000
1!
b1001 %
1'
b1001 +
#322060000000
0!
0'
#322070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#322080000000
0!
0'
#322090000000
1!
1$
b1 %
1'
1*
b1 +
#322100000000
0!
0'
#322110000000
1!
b10 %
1'
b10 +
#322120000000
0!
0'
#322130000000
1!
b11 %
1'
b11 +
#322140000000
0!
0'
#322150000000
1!
b100 %
1'
b100 +
#322160000000
0!
0'
#322170000000
1!
b101 %
1'
b101 +
#322180000000
0!
0'
#322190000000
1!
0$
b110 %
1'
0*
b110 +
#322200000000
0!
0'
#322210000000
1!
b111 %
1'
b111 +
#322220000000
0!
0'
#322230000000
1!
b1000 %
1'
b1000 +
#322240000000
0!
0'
#322250000000
1!
b1001 %
1'
b1001 +
#322260000000
0!
0'
#322270000000
1!
b0 %
1'
b0 +
#322280000000
1"
1(
#322290000000
0!
0"
b100 &
0'
0(
b100 ,
#322300000000
1!
1$
b1 %
1'
1*
b1 +
#322310000000
0!
0'
#322320000000
1!
b10 %
1'
b10 +
#322330000000
0!
0'
#322340000000
1!
b11 %
1'
b11 +
#322350000000
0!
0'
#322360000000
1!
b100 %
1'
b100 +
#322370000000
0!
0'
#322380000000
1!
b101 %
1'
b101 +
#322390000000
0!
0'
#322400000000
1!
b110 %
1'
b110 +
#322410000000
0!
0'
#322420000000
1!
b111 %
1'
b111 +
#322430000000
0!
0'
#322440000000
1!
0$
b1000 %
1'
0*
b1000 +
#322450000000
0!
0'
#322460000000
1!
b1001 %
1'
b1001 +
#322470000000
0!
0'
#322480000000
1!
b0 %
1'
b0 +
#322490000000
0!
0'
#322500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#322510000000
0!
0'
#322520000000
1!
b10 %
1'
b10 +
#322530000000
0!
0'
#322540000000
1!
b11 %
1'
b11 +
#322550000000
0!
0'
#322560000000
1!
b100 %
1'
b100 +
#322570000000
0!
0'
#322580000000
1!
b101 %
1'
b101 +
#322590000000
0!
0'
#322600000000
1!
0$
b110 %
1'
0*
b110 +
#322610000000
0!
0'
#322620000000
1!
b111 %
1'
b111 +
#322630000000
0!
0'
#322640000000
1!
b1000 %
1'
b1000 +
#322650000000
0!
0'
#322660000000
1!
b1001 %
1'
b1001 +
#322670000000
0!
0'
#322680000000
1!
b0 %
1'
b0 +
#322690000000
0!
0'
#322700000000
1!
1$
b1 %
1'
1*
b1 +
#322710000000
1"
1(
#322720000000
0!
0"
b100 &
0'
0(
b100 ,
#322730000000
1!
b10 %
1'
b10 +
#322740000000
0!
0'
#322750000000
1!
b11 %
1'
b11 +
#322760000000
0!
0'
#322770000000
1!
b100 %
1'
b100 +
#322780000000
0!
0'
#322790000000
1!
b101 %
1'
b101 +
#322800000000
0!
0'
#322810000000
1!
b110 %
1'
b110 +
#322820000000
0!
0'
#322830000000
1!
b111 %
1'
b111 +
#322840000000
0!
0'
#322850000000
1!
0$
b1000 %
1'
0*
b1000 +
#322860000000
0!
0'
#322870000000
1!
b1001 %
1'
b1001 +
#322880000000
0!
0'
#322890000000
1!
b0 %
1'
b0 +
#322900000000
0!
0'
#322910000000
1!
1$
b1 %
1'
1*
b1 +
#322920000000
0!
0'
#322930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#322940000000
0!
0'
#322950000000
1!
b11 %
1'
b11 +
#322960000000
0!
0'
#322970000000
1!
b100 %
1'
b100 +
#322980000000
0!
0'
#322990000000
1!
b101 %
1'
b101 +
#323000000000
0!
0'
#323010000000
1!
0$
b110 %
1'
0*
b110 +
#323020000000
0!
0'
#323030000000
1!
b111 %
1'
b111 +
#323040000000
0!
0'
#323050000000
1!
b1000 %
1'
b1000 +
#323060000000
0!
0'
#323070000000
1!
b1001 %
1'
b1001 +
#323080000000
0!
0'
#323090000000
1!
b0 %
1'
b0 +
#323100000000
0!
0'
#323110000000
1!
1$
b1 %
1'
1*
b1 +
#323120000000
0!
0'
#323130000000
1!
b10 %
1'
b10 +
#323140000000
1"
1(
#323150000000
0!
0"
b100 &
0'
0(
b100 ,
#323160000000
1!
b11 %
1'
b11 +
#323170000000
0!
0'
#323180000000
1!
b100 %
1'
b100 +
#323190000000
0!
0'
#323200000000
1!
b101 %
1'
b101 +
#323210000000
0!
0'
#323220000000
1!
b110 %
1'
b110 +
#323230000000
0!
0'
#323240000000
1!
b111 %
1'
b111 +
#323250000000
0!
0'
#323260000000
1!
0$
b1000 %
1'
0*
b1000 +
#323270000000
0!
0'
#323280000000
1!
b1001 %
1'
b1001 +
#323290000000
0!
0'
#323300000000
1!
b0 %
1'
b0 +
#323310000000
0!
0'
#323320000000
1!
1$
b1 %
1'
1*
b1 +
#323330000000
0!
0'
#323340000000
1!
b10 %
1'
b10 +
#323350000000
0!
0'
#323360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#323370000000
0!
0'
#323380000000
1!
b100 %
1'
b100 +
#323390000000
0!
0'
#323400000000
1!
b101 %
1'
b101 +
#323410000000
0!
0'
#323420000000
1!
0$
b110 %
1'
0*
b110 +
#323430000000
0!
0'
#323440000000
1!
b111 %
1'
b111 +
#323450000000
0!
0'
#323460000000
1!
b1000 %
1'
b1000 +
#323470000000
0!
0'
#323480000000
1!
b1001 %
1'
b1001 +
#323490000000
0!
0'
#323500000000
1!
b0 %
1'
b0 +
#323510000000
0!
0'
#323520000000
1!
1$
b1 %
1'
1*
b1 +
#323530000000
0!
0'
#323540000000
1!
b10 %
1'
b10 +
#323550000000
0!
0'
#323560000000
1!
b11 %
1'
b11 +
#323570000000
1"
1(
#323580000000
0!
0"
b100 &
0'
0(
b100 ,
#323590000000
1!
b100 %
1'
b100 +
#323600000000
0!
0'
#323610000000
1!
b101 %
1'
b101 +
#323620000000
0!
0'
#323630000000
1!
b110 %
1'
b110 +
#323640000000
0!
0'
#323650000000
1!
b111 %
1'
b111 +
#323660000000
0!
0'
#323670000000
1!
0$
b1000 %
1'
0*
b1000 +
#323680000000
0!
0'
#323690000000
1!
b1001 %
1'
b1001 +
#323700000000
0!
0'
#323710000000
1!
b0 %
1'
b0 +
#323720000000
0!
0'
#323730000000
1!
1$
b1 %
1'
1*
b1 +
#323740000000
0!
0'
#323750000000
1!
b10 %
1'
b10 +
#323760000000
0!
0'
#323770000000
1!
b11 %
1'
b11 +
#323780000000
0!
0'
#323790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#323800000000
0!
0'
#323810000000
1!
b101 %
1'
b101 +
#323820000000
0!
0'
#323830000000
1!
0$
b110 %
1'
0*
b110 +
#323840000000
0!
0'
#323850000000
1!
b111 %
1'
b111 +
#323860000000
0!
0'
#323870000000
1!
b1000 %
1'
b1000 +
#323880000000
0!
0'
#323890000000
1!
b1001 %
1'
b1001 +
#323900000000
0!
0'
#323910000000
1!
b0 %
1'
b0 +
#323920000000
0!
0'
#323930000000
1!
1$
b1 %
1'
1*
b1 +
#323940000000
0!
0'
#323950000000
1!
b10 %
1'
b10 +
#323960000000
0!
0'
#323970000000
1!
b11 %
1'
b11 +
#323980000000
0!
0'
#323990000000
1!
b100 %
1'
b100 +
#324000000000
1"
1(
#324010000000
0!
0"
b100 &
0'
0(
b100 ,
#324020000000
1!
b101 %
1'
b101 +
#324030000000
0!
0'
#324040000000
1!
b110 %
1'
b110 +
#324050000000
0!
0'
#324060000000
1!
b111 %
1'
b111 +
#324070000000
0!
0'
#324080000000
1!
0$
b1000 %
1'
0*
b1000 +
#324090000000
0!
0'
#324100000000
1!
b1001 %
1'
b1001 +
#324110000000
0!
0'
#324120000000
1!
b0 %
1'
b0 +
#324130000000
0!
0'
#324140000000
1!
1$
b1 %
1'
1*
b1 +
#324150000000
0!
0'
#324160000000
1!
b10 %
1'
b10 +
#324170000000
0!
0'
#324180000000
1!
b11 %
1'
b11 +
#324190000000
0!
0'
#324200000000
1!
b100 %
1'
b100 +
#324210000000
0!
0'
#324220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#324230000000
0!
0'
#324240000000
1!
0$
b110 %
1'
0*
b110 +
#324250000000
0!
0'
#324260000000
1!
b111 %
1'
b111 +
#324270000000
0!
0'
#324280000000
1!
b1000 %
1'
b1000 +
#324290000000
0!
0'
#324300000000
1!
b1001 %
1'
b1001 +
#324310000000
0!
0'
#324320000000
1!
b0 %
1'
b0 +
#324330000000
0!
0'
#324340000000
1!
1$
b1 %
1'
1*
b1 +
#324350000000
0!
0'
#324360000000
1!
b10 %
1'
b10 +
#324370000000
0!
0'
#324380000000
1!
b11 %
1'
b11 +
#324390000000
0!
0'
#324400000000
1!
b100 %
1'
b100 +
#324410000000
0!
0'
#324420000000
1!
b101 %
1'
b101 +
#324430000000
1"
1(
#324440000000
0!
0"
b100 &
0'
0(
b100 ,
#324450000000
1!
b110 %
1'
b110 +
#324460000000
0!
0'
#324470000000
1!
b111 %
1'
b111 +
#324480000000
0!
0'
#324490000000
1!
0$
b1000 %
1'
0*
b1000 +
#324500000000
0!
0'
#324510000000
1!
b1001 %
1'
b1001 +
#324520000000
0!
0'
#324530000000
1!
b0 %
1'
b0 +
#324540000000
0!
0'
#324550000000
1!
1$
b1 %
1'
1*
b1 +
#324560000000
0!
0'
#324570000000
1!
b10 %
1'
b10 +
#324580000000
0!
0'
#324590000000
1!
b11 %
1'
b11 +
#324600000000
0!
0'
#324610000000
1!
b100 %
1'
b100 +
#324620000000
0!
0'
#324630000000
1!
b101 %
1'
b101 +
#324640000000
0!
0'
#324650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#324660000000
0!
0'
#324670000000
1!
b111 %
1'
b111 +
#324680000000
0!
0'
#324690000000
1!
b1000 %
1'
b1000 +
#324700000000
0!
0'
#324710000000
1!
b1001 %
1'
b1001 +
#324720000000
0!
0'
#324730000000
1!
b0 %
1'
b0 +
#324740000000
0!
0'
#324750000000
1!
1$
b1 %
1'
1*
b1 +
#324760000000
0!
0'
#324770000000
1!
b10 %
1'
b10 +
#324780000000
0!
0'
#324790000000
1!
b11 %
1'
b11 +
#324800000000
0!
0'
#324810000000
1!
b100 %
1'
b100 +
#324820000000
0!
0'
#324830000000
1!
b101 %
1'
b101 +
#324840000000
0!
0'
#324850000000
1!
0$
b110 %
1'
0*
b110 +
#324860000000
1"
1(
#324870000000
0!
0"
b100 &
0'
0(
b100 ,
#324880000000
1!
1$
b111 %
1'
1*
b111 +
#324890000000
0!
0'
#324900000000
1!
0$
b1000 %
1'
0*
b1000 +
#324910000000
0!
0'
#324920000000
1!
b1001 %
1'
b1001 +
#324930000000
0!
0'
#324940000000
1!
b0 %
1'
b0 +
#324950000000
0!
0'
#324960000000
1!
1$
b1 %
1'
1*
b1 +
#324970000000
0!
0'
#324980000000
1!
b10 %
1'
b10 +
#324990000000
0!
0'
#325000000000
1!
b11 %
1'
b11 +
#325010000000
0!
0'
#325020000000
1!
b100 %
1'
b100 +
#325030000000
0!
0'
#325040000000
1!
b101 %
1'
b101 +
#325050000000
0!
0'
#325060000000
1!
b110 %
1'
b110 +
#325070000000
0!
0'
#325080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#325090000000
0!
0'
#325100000000
1!
b1000 %
1'
b1000 +
#325110000000
0!
0'
#325120000000
1!
b1001 %
1'
b1001 +
#325130000000
0!
0'
#325140000000
1!
b0 %
1'
b0 +
#325150000000
0!
0'
#325160000000
1!
1$
b1 %
1'
1*
b1 +
#325170000000
0!
0'
#325180000000
1!
b10 %
1'
b10 +
#325190000000
0!
0'
#325200000000
1!
b11 %
1'
b11 +
#325210000000
0!
0'
#325220000000
1!
b100 %
1'
b100 +
#325230000000
0!
0'
#325240000000
1!
b101 %
1'
b101 +
#325250000000
0!
0'
#325260000000
1!
0$
b110 %
1'
0*
b110 +
#325270000000
0!
0'
#325280000000
1!
b111 %
1'
b111 +
#325290000000
1"
1(
#325300000000
0!
0"
b100 &
0'
0(
b100 ,
#325310000000
1!
b1000 %
1'
b1000 +
#325320000000
0!
0'
#325330000000
1!
b1001 %
1'
b1001 +
#325340000000
0!
0'
#325350000000
1!
b0 %
1'
b0 +
#325360000000
0!
0'
#325370000000
1!
1$
b1 %
1'
1*
b1 +
#325380000000
0!
0'
#325390000000
1!
b10 %
1'
b10 +
#325400000000
0!
0'
#325410000000
1!
b11 %
1'
b11 +
#325420000000
0!
0'
#325430000000
1!
b100 %
1'
b100 +
#325440000000
0!
0'
#325450000000
1!
b101 %
1'
b101 +
#325460000000
0!
0'
#325470000000
1!
b110 %
1'
b110 +
#325480000000
0!
0'
#325490000000
1!
b111 %
1'
b111 +
#325500000000
0!
0'
#325510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#325520000000
0!
0'
#325530000000
1!
b1001 %
1'
b1001 +
#325540000000
0!
0'
#325550000000
1!
b0 %
1'
b0 +
#325560000000
0!
0'
#325570000000
1!
1$
b1 %
1'
1*
b1 +
#325580000000
0!
0'
#325590000000
1!
b10 %
1'
b10 +
#325600000000
0!
0'
#325610000000
1!
b11 %
1'
b11 +
#325620000000
0!
0'
#325630000000
1!
b100 %
1'
b100 +
#325640000000
0!
0'
#325650000000
1!
b101 %
1'
b101 +
#325660000000
0!
0'
#325670000000
1!
0$
b110 %
1'
0*
b110 +
#325680000000
0!
0'
#325690000000
1!
b111 %
1'
b111 +
#325700000000
0!
0'
#325710000000
1!
b1000 %
1'
b1000 +
#325720000000
1"
1(
#325730000000
0!
0"
b100 &
0'
0(
b100 ,
#325740000000
1!
b1001 %
1'
b1001 +
#325750000000
0!
0'
#325760000000
1!
b0 %
1'
b0 +
#325770000000
0!
0'
#325780000000
1!
1$
b1 %
1'
1*
b1 +
#325790000000
0!
0'
#325800000000
1!
b10 %
1'
b10 +
#325810000000
0!
0'
#325820000000
1!
b11 %
1'
b11 +
#325830000000
0!
0'
#325840000000
1!
b100 %
1'
b100 +
#325850000000
0!
0'
#325860000000
1!
b101 %
1'
b101 +
#325870000000
0!
0'
#325880000000
1!
b110 %
1'
b110 +
#325890000000
0!
0'
#325900000000
1!
b111 %
1'
b111 +
#325910000000
0!
0'
#325920000000
1!
0$
b1000 %
1'
0*
b1000 +
#325930000000
0!
0'
#325940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#325950000000
0!
0'
#325960000000
1!
b0 %
1'
b0 +
#325970000000
0!
0'
#325980000000
1!
1$
b1 %
1'
1*
b1 +
#325990000000
0!
0'
#326000000000
1!
b10 %
1'
b10 +
#326010000000
0!
0'
#326020000000
1!
b11 %
1'
b11 +
#326030000000
0!
0'
#326040000000
1!
b100 %
1'
b100 +
#326050000000
0!
0'
#326060000000
1!
b101 %
1'
b101 +
#326070000000
0!
0'
#326080000000
1!
0$
b110 %
1'
0*
b110 +
#326090000000
0!
0'
#326100000000
1!
b111 %
1'
b111 +
#326110000000
0!
0'
#326120000000
1!
b1000 %
1'
b1000 +
#326130000000
0!
0'
#326140000000
1!
b1001 %
1'
b1001 +
#326150000000
1"
1(
#326160000000
0!
0"
b100 &
0'
0(
b100 ,
#326170000000
1!
b0 %
1'
b0 +
#326180000000
0!
0'
#326190000000
1!
1$
b1 %
1'
1*
b1 +
#326200000000
0!
0'
#326210000000
1!
b10 %
1'
b10 +
#326220000000
0!
0'
#326230000000
1!
b11 %
1'
b11 +
#326240000000
0!
0'
#326250000000
1!
b100 %
1'
b100 +
#326260000000
0!
0'
#326270000000
1!
b101 %
1'
b101 +
#326280000000
0!
0'
#326290000000
1!
b110 %
1'
b110 +
#326300000000
0!
0'
#326310000000
1!
b111 %
1'
b111 +
#326320000000
0!
0'
#326330000000
1!
0$
b1000 %
1'
0*
b1000 +
#326340000000
0!
0'
#326350000000
1!
b1001 %
1'
b1001 +
#326360000000
0!
0'
#326370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#326380000000
0!
0'
#326390000000
1!
1$
b1 %
1'
1*
b1 +
#326400000000
0!
0'
#326410000000
1!
b10 %
1'
b10 +
#326420000000
0!
0'
#326430000000
1!
b11 %
1'
b11 +
#326440000000
0!
0'
#326450000000
1!
b100 %
1'
b100 +
#326460000000
0!
0'
#326470000000
1!
b101 %
1'
b101 +
#326480000000
0!
0'
#326490000000
1!
0$
b110 %
1'
0*
b110 +
#326500000000
0!
0'
#326510000000
1!
b111 %
1'
b111 +
#326520000000
0!
0'
#326530000000
1!
b1000 %
1'
b1000 +
#326540000000
0!
0'
#326550000000
1!
b1001 %
1'
b1001 +
#326560000000
0!
0'
#326570000000
1!
b0 %
1'
b0 +
#326580000000
1"
1(
#326590000000
0!
0"
b100 &
0'
0(
b100 ,
#326600000000
1!
1$
b1 %
1'
1*
b1 +
#326610000000
0!
0'
#326620000000
1!
b10 %
1'
b10 +
#326630000000
0!
0'
#326640000000
1!
b11 %
1'
b11 +
#326650000000
0!
0'
#326660000000
1!
b100 %
1'
b100 +
#326670000000
0!
0'
#326680000000
1!
b101 %
1'
b101 +
#326690000000
0!
0'
#326700000000
1!
b110 %
1'
b110 +
#326710000000
0!
0'
#326720000000
1!
b111 %
1'
b111 +
#326730000000
0!
0'
#326740000000
1!
0$
b1000 %
1'
0*
b1000 +
#326750000000
0!
0'
#326760000000
1!
b1001 %
1'
b1001 +
#326770000000
0!
0'
#326780000000
1!
b0 %
1'
b0 +
#326790000000
0!
0'
#326800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#326810000000
0!
0'
#326820000000
1!
b10 %
1'
b10 +
#326830000000
0!
0'
#326840000000
1!
b11 %
1'
b11 +
#326850000000
0!
0'
#326860000000
1!
b100 %
1'
b100 +
#326870000000
0!
0'
#326880000000
1!
b101 %
1'
b101 +
#326890000000
0!
0'
#326900000000
1!
0$
b110 %
1'
0*
b110 +
#326910000000
0!
0'
#326920000000
1!
b111 %
1'
b111 +
#326930000000
0!
0'
#326940000000
1!
b1000 %
1'
b1000 +
#326950000000
0!
0'
#326960000000
1!
b1001 %
1'
b1001 +
#326970000000
0!
0'
#326980000000
1!
b0 %
1'
b0 +
#326990000000
0!
0'
#327000000000
1!
1$
b1 %
1'
1*
b1 +
#327010000000
1"
1(
#327020000000
0!
0"
b100 &
0'
0(
b100 ,
#327030000000
1!
b10 %
1'
b10 +
#327040000000
0!
0'
#327050000000
1!
b11 %
1'
b11 +
#327060000000
0!
0'
#327070000000
1!
b100 %
1'
b100 +
#327080000000
0!
0'
#327090000000
1!
b101 %
1'
b101 +
#327100000000
0!
0'
#327110000000
1!
b110 %
1'
b110 +
#327120000000
0!
0'
#327130000000
1!
b111 %
1'
b111 +
#327140000000
0!
0'
#327150000000
1!
0$
b1000 %
1'
0*
b1000 +
#327160000000
0!
0'
#327170000000
1!
b1001 %
1'
b1001 +
#327180000000
0!
0'
#327190000000
1!
b0 %
1'
b0 +
#327200000000
0!
0'
#327210000000
1!
1$
b1 %
1'
1*
b1 +
#327220000000
0!
0'
#327230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#327240000000
0!
0'
#327250000000
1!
b11 %
1'
b11 +
#327260000000
0!
0'
#327270000000
1!
b100 %
1'
b100 +
#327280000000
0!
0'
#327290000000
1!
b101 %
1'
b101 +
#327300000000
0!
0'
#327310000000
1!
0$
b110 %
1'
0*
b110 +
#327320000000
0!
0'
#327330000000
1!
b111 %
1'
b111 +
#327340000000
0!
0'
#327350000000
1!
b1000 %
1'
b1000 +
#327360000000
0!
0'
#327370000000
1!
b1001 %
1'
b1001 +
#327380000000
0!
0'
#327390000000
1!
b0 %
1'
b0 +
#327400000000
0!
0'
#327410000000
1!
1$
b1 %
1'
1*
b1 +
#327420000000
0!
0'
#327430000000
1!
b10 %
1'
b10 +
#327440000000
1"
1(
#327450000000
0!
0"
b100 &
0'
0(
b100 ,
#327460000000
1!
b11 %
1'
b11 +
#327470000000
0!
0'
#327480000000
1!
b100 %
1'
b100 +
#327490000000
0!
0'
#327500000000
1!
b101 %
1'
b101 +
#327510000000
0!
0'
#327520000000
1!
b110 %
1'
b110 +
#327530000000
0!
0'
#327540000000
1!
b111 %
1'
b111 +
#327550000000
0!
0'
#327560000000
1!
0$
b1000 %
1'
0*
b1000 +
#327570000000
0!
0'
#327580000000
1!
b1001 %
1'
b1001 +
#327590000000
0!
0'
#327600000000
1!
b0 %
1'
b0 +
#327610000000
0!
0'
#327620000000
1!
1$
b1 %
1'
1*
b1 +
#327630000000
0!
0'
#327640000000
1!
b10 %
1'
b10 +
#327650000000
0!
0'
#327660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#327670000000
0!
0'
#327680000000
1!
b100 %
1'
b100 +
#327690000000
0!
0'
#327700000000
1!
b101 %
1'
b101 +
#327710000000
0!
0'
#327720000000
1!
0$
b110 %
1'
0*
b110 +
#327730000000
0!
0'
#327740000000
1!
b111 %
1'
b111 +
#327750000000
0!
0'
#327760000000
1!
b1000 %
1'
b1000 +
#327770000000
0!
0'
#327780000000
1!
b1001 %
1'
b1001 +
#327790000000
0!
0'
#327800000000
1!
b0 %
1'
b0 +
#327810000000
0!
0'
#327820000000
1!
1$
b1 %
1'
1*
b1 +
#327830000000
0!
0'
#327840000000
1!
b10 %
1'
b10 +
#327850000000
0!
0'
#327860000000
1!
b11 %
1'
b11 +
#327870000000
1"
1(
#327880000000
0!
0"
b100 &
0'
0(
b100 ,
#327890000000
1!
b100 %
1'
b100 +
#327900000000
0!
0'
#327910000000
1!
b101 %
1'
b101 +
#327920000000
0!
0'
#327930000000
1!
b110 %
1'
b110 +
#327940000000
0!
0'
#327950000000
1!
b111 %
1'
b111 +
#327960000000
0!
0'
#327970000000
1!
0$
b1000 %
1'
0*
b1000 +
#327980000000
0!
0'
#327990000000
1!
b1001 %
1'
b1001 +
#328000000000
0!
0'
#328010000000
1!
b0 %
1'
b0 +
#328020000000
0!
0'
#328030000000
1!
1$
b1 %
1'
1*
b1 +
#328040000000
0!
0'
#328050000000
1!
b10 %
1'
b10 +
#328060000000
0!
0'
#328070000000
1!
b11 %
1'
b11 +
#328080000000
0!
0'
#328090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#328100000000
0!
0'
#328110000000
1!
b101 %
1'
b101 +
#328120000000
0!
0'
#328130000000
1!
0$
b110 %
1'
0*
b110 +
#328140000000
0!
0'
#328150000000
1!
b111 %
1'
b111 +
#328160000000
0!
0'
#328170000000
1!
b1000 %
1'
b1000 +
#328180000000
0!
0'
#328190000000
1!
b1001 %
1'
b1001 +
#328200000000
0!
0'
#328210000000
1!
b0 %
1'
b0 +
#328220000000
0!
0'
#328230000000
1!
1$
b1 %
1'
1*
b1 +
#328240000000
0!
0'
#328250000000
1!
b10 %
1'
b10 +
#328260000000
0!
0'
#328270000000
1!
b11 %
1'
b11 +
#328280000000
0!
0'
#328290000000
1!
b100 %
1'
b100 +
#328300000000
1"
1(
#328310000000
0!
0"
b100 &
0'
0(
b100 ,
#328320000000
1!
b101 %
1'
b101 +
#328330000000
0!
0'
#328340000000
1!
b110 %
1'
b110 +
#328350000000
0!
0'
#328360000000
1!
b111 %
1'
b111 +
#328370000000
0!
0'
#328380000000
1!
0$
b1000 %
1'
0*
b1000 +
#328390000000
0!
0'
#328400000000
1!
b1001 %
1'
b1001 +
#328410000000
0!
0'
#328420000000
1!
b0 %
1'
b0 +
#328430000000
0!
0'
#328440000000
1!
1$
b1 %
1'
1*
b1 +
#328450000000
0!
0'
#328460000000
1!
b10 %
1'
b10 +
#328470000000
0!
0'
#328480000000
1!
b11 %
1'
b11 +
#328490000000
0!
0'
#328500000000
1!
b100 %
1'
b100 +
#328510000000
0!
0'
#328520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#328530000000
0!
0'
#328540000000
1!
0$
b110 %
1'
0*
b110 +
#328550000000
0!
0'
#328560000000
1!
b111 %
1'
b111 +
#328570000000
0!
0'
#328580000000
1!
b1000 %
1'
b1000 +
#328590000000
0!
0'
#328600000000
1!
b1001 %
1'
b1001 +
#328610000000
0!
0'
#328620000000
1!
b0 %
1'
b0 +
#328630000000
0!
0'
#328640000000
1!
1$
b1 %
1'
1*
b1 +
#328650000000
0!
0'
#328660000000
1!
b10 %
1'
b10 +
#328670000000
0!
0'
#328680000000
1!
b11 %
1'
b11 +
#328690000000
0!
0'
#328700000000
1!
b100 %
1'
b100 +
#328710000000
0!
0'
#328720000000
1!
b101 %
1'
b101 +
#328730000000
1"
1(
#328740000000
0!
0"
b100 &
0'
0(
b100 ,
#328750000000
1!
b110 %
1'
b110 +
#328760000000
0!
0'
#328770000000
1!
b111 %
1'
b111 +
#328780000000
0!
0'
#328790000000
1!
0$
b1000 %
1'
0*
b1000 +
#328800000000
0!
0'
#328810000000
1!
b1001 %
1'
b1001 +
#328820000000
0!
0'
#328830000000
1!
b0 %
1'
b0 +
#328840000000
0!
0'
#328850000000
1!
1$
b1 %
1'
1*
b1 +
#328860000000
0!
0'
#328870000000
1!
b10 %
1'
b10 +
#328880000000
0!
0'
#328890000000
1!
b11 %
1'
b11 +
#328900000000
0!
0'
#328910000000
1!
b100 %
1'
b100 +
#328920000000
0!
0'
#328930000000
1!
b101 %
1'
b101 +
#328940000000
0!
0'
#328950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#328960000000
0!
0'
#328970000000
1!
b111 %
1'
b111 +
#328980000000
0!
0'
#328990000000
1!
b1000 %
1'
b1000 +
#329000000000
0!
0'
#329010000000
1!
b1001 %
1'
b1001 +
#329020000000
0!
0'
#329030000000
1!
b0 %
1'
b0 +
#329040000000
0!
0'
#329050000000
1!
1$
b1 %
1'
1*
b1 +
#329060000000
0!
0'
#329070000000
1!
b10 %
1'
b10 +
#329080000000
0!
0'
#329090000000
1!
b11 %
1'
b11 +
#329100000000
0!
0'
#329110000000
1!
b100 %
1'
b100 +
#329120000000
0!
0'
#329130000000
1!
b101 %
1'
b101 +
#329140000000
0!
0'
#329150000000
1!
0$
b110 %
1'
0*
b110 +
#329160000000
1"
1(
#329170000000
0!
0"
b100 &
0'
0(
b100 ,
#329180000000
1!
1$
b111 %
1'
1*
b111 +
#329190000000
0!
0'
#329200000000
1!
0$
b1000 %
1'
0*
b1000 +
#329210000000
0!
0'
#329220000000
1!
b1001 %
1'
b1001 +
#329230000000
0!
0'
#329240000000
1!
b0 %
1'
b0 +
#329250000000
0!
0'
#329260000000
1!
1$
b1 %
1'
1*
b1 +
#329270000000
0!
0'
#329280000000
1!
b10 %
1'
b10 +
#329290000000
0!
0'
#329300000000
1!
b11 %
1'
b11 +
#329310000000
0!
0'
#329320000000
1!
b100 %
1'
b100 +
#329330000000
0!
0'
#329340000000
1!
b101 %
1'
b101 +
#329350000000
0!
0'
#329360000000
1!
b110 %
1'
b110 +
#329370000000
0!
0'
#329380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#329390000000
0!
0'
#329400000000
1!
b1000 %
1'
b1000 +
#329410000000
0!
0'
#329420000000
1!
b1001 %
1'
b1001 +
#329430000000
0!
0'
#329440000000
1!
b0 %
1'
b0 +
#329450000000
0!
0'
#329460000000
1!
1$
b1 %
1'
1*
b1 +
#329470000000
0!
0'
#329480000000
1!
b10 %
1'
b10 +
#329490000000
0!
0'
#329500000000
1!
b11 %
1'
b11 +
#329510000000
0!
0'
#329520000000
1!
b100 %
1'
b100 +
#329530000000
0!
0'
#329540000000
1!
b101 %
1'
b101 +
#329550000000
0!
0'
#329560000000
1!
0$
b110 %
1'
0*
b110 +
#329570000000
0!
0'
#329580000000
1!
b111 %
1'
b111 +
#329590000000
1"
1(
#329600000000
0!
0"
b100 &
0'
0(
b100 ,
#329610000000
1!
b1000 %
1'
b1000 +
#329620000000
0!
0'
#329630000000
1!
b1001 %
1'
b1001 +
#329640000000
0!
0'
#329650000000
1!
b0 %
1'
b0 +
#329660000000
0!
0'
#329670000000
1!
1$
b1 %
1'
1*
b1 +
#329680000000
0!
0'
#329690000000
1!
b10 %
1'
b10 +
#329700000000
0!
0'
#329710000000
1!
b11 %
1'
b11 +
#329720000000
0!
0'
#329730000000
1!
b100 %
1'
b100 +
#329740000000
0!
0'
#329750000000
1!
b101 %
1'
b101 +
#329760000000
0!
0'
#329770000000
1!
b110 %
1'
b110 +
#329780000000
0!
0'
#329790000000
1!
b111 %
1'
b111 +
#329800000000
0!
0'
#329810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#329820000000
0!
0'
#329830000000
1!
b1001 %
1'
b1001 +
#329840000000
0!
0'
#329850000000
1!
b0 %
1'
b0 +
#329860000000
0!
0'
#329870000000
1!
1$
b1 %
1'
1*
b1 +
#329880000000
0!
0'
#329890000000
1!
b10 %
1'
b10 +
#329900000000
0!
0'
#329910000000
1!
b11 %
1'
b11 +
#329920000000
0!
0'
#329930000000
1!
b100 %
1'
b100 +
#329940000000
0!
0'
#329950000000
1!
b101 %
1'
b101 +
#329960000000
0!
0'
#329970000000
1!
0$
b110 %
1'
0*
b110 +
#329980000000
0!
0'
#329990000000
1!
b111 %
1'
b111 +
#330000000000
0!
0'
#330010000000
1!
b1000 %
1'
b1000 +
#330020000000
1"
1(
#330030000000
0!
0"
b100 &
0'
0(
b100 ,
#330040000000
1!
b1001 %
1'
b1001 +
#330050000000
0!
0'
#330060000000
1!
b0 %
1'
b0 +
#330070000000
0!
0'
#330080000000
1!
1$
b1 %
1'
1*
b1 +
#330090000000
0!
0'
#330100000000
1!
b10 %
1'
b10 +
#330110000000
0!
0'
#330120000000
1!
b11 %
1'
b11 +
#330130000000
0!
0'
#330140000000
1!
b100 %
1'
b100 +
#330150000000
0!
0'
#330160000000
1!
b101 %
1'
b101 +
#330170000000
0!
0'
#330180000000
1!
b110 %
1'
b110 +
#330190000000
0!
0'
#330200000000
1!
b111 %
1'
b111 +
#330210000000
0!
0'
#330220000000
1!
0$
b1000 %
1'
0*
b1000 +
#330230000000
0!
0'
#330240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#330250000000
0!
0'
#330260000000
1!
b0 %
1'
b0 +
#330270000000
0!
0'
#330280000000
1!
1$
b1 %
1'
1*
b1 +
#330290000000
0!
0'
#330300000000
1!
b10 %
1'
b10 +
#330310000000
0!
0'
#330320000000
1!
b11 %
1'
b11 +
#330330000000
0!
0'
#330340000000
1!
b100 %
1'
b100 +
#330350000000
0!
0'
#330360000000
1!
b101 %
1'
b101 +
#330370000000
0!
0'
#330380000000
1!
0$
b110 %
1'
0*
b110 +
#330390000000
0!
0'
#330400000000
1!
b111 %
1'
b111 +
#330410000000
0!
0'
#330420000000
1!
b1000 %
1'
b1000 +
#330430000000
0!
0'
#330440000000
1!
b1001 %
1'
b1001 +
#330450000000
1"
1(
#330460000000
0!
0"
b100 &
0'
0(
b100 ,
#330470000000
1!
b0 %
1'
b0 +
#330480000000
0!
0'
#330490000000
1!
1$
b1 %
1'
1*
b1 +
#330500000000
0!
0'
#330510000000
1!
b10 %
1'
b10 +
#330520000000
0!
0'
#330530000000
1!
b11 %
1'
b11 +
#330540000000
0!
0'
#330550000000
1!
b100 %
1'
b100 +
#330560000000
0!
0'
#330570000000
1!
b101 %
1'
b101 +
#330580000000
0!
0'
#330590000000
1!
b110 %
1'
b110 +
#330600000000
0!
0'
#330610000000
1!
b111 %
1'
b111 +
#330620000000
0!
0'
#330630000000
1!
0$
b1000 %
1'
0*
b1000 +
#330640000000
0!
0'
#330650000000
1!
b1001 %
1'
b1001 +
#330660000000
0!
0'
#330670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#330680000000
0!
0'
#330690000000
1!
1$
b1 %
1'
1*
b1 +
#330700000000
0!
0'
#330710000000
1!
b10 %
1'
b10 +
#330720000000
0!
0'
#330730000000
1!
b11 %
1'
b11 +
#330740000000
0!
0'
#330750000000
1!
b100 %
1'
b100 +
#330760000000
0!
0'
#330770000000
1!
b101 %
1'
b101 +
#330780000000
0!
0'
#330790000000
1!
0$
b110 %
1'
0*
b110 +
#330800000000
0!
0'
#330810000000
1!
b111 %
1'
b111 +
#330820000000
0!
0'
#330830000000
1!
b1000 %
1'
b1000 +
#330840000000
0!
0'
#330850000000
1!
b1001 %
1'
b1001 +
#330860000000
0!
0'
#330870000000
1!
b0 %
1'
b0 +
#330880000000
1"
1(
#330890000000
0!
0"
b100 &
0'
0(
b100 ,
#330900000000
1!
1$
b1 %
1'
1*
b1 +
#330910000000
0!
0'
#330920000000
1!
b10 %
1'
b10 +
#330930000000
0!
0'
#330940000000
1!
b11 %
1'
b11 +
#330950000000
0!
0'
#330960000000
1!
b100 %
1'
b100 +
#330970000000
0!
0'
#330980000000
1!
b101 %
1'
b101 +
#330990000000
0!
0'
#331000000000
1!
b110 %
1'
b110 +
#331010000000
0!
0'
#331020000000
1!
b111 %
1'
b111 +
#331030000000
0!
0'
#331040000000
1!
0$
b1000 %
1'
0*
b1000 +
#331050000000
0!
0'
#331060000000
1!
b1001 %
1'
b1001 +
#331070000000
0!
0'
#331080000000
1!
b0 %
1'
b0 +
#331090000000
0!
0'
#331100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#331110000000
0!
0'
#331120000000
1!
b10 %
1'
b10 +
#331130000000
0!
0'
#331140000000
1!
b11 %
1'
b11 +
#331150000000
0!
0'
#331160000000
1!
b100 %
1'
b100 +
#331170000000
0!
0'
#331180000000
1!
b101 %
1'
b101 +
#331190000000
0!
0'
#331200000000
1!
0$
b110 %
1'
0*
b110 +
#331210000000
0!
0'
#331220000000
1!
b111 %
1'
b111 +
#331230000000
0!
0'
#331240000000
1!
b1000 %
1'
b1000 +
#331250000000
0!
0'
#331260000000
1!
b1001 %
1'
b1001 +
#331270000000
0!
0'
#331280000000
1!
b0 %
1'
b0 +
#331290000000
0!
0'
#331300000000
1!
1$
b1 %
1'
1*
b1 +
#331310000000
1"
1(
#331320000000
0!
0"
b100 &
0'
0(
b100 ,
#331330000000
1!
b10 %
1'
b10 +
#331340000000
0!
0'
#331350000000
1!
b11 %
1'
b11 +
#331360000000
0!
0'
#331370000000
1!
b100 %
1'
b100 +
#331380000000
0!
0'
#331390000000
1!
b101 %
1'
b101 +
#331400000000
0!
0'
#331410000000
1!
b110 %
1'
b110 +
#331420000000
0!
0'
#331430000000
1!
b111 %
1'
b111 +
#331440000000
0!
0'
#331450000000
1!
0$
b1000 %
1'
0*
b1000 +
#331460000000
0!
0'
#331470000000
1!
b1001 %
1'
b1001 +
#331480000000
0!
0'
#331490000000
1!
b0 %
1'
b0 +
#331500000000
0!
0'
#331510000000
1!
1$
b1 %
1'
1*
b1 +
#331520000000
0!
0'
#331530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#331540000000
0!
0'
#331550000000
1!
b11 %
1'
b11 +
#331560000000
0!
0'
#331570000000
1!
b100 %
1'
b100 +
#331580000000
0!
0'
#331590000000
1!
b101 %
1'
b101 +
#331600000000
0!
0'
#331610000000
1!
0$
b110 %
1'
0*
b110 +
#331620000000
0!
0'
#331630000000
1!
b111 %
1'
b111 +
#331640000000
0!
0'
#331650000000
1!
b1000 %
1'
b1000 +
#331660000000
0!
0'
#331670000000
1!
b1001 %
1'
b1001 +
#331680000000
0!
0'
#331690000000
1!
b0 %
1'
b0 +
#331700000000
0!
0'
#331710000000
1!
1$
b1 %
1'
1*
b1 +
#331720000000
0!
0'
#331730000000
1!
b10 %
1'
b10 +
#331740000000
1"
1(
#331750000000
0!
0"
b100 &
0'
0(
b100 ,
#331760000000
1!
b11 %
1'
b11 +
#331770000000
0!
0'
#331780000000
1!
b100 %
1'
b100 +
#331790000000
0!
0'
#331800000000
1!
b101 %
1'
b101 +
#331810000000
0!
0'
#331820000000
1!
b110 %
1'
b110 +
#331830000000
0!
0'
#331840000000
1!
b111 %
1'
b111 +
#331850000000
0!
0'
#331860000000
1!
0$
b1000 %
1'
0*
b1000 +
#331870000000
0!
0'
#331880000000
1!
b1001 %
1'
b1001 +
#331890000000
0!
0'
#331900000000
1!
b0 %
1'
b0 +
#331910000000
0!
0'
#331920000000
1!
1$
b1 %
1'
1*
b1 +
#331930000000
0!
0'
#331940000000
1!
b10 %
1'
b10 +
#331950000000
0!
0'
#331960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#331970000000
0!
0'
#331980000000
1!
b100 %
1'
b100 +
#331990000000
0!
0'
#332000000000
1!
b101 %
1'
b101 +
#332010000000
0!
0'
#332020000000
1!
0$
b110 %
1'
0*
b110 +
#332030000000
0!
0'
#332040000000
1!
b111 %
1'
b111 +
#332050000000
0!
0'
#332060000000
1!
b1000 %
1'
b1000 +
#332070000000
0!
0'
#332080000000
1!
b1001 %
1'
b1001 +
#332090000000
0!
0'
#332100000000
1!
b0 %
1'
b0 +
#332110000000
0!
0'
#332120000000
1!
1$
b1 %
1'
1*
b1 +
#332130000000
0!
0'
#332140000000
1!
b10 %
1'
b10 +
#332150000000
0!
0'
#332160000000
1!
b11 %
1'
b11 +
#332170000000
1"
1(
#332180000000
0!
0"
b100 &
0'
0(
b100 ,
#332190000000
1!
b100 %
1'
b100 +
#332200000000
0!
0'
#332210000000
1!
b101 %
1'
b101 +
#332220000000
0!
0'
#332230000000
1!
b110 %
1'
b110 +
#332240000000
0!
0'
#332250000000
1!
b111 %
1'
b111 +
#332260000000
0!
0'
#332270000000
1!
0$
b1000 %
1'
0*
b1000 +
#332280000000
0!
0'
#332290000000
1!
b1001 %
1'
b1001 +
#332300000000
0!
0'
#332310000000
1!
b0 %
1'
b0 +
#332320000000
0!
0'
#332330000000
1!
1$
b1 %
1'
1*
b1 +
#332340000000
0!
0'
#332350000000
1!
b10 %
1'
b10 +
#332360000000
0!
0'
#332370000000
1!
b11 %
1'
b11 +
#332380000000
0!
0'
#332390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#332400000000
0!
0'
#332410000000
1!
b101 %
1'
b101 +
#332420000000
0!
0'
#332430000000
1!
0$
b110 %
1'
0*
b110 +
#332440000000
0!
0'
#332450000000
1!
b111 %
1'
b111 +
#332460000000
0!
0'
#332470000000
1!
b1000 %
1'
b1000 +
#332480000000
0!
0'
#332490000000
1!
b1001 %
1'
b1001 +
#332500000000
0!
0'
#332510000000
1!
b0 %
1'
b0 +
#332520000000
0!
0'
#332530000000
1!
1$
b1 %
1'
1*
b1 +
#332540000000
0!
0'
#332550000000
1!
b10 %
1'
b10 +
#332560000000
0!
0'
#332570000000
1!
b11 %
1'
b11 +
#332580000000
0!
0'
#332590000000
1!
b100 %
1'
b100 +
#332600000000
1"
1(
#332610000000
0!
0"
b100 &
0'
0(
b100 ,
#332620000000
1!
b101 %
1'
b101 +
#332630000000
0!
0'
#332640000000
1!
b110 %
1'
b110 +
#332650000000
0!
0'
#332660000000
1!
b111 %
1'
b111 +
#332670000000
0!
0'
#332680000000
1!
0$
b1000 %
1'
0*
b1000 +
#332690000000
0!
0'
#332700000000
1!
b1001 %
1'
b1001 +
#332710000000
0!
0'
#332720000000
1!
b0 %
1'
b0 +
#332730000000
0!
0'
#332740000000
1!
1$
b1 %
1'
1*
b1 +
#332750000000
0!
0'
#332760000000
1!
b10 %
1'
b10 +
#332770000000
0!
0'
#332780000000
1!
b11 %
1'
b11 +
#332790000000
0!
0'
#332800000000
1!
b100 %
1'
b100 +
#332810000000
0!
0'
#332820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#332830000000
0!
0'
#332840000000
1!
0$
b110 %
1'
0*
b110 +
#332850000000
0!
0'
#332860000000
1!
b111 %
1'
b111 +
#332870000000
0!
0'
#332880000000
1!
b1000 %
1'
b1000 +
#332890000000
0!
0'
#332900000000
1!
b1001 %
1'
b1001 +
#332910000000
0!
0'
#332920000000
1!
b0 %
1'
b0 +
#332930000000
0!
0'
#332940000000
1!
1$
b1 %
1'
1*
b1 +
#332950000000
0!
0'
#332960000000
1!
b10 %
1'
b10 +
#332970000000
0!
0'
#332980000000
1!
b11 %
1'
b11 +
#332990000000
0!
0'
#333000000000
1!
b100 %
1'
b100 +
#333010000000
0!
0'
#333020000000
1!
b101 %
1'
b101 +
#333030000000
1"
1(
#333040000000
0!
0"
b100 &
0'
0(
b100 ,
#333050000000
1!
b110 %
1'
b110 +
#333060000000
0!
0'
#333070000000
1!
b111 %
1'
b111 +
#333080000000
0!
0'
#333090000000
1!
0$
b1000 %
1'
0*
b1000 +
#333100000000
0!
0'
#333110000000
1!
b1001 %
1'
b1001 +
#333120000000
0!
0'
#333130000000
1!
b0 %
1'
b0 +
#333140000000
0!
0'
#333150000000
1!
1$
b1 %
1'
1*
b1 +
#333160000000
0!
0'
#333170000000
1!
b10 %
1'
b10 +
#333180000000
0!
0'
#333190000000
1!
b11 %
1'
b11 +
#333200000000
0!
0'
#333210000000
1!
b100 %
1'
b100 +
#333220000000
0!
0'
#333230000000
1!
b101 %
1'
b101 +
#333240000000
0!
0'
#333250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#333260000000
0!
0'
#333270000000
1!
b111 %
1'
b111 +
#333280000000
0!
0'
#333290000000
1!
b1000 %
1'
b1000 +
#333300000000
0!
0'
#333310000000
1!
b1001 %
1'
b1001 +
#333320000000
0!
0'
#333330000000
1!
b0 %
1'
b0 +
#333340000000
0!
0'
#333350000000
1!
1$
b1 %
1'
1*
b1 +
#333360000000
0!
0'
#333370000000
1!
b10 %
1'
b10 +
#333380000000
0!
0'
#333390000000
1!
b11 %
1'
b11 +
#333400000000
0!
0'
#333410000000
1!
b100 %
1'
b100 +
#333420000000
0!
0'
#333430000000
1!
b101 %
1'
b101 +
#333440000000
0!
0'
#333450000000
1!
0$
b110 %
1'
0*
b110 +
#333460000000
1"
1(
#333470000000
0!
0"
b100 &
0'
0(
b100 ,
#333480000000
1!
1$
b111 %
1'
1*
b111 +
#333490000000
0!
0'
#333500000000
1!
0$
b1000 %
1'
0*
b1000 +
#333510000000
0!
0'
#333520000000
1!
b1001 %
1'
b1001 +
#333530000000
0!
0'
#333540000000
1!
b0 %
1'
b0 +
#333550000000
0!
0'
#333560000000
1!
1$
b1 %
1'
1*
b1 +
#333570000000
0!
0'
#333580000000
1!
b10 %
1'
b10 +
#333590000000
0!
0'
#333600000000
1!
b11 %
1'
b11 +
#333610000000
0!
0'
#333620000000
1!
b100 %
1'
b100 +
#333630000000
0!
0'
#333640000000
1!
b101 %
1'
b101 +
#333650000000
0!
0'
#333660000000
1!
b110 %
1'
b110 +
#333670000000
0!
0'
#333680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#333690000000
0!
0'
#333700000000
1!
b1000 %
1'
b1000 +
#333710000000
0!
0'
#333720000000
1!
b1001 %
1'
b1001 +
#333730000000
0!
0'
#333740000000
1!
b0 %
1'
b0 +
#333750000000
0!
0'
#333760000000
1!
1$
b1 %
1'
1*
b1 +
#333770000000
0!
0'
#333780000000
1!
b10 %
1'
b10 +
#333790000000
0!
0'
#333800000000
1!
b11 %
1'
b11 +
#333810000000
0!
0'
#333820000000
1!
b100 %
1'
b100 +
#333830000000
0!
0'
#333840000000
1!
b101 %
1'
b101 +
#333850000000
0!
0'
#333860000000
1!
0$
b110 %
1'
0*
b110 +
#333870000000
0!
0'
#333880000000
1!
b111 %
1'
b111 +
#333890000000
1"
1(
#333900000000
0!
0"
b100 &
0'
0(
b100 ,
#333910000000
1!
b1000 %
1'
b1000 +
#333920000000
0!
0'
#333930000000
1!
b1001 %
1'
b1001 +
#333940000000
0!
0'
#333950000000
1!
b0 %
1'
b0 +
#333960000000
0!
0'
#333970000000
1!
1$
b1 %
1'
1*
b1 +
#333980000000
0!
0'
#333990000000
1!
b10 %
1'
b10 +
#334000000000
0!
0'
#334010000000
1!
b11 %
1'
b11 +
#334020000000
0!
0'
#334030000000
1!
b100 %
1'
b100 +
#334040000000
0!
0'
#334050000000
1!
b101 %
1'
b101 +
#334060000000
0!
0'
#334070000000
1!
b110 %
1'
b110 +
#334080000000
0!
0'
#334090000000
1!
b111 %
1'
b111 +
#334100000000
0!
0'
#334110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#334120000000
0!
0'
#334130000000
1!
b1001 %
1'
b1001 +
#334140000000
0!
0'
#334150000000
1!
b0 %
1'
b0 +
#334160000000
0!
0'
#334170000000
1!
1$
b1 %
1'
1*
b1 +
#334180000000
0!
0'
#334190000000
1!
b10 %
1'
b10 +
#334200000000
0!
0'
#334210000000
1!
b11 %
1'
b11 +
#334220000000
0!
0'
#334230000000
1!
b100 %
1'
b100 +
#334240000000
0!
0'
#334250000000
1!
b101 %
1'
b101 +
#334260000000
0!
0'
#334270000000
1!
0$
b110 %
1'
0*
b110 +
#334280000000
0!
0'
#334290000000
1!
b111 %
1'
b111 +
#334300000000
0!
0'
#334310000000
1!
b1000 %
1'
b1000 +
#334320000000
1"
1(
#334330000000
0!
0"
b100 &
0'
0(
b100 ,
#334340000000
1!
b1001 %
1'
b1001 +
#334350000000
0!
0'
#334360000000
1!
b0 %
1'
b0 +
#334370000000
0!
0'
#334380000000
1!
1$
b1 %
1'
1*
b1 +
#334390000000
0!
0'
#334400000000
1!
b10 %
1'
b10 +
#334410000000
0!
0'
#334420000000
1!
b11 %
1'
b11 +
#334430000000
0!
0'
#334440000000
1!
b100 %
1'
b100 +
#334450000000
0!
0'
#334460000000
1!
b101 %
1'
b101 +
#334470000000
0!
0'
#334480000000
1!
b110 %
1'
b110 +
#334490000000
0!
0'
#334500000000
1!
b111 %
1'
b111 +
#334510000000
0!
0'
#334520000000
1!
0$
b1000 %
1'
0*
b1000 +
#334530000000
0!
0'
#334540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#334550000000
0!
0'
#334560000000
1!
b0 %
1'
b0 +
#334570000000
0!
0'
#334580000000
1!
1$
b1 %
1'
1*
b1 +
#334590000000
0!
0'
#334600000000
1!
b10 %
1'
b10 +
#334610000000
0!
0'
#334620000000
1!
b11 %
1'
b11 +
#334630000000
0!
0'
#334640000000
1!
b100 %
1'
b100 +
#334650000000
0!
0'
#334660000000
1!
b101 %
1'
b101 +
#334670000000
0!
0'
#334680000000
1!
0$
b110 %
1'
0*
b110 +
#334690000000
0!
0'
#334700000000
1!
b111 %
1'
b111 +
#334710000000
0!
0'
#334720000000
1!
b1000 %
1'
b1000 +
#334730000000
0!
0'
#334740000000
1!
b1001 %
1'
b1001 +
#334750000000
1"
1(
#334760000000
0!
0"
b100 &
0'
0(
b100 ,
#334770000000
1!
b0 %
1'
b0 +
#334780000000
0!
0'
#334790000000
1!
1$
b1 %
1'
1*
b1 +
#334800000000
0!
0'
#334810000000
1!
b10 %
1'
b10 +
#334820000000
0!
0'
#334830000000
1!
b11 %
1'
b11 +
#334840000000
0!
0'
#334850000000
1!
b100 %
1'
b100 +
#334860000000
0!
0'
#334870000000
1!
b101 %
1'
b101 +
#334880000000
0!
0'
#334890000000
1!
b110 %
1'
b110 +
#334900000000
0!
0'
#334910000000
1!
b111 %
1'
b111 +
#334920000000
0!
0'
#334930000000
1!
0$
b1000 %
1'
0*
b1000 +
#334940000000
0!
0'
#334950000000
1!
b1001 %
1'
b1001 +
#334960000000
0!
0'
#334970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#334980000000
0!
0'
#334990000000
1!
1$
b1 %
1'
1*
b1 +
#335000000000
0!
0'
#335010000000
1!
b10 %
1'
b10 +
#335020000000
0!
0'
#335030000000
1!
b11 %
1'
b11 +
#335040000000
0!
0'
#335050000000
1!
b100 %
1'
b100 +
#335060000000
0!
0'
#335070000000
1!
b101 %
1'
b101 +
#335080000000
0!
0'
#335090000000
1!
0$
b110 %
1'
0*
b110 +
#335100000000
0!
0'
#335110000000
1!
b111 %
1'
b111 +
#335120000000
0!
0'
#335130000000
1!
b1000 %
1'
b1000 +
#335140000000
0!
0'
#335150000000
1!
b1001 %
1'
b1001 +
#335160000000
0!
0'
#335170000000
1!
b0 %
1'
b0 +
#335180000000
1"
1(
#335190000000
0!
0"
b100 &
0'
0(
b100 ,
#335200000000
1!
1$
b1 %
1'
1*
b1 +
#335210000000
0!
0'
#335220000000
1!
b10 %
1'
b10 +
#335230000000
0!
0'
#335240000000
1!
b11 %
1'
b11 +
#335250000000
0!
0'
#335260000000
1!
b100 %
1'
b100 +
#335270000000
0!
0'
#335280000000
1!
b101 %
1'
b101 +
#335290000000
0!
0'
#335300000000
1!
b110 %
1'
b110 +
#335310000000
0!
0'
#335320000000
1!
b111 %
1'
b111 +
#335330000000
0!
0'
#335340000000
1!
0$
b1000 %
1'
0*
b1000 +
#335350000000
0!
0'
#335360000000
1!
b1001 %
1'
b1001 +
#335370000000
0!
0'
#335380000000
1!
b0 %
1'
b0 +
#335390000000
0!
0'
#335400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#335410000000
0!
0'
#335420000000
1!
b10 %
1'
b10 +
#335430000000
0!
0'
#335440000000
1!
b11 %
1'
b11 +
#335450000000
0!
0'
#335460000000
1!
b100 %
1'
b100 +
#335470000000
0!
0'
#335480000000
1!
b101 %
1'
b101 +
#335490000000
0!
0'
#335500000000
1!
0$
b110 %
1'
0*
b110 +
#335510000000
0!
0'
#335520000000
1!
b111 %
1'
b111 +
#335530000000
0!
0'
#335540000000
1!
b1000 %
1'
b1000 +
#335550000000
0!
0'
#335560000000
1!
b1001 %
1'
b1001 +
#335570000000
0!
0'
#335580000000
1!
b0 %
1'
b0 +
#335590000000
0!
0'
#335600000000
1!
1$
b1 %
1'
1*
b1 +
#335610000000
1"
1(
#335620000000
0!
0"
b100 &
0'
0(
b100 ,
#335630000000
1!
b10 %
1'
b10 +
#335640000000
0!
0'
#335650000000
1!
b11 %
1'
b11 +
#335660000000
0!
0'
#335670000000
1!
b100 %
1'
b100 +
#335680000000
0!
0'
#335690000000
1!
b101 %
1'
b101 +
#335700000000
0!
0'
#335710000000
1!
b110 %
1'
b110 +
#335720000000
0!
0'
#335730000000
1!
b111 %
1'
b111 +
#335740000000
0!
0'
#335750000000
1!
0$
b1000 %
1'
0*
b1000 +
#335760000000
0!
0'
#335770000000
1!
b1001 %
1'
b1001 +
#335780000000
0!
0'
#335790000000
1!
b0 %
1'
b0 +
#335800000000
0!
0'
#335810000000
1!
1$
b1 %
1'
1*
b1 +
#335820000000
0!
0'
#335830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#335840000000
0!
0'
#335850000000
1!
b11 %
1'
b11 +
#335860000000
0!
0'
#335870000000
1!
b100 %
1'
b100 +
#335880000000
0!
0'
#335890000000
1!
b101 %
1'
b101 +
#335900000000
0!
0'
#335910000000
1!
0$
b110 %
1'
0*
b110 +
#335920000000
0!
0'
#335930000000
1!
b111 %
1'
b111 +
#335940000000
0!
0'
#335950000000
1!
b1000 %
1'
b1000 +
#335960000000
0!
0'
#335970000000
1!
b1001 %
1'
b1001 +
#335980000000
0!
0'
#335990000000
1!
b0 %
1'
b0 +
#336000000000
0!
0'
#336010000000
1!
1$
b1 %
1'
1*
b1 +
#336020000000
0!
0'
#336030000000
1!
b10 %
1'
b10 +
#336040000000
1"
1(
#336050000000
0!
0"
b100 &
0'
0(
b100 ,
#336060000000
1!
b11 %
1'
b11 +
#336070000000
0!
0'
#336080000000
1!
b100 %
1'
b100 +
#336090000000
0!
0'
#336100000000
1!
b101 %
1'
b101 +
#336110000000
0!
0'
#336120000000
1!
b110 %
1'
b110 +
#336130000000
0!
0'
#336140000000
1!
b111 %
1'
b111 +
#336150000000
0!
0'
#336160000000
1!
0$
b1000 %
1'
0*
b1000 +
#336170000000
0!
0'
#336180000000
1!
b1001 %
1'
b1001 +
#336190000000
0!
0'
#336200000000
1!
b0 %
1'
b0 +
#336210000000
0!
0'
#336220000000
1!
1$
b1 %
1'
1*
b1 +
#336230000000
0!
0'
#336240000000
1!
b10 %
1'
b10 +
#336250000000
0!
0'
#336260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#336270000000
0!
0'
#336280000000
1!
b100 %
1'
b100 +
#336290000000
0!
0'
#336300000000
1!
b101 %
1'
b101 +
#336310000000
0!
0'
#336320000000
1!
0$
b110 %
1'
0*
b110 +
#336330000000
0!
0'
#336340000000
1!
b111 %
1'
b111 +
#336350000000
0!
0'
#336360000000
1!
b1000 %
1'
b1000 +
#336370000000
0!
0'
#336380000000
1!
b1001 %
1'
b1001 +
#336390000000
0!
0'
#336400000000
1!
b0 %
1'
b0 +
#336410000000
0!
0'
#336420000000
1!
1$
b1 %
1'
1*
b1 +
#336430000000
0!
0'
#336440000000
1!
b10 %
1'
b10 +
#336450000000
0!
0'
#336460000000
1!
b11 %
1'
b11 +
#336470000000
1"
1(
#336480000000
0!
0"
b100 &
0'
0(
b100 ,
#336490000000
1!
b100 %
1'
b100 +
#336500000000
0!
0'
#336510000000
1!
b101 %
1'
b101 +
#336520000000
0!
0'
#336530000000
1!
b110 %
1'
b110 +
#336540000000
0!
0'
#336550000000
1!
b111 %
1'
b111 +
#336560000000
0!
0'
#336570000000
1!
0$
b1000 %
1'
0*
b1000 +
#336580000000
0!
0'
#336590000000
1!
b1001 %
1'
b1001 +
#336600000000
0!
0'
#336610000000
1!
b0 %
1'
b0 +
#336620000000
0!
0'
#336630000000
1!
1$
b1 %
1'
1*
b1 +
#336640000000
0!
0'
#336650000000
1!
b10 %
1'
b10 +
#336660000000
0!
0'
#336670000000
1!
b11 %
1'
b11 +
#336680000000
0!
0'
#336690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#336700000000
0!
0'
#336710000000
1!
b101 %
1'
b101 +
#336720000000
0!
0'
#336730000000
1!
0$
b110 %
1'
0*
b110 +
#336740000000
0!
0'
#336750000000
1!
b111 %
1'
b111 +
#336760000000
0!
0'
#336770000000
1!
b1000 %
1'
b1000 +
#336780000000
0!
0'
#336790000000
1!
b1001 %
1'
b1001 +
#336800000000
0!
0'
#336810000000
1!
b0 %
1'
b0 +
#336820000000
0!
0'
#336830000000
1!
1$
b1 %
1'
1*
b1 +
#336840000000
0!
0'
#336850000000
1!
b10 %
1'
b10 +
#336860000000
0!
0'
#336870000000
1!
b11 %
1'
b11 +
#336880000000
0!
0'
#336890000000
1!
b100 %
1'
b100 +
#336900000000
1"
1(
#336910000000
0!
0"
b100 &
0'
0(
b100 ,
#336920000000
1!
b101 %
1'
b101 +
#336930000000
0!
0'
#336940000000
1!
b110 %
1'
b110 +
#336950000000
0!
0'
#336960000000
1!
b111 %
1'
b111 +
#336970000000
0!
0'
#336980000000
1!
0$
b1000 %
1'
0*
b1000 +
#336990000000
0!
0'
#337000000000
1!
b1001 %
1'
b1001 +
#337010000000
0!
0'
#337020000000
1!
b0 %
1'
b0 +
#337030000000
0!
0'
#337040000000
1!
1$
b1 %
1'
1*
b1 +
#337050000000
0!
0'
#337060000000
1!
b10 %
1'
b10 +
#337070000000
0!
0'
#337080000000
1!
b11 %
1'
b11 +
#337090000000
0!
0'
#337100000000
1!
b100 %
1'
b100 +
#337110000000
0!
0'
#337120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#337130000000
0!
0'
#337140000000
1!
0$
b110 %
1'
0*
b110 +
#337150000000
0!
0'
#337160000000
1!
b111 %
1'
b111 +
#337170000000
0!
0'
#337180000000
1!
b1000 %
1'
b1000 +
#337190000000
0!
0'
#337200000000
1!
b1001 %
1'
b1001 +
#337210000000
0!
0'
#337220000000
1!
b0 %
1'
b0 +
#337230000000
0!
0'
#337240000000
1!
1$
b1 %
1'
1*
b1 +
#337250000000
0!
0'
#337260000000
1!
b10 %
1'
b10 +
#337270000000
0!
0'
#337280000000
1!
b11 %
1'
b11 +
#337290000000
0!
0'
#337300000000
1!
b100 %
1'
b100 +
#337310000000
0!
0'
#337320000000
1!
b101 %
1'
b101 +
#337330000000
1"
1(
#337340000000
0!
0"
b100 &
0'
0(
b100 ,
#337350000000
1!
b110 %
1'
b110 +
#337360000000
0!
0'
#337370000000
1!
b111 %
1'
b111 +
#337380000000
0!
0'
#337390000000
1!
0$
b1000 %
1'
0*
b1000 +
#337400000000
0!
0'
#337410000000
1!
b1001 %
1'
b1001 +
#337420000000
0!
0'
#337430000000
1!
b0 %
1'
b0 +
#337440000000
0!
0'
#337450000000
1!
1$
b1 %
1'
1*
b1 +
#337460000000
0!
0'
#337470000000
1!
b10 %
1'
b10 +
#337480000000
0!
0'
#337490000000
1!
b11 %
1'
b11 +
#337500000000
0!
0'
#337510000000
1!
b100 %
1'
b100 +
#337520000000
0!
0'
#337530000000
1!
b101 %
1'
b101 +
#337540000000
0!
0'
#337550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#337560000000
0!
0'
#337570000000
1!
b111 %
1'
b111 +
#337580000000
0!
0'
#337590000000
1!
b1000 %
1'
b1000 +
#337600000000
0!
0'
#337610000000
1!
b1001 %
1'
b1001 +
#337620000000
0!
0'
#337630000000
1!
b0 %
1'
b0 +
#337640000000
0!
0'
#337650000000
1!
1$
b1 %
1'
1*
b1 +
#337660000000
0!
0'
#337670000000
1!
b10 %
1'
b10 +
#337680000000
0!
0'
#337690000000
1!
b11 %
1'
b11 +
#337700000000
0!
0'
#337710000000
1!
b100 %
1'
b100 +
#337720000000
0!
0'
#337730000000
1!
b101 %
1'
b101 +
#337740000000
0!
0'
#337750000000
1!
0$
b110 %
1'
0*
b110 +
#337760000000
1"
1(
#337770000000
0!
0"
b100 &
0'
0(
b100 ,
#337780000000
1!
1$
b111 %
1'
1*
b111 +
#337790000000
0!
0'
#337800000000
1!
0$
b1000 %
1'
0*
b1000 +
#337810000000
0!
0'
#337820000000
1!
b1001 %
1'
b1001 +
#337830000000
0!
0'
#337840000000
1!
b0 %
1'
b0 +
#337850000000
0!
0'
#337860000000
1!
1$
b1 %
1'
1*
b1 +
#337870000000
0!
0'
#337880000000
1!
b10 %
1'
b10 +
#337890000000
0!
0'
#337900000000
1!
b11 %
1'
b11 +
#337910000000
0!
0'
#337920000000
1!
b100 %
1'
b100 +
#337930000000
0!
0'
#337940000000
1!
b101 %
1'
b101 +
#337950000000
0!
0'
#337960000000
1!
b110 %
1'
b110 +
#337970000000
0!
0'
#337980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#337990000000
0!
0'
#338000000000
1!
b1000 %
1'
b1000 +
#338010000000
0!
0'
#338020000000
1!
b1001 %
1'
b1001 +
#338030000000
0!
0'
#338040000000
1!
b0 %
1'
b0 +
#338050000000
0!
0'
#338060000000
1!
1$
b1 %
1'
1*
b1 +
#338070000000
0!
0'
#338080000000
1!
b10 %
1'
b10 +
#338090000000
0!
0'
#338100000000
1!
b11 %
1'
b11 +
#338110000000
0!
0'
#338120000000
1!
b100 %
1'
b100 +
#338130000000
0!
0'
#338140000000
1!
b101 %
1'
b101 +
#338150000000
0!
0'
#338160000000
1!
0$
b110 %
1'
0*
b110 +
#338170000000
0!
0'
#338180000000
1!
b111 %
1'
b111 +
#338190000000
1"
1(
#338200000000
0!
0"
b100 &
0'
0(
b100 ,
#338210000000
1!
b1000 %
1'
b1000 +
#338220000000
0!
0'
#338230000000
1!
b1001 %
1'
b1001 +
#338240000000
0!
0'
#338250000000
1!
b0 %
1'
b0 +
#338260000000
0!
0'
#338270000000
1!
1$
b1 %
1'
1*
b1 +
#338280000000
0!
0'
#338290000000
1!
b10 %
1'
b10 +
#338300000000
0!
0'
#338310000000
1!
b11 %
1'
b11 +
#338320000000
0!
0'
#338330000000
1!
b100 %
1'
b100 +
#338340000000
0!
0'
#338350000000
1!
b101 %
1'
b101 +
#338360000000
0!
0'
#338370000000
1!
b110 %
1'
b110 +
#338380000000
0!
0'
#338390000000
1!
b111 %
1'
b111 +
#338400000000
0!
0'
#338410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#338420000000
0!
0'
#338430000000
1!
b1001 %
1'
b1001 +
#338440000000
0!
0'
#338450000000
1!
b0 %
1'
b0 +
#338460000000
0!
0'
#338470000000
1!
1$
b1 %
1'
1*
b1 +
#338480000000
0!
0'
#338490000000
1!
b10 %
1'
b10 +
#338500000000
0!
0'
#338510000000
1!
b11 %
1'
b11 +
#338520000000
0!
0'
#338530000000
1!
b100 %
1'
b100 +
#338540000000
0!
0'
#338550000000
1!
b101 %
1'
b101 +
#338560000000
0!
0'
#338570000000
1!
0$
b110 %
1'
0*
b110 +
#338580000000
0!
0'
#338590000000
1!
b111 %
1'
b111 +
#338600000000
0!
0'
#338610000000
1!
b1000 %
1'
b1000 +
#338620000000
1"
1(
#338630000000
0!
0"
b100 &
0'
0(
b100 ,
#338640000000
1!
b1001 %
1'
b1001 +
#338650000000
0!
0'
#338660000000
1!
b0 %
1'
b0 +
#338670000000
0!
0'
#338680000000
1!
1$
b1 %
1'
1*
b1 +
#338690000000
0!
0'
#338700000000
1!
b10 %
1'
b10 +
#338710000000
0!
0'
#338720000000
1!
b11 %
1'
b11 +
#338730000000
0!
0'
#338740000000
1!
b100 %
1'
b100 +
#338750000000
0!
0'
#338760000000
1!
b101 %
1'
b101 +
#338770000000
0!
0'
#338780000000
1!
b110 %
1'
b110 +
#338790000000
0!
0'
#338800000000
1!
b111 %
1'
b111 +
#338810000000
0!
0'
#338820000000
1!
0$
b1000 %
1'
0*
b1000 +
#338830000000
0!
0'
#338840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#338850000000
0!
0'
#338860000000
1!
b0 %
1'
b0 +
#338870000000
0!
0'
#338880000000
1!
1$
b1 %
1'
1*
b1 +
#338890000000
0!
0'
#338900000000
1!
b10 %
1'
b10 +
#338910000000
0!
0'
#338920000000
1!
b11 %
1'
b11 +
#338930000000
0!
0'
#338940000000
1!
b100 %
1'
b100 +
#338950000000
0!
0'
#338960000000
1!
b101 %
1'
b101 +
#338970000000
0!
0'
#338980000000
1!
0$
b110 %
1'
0*
b110 +
#338990000000
0!
0'
#339000000000
1!
b111 %
1'
b111 +
#339010000000
0!
0'
#339020000000
1!
b1000 %
1'
b1000 +
#339030000000
0!
0'
#339040000000
1!
b1001 %
1'
b1001 +
#339050000000
1"
1(
#339060000000
0!
0"
b100 &
0'
0(
b100 ,
#339070000000
1!
b0 %
1'
b0 +
#339080000000
0!
0'
#339090000000
1!
1$
b1 %
1'
1*
b1 +
#339100000000
0!
0'
#339110000000
1!
b10 %
1'
b10 +
#339120000000
0!
0'
#339130000000
1!
b11 %
1'
b11 +
#339140000000
0!
0'
#339150000000
1!
b100 %
1'
b100 +
#339160000000
0!
0'
#339170000000
1!
b101 %
1'
b101 +
#339180000000
0!
0'
#339190000000
1!
b110 %
1'
b110 +
#339200000000
0!
0'
#339210000000
1!
b111 %
1'
b111 +
#339220000000
0!
0'
#339230000000
1!
0$
b1000 %
1'
0*
b1000 +
#339240000000
0!
0'
#339250000000
1!
b1001 %
1'
b1001 +
#339260000000
0!
0'
#339270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#339280000000
0!
0'
#339290000000
1!
1$
b1 %
1'
1*
b1 +
#339300000000
0!
0'
#339310000000
1!
b10 %
1'
b10 +
#339320000000
0!
0'
#339330000000
1!
b11 %
1'
b11 +
#339340000000
0!
0'
#339350000000
1!
b100 %
1'
b100 +
#339360000000
0!
0'
#339370000000
1!
b101 %
1'
b101 +
#339380000000
0!
0'
#339390000000
1!
0$
b110 %
1'
0*
b110 +
#339400000000
0!
0'
#339410000000
1!
b111 %
1'
b111 +
#339420000000
0!
0'
#339430000000
1!
b1000 %
1'
b1000 +
#339440000000
0!
0'
#339450000000
1!
b1001 %
1'
b1001 +
#339460000000
0!
0'
#339470000000
1!
b0 %
1'
b0 +
#339480000000
1"
1(
#339490000000
0!
0"
b100 &
0'
0(
b100 ,
#339500000000
1!
1$
b1 %
1'
1*
b1 +
#339510000000
0!
0'
#339520000000
1!
b10 %
1'
b10 +
#339530000000
0!
0'
#339540000000
1!
b11 %
1'
b11 +
#339550000000
0!
0'
#339560000000
1!
b100 %
1'
b100 +
#339570000000
0!
0'
#339580000000
1!
b101 %
1'
b101 +
#339590000000
0!
0'
#339600000000
1!
b110 %
1'
b110 +
#339610000000
0!
0'
#339620000000
1!
b111 %
1'
b111 +
#339630000000
0!
0'
#339640000000
1!
0$
b1000 %
1'
0*
b1000 +
#339650000000
0!
0'
#339660000000
1!
b1001 %
1'
b1001 +
#339670000000
0!
0'
#339680000000
1!
b0 %
1'
b0 +
#339690000000
0!
0'
#339700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#339710000000
0!
0'
#339720000000
1!
b10 %
1'
b10 +
#339730000000
0!
0'
#339740000000
1!
b11 %
1'
b11 +
#339750000000
0!
0'
#339760000000
1!
b100 %
1'
b100 +
#339770000000
0!
0'
#339780000000
1!
b101 %
1'
b101 +
#339790000000
0!
0'
#339800000000
1!
0$
b110 %
1'
0*
b110 +
#339810000000
0!
0'
#339820000000
1!
b111 %
1'
b111 +
#339830000000
0!
0'
#339840000000
1!
b1000 %
1'
b1000 +
#339850000000
0!
0'
#339860000000
1!
b1001 %
1'
b1001 +
#339870000000
0!
0'
#339880000000
1!
b0 %
1'
b0 +
#339890000000
0!
0'
#339900000000
1!
1$
b1 %
1'
1*
b1 +
#339910000000
1"
1(
#339920000000
0!
0"
b100 &
0'
0(
b100 ,
#339930000000
1!
b10 %
1'
b10 +
#339940000000
0!
0'
#339950000000
1!
b11 %
1'
b11 +
#339960000000
0!
0'
#339970000000
1!
b100 %
1'
b100 +
#339980000000
0!
0'
#339990000000
1!
b101 %
1'
b101 +
#340000000000
0!
0'
#340010000000
1!
b110 %
1'
b110 +
#340020000000
0!
0'
#340030000000
1!
b111 %
1'
b111 +
#340040000000
0!
0'
#340050000000
1!
0$
b1000 %
1'
0*
b1000 +
#340060000000
0!
0'
#340070000000
1!
b1001 %
1'
b1001 +
#340080000000
0!
0'
#340090000000
1!
b0 %
1'
b0 +
#340100000000
0!
0'
#340110000000
1!
1$
b1 %
1'
1*
b1 +
#340120000000
0!
0'
#340130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#340140000000
0!
0'
#340150000000
1!
b11 %
1'
b11 +
#340160000000
0!
0'
#340170000000
1!
b100 %
1'
b100 +
#340180000000
0!
0'
#340190000000
1!
b101 %
1'
b101 +
#340200000000
0!
0'
#340210000000
1!
0$
b110 %
1'
0*
b110 +
#340220000000
0!
0'
#340230000000
1!
b111 %
1'
b111 +
#340240000000
0!
0'
#340250000000
1!
b1000 %
1'
b1000 +
#340260000000
0!
0'
#340270000000
1!
b1001 %
1'
b1001 +
#340280000000
0!
0'
#340290000000
1!
b0 %
1'
b0 +
#340300000000
0!
0'
#340310000000
1!
1$
b1 %
1'
1*
b1 +
#340320000000
0!
0'
#340330000000
1!
b10 %
1'
b10 +
#340340000000
1"
1(
#340350000000
0!
0"
b100 &
0'
0(
b100 ,
#340360000000
1!
b11 %
1'
b11 +
#340370000000
0!
0'
#340380000000
1!
b100 %
1'
b100 +
#340390000000
0!
0'
#340400000000
1!
b101 %
1'
b101 +
#340410000000
0!
0'
#340420000000
1!
b110 %
1'
b110 +
#340430000000
0!
0'
#340440000000
1!
b111 %
1'
b111 +
#340450000000
0!
0'
#340460000000
1!
0$
b1000 %
1'
0*
b1000 +
#340470000000
0!
0'
#340480000000
1!
b1001 %
1'
b1001 +
#340490000000
0!
0'
#340500000000
1!
b0 %
1'
b0 +
#340510000000
0!
0'
#340520000000
1!
1$
b1 %
1'
1*
b1 +
#340530000000
0!
0'
#340540000000
1!
b10 %
1'
b10 +
#340550000000
0!
0'
#340560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#340570000000
0!
0'
#340580000000
1!
b100 %
1'
b100 +
#340590000000
0!
0'
#340600000000
1!
b101 %
1'
b101 +
#340610000000
0!
0'
#340620000000
1!
0$
b110 %
1'
0*
b110 +
#340630000000
0!
0'
#340640000000
1!
b111 %
1'
b111 +
#340650000000
0!
0'
#340660000000
1!
b1000 %
1'
b1000 +
#340670000000
0!
0'
#340680000000
1!
b1001 %
1'
b1001 +
#340690000000
0!
0'
#340700000000
1!
b0 %
1'
b0 +
#340710000000
0!
0'
#340720000000
1!
1$
b1 %
1'
1*
b1 +
#340730000000
0!
0'
#340740000000
1!
b10 %
1'
b10 +
#340750000000
0!
0'
#340760000000
1!
b11 %
1'
b11 +
#340770000000
1"
1(
#340780000000
0!
0"
b100 &
0'
0(
b100 ,
#340790000000
1!
b100 %
1'
b100 +
#340800000000
0!
0'
#340810000000
1!
b101 %
1'
b101 +
#340820000000
0!
0'
#340830000000
1!
b110 %
1'
b110 +
#340840000000
0!
0'
#340850000000
1!
b111 %
1'
b111 +
#340860000000
0!
0'
#340870000000
1!
0$
b1000 %
1'
0*
b1000 +
#340880000000
0!
0'
#340890000000
1!
b1001 %
1'
b1001 +
#340900000000
0!
0'
#340910000000
1!
b0 %
1'
b0 +
#340920000000
0!
0'
#340930000000
1!
1$
b1 %
1'
1*
b1 +
#340940000000
0!
0'
#340950000000
1!
b10 %
1'
b10 +
#340960000000
0!
0'
#340970000000
1!
b11 %
1'
b11 +
#340980000000
0!
0'
#340990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#341000000000
0!
0'
#341010000000
1!
b101 %
1'
b101 +
#341020000000
0!
0'
#341030000000
1!
0$
b110 %
1'
0*
b110 +
#341040000000
0!
0'
#341050000000
1!
b111 %
1'
b111 +
#341060000000
0!
0'
#341070000000
1!
b1000 %
1'
b1000 +
#341080000000
0!
0'
#341090000000
1!
b1001 %
1'
b1001 +
#341100000000
0!
0'
#341110000000
1!
b0 %
1'
b0 +
#341120000000
0!
0'
#341130000000
1!
1$
b1 %
1'
1*
b1 +
#341140000000
0!
0'
#341150000000
1!
b10 %
1'
b10 +
#341160000000
0!
0'
#341170000000
1!
b11 %
1'
b11 +
#341180000000
0!
0'
#341190000000
1!
b100 %
1'
b100 +
#341200000000
1"
1(
#341210000000
0!
0"
b100 &
0'
0(
b100 ,
#341220000000
1!
b101 %
1'
b101 +
#341230000000
0!
0'
#341240000000
1!
b110 %
1'
b110 +
#341250000000
0!
0'
#341260000000
1!
b111 %
1'
b111 +
#341270000000
0!
0'
#341280000000
1!
0$
b1000 %
1'
0*
b1000 +
#341290000000
0!
0'
#341300000000
1!
b1001 %
1'
b1001 +
#341310000000
0!
0'
#341320000000
1!
b0 %
1'
b0 +
#341330000000
0!
0'
#341340000000
1!
1$
b1 %
1'
1*
b1 +
#341350000000
0!
0'
#341360000000
1!
b10 %
1'
b10 +
#341370000000
0!
0'
#341380000000
1!
b11 %
1'
b11 +
#341390000000
0!
0'
#341400000000
1!
b100 %
1'
b100 +
#341410000000
0!
0'
#341420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#341430000000
0!
0'
#341440000000
1!
0$
b110 %
1'
0*
b110 +
#341450000000
0!
0'
#341460000000
1!
b111 %
1'
b111 +
#341470000000
0!
0'
#341480000000
1!
b1000 %
1'
b1000 +
#341490000000
0!
0'
#341500000000
1!
b1001 %
1'
b1001 +
#341510000000
0!
0'
#341520000000
1!
b0 %
1'
b0 +
#341530000000
0!
0'
#341540000000
1!
1$
b1 %
1'
1*
b1 +
#341550000000
0!
0'
#341560000000
1!
b10 %
1'
b10 +
#341570000000
0!
0'
#341580000000
1!
b11 %
1'
b11 +
#341590000000
0!
0'
#341600000000
1!
b100 %
1'
b100 +
#341610000000
0!
0'
#341620000000
1!
b101 %
1'
b101 +
#341630000000
1"
1(
#341640000000
0!
0"
b100 &
0'
0(
b100 ,
#341650000000
1!
b110 %
1'
b110 +
#341660000000
0!
0'
#341670000000
1!
b111 %
1'
b111 +
#341680000000
0!
0'
#341690000000
1!
0$
b1000 %
1'
0*
b1000 +
#341700000000
0!
0'
#341710000000
1!
b1001 %
1'
b1001 +
#341720000000
0!
0'
#341730000000
1!
b0 %
1'
b0 +
#341740000000
0!
0'
#341750000000
1!
1$
b1 %
1'
1*
b1 +
#341760000000
0!
0'
#341770000000
1!
b10 %
1'
b10 +
#341780000000
0!
0'
#341790000000
1!
b11 %
1'
b11 +
#341800000000
0!
0'
#341810000000
1!
b100 %
1'
b100 +
#341820000000
0!
0'
#341830000000
1!
b101 %
1'
b101 +
#341840000000
0!
0'
#341850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#341860000000
0!
0'
#341870000000
1!
b111 %
1'
b111 +
#341880000000
0!
0'
#341890000000
1!
b1000 %
1'
b1000 +
#341900000000
0!
0'
#341910000000
1!
b1001 %
1'
b1001 +
#341920000000
0!
0'
#341930000000
1!
b0 %
1'
b0 +
#341940000000
0!
0'
#341950000000
1!
1$
b1 %
1'
1*
b1 +
#341960000000
0!
0'
#341970000000
1!
b10 %
1'
b10 +
#341980000000
0!
0'
#341990000000
1!
b11 %
1'
b11 +
#342000000000
0!
0'
#342010000000
1!
b100 %
1'
b100 +
#342020000000
0!
0'
#342030000000
1!
b101 %
1'
b101 +
#342040000000
0!
0'
#342050000000
1!
0$
b110 %
1'
0*
b110 +
#342060000000
1"
1(
#342070000000
0!
0"
b100 &
0'
0(
b100 ,
#342080000000
1!
1$
b111 %
1'
1*
b111 +
#342090000000
0!
0'
#342100000000
1!
0$
b1000 %
1'
0*
b1000 +
#342110000000
0!
0'
#342120000000
1!
b1001 %
1'
b1001 +
#342130000000
0!
0'
#342140000000
1!
b0 %
1'
b0 +
#342150000000
0!
0'
#342160000000
1!
1$
b1 %
1'
1*
b1 +
#342170000000
0!
0'
#342180000000
1!
b10 %
1'
b10 +
#342190000000
0!
0'
#342200000000
1!
b11 %
1'
b11 +
#342210000000
0!
0'
#342220000000
1!
b100 %
1'
b100 +
#342230000000
0!
0'
#342240000000
1!
b101 %
1'
b101 +
#342250000000
0!
0'
#342260000000
1!
b110 %
1'
b110 +
#342270000000
0!
0'
#342280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#342290000000
0!
0'
#342300000000
1!
b1000 %
1'
b1000 +
#342310000000
0!
0'
#342320000000
1!
b1001 %
1'
b1001 +
#342330000000
0!
0'
#342340000000
1!
b0 %
1'
b0 +
#342350000000
0!
0'
#342360000000
1!
1$
b1 %
1'
1*
b1 +
#342370000000
0!
0'
#342380000000
1!
b10 %
1'
b10 +
#342390000000
0!
0'
#342400000000
1!
b11 %
1'
b11 +
#342410000000
0!
0'
#342420000000
1!
b100 %
1'
b100 +
#342430000000
0!
0'
#342440000000
1!
b101 %
1'
b101 +
#342450000000
0!
0'
#342460000000
1!
0$
b110 %
1'
0*
b110 +
#342470000000
0!
0'
#342480000000
1!
b111 %
1'
b111 +
#342490000000
1"
1(
#342500000000
0!
0"
b100 &
0'
0(
b100 ,
#342510000000
1!
b1000 %
1'
b1000 +
#342520000000
0!
0'
#342530000000
1!
b1001 %
1'
b1001 +
#342540000000
0!
0'
#342550000000
1!
b0 %
1'
b0 +
#342560000000
0!
0'
#342570000000
1!
1$
b1 %
1'
1*
b1 +
#342580000000
0!
0'
#342590000000
1!
b10 %
1'
b10 +
#342600000000
0!
0'
#342610000000
1!
b11 %
1'
b11 +
#342620000000
0!
0'
#342630000000
1!
b100 %
1'
b100 +
#342640000000
0!
0'
#342650000000
1!
b101 %
1'
b101 +
#342660000000
0!
0'
#342670000000
1!
b110 %
1'
b110 +
#342680000000
0!
0'
#342690000000
1!
b111 %
1'
b111 +
#342700000000
0!
0'
#342710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#342720000000
0!
0'
#342730000000
1!
b1001 %
1'
b1001 +
#342740000000
0!
0'
#342750000000
1!
b0 %
1'
b0 +
#342760000000
0!
0'
#342770000000
1!
1$
b1 %
1'
1*
b1 +
#342780000000
0!
0'
#342790000000
1!
b10 %
1'
b10 +
#342800000000
0!
0'
#342810000000
1!
b11 %
1'
b11 +
#342820000000
0!
0'
#342830000000
1!
b100 %
1'
b100 +
#342840000000
0!
0'
#342850000000
1!
b101 %
1'
b101 +
#342860000000
0!
0'
#342870000000
1!
0$
b110 %
1'
0*
b110 +
#342880000000
0!
0'
#342890000000
1!
b111 %
1'
b111 +
#342900000000
0!
0'
#342910000000
1!
b1000 %
1'
b1000 +
#342920000000
1"
1(
#342930000000
0!
0"
b100 &
0'
0(
b100 ,
#342940000000
1!
b1001 %
1'
b1001 +
#342950000000
0!
0'
#342960000000
1!
b0 %
1'
b0 +
#342970000000
0!
0'
#342980000000
1!
1$
b1 %
1'
1*
b1 +
#342990000000
0!
0'
#343000000000
1!
b10 %
1'
b10 +
#343010000000
0!
0'
#343020000000
1!
b11 %
1'
b11 +
#343030000000
0!
0'
#343040000000
1!
b100 %
1'
b100 +
#343050000000
0!
0'
#343060000000
1!
b101 %
1'
b101 +
#343070000000
0!
0'
#343080000000
1!
b110 %
1'
b110 +
#343090000000
0!
0'
#343100000000
1!
b111 %
1'
b111 +
#343110000000
0!
0'
#343120000000
1!
0$
b1000 %
1'
0*
b1000 +
#343130000000
0!
0'
#343140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#343150000000
0!
0'
#343160000000
1!
b0 %
1'
b0 +
#343170000000
0!
0'
#343180000000
1!
1$
b1 %
1'
1*
b1 +
#343190000000
0!
0'
#343200000000
1!
b10 %
1'
b10 +
#343210000000
0!
0'
#343220000000
1!
b11 %
1'
b11 +
#343230000000
0!
0'
#343240000000
1!
b100 %
1'
b100 +
#343250000000
0!
0'
#343260000000
1!
b101 %
1'
b101 +
#343270000000
0!
0'
#343280000000
1!
0$
b110 %
1'
0*
b110 +
#343290000000
0!
0'
#343300000000
1!
b111 %
1'
b111 +
#343310000000
0!
0'
#343320000000
1!
b1000 %
1'
b1000 +
#343330000000
0!
0'
#343340000000
1!
b1001 %
1'
b1001 +
#343350000000
1"
1(
#343360000000
0!
0"
b100 &
0'
0(
b100 ,
#343370000000
1!
b0 %
1'
b0 +
#343380000000
0!
0'
#343390000000
1!
1$
b1 %
1'
1*
b1 +
#343400000000
0!
0'
#343410000000
1!
b10 %
1'
b10 +
#343420000000
0!
0'
#343430000000
1!
b11 %
1'
b11 +
#343440000000
0!
0'
#343450000000
1!
b100 %
1'
b100 +
#343460000000
0!
0'
#343470000000
1!
b101 %
1'
b101 +
#343480000000
0!
0'
#343490000000
1!
b110 %
1'
b110 +
#343500000000
0!
0'
#343510000000
1!
b111 %
1'
b111 +
#343520000000
0!
0'
#343530000000
1!
0$
b1000 %
1'
0*
b1000 +
#343540000000
0!
0'
#343550000000
1!
b1001 %
1'
b1001 +
#343560000000
0!
0'
#343570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#343580000000
0!
0'
#343590000000
1!
1$
b1 %
1'
1*
b1 +
#343600000000
0!
0'
#343610000000
1!
b10 %
1'
b10 +
#343620000000
0!
0'
#343630000000
1!
b11 %
1'
b11 +
#343640000000
0!
0'
#343650000000
1!
b100 %
1'
b100 +
#343660000000
0!
0'
#343670000000
1!
b101 %
1'
b101 +
#343680000000
0!
0'
#343690000000
1!
0$
b110 %
1'
0*
b110 +
#343700000000
0!
0'
#343710000000
1!
b111 %
1'
b111 +
#343720000000
0!
0'
#343730000000
1!
b1000 %
1'
b1000 +
#343740000000
0!
0'
#343750000000
1!
b1001 %
1'
b1001 +
#343760000000
0!
0'
#343770000000
1!
b0 %
1'
b0 +
#343780000000
1"
1(
#343790000000
0!
0"
b100 &
0'
0(
b100 ,
#343800000000
1!
1$
b1 %
1'
1*
b1 +
#343810000000
0!
0'
#343820000000
1!
b10 %
1'
b10 +
#343830000000
0!
0'
#343840000000
1!
b11 %
1'
b11 +
#343850000000
0!
0'
#343860000000
1!
b100 %
1'
b100 +
#343870000000
0!
0'
#343880000000
1!
b101 %
1'
b101 +
#343890000000
0!
0'
#343900000000
1!
b110 %
1'
b110 +
#343910000000
0!
0'
#343920000000
1!
b111 %
1'
b111 +
#343930000000
0!
0'
#343940000000
1!
0$
b1000 %
1'
0*
b1000 +
#343950000000
0!
0'
#343960000000
1!
b1001 %
1'
b1001 +
#343970000000
0!
0'
#343980000000
1!
b0 %
1'
b0 +
#343990000000
0!
0'
#344000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#344010000000
0!
0'
#344020000000
1!
b10 %
1'
b10 +
#344030000000
0!
0'
#344040000000
1!
b11 %
1'
b11 +
#344050000000
0!
0'
#344060000000
1!
b100 %
1'
b100 +
#344070000000
0!
0'
#344080000000
1!
b101 %
1'
b101 +
#344090000000
0!
0'
#344100000000
1!
0$
b110 %
1'
0*
b110 +
#344110000000
0!
0'
#344120000000
1!
b111 %
1'
b111 +
#344130000000
0!
0'
#344140000000
1!
b1000 %
1'
b1000 +
#344150000000
0!
0'
#344160000000
1!
b1001 %
1'
b1001 +
#344170000000
0!
0'
#344180000000
1!
b0 %
1'
b0 +
#344190000000
0!
0'
#344200000000
1!
1$
b1 %
1'
1*
b1 +
#344210000000
1"
1(
#344220000000
0!
0"
b100 &
0'
0(
b100 ,
#344230000000
1!
b10 %
1'
b10 +
#344240000000
0!
0'
#344250000000
1!
b11 %
1'
b11 +
#344260000000
0!
0'
#344270000000
1!
b100 %
1'
b100 +
#344280000000
0!
0'
#344290000000
1!
b101 %
1'
b101 +
#344300000000
0!
0'
#344310000000
1!
b110 %
1'
b110 +
#344320000000
0!
0'
#344330000000
1!
b111 %
1'
b111 +
#344340000000
0!
0'
#344350000000
1!
0$
b1000 %
1'
0*
b1000 +
#344360000000
0!
0'
#344370000000
1!
b1001 %
1'
b1001 +
#344380000000
0!
0'
#344390000000
1!
b0 %
1'
b0 +
#344400000000
0!
0'
#344410000000
1!
1$
b1 %
1'
1*
b1 +
#344420000000
0!
0'
#344430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#344440000000
0!
0'
#344450000000
1!
b11 %
1'
b11 +
#344460000000
0!
0'
#344470000000
1!
b100 %
1'
b100 +
#344480000000
0!
0'
#344490000000
1!
b101 %
1'
b101 +
#344500000000
0!
0'
#344510000000
1!
0$
b110 %
1'
0*
b110 +
#344520000000
0!
0'
#344530000000
1!
b111 %
1'
b111 +
#344540000000
0!
0'
#344550000000
1!
b1000 %
1'
b1000 +
#344560000000
0!
0'
#344570000000
1!
b1001 %
1'
b1001 +
#344580000000
0!
0'
#344590000000
1!
b0 %
1'
b0 +
#344600000000
0!
0'
#344610000000
1!
1$
b1 %
1'
1*
b1 +
#344620000000
0!
0'
#344630000000
1!
b10 %
1'
b10 +
#344640000000
1"
1(
#344650000000
0!
0"
b100 &
0'
0(
b100 ,
#344660000000
1!
b11 %
1'
b11 +
#344670000000
0!
0'
#344680000000
1!
b100 %
1'
b100 +
#344690000000
0!
0'
#344700000000
1!
b101 %
1'
b101 +
#344710000000
0!
0'
#344720000000
1!
b110 %
1'
b110 +
#344730000000
0!
0'
#344740000000
1!
b111 %
1'
b111 +
#344750000000
0!
0'
#344760000000
1!
0$
b1000 %
1'
0*
b1000 +
#344770000000
0!
0'
#344780000000
1!
b1001 %
1'
b1001 +
#344790000000
0!
0'
#344800000000
1!
b0 %
1'
b0 +
#344810000000
0!
0'
#344820000000
1!
1$
b1 %
1'
1*
b1 +
#344830000000
0!
0'
#344840000000
1!
b10 %
1'
b10 +
#344850000000
0!
0'
#344860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#344870000000
0!
0'
#344880000000
1!
b100 %
1'
b100 +
#344890000000
0!
0'
#344900000000
1!
b101 %
1'
b101 +
#344910000000
0!
0'
#344920000000
1!
0$
b110 %
1'
0*
b110 +
#344930000000
0!
0'
#344940000000
1!
b111 %
1'
b111 +
#344950000000
0!
0'
#344960000000
1!
b1000 %
1'
b1000 +
#344970000000
0!
0'
#344980000000
1!
b1001 %
1'
b1001 +
#344990000000
0!
0'
#345000000000
1!
b0 %
1'
b0 +
#345010000000
0!
0'
#345020000000
1!
1$
b1 %
1'
1*
b1 +
#345030000000
0!
0'
#345040000000
1!
b10 %
1'
b10 +
#345050000000
0!
0'
#345060000000
1!
b11 %
1'
b11 +
#345070000000
1"
1(
#345080000000
0!
0"
b100 &
0'
0(
b100 ,
#345090000000
1!
b100 %
1'
b100 +
#345100000000
0!
0'
#345110000000
1!
b101 %
1'
b101 +
#345120000000
0!
0'
#345130000000
1!
b110 %
1'
b110 +
#345140000000
0!
0'
#345150000000
1!
b111 %
1'
b111 +
#345160000000
0!
0'
#345170000000
1!
0$
b1000 %
1'
0*
b1000 +
#345180000000
0!
0'
#345190000000
1!
b1001 %
1'
b1001 +
#345200000000
0!
0'
#345210000000
1!
b0 %
1'
b0 +
#345220000000
0!
0'
#345230000000
1!
1$
b1 %
1'
1*
b1 +
#345240000000
0!
0'
#345250000000
1!
b10 %
1'
b10 +
#345260000000
0!
0'
#345270000000
1!
b11 %
1'
b11 +
#345280000000
0!
0'
#345290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#345300000000
0!
0'
#345310000000
1!
b101 %
1'
b101 +
#345320000000
0!
0'
#345330000000
1!
0$
b110 %
1'
0*
b110 +
#345340000000
0!
0'
#345350000000
1!
b111 %
1'
b111 +
#345360000000
0!
0'
#345370000000
1!
b1000 %
1'
b1000 +
#345380000000
0!
0'
#345390000000
1!
b1001 %
1'
b1001 +
#345400000000
0!
0'
#345410000000
1!
b0 %
1'
b0 +
#345420000000
0!
0'
#345430000000
1!
1$
b1 %
1'
1*
b1 +
#345440000000
0!
0'
#345450000000
1!
b10 %
1'
b10 +
#345460000000
0!
0'
#345470000000
1!
b11 %
1'
b11 +
#345480000000
0!
0'
#345490000000
1!
b100 %
1'
b100 +
#345500000000
1"
1(
#345510000000
0!
0"
b100 &
0'
0(
b100 ,
#345520000000
1!
b101 %
1'
b101 +
#345530000000
0!
0'
#345540000000
1!
b110 %
1'
b110 +
#345550000000
0!
0'
#345560000000
1!
b111 %
1'
b111 +
#345570000000
0!
0'
#345580000000
1!
0$
b1000 %
1'
0*
b1000 +
#345590000000
0!
0'
#345600000000
1!
b1001 %
1'
b1001 +
#345610000000
0!
0'
#345620000000
1!
b0 %
1'
b0 +
#345630000000
0!
0'
#345640000000
1!
1$
b1 %
1'
1*
b1 +
#345650000000
0!
0'
#345660000000
1!
b10 %
1'
b10 +
#345670000000
0!
0'
#345680000000
1!
b11 %
1'
b11 +
#345690000000
0!
0'
#345700000000
1!
b100 %
1'
b100 +
#345710000000
0!
0'
#345720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#345730000000
0!
0'
#345740000000
1!
0$
b110 %
1'
0*
b110 +
#345750000000
0!
0'
#345760000000
1!
b111 %
1'
b111 +
#345770000000
0!
0'
#345780000000
1!
b1000 %
1'
b1000 +
#345790000000
0!
0'
#345800000000
1!
b1001 %
1'
b1001 +
#345810000000
0!
0'
#345820000000
1!
b0 %
1'
b0 +
#345830000000
0!
0'
#345840000000
1!
1$
b1 %
1'
1*
b1 +
#345850000000
0!
0'
#345860000000
1!
b10 %
1'
b10 +
#345870000000
0!
0'
#345880000000
1!
b11 %
1'
b11 +
#345890000000
0!
0'
#345900000000
1!
b100 %
1'
b100 +
#345910000000
0!
0'
#345920000000
1!
b101 %
1'
b101 +
#345930000000
1"
1(
#345940000000
0!
0"
b100 &
0'
0(
b100 ,
#345950000000
1!
b110 %
1'
b110 +
#345960000000
0!
0'
#345970000000
1!
b111 %
1'
b111 +
#345980000000
0!
0'
#345990000000
1!
0$
b1000 %
1'
0*
b1000 +
#346000000000
0!
0'
#346010000000
1!
b1001 %
1'
b1001 +
#346020000000
0!
0'
#346030000000
1!
b0 %
1'
b0 +
#346040000000
0!
0'
#346050000000
1!
1$
b1 %
1'
1*
b1 +
#346060000000
0!
0'
#346070000000
1!
b10 %
1'
b10 +
#346080000000
0!
0'
#346090000000
1!
b11 %
1'
b11 +
#346100000000
0!
0'
#346110000000
1!
b100 %
1'
b100 +
#346120000000
0!
0'
#346130000000
1!
b101 %
1'
b101 +
#346140000000
0!
0'
#346150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#346160000000
0!
0'
#346170000000
1!
b111 %
1'
b111 +
#346180000000
0!
0'
#346190000000
1!
b1000 %
1'
b1000 +
#346200000000
0!
0'
#346210000000
1!
b1001 %
1'
b1001 +
#346220000000
0!
0'
#346230000000
1!
b0 %
1'
b0 +
#346240000000
0!
0'
#346250000000
1!
1$
b1 %
1'
1*
b1 +
#346260000000
0!
0'
#346270000000
1!
b10 %
1'
b10 +
#346280000000
0!
0'
#346290000000
1!
b11 %
1'
b11 +
#346300000000
0!
0'
#346310000000
1!
b100 %
1'
b100 +
#346320000000
0!
0'
#346330000000
1!
b101 %
1'
b101 +
#346340000000
0!
0'
#346350000000
1!
0$
b110 %
1'
0*
b110 +
#346360000000
1"
1(
#346370000000
0!
0"
b100 &
0'
0(
b100 ,
#346380000000
1!
1$
b111 %
1'
1*
b111 +
#346390000000
0!
0'
#346400000000
1!
0$
b1000 %
1'
0*
b1000 +
#346410000000
0!
0'
#346420000000
1!
b1001 %
1'
b1001 +
#346430000000
0!
0'
#346440000000
1!
b0 %
1'
b0 +
#346450000000
0!
0'
#346460000000
1!
1$
b1 %
1'
1*
b1 +
#346470000000
0!
0'
#346480000000
1!
b10 %
1'
b10 +
#346490000000
0!
0'
#346500000000
1!
b11 %
1'
b11 +
#346510000000
0!
0'
#346520000000
1!
b100 %
1'
b100 +
#346530000000
0!
0'
#346540000000
1!
b101 %
1'
b101 +
#346550000000
0!
0'
#346560000000
1!
b110 %
1'
b110 +
#346570000000
0!
0'
#346580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#346590000000
0!
0'
#346600000000
1!
b1000 %
1'
b1000 +
#346610000000
0!
0'
#346620000000
1!
b1001 %
1'
b1001 +
#346630000000
0!
0'
#346640000000
1!
b0 %
1'
b0 +
#346650000000
0!
0'
#346660000000
1!
1$
b1 %
1'
1*
b1 +
#346670000000
0!
0'
#346680000000
1!
b10 %
1'
b10 +
#346690000000
0!
0'
#346700000000
1!
b11 %
1'
b11 +
#346710000000
0!
0'
#346720000000
1!
b100 %
1'
b100 +
#346730000000
0!
0'
#346740000000
1!
b101 %
1'
b101 +
#346750000000
0!
0'
#346760000000
1!
0$
b110 %
1'
0*
b110 +
#346770000000
0!
0'
#346780000000
1!
b111 %
1'
b111 +
#346790000000
1"
1(
#346800000000
0!
0"
b100 &
0'
0(
b100 ,
#346810000000
1!
b1000 %
1'
b1000 +
#346820000000
0!
0'
#346830000000
1!
b1001 %
1'
b1001 +
#346840000000
0!
0'
#346850000000
1!
b0 %
1'
b0 +
#346860000000
0!
0'
#346870000000
1!
1$
b1 %
1'
1*
b1 +
#346880000000
0!
0'
#346890000000
1!
b10 %
1'
b10 +
#346900000000
0!
0'
#346910000000
1!
b11 %
1'
b11 +
#346920000000
0!
0'
#346930000000
1!
b100 %
1'
b100 +
#346940000000
0!
0'
#346950000000
1!
b101 %
1'
b101 +
#346960000000
0!
0'
#346970000000
1!
b110 %
1'
b110 +
#346980000000
0!
0'
#346990000000
1!
b111 %
1'
b111 +
#347000000000
0!
0'
#347010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#347020000000
0!
0'
#347030000000
1!
b1001 %
1'
b1001 +
#347040000000
0!
0'
#347050000000
1!
b0 %
1'
b0 +
#347060000000
0!
0'
#347070000000
1!
1$
b1 %
1'
1*
b1 +
#347080000000
0!
0'
#347090000000
1!
b10 %
1'
b10 +
#347100000000
0!
0'
#347110000000
1!
b11 %
1'
b11 +
#347120000000
0!
0'
#347130000000
1!
b100 %
1'
b100 +
#347140000000
0!
0'
#347150000000
1!
b101 %
1'
b101 +
#347160000000
0!
0'
#347170000000
1!
0$
b110 %
1'
0*
b110 +
#347180000000
0!
0'
#347190000000
1!
b111 %
1'
b111 +
#347200000000
0!
0'
#347210000000
1!
b1000 %
1'
b1000 +
#347220000000
1"
1(
#347230000000
0!
0"
b100 &
0'
0(
b100 ,
#347240000000
1!
b1001 %
1'
b1001 +
#347250000000
0!
0'
#347260000000
1!
b0 %
1'
b0 +
#347270000000
0!
0'
#347280000000
1!
1$
b1 %
1'
1*
b1 +
#347290000000
0!
0'
#347300000000
1!
b10 %
1'
b10 +
#347310000000
0!
0'
#347320000000
1!
b11 %
1'
b11 +
#347330000000
0!
0'
#347340000000
1!
b100 %
1'
b100 +
#347350000000
0!
0'
#347360000000
1!
b101 %
1'
b101 +
#347370000000
0!
0'
#347380000000
1!
b110 %
1'
b110 +
#347390000000
0!
0'
#347400000000
1!
b111 %
1'
b111 +
#347410000000
0!
0'
#347420000000
1!
0$
b1000 %
1'
0*
b1000 +
#347430000000
0!
0'
#347440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#347450000000
0!
0'
#347460000000
1!
b0 %
1'
b0 +
#347470000000
0!
0'
#347480000000
1!
1$
b1 %
1'
1*
b1 +
#347490000000
0!
0'
#347500000000
1!
b10 %
1'
b10 +
#347510000000
0!
0'
#347520000000
1!
b11 %
1'
b11 +
#347530000000
0!
0'
#347540000000
1!
b100 %
1'
b100 +
#347550000000
0!
0'
#347560000000
1!
b101 %
1'
b101 +
#347570000000
0!
0'
#347580000000
1!
0$
b110 %
1'
0*
b110 +
#347590000000
0!
0'
#347600000000
1!
b111 %
1'
b111 +
#347610000000
0!
0'
#347620000000
1!
b1000 %
1'
b1000 +
#347630000000
0!
0'
#347640000000
1!
b1001 %
1'
b1001 +
#347650000000
1"
1(
#347660000000
0!
0"
b100 &
0'
0(
b100 ,
#347670000000
1!
b0 %
1'
b0 +
#347680000000
0!
0'
#347690000000
1!
1$
b1 %
1'
1*
b1 +
#347700000000
0!
0'
#347710000000
1!
b10 %
1'
b10 +
#347720000000
0!
0'
#347730000000
1!
b11 %
1'
b11 +
#347740000000
0!
0'
#347750000000
1!
b100 %
1'
b100 +
#347760000000
0!
0'
#347770000000
1!
b101 %
1'
b101 +
#347780000000
0!
0'
#347790000000
1!
b110 %
1'
b110 +
#347800000000
0!
0'
#347810000000
1!
b111 %
1'
b111 +
#347820000000
0!
0'
#347830000000
1!
0$
b1000 %
1'
0*
b1000 +
#347840000000
0!
0'
#347850000000
1!
b1001 %
1'
b1001 +
#347860000000
0!
0'
#347870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#347880000000
0!
0'
#347890000000
1!
1$
b1 %
1'
1*
b1 +
#347900000000
0!
0'
#347910000000
1!
b10 %
1'
b10 +
#347920000000
0!
0'
#347930000000
1!
b11 %
1'
b11 +
#347940000000
0!
0'
#347950000000
1!
b100 %
1'
b100 +
#347960000000
0!
0'
#347970000000
1!
b101 %
1'
b101 +
#347980000000
0!
0'
#347990000000
1!
0$
b110 %
1'
0*
b110 +
#348000000000
0!
0'
#348010000000
1!
b111 %
1'
b111 +
#348020000000
0!
0'
#348030000000
1!
b1000 %
1'
b1000 +
#348040000000
0!
0'
#348050000000
1!
b1001 %
1'
b1001 +
#348060000000
0!
0'
#348070000000
1!
b0 %
1'
b0 +
#348080000000
1"
1(
#348090000000
0!
0"
b100 &
0'
0(
b100 ,
#348100000000
1!
1$
b1 %
1'
1*
b1 +
#348110000000
0!
0'
#348120000000
1!
b10 %
1'
b10 +
#348130000000
0!
0'
#348140000000
1!
b11 %
1'
b11 +
#348150000000
0!
0'
#348160000000
1!
b100 %
1'
b100 +
#348170000000
0!
0'
#348180000000
1!
b101 %
1'
b101 +
#348190000000
0!
0'
#348200000000
1!
b110 %
1'
b110 +
#348210000000
0!
0'
#348220000000
1!
b111 %
1'
b111 +
#348230000000
0!
0'
#348240000000
1!
0$
b1000 %
1'
0*
b1000 +
#348250000000
0!
0'
#348260000000
1!
b1001 %
1'
b1001 +
#348270000000
0!
0'
#348280000000
1!
b0 %
1'
b0 +
#348290000000
0!
0'
#348300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#348310000000
0!
0'
#348320000000
1!
b10 %
1'
b10 +
#348330000000
0!
0'
#348340000000
1!
b11 %
1'
b11 +
#348350000000
0!
0'
#348360000000
1!
b100 %
1'
b100 +
#348370000000
0!
0'
#348380000000
1!
b101 %
1'
b101 +
#348390000000
0!
0'
#348400000000
1!
0$
b110 %
1'
0*
b110 +
#348410000000
0!
0'
#348420000000
1!
b111 %
1'
b111 +
#348430000000
0!
0'
#348440000000
1!
b1000 %
1'
b1000 +
#348450000000
0!
0'
#348460000000
1!
b1001 %
1'
b1001 +
#348470000000
0!
0'
#348480000000
1!
b0 %
1'
b0 +
#348490000000
0!
0'
#348500000000
1!
1$
b1 %
1'
1*
b1 +
#348510000000
1"
1(
#348520000000
0!
0"
b100 &
0'
0(
b100 ,
#348530000000
1!
b10 %
1'
b10 +
#348540000000
0!
0'
#348550000000
1!
b11 %
1'
b11 +
#348560000000
0!
0'
#348570000000
1!
b100 %
1'
b100 +
#348580000000
0!
0'
#348590000000
1!
b101 %
1'
b101 +
#348600000000
0!
0'
#348610000000
1!
b110 %
1'
b110 +
#348620000000
0!
0'
#348630000000
1!
b111 %
1'
b111 +
#348640000000
0!
0'
#348650000000
1!
0$
b1000 %
1'
0*
b1000 +
#348660000000
0!
0'
#348670000000
1!
b1001 %
1'
b1001 +
#348680000000
0!
0'
#348690000000
1!
b0 %
1'
b0 +
#348700000000
0!
0'
#348710000000
1!
1$
b1 %
1'
1*
b1 +
#348720000000
0!
0'
#348730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#348740000000
0!
0'
#348750000000
1!
b11 %
1'
b11 +
#348760000000
0!
0'
#348770000000
1!
b100 %
1'
b100 +
#348780000000
0!
0'
#348790000000
1!
b101 %
1'
b101 +
#348800000000
0!
0'
#348810000000
1!
0$
b110 %
1'
0*
b110 +
#348820000000
0!
0'
#348830000000
1!
b111 %
1'
b111 +
#348840000000
0!
0'
#348850000000
1!
b1000 %
1'
b1000 +
#348860000000
0!
0'
#348870000000
1!
b1001 %
1'
b1001 +
#348880000000
0!
0'
#348890000000
1!
b0 %
1'
b0 +
#348900000000
0!
0'
#348910000000
1!
1$
b1 %
1'
1*
b1 +
#348920000000
0!
0'
#348930000000
1!
b10 %
1'
b10 +
#348940000000
1"
1(
#348950000000
0!
0"
b100 &
0'
0(
b100 ,
#348960000000
1!
b11 %
1'
b11 +
#348970000000
0!
0'
#348980000000
1!
b100 %
1'
b100 +
#348990000000
0!
0'
#349000000000
1!
b101 %
1'
b101 +
#349010000000
0!
0'
#349020000000
1!
b110 %
1'
b110 +
#349030000000
0!
0'
#349040000000
1!
b111 %
1'
b111 +
#349050000000
0!
0'
#349060000000
1!
0$
b1000 %
1'
0*
b1000 +
#349070000000
0!
0'
#349080000000
1!
b1001 %
1'
b1001 +
#349090000000
0!
0'
#349100000000
1!
b0 %
1'
b0 +
#349110000000
0!
0'
#349120000000
1!
1$
b1 %
1'
1*
b1 +
#349130000000
0!
0'
#349140000000
1!
b10 %
1'
b10 +
#349150000000
0!
0'
#349160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#349170000000
0!
0'
#349180000000
1!
b100 %
1'
b100 +
#349190000000
0!
0'
#349200000000
1!
b101 %
1'
b101 +
#349210000000
0!
0'
#349220000000
1!
0$
b110 %
1'
0*
b110 +
#349230000000
0!
0'
#349240000000
1!
b111 %
1'
b111 +
#349250000000
0!
0'
#349260000000
1!
b1000 %
1'
b1000 +
#349270000000
0!
0'
#349280000000
1!
b1001 %
1'
b1001 +
#349290000000
0!
0'
#349300000000
1!
b0 %
1'
b0 +
#349310000000
0!
0'
#349320000000
1!
1$
b1 %
1'
1*
b1 +
#349330000000
0!
0'
#349340000000
1!
b10 %
1'
b10 +
#349350000000
0!
0'
#349360000000
1!
b11 %
1'
b11 +
#349370000000
1"
1(
#349380000000
0!
0"
b100 &
0'
0(
b100 ,
#349390000000
1!
b100 %
1'
b100 +
#349400000000
0!
0'
#349410000000
1!
b101 %
1'
b101 +
#349420000000
0!
0'
#349430000000
1!
b110 %
1'
b110 +
#349440000000
0!
0'
#349450000000
1!
b111 %
1'
b111 +
#349460000000
0!
0'
#349470000000
1!
0$
b1000 %
1'
0*
b1000 +
#349480000000
0!
0'
#349490000000
1!
b1001 %
1'
b1001 +
#349500000000
0!
0'
#349510000000
1!
b0 %
1'
b0 +
#349520000000
0!
0'
#349530000000
1!
1$
b1 %
1'
1*
b1 +
#349540000000
0!
0'
#349550000000
1!
b10 %
1'
b10 +
#349560000000
0!
0'
#349570000000
1!
b11 %
1'
b11 +
#349580000000
0!
0'
#349590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#349600000000
0!
0'
#349610000000
1!
b101 %
1'
b101 +
#349620000000
0!
0'
#349630000000
1!
0$
b110 %
1'
0*
b110 +
#349640000000
0!
0'
#349650000000
1!
b111 %
1'
b111 +
#349660000000
0!
0'
#349670000000
1!
b1000 %
1'
b1000 +
#349680000000
0!
0'
#349690000000
1!
b1001 %
1'
b1001 +
#349700000000
0!
0'
#349710000000
1!
b0 %
1'
b0 +
#349720000000
0!
0'
#349730000000
1!
1$
b1 %
1'
1*
b1 +
#349740000000
0!
0'
#349750000000
1!
b10 %
1'
b10 +
#349760000000
0!
0'
#349770000000
1!
b11 %
1'
b11 +
#349780000000
0!
0'
#349790000000
1!
b100 %
1'
b100 +
#349800000000
1"
1(
#349810000000
0!
0"
b100 &
0'
0(
b100 ,
#349820000000
1!
b101 %
1'
b101 +
#349830000000
0!
0'
#349840000000
1!
b110 %
1'
b110 +
#349850000000
0!
0'
#349860000000
1!
b111 %
1'
b111 +
#349870000000
0!
0'
#349880000000
1!
0$
b1000 %
1'
0*
b1000 +
#349890000000
0!
0'
#349900000000
1!
b1001 %
1'
b1001 +
#349910000000
0!
0'
#349920000000
1!
b0 %
1'
b0 +
#349930000000
0!
0'
#349940000000
1!
1$
b1 %
1'
1*
b1 +
#349950000000
0!
0'
#349960000000
1!
b10 %
1'
b10 +
#349970000000
0!
0'
#349980000000
1!
b11 %
1'
b11 +
#349990000000
0!
0'
#350000000000
1!
b100 %
1'
b100 +
#350010000000
0!
0'
#350020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#350030000000
0!
0'
#350040000000
1!
0$
b110 %
1'
0*
b110 +
#350050000000
0!
0'
#350060000000
1!
b111 %
1'
b111 +
#350070000000
0!
0'
#350080000000
1!
b1000 %
1'
b1000 +
#350090000000
0!
0'
#350100000000
1!
b1001 %
1'
b1001 +
#350110000000
0!
0'
#350120000000
1!
b0 %
1'
b0 +
#350130000000
0!
0'
#350140000000
1!
1$
b1 %
1'
1*
b1 +
#350150000000
0!
0'
#350160000000
1!
b10 %
1'
b10 +
#350170000000
0!
0'
#350180000000
1!
b11 %
1'
b11 +
#350190000000
0!
0'
#350200000000
1!
b100 %
1'
b100 +
#350210000000
0!
0'
#350220000000
1!
b101 %
1'
b101 +
#350230000000
1"
1(
#350240000000
0!
0"
b100 &
0'
0(
b100 ,
#350250000000
1!
b110 %
1'
b110 +
#350260000000
0!
0'
#350270000000
1!
b111 %
1'
b111 +
#350280000000
0!
0'
#350290000000
1!
0$
b1000 %
1'
0*
b1000 +
#350300000000
0!
0'
#350310000000
1!
b1001 %
1'
b1001 +
#350320000000
0!
0'
#350330000000
1!
b0 %
1'
b0 +
#350340000000
0!
0'
#350350000000
1!
1$
b1 %
1'
1*
b1 +
#350360000000
0!
0'
#350370000000
1!
b10 %
1'
b10 +
#350380000000
0!
0'
#350390000000
1!
b11 %
1'
b11 +
#350400000000
0!
0'
#350410000000
1!
b100 %
1'
b100 +
#350420000000
0!
0'
#350430000000
1!
b101 %
1'
b101 +
#350440000000
0!
0'
#350450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#350460000000
0!
0'
#350470000000
1!
b111 %
1'
b111 +
#350480000000
0!
0'
#350490000000
1!
b1000 %
1'
b1000 +
#350500000000
0!
0'
#350510000000
1!
b1001 %
1'
b1001 +
#350520000000
0!
0'
#350530000000
1!
b0 %
1'
b0 +
#350540000000
0!
0'
#350550000000
1!
1$
b1 %
1'
1*
b1 +
#350560000000
0!
0'
#350570000000
1!
b10 %
1'
b10 +
#350580000000
0!
0'
#350590000000
1!
b11 %
1'
b11 +
#350600000000
0!
0'
#350610000000
1!
b100 %
1'
b100 +
#350620000000
0!
0'
#350630000000
1!
b101 %
1'
b101 +
#350640000000
0!
0'
#350650000000
1!
0$
b110 %
1'
0*
b110 +
#350660000000
1"
1(
#350670000000
0!
0"
b100 &
0'
0(
b100 ,
#350680000000
1!
1$
b111 %
1'
1*
b111 +
#350690000000
0!
0'
#350700000000
1!
0$
b1000 %
1'
0*
b1000 +
#350710000000
0!
0'
#350720000000
1!
b1001 %
1'
b1001 +
#350730000000
0!
0'
#350740000000
1!
b0 %
1'
b0 +
#350750000000
0!
0'
#350760000000
1!
1$
b1 %
1'
1*
b1 +
#350770000000
0!
0'
#350780000000
1!
b10 %
1'
b10 +
#350790000000
0!
0'
#350800000000
1!
b11 %
1'
b11 +
#350810000000
0!
0'
#350820000000
1!
b100 %
1'
b100 +
#350830000000
0!
0'
#350840000000
1!
b101 %
1'
b101 +
#350850000000
0!
0'
#350860000000
1!
b110 %
1'
b110 +
#350870000000
0!
0'
#350880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#350890000000
0!
0'
#350900000000
1!
b1000 %
1'
b1000 +
#350910000000
0!
0'
#350920000000
1!
b1001 %
1'
b1001 +
#350930000000
0!
0'
#350940000000
1!
b0 %
1'
b0 +
#350950000000
0!
0'
#350960000000
1!
1$
b1 %
1'
1*
b1 +
#350970000000
0!
0'
#350980000000
1!
b10 %
1'
b10 +
#350990000000
0!
0'
#351000000000
1!
b11 %
1'
b11 +
#351010000000
0!
0'
#351020000000
1!
b100 %
1'
b100 +
#351030000000
0!
0'
#351040000000
1!
b101 %
1'
b101 +
#351050000000
0!
0'
#351060000000
1!
0$
b110 %
1'
0*
b110 +
#351070000000
0!
0'
#351080000000
1!
b111 %
1'
b111 +
#351090000000
1"
1(
#351100000000
0!
0"
b100 &
0'
0(
b100 ,
#351110000000
1!
b1000 %
1'
b1000 +
#351120000000
0!
0'
#351130000000
1!
b1001 %
1'
b1001 +
#351140000000
0!
0'
#351150000000
1!
b0 %
1'
b0 +
#351160000000
0!
0'
#351170000000
1!
1$
b1 %
1'
1*
b1 +
#351180000000
0!
0'
#351190000000
1!
b10 %
1'
b10 +
#351200000000
0!
0'
#351210000000
1!
b11 %
1'
b11 +
#351220000000
0!
0'
#351230000000
1!
b100 %
1'
b100 +
#351240000000
0!
0'
#351250000000
1!
b101 %
1'
b101 +
#351260000000
0!
0'
#351270000000
1!
b110 %
1'
b110 +
#351280000000
0!
0'
#351290000000
1!
b111 %
1'
b111 +
#351300000000
0!
0'
#351310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#351320000000
0!
0'
#351330000000
1!
b1001 %
1'
b1001 +
#351340000000
0!
0'
#351350000000
1!
b0 %
1'
b0 +
#351360000000
0!
0'
#351370000000
1!
1$
b1 %
1'
1*
b1 +
#351380000000
0!
0'
#351390000000
1!
b10 %
1'
b10 +
#351400000000
0!
0'
#351410000000
1!
b11 %
1'
b11 +
#351420000000
0!
0'
#351430000000
1!
b100 %
1'
b100 +
#351440000000
0!
0'
#351450000000
1!
b101 %
1'
b101 +
#351460000000
0!
0'
#351470000000
1!
0$
b110 %
1'
0*
b110 +
#351480000000
0!
0'
#351490000000
1!
b111 %
1'
b111 +
#351500000000
0!
0'
#351510000000
1!
b1000 %
1'
b1000 +
#351520000000
1"
1(
#351530000000
0!
0"
b100 &
0'
0(
b100 ,
#351540000000
1!
b1001 %
1'
b1001 +
#351550000000
0!
0'
#351560000000
1!
b0 %
1'
b0 +
#351570000000
0!
0'
#351580000000
1!
1$
b1 %
1'
1*
b1 +
#351590000000
0!
0'
#351600000000
1!
b10 %
1'
b10 +
#351610000000
0!
0'
#351620000000
1!
b11 %
1'
b11 +
#351630000000
0!
0'
#351640000000
1!
b100 %
1'
b100 +
#351650000000
0!
0'
#351660000000
1!
b101 %
1'
b101 +
#351670000000
0!
0'
#351680000000
1!
b110 %
1'
b110 +
#351690000000
0!
0'
#351700000000
1!
b111 %
1'
b111 +
#351710000000
0!
0'
#351720000000
1!
0$
b1000 %
1'
0*
b1000 +
#351730000000
0!
0'
#351740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#351750000000
0!
0'
#351760000000
1!
b0 %
1'
b0 +
#351770000000
0!
0'
#351780000000
1!
1$
b1 %
1'
1*
b1 +
#351790000000
0!
0'
#351800000000
1!
b10 %
1'
b10 +
#351810000000
0!
0'
#351820000000
1!
b11 %
1'
b11 +
#351830000000
0!
0'
#351840000000
1!
b100 %
1'
b100 +
#351850000000
0!
0'
#351860000000
1!
b101 %
1'
b101 +
#351870000000
0!
0'
#351880000000
1!
0$
b110 %
1'
0*
b110 +
#351890000000
0!
0'
#351900000000
1!
b111 %
1'
b111 +
#351910000000
0!
0'
#351920000000
1!
b1000 %
1'
b1000 +
#351930000000
0!
0'
#351940000000
1!
b1001 %
1'
b1001 +
#351950000000
1"
1(
#351960000000
0!
0"
b100 &
0'
0(
b100 ,
#351970000000
1!
b0 %
1'
b0 +
#351980000000
0!
0'
#351990000000
1!
1$
b1 %
1'
1*
b1 +
#352000000000
0!
0'
#352010000000
1!
b10 %
1'
b10 +
#352020000000
0!
0'
#352030000000
1!
b11 %
1'
b11 +
#352040000000
0!
0'
#352050000000
1!
b100 %
1'
b100 +
#352060000000
0!
0'
#352070000000
1!
b101 %
1'
b101 +
#352080000000
0!
0'
#352090000000
1!
b110 %
1'
b110 +
#352100000000
0!
0'
#352110000000
1!
b111 %
1'
b111 +
#352120000000
0!
0'
#352130000000
1!
0$
b1000 %
1'
0*
b1000 +
#352140000000
0!
0'
#352150000000
1!
b1001 %
1'
b1001 +
#352160000000
0!
0'
#352170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#352180000000
0!
0'
#352190000000
1!
1$
b1 %
1'
1*
b1 +
#352200000000
0!
0'
#352210000000
1!
b10 %
1'
b10 +
#352220000000
0!
0'
#352230000000
1!
b11 %
1'
b11 +
#352240000000
0!
0'
#352250000000
1!
b100 %
1'
b100 +
#352260000000
0!
0'
#352270000000
1!
b101 %
1'
b101 +
#352280000000
0!
0'
#352290000000
1!
0$
b110 %
1'
0*
b110 +
#352300000000
0!
0'
#352310000000
1!
b111 %
1'
b111 +
#352320000000
0!
0'
#352330000000
1!
b1000 %
1'
b1000 +
#352340000000
0!
0'
#352350000000
1!
b1001 %
1'
b1001 +
#352360000000
0!
0'
#352370000000
1!
b0 %
1'
b0 +
#352380000000
1"
1(
#352390000000
0!
0"
b100 &
0'
0(
b100 ,
#352400000000
1!
1$
b1 %
1'
1*
b1 +
#352410000000
0!
0'
#352420000000
1!
b10 %
1'
b10 +
#352430000000
0!
0'
#352440000000
1!
b11 %
1'
b11 +
#352450000000
0!
0'
#352460000000
1!
b100 %
1'
b100 +
#352470000000
0!
0'
#352480000000
1!
b101 %
1'
b101 +
#352490000000
0!
0'
#352500000000
1!
b110 %
1'
b110 +
#352510000000
0!
0'
#352520000000
1!
b111 %
1'
b111 +
#352530000000
0!
0'
#352540000000
1!
0$
b1000 %
1'
0*
b1000 +
#352550000000
0!
0'
#352560000000
1!
b1001 %
1'
b1001 +
#352570000000
0!
0'
#352580000000
1!
b0 %
1'
b0 +
#352590000000
0!
0'
#352600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#352610000000
0!
0'
#352620000000
1!
b10 %
1'
b10 +
#352630000000
0!
0'
#352640000000
1!
b11 %
1'
b11 +
#352650000000
0!
0'
#352660000000
1!
b100 %
1'
b100 +
#352670000000
0!
0'
#352680000000
1!
b101 %
1'
b101 +
#352690000000
0!
0'
#352700000000
1!
0$
b110 %
1'
0*
b110 +
#352710000000
0!
0'
#352720000000
1!
b111 %
1'
b111 +
#352730000000
0!
0'
#352740000000
1!
b1000 %
1'
b1000 +
#352750000000
0!
0'
#352760000000
1!
b1001 %
1'
b1001 +
#352770000000
0!
0'
#352780000000
1!
b0 %
1'
b0 +
#352790000000
0!
0'
#352800000000
1!
1$
b1 %
1'
1*
b1 +
#352810000000
1"
1(
#352820000000
0!
0"
b100 &
0'
0(
b100 ,
#352830000000
1!
b10 %
1'
b10 +
#352840000000
0!
0'
#352850000000
1!
b11 %
1'
b11 +
#352860000000
0!
0'
#352870000000
1!
b100 %
1'
b100 +
#352880000000
0!
0'
#352890000000
1!
b101 %
1'
b101 +
#352900000000
0!
0'
#352910000000
1!
b110 %
1'
b110 +
#352920000000
0!
0'
#352930000000
1!
b111 %
1'
b111 +
#352940000000
0!
0'
#352950000000
1!
0$
b1000 %
1'
0*
b1000 +
#352960000000
0!
0'
#352970000000
1!
b1001 %
1'
b1001 +
#352980000000
0!
0'
#352990000000
1!
b0 %
1'
b0 +
#353000000000
0!
0'
#353010000000
1!
1$
b1 %
1'
1*
b1 +
#353020000000
0!
0'
#353030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#353040000000
0!
0'
#353050000000
1!
b11 %
1'
b11 +
#353060000000
0!
0'
#353070000000
1!
b100 %
1'
b100 +
#353080000000
0!
0'
#353090000000
1!
b101 %
1'
b101 +
#353100000000
0!
0'
#353110000000
1!
0$
b110 %
1'
0*
b110 +
#353120000000
0!
0'
#353130000000
1!
b111 %
1'
b111 +
#353140000000
0!
0'
#353150000000
1!
b1000 %
1'
b1000 +
#353160000000
0!
0'
#353170000000
1!
b1001 %
1'
b1001 +
#353180000000
0!
0'
#353190000000
1!
b0 %
1'
b0 +
#353200000000
0!
0'
#353210000000
1!
1$
b1 %
1'
1*
b1 +
#353220000000
0!
0'
#353230000000
1!
b10 %
1'
b10 +
#353240000000
1"
1(
#353250000000
0!
0"
b100 &
0'
0(
b100 ,
#353260000000
1!
b11 %
1'
b11 +
#353270000000
0!
0'
#353280000000
1!
b100 %
1'
b100 +
#353290000000
0!
0'
#353300000000
1!
b101 %
1'
b101 +
#353310000000
0!
0'
#353320000000
1!
b110 %
1'
b110 +
#353330000000
0!
0'
#353340000000
1!
b111 %
1'
b111 +
#353350000000
0!
0'
#353360000000
1!
0$
b1000 %
1'
0*
b1000 +
#353370000000
0!
0'
#353380000000
1!
b1001 %
1'
b1001 +
#353390000000
0!
0'
#353400000000
1!
b0 %
1'
b0 +
#353410000000
0!
0'
#353420000000
1!
1$
b1 %
1'
1*
b1 +
#353430000000
0!
0'
#353440000000
1!
b10 %
1'
b10 +
#353450000000
0!
0'
#353460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#353470000000
0!
0'
#353480000000
1!
b100 %
1'
b100 +
#353490000000
0!
0'
#353500000000
1!
b101 %
1'
b101 +
#353510000000
0!
0'
#353520000000
1!
0$
b110 %
1'
0*
b110 +
#353530000000
0!
0'
#353540000000
1!
b111 %
1'
b111 +
#353550000000
0!
0'
#353560000000
1!
b1000 %
1'
b1000 +
#353570000000
0!
0'
#353580000000
1!
b1001 %
1'
b1001 +
#353590000000
0!
0'
#353600000000
1!
b0 %
1'
b0 +
#353610000000
0!
0'
#353620000000
1!
1$
b1 %
1'
1*
b1 +
#353630000000
0!
0'
#353640000000
1!
b10 %
1'
b10 +
#353650000000
0!
0'
#353660000000
1!
b11 %
1'
b11 +
#353670000000
1"
1(
#353680000000
0!
0"
b100 &
0'
0(
b100 ,
#353690000000
1!
b100 %
1'
b100 +
#353700000000
0!
0'
#353710000000
1!
b101 %
1'
b101 +
#353720000000
0!
0'
#353730000000
1!
b110 %
1'
b110 +
#353740000000
0!
0'
#353750000000
1!
b111 %
1'
b111 +
#353760000000
0!
0'
#353770000000
1!
0$
b1000 %
1'
0*
b1000 +
#353780000000
0!
0'
#353790000000
1!
b1001 %
1'
b1001 +
#353800000000
0!
0'
#353810000000
1!
b0 %
1'
b0 +
#353820000000
0!
0'
#353830000000
1!
1$
b1 %
1'
1*
b1 +
#353840000000
0!
0'
#353850000000
1!
b10 %
1'
b10 +
#353860000000
0!
0'
#353870000000
1!
b11 %
1'
b11 +
#353880000000
0!
0'
#353890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#353900000000
0!
0'
#353910000000
1!
b101 %
1'
b101 +
#353920000000
0!
0'
#353930000000
1!
0$
b110 %
1'
0*
b110 +
#353940000000
0!
0'
#353950000000
1!
b111 %
1'
b111 +
#353960000000
0!
0'
#353970000000
1!
b1000 %
1'
b1000 +
#353980000000
0!
0'
#353990000000
1!
b1001 %
1'
b1001 +
#354000000000
0!
0'
#354010000000
1!
b0 %
1'
b0 +
#354020000000
0!
0'
#354030000000
1!
1$
b1 %
1'
1*
b1 +
#354040000000
0!
0'
#354050000000
1!
b10 %
1'
b10 +
#354060000000
0!
0'
#354070000000
1!
b11 %
1'
b11 +
#354080000000
0!
0'
#354090000000
1!
b100 %
1'
b100 +
#354100000000
1"
1(
#354110000000
0!
0"
b100 &
0'
0(
b100 ,
#354120000000
1!
b101 %
1'
b101 +
#354130000000
0!
0'
#354140000000
1!
b110 %
1'
b110 +
#354150000000
0!
0'
#354160000000
1!
b111 %
1'
b111 +
#354170000000
0!
0'
#354180000000
1!
0$
b1000 %
1'
0*
b1000 +
#354190000000
0!
0'
#354200000000
1!
b1001 %
1'
b1001 +
#354210000000
0!
0'
#354220000000
1!
b0 %
1'
b0 +
#354230000000
0!
0'
#354240000000
1!
1$
b1 %
1'
1*
b1 +
#354250000000
0!
0'
#354260000000
1!
b10 %
1'
b10 +
#354270000000
0!
0'
#354280000000
1!
b11 %
1'
b11 +
#354290000000
0!
0'
#354300000000
1!
b100 %
1'
b100 +
#354310000000
0!
0'
#354320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#354330000000
0!
0'
#354340000000
1!
0$
b110 %
1'
0*
b110 +
#354350000000
0!
0'
#354360000000
1!
b111 %
1'
b111 +
#354370000000
0!
0'
#354380000000
1!
b1000 %
1'
b1000 +
#354390000000
0!
0'
#354400000000
1!
b1001 %
1'
b1001 +
#354410000000
0!
0'
#354420000000
1!
b0 %
1'
b0 +
#354430000000
0!
0'
#354440000000
1!
1$
b1 %
1'
1*
b1 +
#354450000000
0!
0'
#354460000000
1!
b10 %
1'
b10 +
#354470000000
0!
0'
#354480000000
1!
b11 %
1'
b11 +
#354490000000
0!
0'
#354500000000
1!
b100 %
1'
b100 +
#354510000000
0!
0'
#354520000000
1!
b101 %
1'
b101 +
#354530000000
1"
1(
#354540000000
0!
0"
b100 &
0'
0(
b100 ,
#354550000000
1!
b110 %
1'
b110 +
#354560000000
0!
0'
#354570000000
1!
b111 %
1'
b111 +
#354580000000
0!
0'
#354590000000
1!
0$
b1000 %
1'
0*
b1000 +
#354600000000
0!
0'
#354610000000
1!
b1001 %
1'
b1001 +
#354620000000
0!
0'
#354630000000
1!
b0 %
1'
b0 +
#354640000000
0!
0'
#354650000000
1!
1$
b1 %
1'
1*
b1 +
#354660000000
0!
0'
#354670000000
1!
b10 %
1'
b10 +
#354680000000
0!
0'
#354690000000
1!
b11 %
1'
b11 +
#354700000000
0!
0'
#354710000000
1!
b100 %
1'
b100 +
#354720000000
0!
0'
#354730000000
1!
b101 %
1'
b101 +
#354740000000
0!
0'
#354750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#354760000000
0!
0'
#354770000000
1!
b111 %
1'
b111 +
#354780000000
0!
0'
#354790000000
1!
b1000 %
1'
b1000 +
#354800000000
0!
0'
#354810000000
1!
b1001 %
1'
b1001 +
#354820000000
0!
0'
#354830000000
1!
b0 %
1'
b0 +
#354840000000
0!
0'
#354850000000
1!
1$
b1 %
1'
1*
b1 +
#354860000000
0!
0'
#354870000000
1!
b10 %
1'
b10 +
#354880000000
0!
0'
#354890000000
1!
b11 %
1'
b11 +
#354900000000
0!
0'
#354910000000
1!
b100 %
1'
b100 +
#354920000000
0!
0'
#354930000000
1!
b101 %
1'
b101 +
#354940000000
0!
0'
#354950000000
1!
0$
b110 %
1'
0*
b110 +
#354960000000
1"
1(
#354970000000
0!
0"
b100 &
0'
0(
b100 ,
#354980000000
1!
1$
b111 %
1'
1*
b111 +
#354990000000
0!
0'
#355000000000
1!
0$
b1000 %
1'
0*
b1000 +
#355010000000
0!
0'
#355020000000
1!
b1001 %
1'
b1001 +
#355030000000
0!
0'
#355040000000
1!
b0 %
1'
b0 +
#355050000000
0!
0'
#355060000000
1!
1$
b1 %
1'
1*
b1 +
#355070000000
0!
0'
#355080000000
1!
b10 %
1'
b10 +
#355090000000
0!
0'
#355100000000
1!
b11 %
1'
b11 +
#355110000000
0!
0'
#355120000000
1!
b100 %
1'
b100 +
#355130000000
0!
0'
#355140000000
1!
b101 %
1'
b101 +
#355150000000
0!
0'
#355160000000
1!
b110 %
1'
b110 +
#355170000000
0!
0'
#355180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#355190000000
0!
0'
#355200000000
1!
b1000 %
1'
b1000 +
#355210000000
0!
0'
#355220000000
1!
b1001 %
1'
b1001 +
#355230000000
0!
0'
#355240000000
1!
b0 %
1'
b0 +
#355250000000
0!
0'
#355260000000
1!
1$
b1 %
1'
1*
b1 +
#355270000000
0!
0'
#355280000000
1!
b10 %
1'
b10 +
#355290000000
0!
0'
#355300000000
1!
b11 %
1'
b11 +
#355310000000
0!
0'
#355320000000
1!
b100 %
1'
b100 +
#355330000000
0!
0'
#355340000000
1!
b101 %
1'
b101 +
#355350000000
0!
0'
#355360000000
1!
0$
b110 %
1'
0*
b110 +
#355370000000
0!
0'
#355380000000
1!
b111 %
1'
b111 +
#355390000000
1"
1(
#355400000000
0!
0"
b100 &
0'
0(
b100 ,
#355410000000
1!
b1000 %
1'
b1000 +
#355420000000
0!
0'
#355430000000
1!
b1001 %
1'
b1001 +
#355440000000
0!
0'
#355450000000
1!
b0 %
1'
b0 +
#355460000000
0!
0'
#355470000000
1!
1$
b1 %
1'
1*
b1 +
#355480000000
0!
0'
#355490000000
1!
b10 %
1'
b10 +
#355500000000
0!
0'
#355510000000
1!
b11 %
1'
b11 +
#355520000000
0!
0'
#355530000000
1!
b100 %
1'
b100 +
#355540000000
0!
0'
#355550000000
1!
b101 %
1'
b101 +
#355560000000
0!
0'
#355570000000
1!
b110 %
1'
b110 +
#355580000000
0!
0'
#355590000000
1!
b111 %
1'
b111 +
#355600000000
0!
0'
#355610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#355620000000
0!
0'
#355630000000
1!
b1001 %
1'
b1001 +
#355640000000
0!
0'
#355650000000
1!
b0 %
1'
b0 +
#355660000000
0!
0'
#355670000000
1!
1$
b1 %
1'
1*
b1 +
#355680000000
0!
0'
#355690000000
1!
b10 %
1'
b10 +
#355700000000
0!
0'
#355710000000
1!
b11 %
1'
b11 +
#355720000000
0!
0'
#355730000000
1!
b100 %
1'
b100 +
#355740000000
0!
0'
#355750000000
1!
b101 %
1'
b101 +
#355760000000
0!
0'
#355770000000
1!
0$
b110 %
1'
0*
b110 +
#355780000000
0!
0'
#355790000000
1!
b111 %
1'
b111 +
#355800000000
0!
0'
#355810000000
1!
b1000 %
1'
b1000 +
#355820000000
1"
1(
#355830000000
0!
0"
b100 &
0'
0(
b100 ,
#355840000000
1!
b1001 %
1'
b1001 +
#355850000000
0!
0'
#355860000000
1!
b0 %
1'
b0 +
#355870000000
0!
0'
#355880000000
1!
1$
b1 %
1'
1*
b1 +
#355890000000
0!
0'
#355900000000
1!
b10 %
1'
b10 +
#355910000000
0!
0'
#355920000000
1!
b11 %
1'
b11 +
#355930000000
0!
0'
#355940000000
1!
b100 %
1'
b100 +
#355950000000
0!
0'
#355960000000
1!
b101 %
1'
b101 +
#355970000000
0!
0'
#355980000000
1!
b110 %
1'
b110 +
#355990000000
0!
0'
#356000000000
1!
b111 %
1'
b111 +
#356010000000
0!
0'
#356020000000
1!
0$
b1000 %
1'
0*
b1000 +
#356030000000
0!
0'
#356040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#356050000000
0!
0'
#356060000000
1!
b0 %
1'
b0 +
#356070000000
0!
0'
#356080000000
1!
1$
b1 %
1'
1*
b1 +
#356090000000
0!
0'
#356100000000
1!
b10 %
1'
b10 +
#356110000000
0!
0'
#356120000000
1!
b11 %
1'
b11 +
#356130000000
0!
0'
#356140000000
1!
b100 %
1'
b100 +
#356150000000
0!
0'
#356160000000
1!
b101 %
1'
b101 +
#356170000000
0!
0'
#356180000000
1!
0$
b110 %
1'
0*
b110 +
#356190000000
0!
0'
#356200000000
1!
b111 %
1'
b111 +
#356210000000
0!
0'
#356220000000
1!
b1000 %
1'
b1000 +
#356230000000
0!
0'
#356240000000
1!
b1001 %
1'
b1001 +
#356250000000
1"
1(
#356260000000
0!
0"
b100 &
0'
0(
b100 ,
#356270000000
1!
b0 %
1'
b0 +
#356280000000
0!
0'
#356290000000
1!
1$
b1 %
1'
1*
b1 +
#356300000000
0!
0'
#356310000000
1!
b10 %
1'
b10 +
#356320000000
0!
0'
#356330000000
1!
b11 %
1'
b11 +
#356340000000
0!
0'
#356350000000
1!
b100 %
1'
b100 +
#356360000000
0!
0'
#356370000000
1!
b101 %
1'
b101 +
#356380000000
0!
0'
#356390000000
1!
b110 %
1'
b110 +
#356400000000
0!
0'
#356410000000
1!
b111 %
1'
b111 +
#356420000000
0!
0'
#356430000000
1!
0$
b1000 %
1'
0*
b1000 +
#356440000000
0!
0'
#356450000000
1!
b1001 %
1'
b1001 +
#356460000000
0!
0'
#356470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#356480000000
0!
0'
#356490000000
1!
1$
b1 %
1'
1*
b1 +
#356500000000
0!
0'
#356510000000
1!
b10 %
1'
b10 +
#356520000000
0!
0'
#356530000000
1!
b11 %
1'
b11 +
#356540000000
0!
0'
#356550000000
1!
b100 %
1'
b100 +
#356560000000
0!
0'
#356570000000
1!
b101 %
1'
b101 +
#356580000000
0!
0'
#356590000000
1!
0$
b110 %
1'
0*
b110 +
#356600000000
0!
0'
#356610000000
1!
b111 %
1'
b111 +
#356620000000
0!
0'
#356630000000
1!
b1000 %
1'
b1000 +
#356640000000
0!
0'
#356650000000
1!
b1001 %
1'
b1001 +
#356660000000
0!
0'
#356670000000
1!
b0 %
1'
b0 +
#356680000000
1"
1(
#356690000000
0!
0"
b100 &
0'
0(
b100 ,
#356700000000
1!
1$
b1 %
1'
1*
b1 +
#356710000000
0!
0'
#356720000000
1!
b10 %
1'
b10 +
#356730000000
0!
0'
#356740000000
1!
b11 %
1'
b11 +
#356750000000
0!
0'
#356760000000
1!
b100 %
1'
b100 +
#356770000000
0!
0'
#356780000000
1!
b101 %
1'
b101 +
#356790000000
0!
0'
#356800000000
1!
b110 %
1'
b110 +
#356810000000
0!
0'
#356820000000
1!
b111 %
1'
b111 +
#356830000000
0!
0'
#356840000000
1!
0$
b1000 %
1'
0*
b1000 +
#356850000000
0!
0'
#356860000000
1!
b1001 %
1'
b1001 +
#356870000000
0!
0'
#356880000000
1!
b0 %
1'
b0 +
#356890000000
0!
0'
#356900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#356910000000
0!
0'
#356920000000
1!
b10 %
1'
b10 +
#356930000000
0!
0'
#356940000000
1!
b11 %
1'
b11 +
#356950000000
0!
0'
#356960000000
1!
b100 %
1'
b100 +
#356970000000
0!
0'
#356980000000
1!
b101 %
1'
b101 +
#356990000000
0!
0'
#357000000000
1!
0$
b110 %
1'
0*
b110 +
#357010000000
0!
0'
#357020000000
1!
b111 %
1'
b111 +
#357030000000
0!
0'
#357040000000
1!
b1000 %
1'
b1000 +
#357050000000
0!
0'
#357060000000
1!
b1001 %
1'
b1001 +
#357070000000
0!
0'
#357080000000
1!
b0 %
1'
b0 +
#357090000000
0!
0'
#357100000000
1!
1$
b1 %
1'
1*
b1 +
#357110000000
1"
1(
#357120000000
0!
0"
b100 &
0'
0(
b100 ,
#357130000000
1!
b10 %
1'
b10 +
#357140000000
0!
0'
#357150000000
1!
b11 %
1'
b11 +
#357160000000
0!
0'
#357170000000
1!
b100 %
1'
b100 +
#357180000000
0!
0'
#357190000000
1!
b101 %
1'
b101 +
#357200000000
0!
0'
#357210000000
1!
b110 %
1'
b110 +
#357220000000
0!
0'
#357230000000
1!
b111 %
1'
b111 +
#357240000000
0!
0'
#357250000000
1!
0$
b1000 %
1'
0*
b1000 +
#357260000000
0!
0'
#357270000000
1!
b1001 %
1'
b1001 +
#357280000000
0!
0'
#357290000000
1!
b0 %
1'
b0 +
#357300000000
0!
0'
#357310000000
1!
1$
b1 %
1'
1*
b1 +
#357320000000
0!
0'
#357330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#357340000000
0!
0'
#357350000000
1!
b11 %
1'
b11 +
#357360000000
0!
0'
#357370000000
1!
b100 %
1'
b100 +
#357380000000
0!
0'
#357390000000
1!
b101 %
1'
b101 +
#357400000000
0!
0'
#357410000000
1!
0$
b110 %
1'
0*
b110 +
#357420000000
0!
0'
#357430000000
1!
b111 %
1'
b111 +
#357440000000
0!
0'
#357450000000
1!
b1000 %
1'
b1000 +
#357460000000
0!
0'
#357470000000
1!
b1001 %
1'
b1001 +
#357480000000
0!
0'
#357490000000
1!
b0 %
1'
b0 +
#357500000000
0!
0'
#357510000000
1!
1$
b1 %
1'
1*
b1 +
#357520000000
0!
0'
#357530000000
1!
b10 %
1'
b10 +
#357540000000
1"
1(
#357550000000
0!
0"
b100 &
0'
0(
b100 ,
#357560000000
1!
b11 %
1'
b11 +
#357570000000
0!
0'
#357580000000
1!
b100 %
1'
b100 +
#357590000000
0!
0'
#357600000000
1!
b101 %
1'
b101 +
#357610000000
0!
0'
#357620000000
1!
b110 %
1'
b110 +
#357630000000
0!
0'
#357640000000
1!
b111 %
1'
b111 +
#357650000000
0!
0'
#357660000000
1!
0$
b1000 %
1'
0*
b1000 +
#357670000000
0!
0'
#357680000000
1!
b1001 %
1'
b1001 +
#357690000000
0!
0'
#357700000000
1!
b0 %
1'
b0 +
#357710000000
0!
0'
#357720000000
1!
1$
b1 %
1'
1*
b1 +
#357730000000
0!
0'
#357740000000
1!
b10 %
1'
b10 +
#357750000000
0!
0'
#357760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#357770000000
0!
0'
#357780000000
1!
b100 %
1'
b100 +
#357790000000
0!
0'
#357800000000
1!
b101 %
1'
b101 +
#357810000000
0!
0'
#357820000000
1!
0$
b110 %
1'
0*
b110 +
#357830000000
0!
0'
#357840000000
1!
b111 %
1'
b111 +
#357850000000
0!
0'
#357860000000
1!
b1000 %
1'
b1000 +
#357870000000
0!
0'
#357880000000
1!
b1001 %
1'
b1001 +
#357890000000
0!
0'
#357900000000
1!
b0 %
1'
b0 +
#357910000000
0!
0'
#357920000000
1!
1$
b1 %
1'
1*
b1 +
#357930000000
0!
0'
#357940000000
1!
b10 %
1'
b10 +
#357950000000
0!
0'
#357960000000
1!
b11 %
1'
b11 +
#357970000000
1"
1(
#357980000000
0!
0"
b100 &
0'
0(
b100 ,
#357990000000
1!
b100 %
1'
b100 +
#358000000000
0!
0'
#358010000000
1!
b101 %
1'
b101 +
#358020000000
0!
0'
#358030000000
1!
b110 %
1'
b110 +
#358040000000
0!
0'
#358050000000
1!
b111 %
1'
b111 +
#358060000000
0!
0'
#358070000000
1!
0$
b1000 %
1'
0*
b1000 +
#358080000000
0!
0'
#358090000000
1!
b1001 %
1'
b1001 +
#358100000000
0!
0'
#358110000000
1!
b0 %
1'
b0 +
#358120000000
0!
0'
#358130000000
1!
1$
b1 %
1'
1*
b1 +
#358140000000
0!
0'
#358150000000
1!
b10 %
1'
b10 +
#358160000000
0!
0'
#358170000000
1!
b11 %
1'
b11 +
#358180000000
0!
0'
#358190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#358200000000
0!
0'
#358210000000
1!
b101 %
1'
b101 +
#358220000000
0!
0'
#358230000000
1!
0$
b110 %
1'
0*
b110 +
#358240000000
0!
0'
#358250000000
1!
b111 %
1'
b111 +
#358260000000
0!
0'
#358270000000
1!
b1000 %
1'
b1000 +
#358280000000
0!
0'
#358290000000
1!
b1001 %
1'
b1001 +
#358300000000
0!
0'
#358310000000
1!
b0 %
1'
b0 +
#358320000000
0!
0'
#358330000000
1!
1$
b1 %
1'
1*
b1 +
#358340000000
0!
0'
#358350000000
1!
b10 %
1'
b10 +
#358360000000
0!
0'
#358370000000
1!
b11 %
1'
b11 +
#358380000000
0!
0'
#358390000000
1!
b100 %
1'
b100 +
#358400000000
1"
1(
#358410000000
0!
0"
b100 &
0'
0(
b100 ,
#358420000000
1!
b101 %
1'
b101 +
#358430000000
0!
0'
#358440000000
1!
b110 %
1'
b110 +
#358450000000
0!
0'
#358460000000
1!
b111 %
1'
b111 +
#358470000000
0!
0'
#358480000000
1!
0$
b1000 %
1'
0*
b1000 +
#358490000000
0!
0'
#358500000000
1!
b1001 %
1'
b1001 +
#358510000000
0!
0'
#358520000000
1!
b0 %
1'
b0 +
#358530000000
0!
0'
#358540000000
1!
1$
b1 %
1'
1*
b1 +
#358550000000
0!
0'
#358560000000
1!
b10 %
1'
b10 +
#358570000000
0!
0'
#358580000000
1!
b11 %
1'
b11 +
#358590000000
0!
0'
#358600000000
1!
b100 %
1'
b100 +
#358610000000
0!
0'
#358620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#358630000000
0!
0'
#358640000000
1!
0$
b110 %
1'
0*
b110 +
#358650000000
0!
0'
#358660000000
1!
b111 %
1'
b111 +
#358670000000
0!
0'
#358680000000
1!
b1000 %
1'
b1000 +
#358690000000
0!
0'
#358700000000
1!
b1001 %
1'
b1001 +
#358710000000
0!
0'
#358720000000
1!
b0 %
1'
b0 +
#358730000000
0!
0'
#358740000000
1!
1$
b1 %
1'
1*
b1 +
#358750000000
0!
0'
#358760000000
1!
b10 %
1'
b10 +
#358770000000
0!
0'
#358780000000
1!
b11 %
1'
b11 +
#358790000000
0!
0'
#358800000000
1!
b100 %
1'
b100 +
#358810000000
0!
0'
#358820000000
1!
b101 %
1'
b101 +
#358830000000
1"
1(
#358840000000
0!
0"
b100 &
0'
0(
b100 ,
#358850000000
1!
b110 %
1'
b110 +
#358860000000
0!
0'
#358870000000
1!
b111 %
1'
b111 +
#358880000000
0!
0'
#358890000000
1!
0$
b1000 %
1'
0*
b1000 +
#358900000000
0!
0'
#358910000000
1!
b1001 %
1'
b1001 +
#358920000000
0!
0'
#358930000000
1!
b0 %
1'
b0 +
#358940000000
0!
0'
#358950000000
1!
1$
b1 %
1'
1*
b1 +
#358960000000
0!
0'
#358970000000
1!
b10 %
1'
b10 +
#358980000000
0!
0'
#358990000000
1!
b11 %
1'
b11 +
#359000000000
0!
0'
#359010000000
1!
b100 %
1'
b100 +
#359020000000
0!
0'
#359030000000
1!
b101 %
1'
b101 +
#359040000000
0!
0'
#359050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#359060000000
0!
0'
#359070000000
1!
b111 %
1'
b111 +
#359080000000
0!
0'
#359090000000
1!
b1000 %
1'
b1000 +
#359100000000
0!
0'
#359110000000
1!
b1001 %
1'
b1001 +
#359120000000
0!
0'
#359130000000
1!
b0 %
1'
b0 +
#359140000000
0!
0'
#359150000000
1!
1$
b1 %
1'
1*
b1 +
#359160000000
0!
0'
#359170000000
1!
b10 %
1'
b10 +
#359180000000
0!
0'
#359190000000
1!
b11 %
1'
b11 +
#359200000000
0!
0'
#359210000000
1!
b100 %
1'
b100 +
#359220000000
0!
0'
#359230000000
1!
b101 %
1'
b101 +
#359240000000
0!
0'
#359250000000
1!
0$
b110 %
1'
0*
b110 +
#359260000000
1"
1(
#359270000000
0!
0"
b100 &
0'
0(
b100 ,
#359280000000
1!
1$
b111 %
1'
1*
b111 +
#359290000000
0!
0'
#359300000000
1!
0$
b1000 %
1'
0*
b1000 +
#359310000000
0!
0'
#359320000000
1!
b1001 %
1'
b1001 +
#359330000000
0!
0'
#359340000000
1!
b0 %
1'
b0 +
#359350000000
0!
0'
#359360000000
1!
1$
b1 %
1'
1*
b1 +
#359370000000
0!
0'
#359380000000
1!
b10 %
1'
b10 +
#359390000000
0!
0'
#359400000000
1!
b11 %
1'
b11 +
#359410000000
0!
0'
#359420000000
1!
b100 %
1'
b100 +
#359430000000
0!
0'
#359440000000
1!
b101 %
1'
b101 +
#359450000000
0!
0'
#359460000000
1!
b110 %
1'
b110 +
#359470000000
0!
0'
#359480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#359490000000
0!
0'
#359500000000
1!
b1000 %
1'
b1000 +
#359510000000
0!
0'
#359520000000
1!
b1001 %
1'
b1001 +
#359530000000
0!
0'
#359540000000
1!
b0 %
1'
b0 +
#359550000000
0!
0'
#359560000000
1!
1$
b1 %
1'
1*
b1 +
#359570000000
0!
0'
#359580000000
1!
b10 %
1'
b10 +
#359590000000
0!
0'
#359600000000
1!
b11 %
1'
b11 +
#359610000000
0!
0'
#359620000000
1!
b100 %
1'
b100 +
#359630000000
0!
0'
#359640000000
1!
b101 %
1'
b101 +
#359650000000
0!
0'
#359660000000
1!
0$
b110 %
1'
0*
b110 +
#359670000000
0!
0'
#359680000000
1!
b111 %
1'
b111 +
#359690000000
1"
1(
#359700000000
0!
0"
b100 &
0'
0(
b100 ,
#359710000000
1!
b1000 %
1'
b1000 +
#359720000000
0!
0'
#359730000000
1!
b1001 %
1'
b1001 +
#359740000000
0!
0'
#359750000000
1!
b0 %
1'
b0 +
#359760000000
0!
0'
#359770000000
1!
1$
b1 %
1'
1*
b1 +
#359780000000
0!
0'
#359790000000
1!
b10 %
1'
b10 +
#359800000000
0!
0'
#359810000000
1!
b11 %
1'
b11 +
#359820000000
0!
0'
#359830000000
1!
b100 %
1'
b100 +
#359840000000
0!
0'
#359850000000
1!
b101 %
1'
b101 +
#359860000000
0!
0'
#359870000000
1!
b110 %
1'
b110 +
#359880000000
0!
0'
#359890000000
1!
b111 %
1'
b111 +
#359900000000
0!
0'
#359910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#359920000000
0!
0'
#359930000000
1!
b1001 %
1'
b1001 +
#359940000000
0!
0'
#359950000000
1!
b0 %
1'
b0 +
#359960000000
0!
0'
#359970000000
1!
1$
b1 %
1'
1*
b1 +
#359980000000
0!
0'
#359990000000
1!
b10 %
1'
b10 +
#360000000000
0!
0'
#360010000000
1!
b11 %
1'
b11 +
#360020000000
0!
0'
#360030000000
1!
b100 %
1'
b100 +
#360040000000
0!
0'
#360050000000
1!
b101 %
1'
b101 +
#360060000000
0!
0'
#360070000000
1!
0$
b110 %
1'
0*
b110 +
#360080000000
0!
0'
#360090000000
1!
b111 %
1'
b111 +
#360100000000
0!
0'
#360110000000
1!
b1000 %
1'
b1000 +
#360120000000
1"
1(
#360130000000
0!
0"
b100 &
0'
0(
b100 ,
#360140000000
1!
b1001 %
1'
b1001 +
#360150000000
0!
0'
#360160000000
1!
b0 %
1'
b0 +
#360170000000
0!
0'
#360180000000
1!
1$
b1 %
1'
1*
b1 +
#360190000000
0!
0'
#360200000000
1!
b10 %
1'
b10 +
#360210000000
0!
0'
#360220000000
1!
b11 %
1'
b11 +
#360230000000
0!
0'
#360240000000
1!
b100 %
1'
b100 +
#360250000000
0!
0'
#360260000000
1!
b101 %
1'
b101 +
#360270000000
0!
0'
#360280000000
1!
b110 %
1'
b110 +
#360290000000
0!
0'
#360300000000
1!
b111 %
1'
b111 +
#360310000000
0!
0'
#360320000000
1!
0$
b1000 %
1'
0*
b1000 +
#360330000000
0!
0'
#360340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#360350000000
0!
0'
#360360000000
1!
b0 %
1'
b0 +
#360370000000
0!
0'
#360380000000
1!
1$
b1 %
1'
1*
b1 +
#360390000000
0!
0'
#360400000000
1!
b10 %
1'
b10 +
#360410000000
0!
0'
#360420000000
1!
b11 %
1'
b11 +
#360430000000
0!
0'
#360440000000
1!
b100 %
1'
b100 +
#360450000000
0!
0'
#360460000000
1!
b101 %
1'
b101 +
#360470000000
0!
0'
#360480000000
1!
0$
b110 %
1'
0*
b110 +
#360490000000
0!
0'
#360500000000
1!
b111 %
1'
b111 +
#360510000000
0!
0'
#360520000000
1!
b1000 %
1'
b1000 +
#360530000000
0!
0'
#360540000000
1!
b1001 %
1'
b1001 +
#360550000000
1"
1(
#360560000000
0!
0"
b100 &
0'
0(
b100 ,
#360570000000
1!
b0 %
1'
b0 +
#360580000000
0!
0'
#360590000000
1!
1$
b1 %
1'
1*
b1 +
#360600000000
0!
0'
#360610000000
1!
b10 %
1'
b10 +
#360620000000
0!
0'
#360630000000
1!
b11 %
1'
b11 +
#360640000000
0!
0'
#360650000000
1!
b100 %
1'
b100 +
#360660000000
0!
0'
#360670000000
1!
b101 %
1'
b101 +
#360680000000
0!
0'
#360690000000
1!
b110 %
1'
b110 +
#360700000000
0!
0'
#360710000000
1!
b111 %
1'
b111 +
#360720000000
0!
0'
#360730000000
1!
0$
b1000 %
1'
0*
b1000 +
#360740000000
0!
0'
#360750000000
1!
b1001 %
1'
b1001 +
#360760000000
0!
0'
#360770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#360780000000
0!
0'
#360790000000
1!
1$
b1 %
1'
1*
b1 +
#360800000000
0!
0'
#360810000000
1!
b10 %
1'
b10 +
#360820000000
0!
0'
#360830000000
1!
b11 %
1'
b11 +
#360840000000
0!
0'
#360850000000
1!
b100 %
1'
b100 +
#360860000000
0!
0'
#360870000000
1!
b101 %
1'
b101 +
#360880000000
0!
0'
#360890000000
1!
0$
b110 %
1'
0*
b110 +
#360900000000
0!
0'
#360910000000
1!
b111 %
1'
b111 +
#360920000000
0!
0'
#360930000000
1!
b1000 %
1'
b1000 +
#360940000000
0!
0'
#360950000000
1!
b1001 %
1'
b1001 +
#360960000000
0!
0'
#360970000000
1!
b0 %
1'
b0 +
#360980000000
1"
1(
#360990000000
0!
0"
b100 &
0'
0(
b100 ,
#361000000000
1!
1$
b1 %
1'
1*
b1 +
#361010000000
0!
0'
#361020000000
1!
b10 %
1'
b10 +
#361030000000
0!
0'
#361040000000
1!
b11 %
1'
b11 +
#361050000000
0!
0'
#361060000000
1!
b100 %
1'
b100 +
#361070000000
0!
0'
#361080000000
1!
b101 %
1'
b101 +
#361090000000
0!
0'
#361100000000
1!
b110 %
1'
b110 +
#361110000000
0!
0'
#361120000000
1!
b111 %
1'
b111 +
#361130000000
0!
0'
#361140000000
1!
0$
b1000 %
1'
0*
b1000 +
#361150000000
0!
0'
#361160000000
1!
b1001 %
1'
b1001 +
#361170000000
0!
0'
#361180000000
1!
b0 %
1'
b0 +
#361190000000
0!
0'
#361200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#361210000000
0!
0'
#361220000000
1!
b10 %
1'
b10 +
#361230000000
0!
0'
#361240000000
1!
b11 %
1'
b11 +
#361250000000
0!
0'
#361260000000
1!
b100 %
1'
b100 +
#361270000000
0!
0'
#361280000000
1!
b101 %
1'
b101 +
#361290000000
0!
0'
#361300000000
1!
0$
b110 %
1'
0*
b110 +
#361310000000
0!
0'
#361320000000
1!
b111 %
1'
b111 +
#361330000000
0!
0'
#361340000000
1!
b1000 %
1'
b1000 +
#361350000000
0!
0'
#361360000000
1!
b1001 %
1'
b1001 +
#361370000000
0!
0'
#361380000000
1!
b0 %
1'
b0 +
#361390000000
0!
0'
#361400000000
1!
1$
b1 %
1'
1*
b1 +
#361410000000
1"
1(
#361420000000
0!
0"
b100 &
0'
0(
b100 ,
#361430000000
1!
b10 %
1'
b10 +
#361440000000
0!
0'
#361450000000
1!
b11 %
1'
b11 +
#361460000000
0!
0'
#361470000000
1!
b100 %
1'
b100 +
#361480000000
0!
0'
#361490000000
1!
b101 %
1'
b101 +
#361500000000
0!
0'
#361510000000
1!
b110 %
1'
b110 +
#361520000000
0!
0'
#361530000000
1!
b111 %
1'
b111 +
#361540000000
0!
0'
#361550000000
1!
0$
b1000 %
1'
0*
b1000 +
#361560000000
0!
0'
#361570000000
1!
b1001 %
1'
b1001 +
#361580000000
0!
0'
#361590000000
1!
b0 %
1'
b0 +
#361600000000
0!
0'
#361610000000
1!
1$
b1 %
1'
1*
b1 +
#361620000000
0!
0'
#361630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#361640000000
0!
0'
#361650000000
1!
b11 %
1'
b11 +
#361660000000
0!
0'
#361670000000
1!
b100 %
1'
b100 +
#361680000000
0!
0'
#361690000000
1!
b101 %
1'
b101 +
#361700000000
0!
0'
#361710000000
1!
0$
b110 %
1'
0*
b110 +
#361720000000
0!
0'
#361730000000
1!
b111 %
1'
b111 +
#361740000000
0!
0'
#361750000000
1!
b1000 %
1'
b1000 +
#361760000000
0!
0'
#361770000000
1!
b1001 %
1'
b1001 +
#361780000000
0!
0'
#361790000000
1!
b0 %
1'
b0 +
#361800000000
0!
0'
#361810000000
1!
1$
b1 %
1'
1*
b1 +
#361820000000
0!
0'
#361830000000
1!
b10 %
1'
b10 +
#361840000000
1"
1(
#361850000000
0!
0"
b100 &
0'
0(
b100 ,
#361860000000
1!
b11 %
1'
b11 +
#361870000000
0!
0'
#361880000000
1!
b100 %
1'
b100 +
#361890000000
0!
0'
#361900000000
1!
b101 %
1'
b101 +
#361910000000
0!
0'
#361920000000
1!
b110 %
1'
b110 +
#361930000000
0!
0'
#361940000000
1!
b111 %
1'
b111 +
#361950000000
0!
0'
#361960000000
1!
0$
b1000 %
1'
0*
b1000 +
#361970000000
0!
0'
#361980000000
1!
b1001 %
1'
b1001 +
#361990000000
0!
0'
#362000000000
1!
b0 %
1'
b0 +
#362010000000
0!
0'
#362020000000
1!
1$
b1 %
1'
1*
b1 +
#362030000000
0!
0'
#362040000000
1!
b10 %
1'
b10 +
#362050000000
0!
0'
#362060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#362070000000
0!
0'
#362080000000
1!
b100 %
1'
b100 +
#362090000000
0!
0'
#362100000000
1!
b101 %
1'
b101 +
#362110000000
0!
0'
#362120000000
1!
0$
b110 %
1'
0*
b110 +
#362130000000
0!
0'
#362140000000
1!
b111 %
1'
b111 +
#362150000000
0!
0'
#362160000000
1!
b1000 %
1'
b1000 +
#362170000000
0!
0'
#362180000000
1!
b1001 %
1'
b1001 +
#362190000000
0!
0'
#362200000000
1!
b0 %
1'
b0 +
#362210000000
0!
0'
#362220000000
1!
1$
b1 %
1'
1*
b1 +
#362230000000
0!
0'
#362240000000
1!
b10 %
1'
b10 +
#362250000000
0!
0'
#362260000000
1!
b11 %
1'
b11 +
#362270000000
1"
1(
#362280000000
0!
0"
b100 &
0'
0(
b100 ,
#362290000000
1!
b100 %
1'
b100 +
#362300000000
0!
0'
#362310000000
1!
b101 %
1'
b101 +
#362320000000
0!
0'
#362330000000
1!
b110 %
1'
b110 +
#362340000000
0!
0'
#362350000000
1!
b111 %
1'
b111 +
#362360000000
0!
0'
#362370000000
1!
0$
b1000 %
1'
0*
b1000 +
#362380000000
0!
0'
#362390000000
1!
b1001 %
1'
b1001 +
#362400000000
0!
0'
#362410000000
1!
b0 %
1'
b0 +
#362420000000
0!
0'
#362430000000
1!
1$
b1 %
1'
1*
b1 +
#362440000000
0!
0'
#362450000000
1!
b10 %
1'
b10 +
#362460000000
0!
0'
#362470000000
1!
b11 %
1'
b11 +
#362480000000
0!
0'
#362490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#362500000000
0!
0'
#362510000000
1!
b101 %
1'
b101 +
#362520000000
0!
0'
#362530000000
1!
0$
b110 %
1'
0*
b110 +
#362540000000
0!
0'
#362550000000
1!
b111 %
1'
b111 +
#362560000000
0!
0'
#362570000000
1!
b1000 %
1'
b1000 +
#362580000000
0!
0'
#362590000000
1!
b1001 %
1'
b1001 +
#362600000000
0!
0'
#362610000000
1!
b0 %
1'
b0 +
#362620000000
0!
0'
#362630000000
1!
1$
b1 %
1'
1*
b1 +
#362640000000
0!
0'
#362650000000
1!
b10 %
1'
b10 +
#362660000000
0!
0'
#362670000000
1!
b11 %
1'
b11 +
#362680000000
0!
0'
#362690000000
1!
b100 %
1'
b100 +
#362700000000
1"
1(
#362710000000
0!
0"
b100 &
0'
0(
b100 ,
#362720000000
1!
b101 %
1'
b101 +
#362730000000
0!
0'
#362740000000
1!
b110 %
1'
b110 +
#362750000000
0!
0'
#362760000000
1!
b111 %
1'
b111 +
#362770000000
0!
0'
#362780000000
1!
0$
b1000 %
1'
0*
b1000 +
#362790000000
0!
0'
#362800000000
1!
b1001 %
1'
b1001 +
#362810000000
0!
0'
#362820000000
1!
b0 %
1'
b0 +
#362830000000
0!
0'
#362840000000
1!
1$
b1 %
1'
1*
b1 +
#362850000000
0!
0'
#362860000000
1!
b10 %
1'
b10 +
#362870000000
0!
0'
#362880000000
1!
b11 %
1'
b11 +
#362890000000
0!
0'
#362900000000
1!
b100 %
1'
b100 +
#362910000000
0!
0'
#362920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#362930000000
0!
0'
#362940000000
1!
0$
b110 %
1'
0*
b110 +
#362950000000
0!
0'
#362960000000
1!
b111 %
1'
b111 +
#362970000000
0!
0'
#362980000000
1!
b1000 %
1'
b1000 +
#362990000000
0!
0'
#363000000000
1!
b1001 %
1'
b1001 +
#363010000000
0!
0'
#363020000000
1!
b0 %
1'
b0 +
#363030000000
0!
0'
#363040000000
1!
1$
b1 %
1'
1*
b1 +
#363050000000
0!
0'
#363060000000
1!
b10 %
1'
b10 +
#363070000000
0!
0'
#363080000000
1!
b11 %
1'
b11 +
#363090000000
0!
0'
#363100000000
1!
b100 %
1'
b100 +
#363110000000
0!
0'
#363120000000
1!
b101 %
1'
b101 +
#363130000000
1"
1(
#363140000000
0!
0"
b100 &
0'
0(
b100 ,
#363150000000
1!
b110 %
1'
b110 +
#363160000000
0!
0'
#363170000000
1!
b111 %
1'
b111 +
#363180000000
0!
0'
#363190000000
1!
0$
b1000 %
1'
0*
b1000 +
#363200000000
0!
0'
#363210000000
1!
b1001 %
1'
b1001 +
#363220000000
0!
0'
#363230000000
1!
b0 %
1'
b0 +
#363240000000
0!
0'
#363250000000
1!
1$
b1 %
1'
1*
b1 +
#363260000000
0!
0'
#363270000000
1!
b10 %
1'
b10 +
#363280000000
0!
0'
#363290000000
1!
b11 %
1'
b11 +
#363300000000
0!
0'
#363310000000
1!
b100 %
1'
b100 +
#363320000000
0!
0'
#363330000000
1!
b101 %
1'
b101 +
#363340000000
0!
0'
#363350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#363360000000
0!
0'
#363370000000
1!
b111 %
1'
b111 +
#363380000000
0!
0'
#363390000000
1!
b1000 %
1'
b1000 +
#363400000000
0!
0'
#363410000000
1!
b1001 %
1'
b1001 +
#363420000000
0!
0'
#363430000000
1!
b0 %
1'
b0 +
#363440000000
0!
0'
#363450000000
1!
1$
b1 %
1'
1*
b1 +
#363460000000
0!
0'
#363470000000
1!
b10 %
1'
b10 +
#363480000000
0!
0'
#363490000000
1!
b11 %
1'
b11 +
#363500000000
0!
0'
#363510000000
1!
b100 %
1'
b100 +
#363520000000
0!
0'
#363530000000
1!
b101 %
1'
b101 +
#363540000000
0!
0'
#363550000000
1!
0$
b110 %
1'
0*
b110 +
#363560000000
1"
1(
#363570000000
0!
0"
b100 &
0'
0(
b100 ,
#363580000000
1!
1$
b111 %
1'
1*
b111 +
#363590000000
0!
0'
#363600000000
1!
0$
b1000 %
1'
0*
b1000 +
#363610000000
0!
0'
#363620000000
1!
b1001 %
1'
b1001 +
#363630000000
0!
0'
#363640000000
1!
b0 %
1'
b0 +
#363650000000
0!
0'
#363660000000
1!
1$
b1 %
1'
1*
b1 +
#363670000000
0!
0'
#363680000000
1!
b10 %
1'
b10 +
#363690000000
0!
0'
#363700000000
1!
b11 %
1'
b11 +
#363710000000
0!
0'
#363720000000
1!
b100 %
1'
b100 +
#363730000000
0!
0'
#363740000000
1!
b101 %
1'
b101 +
#363750000000
0!
0'
#363760000000
1!
b110 %
1'
b110 +
#363770000000
0!
0'
#363780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#363790000000
0!
0'
#363800000000
1!
b1000 %
1'
b1000 +
#363810000000
0!
0'
#363820000000
1!
b1001 %
1'
b1001 +
#363830000000
0!
0'
#363840000000
1!
b0 %
1'
b0 +
#363850000000
0!
0'
#363860000000
1!
1$
b1 %
1'
1*
b1 +
#363870000000
0!
0'
#363880000000
1!
b10 %
1'
b10 +
#363890000000
0!
0'
#363900000000
1!
b11 %
1'
b11 +
#363910000000
0!
0'
#363920000000
1!
b100 %
1'
b100 +
#363930000000
0!
0'
#363940000000
1!
b101 %
1'
b101 +
#363950000000
0!
0'
#363960000000
1!
0$
b110 %
1'
0*
b110 +
#363970000000
0!
0'
#363980000000
1!
b111 %
1'
b111 +
#363990000000
1"
1(
#364000000000
0!
0"
b100 &
0'
0(
b100 ,
#364010000000
1!
b1000 %
1'
b1000 +
#364020000000
0!
0'
#364030000000
1!
b1001 %
1'
b1001 +
#364040000000
0!
0'
#364050000000
1!
b0 %
1'
b0 +
#364060000000
0!
0'
#364070000000
1!
1$
b1 %
1'
1*
b1 +
#364080000000
0!
0'
#364090000000
1!
b10 %
1'
b10 +
#364100000000
0!
0'
#364110000000
1!
b11 %
1'
b11 +
#364120000000
0!
0'
#364130000000
1!
b100 %
1'
b100 +
#364140000000
0!
0'
#364150000000
1!
b101 %
1'
b101 +
#364160000000
0!
0'
#364170000000
1!
b110 %
1'
b110 +
#364180000000
0!
0'
#364190000000
1!
b111 %
1'
b111 +
#364200000000
0!
0'
#364210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#364220000000
0!
0'
#364230000000
1!
b1001 %
1'
b1001 +
#364240000000
0!
0'
#364250000000
1!
b0 %
1'
b0 +
#364260000000
0!
0'
#364270000000
1!
1$
b1 %
1'
1*
b1 +
#364280000000
0!
0'
#364290000000
1!
b10 %
1'
b10 +
#364300000000
0!
0'
#364310000000
1!
b11 %
1'
b11 +
#364320000000
0!
0'
#364330000000
1!
b100 %
1'
b100 +
#364340000000
0!
0'
#364350000000
1!
b101 %
1'
b101 +
#364360000000
0!
0'
#364370000000
1!
0$
b110 %
1'
0*
b110 +
#364380000000
0!
0'
#364390000000
1!
b111 %
1'
b111 +
#364400000000
0!
0'
#364410000000
1!
b1000 %
1'
b1000 +
#364420000000
1"
1(
#364430000000
0!
0"
b100 &
0'
0(
b100 ,
#364440000000
1!
b1001 %
1'
b1001 +
#364450000000
0!
0'
#364460000000
1!
b0 %
1'
b0 +
#364470000000
0!
0'
#364480000000
1!
1$
b1 %
1'
1*
b1 +
#364490000000
0!
0'
#364500000000
1!
b10 %
1'
b10 +
#364510000000
0!
0'
#364520000000
1!
b11 %
1'
b11 +
#364530000000
0!
0'
#364540000000
1!
b100 %
1'
b100 +
#364550000000
0!
0'
#364560000000
1!
b101 %
1'
b101 +
#364570000000
0!
0'
#364580000000
1!
b110 %
1'
b110 +
#364590000000
0!
0'
#364600000000
1!
b111 %
1'
b111 +
#364610000000
0!
0'
#364620000000
1!
0$
b1000 %
1'
0*
b1000 +
#364630000000
0!
0'
#364640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#364650000000
0!
0'
#364660000000
1!
b0 %
1'
b0 +
#364670000000
0!
0'
#364680000000
1!
1$
b1 %
1'
1*
b1 +
#364690000000
0!
0'
#364700000000
1!
b10 %
1'
b10 +
#364710000000
0!
0'
#364720000000
1!
b11 %
1'
b11 +
#364730000000
0!
0'
#364740000000
1!
b100 %
1'
b100 +
#364750000000
0!
0'
#364760000000
1!
b101 %
1'
b101 +
#364770000000
0!
0'
#364780000000
1!
0$
b110 %
1'
0*
b110 +
#364790000000
0!
0'
#364800000000
1!
b111 %
1'
b111 +
#364810000000
0!
0'
#364820000000
1!
b1000 %
1'
b1000 +
#364830000000
0!
0'
#364840000000
1!
b1001 %
1'
b1001 +
#364850000000
1"
1(
#364860000000
0!
0"
b100 &
0'
0(
b100 ,
#364870000000
1!
b0 %
1'
b0 +
#364880000000
0!
0'
#364890000000
1!
1$
b1 %
1'
1*
b1 +
#364900000000
0!
0'
#364910000000
1!
b10 %
1'
b10 +
#364920000000
0!
0'
#364930000000
1!
b11 %
1'
b11 +
#364940000000
0!
0'
#364950000000
1!
b100 %
1'
b100 +
#364960000000
0!
0'
#364970000000
1!
b101 %
1'
b101 +
#364980000000
0!
0'
#364990000000
1!
b110 %
1'
b110 +
#365000000000
0!
0'
#365010000000
1!
b111 %
1'
b111 +
#365020000000
0!
0'
#365030000000
1!
0$
b1000 %
1'
0*
b1000 +
#365040000000
0!
0'
#365050000000
1!
b1001 %
1'
b1001 +
#365060000000
0!
0'
#365070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#365080000000
0!
0'
#365090000000
1!
1$
b1 %
1'
1*
b1 +
#365100000000
0!
0'
#365110000000
1!
b10 %
1'
b10 +
#365120000000
0!
0'
#365130000000
1!
b11 %
1'
b11 +
#365140000000
0!
0'
#365150000000
1!
b100 %
1'
b100 +
#365160000000
0!
0'
#365170000000
1!
b101 %
1'
b101 +
#365180000000
0!
0'
#365190000000
1!
0$
b110 %
1'
0*
b110 +
#365200000000
0!
0'
#365210000000
1!
b111 %
1'
b111 +
#365220000000
0!
0'
#365230000000
1!
b1000 %
1'
b1000 +
#365240000000
0!
0'
#365250000000
1!
b1001 %
1'
b1001 +
#365260000000
0!
0'
#365270000000
1!
b0 %
1'
b0 +
#365280000000
1"
1(
#365290000000
0!
0"
b100 &
0'
0(
b100 ,
#365300000000
1!
1$
b1 %
1'
1*
b1 +
#365310000000
0!
0'
#365320000000
1!
b10 %
1'
b10 +
#365330000000
0!
0'
#365340000000
1!
b11 %
1'
b11 +
#365350000000
0!
0'
#365360000000
1!
b100 %
1'
b100 +
#365370000000
0!
0'
#365380000000
1!
b101 %
1'
b101 +
#365390000000
0!
0'
#365400000000
1!
b110 %
1'
b110 +
#365410000000
0!
0'
#365420000000
1!
b111 %
1'
b111 +
#365430000000
0!
0'
#365440000000
1!
0$
b1000 %
1'
0*
b1000 +
#365450000000
0!
0'
#365460000000
1!
b1001 %
1'
b1001 +
#365470000000
0!
0'
#365480000000
1!
b0 %
1'
b0 +
#365490000000
0!
0'
#365500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#365510000000
0!
0'
#365520000000
1!
b10 %
1'
b10 +
#365530000000
0!
0'
#365540000000
1!
b11 %
1'
b11 +
#365550000000
0!
0'
#365560000000
1!
b100 %
1'
b100 +
#365570000000
0!
0'
#365580000000
1!
b101 %
1'
b101 +
#365590000000
0!
0'
#365600000000
1!
0$
b110 %
1'
0*
b110 +
#365610000000
0!
0'
#365620000000
1!
b111 %
1'
b111 +
#365630000000
0!
0'
#365640000000
1!
b1000 %
1'
b1000 +
#365650000000
0!
0'
#365660000000
1!
b1001 %
1'
b1001 +
#365670000000
0!
0'
#365680000000
1!
b0 %
1'
b0 +
#365690000000
0!
0'
#365700000000
1!
1$
b1 %
1'
1*
b1 +
#365710000000
1"
1(
#365720000000
0!
0"
b100 &
0'
0(
b100 ,
#365730000000
1!
b10 %
1'
b10 +
#365740000000
0!
0'
#365750000000
1!
b11 %
1'
b11 +
#365760000000
0!
0'
#365770000000
1!
b100 %
1'
b100 +
#365780000000
0!
0'
#365790000000
1!
b101 %
1'
b101 +
#365800000000
0!
0'
#365810000000
1!
b110 %
1'
b110 +
#365820000000
0!
0'
#365830000000
1!
b111 %
1'
b111 +
#365840000000
0!
0'
#365850000000
1!
0$
b1000 %
1'
0*
b1000 +
#365860000000
0!
0'
#365870000000
1!
b1001 %
1'
b1001 +
#365880000000
0!
0'
#365890000000
1!
b0 %
1'
b0 +
#365900000000
0!
0'
#365910000000
1!
1$
b1 %
1'
1*
b1 +
#365920000000
0!
0'
#365930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#365940000000
0!
0'
#365950000000
1!
b11 %
1'
b11 +
#365960000000
0!
0'
#365970000000
1!
b100 %
1'
b100 +
#365980000000
0!
0'
#365990000000
1!
b101 %
1'
b101 +
#366000000000
0!
0'
#366010000000
1!
0$
b110 %
1'
0*
b110 +
#366020000000
0!
0'
#366030000000
1!
b111 %
1'
b111 +
#366040000000
0!
0'
#366050000000
1!
b1000 %
1'
b1000 +
#366060000000
0!
0'
#366070000000
1!
b1001 %
1'
b1001 +
#366080000000
0!
0'
#366090000000
1!
b0 %
1'
b0 +
#366100000000
0!
0'
#366110000000
1!
1$
b1 %
1'
1*
b1 +
#366120000000
0!
0'
#366130000000
1!
b10 %
1'
b10 +
#366140000000
1"
1(
#366150000000
0!
0"
b100 &
0'
0(
b100 ,
#366160000000
1!
b11 %
1'
b11 +
#366170000000
0!
0'
#366180000000
1!
b100 %
1'
b100 +
#366190000000
0!
0'
#366200000000
1!
b101 %
1'
b101 +
#366210000000
0!
0'
#366220000000
1!
b110 %
1'
b110 +
#366230000000
0!
0'
#366240000000
1!
b111 %
1'
b111 +
#366250000000
0!
0'
#366260000000
1!
0$
b1000 %
1'
0*
b1000 +
#366270000000
0!
0'
#366280000000
1!
b1001 %
1'
b1001 +
#366290000000
0!
0'
#366300000000
1!
b0 %
1'
b0 +
#366310000000
0!
0'
#366320000000
1!
1$
b1 %
1'
1*
b1 +
#366330000000
0!
0'
#366340000000
1!
b10 %
1'
b10 +
#366350000000
0!
0'
#366360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#366370000000
0!
0'
#366380000000
1!
b100 %
1'
b100 +
#366390000000
0!
0'
#366400000000
1!
b101 %
1'
b101 +
#366410000000
0!
0'
#366420000000
1!
0$
b110 %
1'
0*
b110 +
#366430000000
0!
0'
#366440000000
1!
b111 %
1'
b111 +
#366450000000
0!
0'
#366460000000
1!
b1000 %
1'
b1000 +
#366470000000
0!
0'
#366480000000
1!
b1001 %
1'
b1001 +
#366490000000
0!
0'
#366500000000
1!
b0 %
1'
b0 +
#366510000000
0!
0'
#366520000000
1!
1$
b1 %
1'
1*
b1 +
#366530000000
0!
0'
#366540000000
1!
b10 %
1'
b10 +
#366550000000
0!
0'
#366560000000
1!
b11 %
1'
b11 +
#366570000000
1"
1(
#366580000000
0!
0"
b100 &
0'
0(
b100 ,
#366590000000
1!
b100 %
1'
b100 +
#366600000000
0!
0'
#366610000000
1!
b101 %
1'
b101 +
#366620000000
0!
0'
#366630000000
1!
b110 %
1'
b110 +
#366640000000
0!
0'
#366650000000
1!
b111 %
1'
b111 +
#366660000000
0!
0'
#366670000000
1!
0$
b1000 %
1'
0*
b1000 +
#366680000000
0!
0'
#366690000000
1!
b1001 %
1'
b1001 +
#366700000000
0!
0'
#366710000000
1!
b0 %
1'
b0 +
#366720000000
0!
0'
#366730000000
1!
1$
b1 %
1'
1*
b1 +
#366740000000
0!
0'
#366750000000
1!
b10 %
1'
b10 +
#366760000000
0!
0'
#366770000000
1!
b11 %
1'
b11 +
#366780000000
0!
0'
#366790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#366800000000
0!
0'
#366810000000
1!
b101 %
1'
b101 +
#366820000000
0!
0'
#366830000000
1!
0$
b110 %
1'
0*
b110 +
#366840000000
0!
0'
#366850000000
1!
b111 %
1'
b111 +
#366860000000
0!
0'
#366870000000
1!
b1000 %
1'
b1000 +
#366880000000
0!
0'
#366890000000
1!
b1001 %
1'
b1001 +
#366900000000
0!
0'
#366910000000
1!
b0 %
1'
b0 +
#366920000000
0!
0'
#366930000000
1!
1$
b1 %
1'
1*
b1 +
#366940000000
0!
0'
#366950000000
1!
b10 %
1'
b10 +
#366960000000
0!
0'
#366970000000
1!
b11 %
1'
b11 +
#366980000000
0!
0'
#366990000000
1!
b100 %
1'
b100 +
#367000000000
1"
1(
#367010000000
0!
0"
b100 &
0'
0(
b100 ,
#367020000000
1!
b101 %
1'
b101 +
#367030000000
0!
0'
#367040000000
1!
b110 %
1'
b110 +
#367050000000
0!
0'
#367060000000
1!
b111 %
1'
b111 +
#367070000000
0!
0'
#367080000000
1!
0$
b1000 %
1'
0*
b1000 +
#367090000000
0!
0'
#367100000000
1!
b1001 %
1'
b1001 +
#367110000000
0!
0'
#367120000000
1!
b0 %
1'
b0 +
#367130000000
0!
0'
#367140000000
1!
1$
b1 %
1'
1*
b1 +
#367150000000
0!
0'
#367160000000
1!
b10 %
1'
b10 +
#367170000000
0!
0'
#367180000000
1!
b11 %
1'
b11 +
#367190000000
0!
0'
#367200000000
1!
b100 %
1'
b100 +
#367210000000
0!
0'
#367220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#367230000000
0!
0'
#367240000000
1!
0$
b110 %
1'
0*
b110 +
#367250000000
0!
0'
#367260000000
1!
b111 %
1'
b111 +
#367270000000
0!
0'
#367280000000
1!
b1000 %
1'
b1000 +
#367290000000
0!
0'
#367300000000
1!
b1001 %
1'
b1001 +
#367310000000
0!
0'
#367320000000
1!
b0 %
1'
b0 +
#367330000000
0!
0'
#367340000000
1!
1$
b1 %
1'
1*
b1 +
#367350000000
0!
0'
#367360000000
1!
b10 %
1'
b10 +
#367370000000
0!
0'
#367380000000
1!
b11 %
1'
b11 +
#367390000000
0!
0'
#367400000000
1!
b100 %
1'
b100 +
#367410000000
0!
0'
#367420000000
1!
b101 %
1'
b101 +
#367430000000
1"
1(
#367440000000
0!
0"
b100 &
0'
0(
b100 ,
#367450000000
1!
b110 %
1'
b110 +
#367460000000
0!
0'
#367470000000
1!
b111 %
1'
b111 +
#367480000000
0!
0'
#367490000000
1!
0$
b1000 %
1'
0*
b1000 +
#367500000000
0!
0'
#367510000000
1!
b1001 %
1'
b1001 +
#367520000000
0!
0'
#367530000000
1!
b0 %
1'
b0 +
#367540000000
0!
0'
#367550000000
1!
1$
b1 %
1'
1*
b1 +
#367560000000
0!
0'
#367570000000
1!
b10 %
1'
b10 +
#367580000000
0!
0'
#367590000000
1!
b11 %
1'
b11 +
#367600000000
0!
0'
#367610000000
1!
b100 %
1'
b100 +
#367620000000
0!
0'
#367630000000
1!
b101 %
1'
b101 +
#367640000000
0!
0'
#367650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#367660000000
0!
0'
#367670000000
1!
b111 %
1'
b111 +
#367680000000
0!
0'
#367690000000
1!
b1000 %
1'
b1000 +
#367700000000
0!
0'
#367710000000
1!
b1001 %
1'
b1001 +
#367720000000
0!
0'
#367730000000
1!
b0 %
1'
b0 +
#367740000000
0!
0'
#367750000000
1!
1$
b1 %
1'
1*
b1 +
#367760000000
0!
0'
#367770000000
1!
b10 %
1'
b10 +
#367780000000
0!
0'
#367790000000
1!
b11 %
1'
b11 +
#367800000000
0!
0'
#367810000000
1!
b100 %
1'
b100 +
#367820000000
0!
0'
#367830000000
1!
b101 %
1'
b101 +
#367840000000
0!
0'
#367850000000
1!
0$
b110 %
1'
0*
b110 +
#367860000000
1"
1(
#367870000000
0!
0"
b100 &
0'
0(
b100 ,
#367880000000
1!
1$
b111 %
1'
1*
b111 +
#367890000000
0!
0'
#367900000000
1!
0$
b1000 %
1'
0*
b1000 +
#367910000000
0!
0'
#367920000000
1!
b1001 %
1'
b1001 +
#367930000000
0!
0'
#367940000000
1!
b0 %
1'
b0 +
#367950000000
0!
0'
#367960000000
1!
1$
b1 %
1'
1*
b1 +
#367970000000
0!
0'
#367980000000
1!
b10 %
1'
b10 +
#367990000000
0!
0'
#368000000000
1!
b11 %
1'
b11 +
#368010000000
0!
0'
#368020000000
1!
b100 %
1'
b100 +
#368030000000
0!
0'
#368040000000
1!
b101 %
1'
b101 +
#368050000000
0!
0'
#368060000000
1!
b110 %
1'
b110 +
#368070000000
0!
0'
#368080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#368090000000
0!
0'
#368100000000
1!
b1000 %
1'
b1000 +
#368110000000
0!
0'
#368120000000
1!
b1001 %
1'
b1001 +
#368130000000
0!
0'
#368140000000
1!
b0 %
1'
b0 +
#368150000000
0!
0'
#368160000000
1!
1$
b1 %
1'
1*
b1 +
#368170000000
0!
0'
#368180000000
1!
b10 %
1'
b10 +
#368190000000
0!
0'
#368200000000
1!
b11 %
1'
b11 +
#368210000000
0!
0'
#368220000000
1!
b100 %
1'
b100 +
#368230000000
0!
0'
#368240000000
1!
b101 %
1'
b101 +
#368250000000
0!
0'
#368260000000
1!
0$
b110 %
1'
0*
b110 +
#368270000000
0!
0'
#368280000000
1!
b111 %
1'
b111 +
#368290000000
1"
1(
#368300000000
0!
0"
b100 &
0'
0(
b100 ,
#368310000000
1!
b1000 %
1'
b1000 +
#368320000000
0!
0'
#368330000000
1!
b1001 %
1'
b1001 +
#368340000000
0!
0'
#368350000000
1!
b0 %
1'
b0 +
#368360000000
0!
0'
#368370000000
1!
1$
b1 %
1'
1*
b1 +
#368380000000
0!
0'
#368390000000
1!
b10 %
1'
b10 +
#368400000000
0!
0'
#368410000000
1!
b11 %
1'
b11 +
#368420000000
0!
0'
#368430000000
1!
b100 %
1'
b100 +
#368440000000
0!
0'
#368450000000
1!
b101 %
1'
b101 +
#368460000000
0!
0'
#368470000000
1!
b110 %
1'
b110 +
#368480000000
0!
0'
#368490000000
1!
b111 %
1'
b111 +
#368500000000
0!
0'
#368510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#368520000000
0!
0'
#368530000000
1!
b1001 %
1'
b1001 +
#368540000000
0!
0'
#368550000000
1!
b0 %
1'
b0 +
#368560000000
0!
0'
#368570000000
1!
1$
b1 %
1'
1*
b1 +
#368580000000
0!
0'
#368590000000
1!
b10 %
1'
b10 +
#368600000000
0!
0'
#368610000000
1!
b11 %
1'
b11 +
#368620000000
0!
0'
#368630000000
1!
b100 %
1'
b100 +
#368640000000
0!
0'
#368650000000
1!
b101 %
1'
b101 +
#368660000000
0!
0'
#368670000000
1!
0$
b110 %
1'
0*
b110 +
#368680000000
0!
0'
#368690000000
1!
b111 %
1'
b111 +
#368700000000
0!
0'
#368710000000
1!
b1000 %
1'
b1000 +
#368720000000
1"
1(
#368730000000
0!
0"
b100 &
0'
0(
b100 ,
#368740000000
1!
b1001 %
1'
b1001 +
#368750000000
0!
0'
#368760000000
1!
b0 %
1'
b0 +
#368770000000
0!
0'
#368780000000
1!
1$
b1 %
1'
1*
b1 +
#368790000000
0!
0'
#368800000000
1!
b10 %
1'
b10 +
#368810000000
0!
0'
#368820000000
1!
b11 %
1'
b11 +
#368830000000
0!
0'
#368840000000
1!
b100 %
1'
b100 +
#368850000000
0!
0'
#368860000000
1!
b101 %
1'
b101 +
#368870000000
0!
0'
#368880000000
1!
b110 %
1'
b110 +
#368890000000
0!
0'
#368900000000
1!
b111 %
1'
b111 +
#368910000000
0!
0'
#368920000000
1!
0$
b1000 %
1'
0*
b1000 +
#368930000000
0!
0'
#368940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#368950000000
0!
0'
#368960000000
1!
b0 %
1'
b0 +
#368970000000
0!
0'
#368980000000
1!
1$
b1 %
1'
1*
b1 +
#368990000000
0!
0'
#369000000000
1!
b10 %
1'
b10 +
#369010000000
0!
0'
#369020000000
1!
b11 %
1'
b11 +
#369030000000
0!
0'
#369040000000
1!
b100 %
1'
b100 +
#369050000000
0!
0'
#369060000000
1!
b101 %
1'
b101 +
#369070000000
0!
0'
#369080000000
1!
0$
b110 %
1'
0*
b110 +
#369090000000
0!
0'
#369100000000
1!
b111 %
1'
b111 +
#369110000000
0!
0'
#369120000000
1!
b1000 %
1'
b1000 +
#369130000000
0!
0'
#369140000000
1!
b1001 %
1'
b1001 +
#369150000000
1"
1(
#369160000000
0!
0"
b100 &
0'
0(
b100 ,
#369170000000
1!
b0 %
1'
b0 +
#369180000000
0!
0'
#369190000000
1!
1$
b1 %
1'
1*
b1 +
#369200000000
0!
0'
#369210000000
1!
b10 %
1'
b10 +
#369220000000
0!
0'
#369230000000
1!
b11 %
1'
b11 +
#369240000000
0!
0'
#369250000000
1!
b100 %
1'
b100 +
#369260000000
0!
0'
#369270000000
1!
b101 %
1'
b101 +
#369280000000
0!
0'
#369290000000
1!
b110 %
1'
b110 +
#369300000000
0!
0'
#369310000000
1!
b111 %
1'
b111 +
#369320000000
0!
0'
#369330000000
1!
0$
b1000 %
1'
0*
b1000 +
#369340000000
0!
0'
#369350000000
1!
b1001 %
1'
b1001 +
#369360000000
0!
0'
#369370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#369380000000
0!
0'
#369390000000
1!
1$
b1 %
1'
1*
b1 +
#369400000000
0!
0'
#369410000000
1!
b10 %
1'
b10 +
#369420000000
0!
0'
#369430000000
1!
b11 %
1'
b11 +
#369440000000
0!
0'
#369450000000
1!
b100 %
1'
b100 +
#369460000000
0!
0'
#369470000000
1!
b101 %
1'
b101 +
#369480000000
0!
0'
#369490000000
1!
0$
b110 %
1'
0*
b110 +
#369500000000
0!
0'
#369510000000
1!
b111 %
1'
b111 +
#369520000000
0!
0'
#369530000000
1!
b1000 %
1'
b1000 +
#369540000000
0!
0'
#369550000000
1!
b1001 %
1'
b1001 +
#369560000000
0!
0'
#369570000000
1!
b0 %
1'
b0 +
#369580000000
1"
1(
#369590000000
0!
0"
b100 &
0'
0(
b100 ,
#369600000000
1!
1$
b1 %
1'
1*
b1 +
#369610000000
0!
0'
#369620000000
1!
b10 %
1'
b10 +
#369630000000
0!
0'
#369640000000
1!
b11 %
1'
b11 +
#369650000000
0!
0'
#369660000000
1!
b100 %
1'
b100 +
#369670000000
0!
0'
#369680000000
1!
b101 %
1'
b101 +
#369690000000
0!
0'
#369700000000
1!
b110 %
1'
b110 +
#369710000000
0!
0'
#369720000000
1!
b111 %
1'
b111 +
#369730000000
0!
0'
#369740000000
1!
0$
b1000 %
1'
0*
b1000 +
#369750000000
0!
0'
#369760000000
1!
b1001 %
1'
b1001 +
#369770000000
0!
0'
#369780000000
1!
b0 %
1'
b0 +
#369790000000
0!
0'
#369800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#369810000000
0!
0'
#369820000000
1!
b10 %
1'
b10 +
#369830000000
0!
0'
#369840000000
1!
b11 %
1'
b11 +
#369850000000
0!
0'
#369860000000
1!
b100 %
1'
b100 +
#369870000000
0!
0'
#369880000000
1!
b101 %
1'
b101 +
#369890000000
0!
0'
#369900000000
1!
0$
b110 %
1'
0*
b110 +
#369910000000
0!
0'
#369920000000
1!
b111 %
1'
b111 +
#369930000000
0!
0'
#369940000000
1!
b1000 %
1'
b1000 +
#369950000000
0!
0'
#369960000000
1!
b1001 %
1'
b1001 +
#369970000000
0!
0'
#369980000000
1!
b0 %
1'
b0 +
#369990000000
0!
0'
#370000000000
1!
1$
b1 %
1'
1*
b1 +
#370010000000
1"
1(
#370020000000
0!
0"
b100 &
0'
0(
b100 ,
#370030000000
1!
b10 %
1'
b10 +
#370040000000
0!
0'
#370050000000
1!
b11 %
1'
b11 +
#370060000000
0!
0'
#370070000000
1!
b100 %
1'
b100 +
#370080000000
0!
0'
#370090000000
1!
b101 %
1'
b101 +
#370100000000
0!
0'
#370110000000
1!
b110 %
1'
b110 +
#370120000000
0!
0'
#370130000000
1!
b111 %
1'
b111 +
#370140000000
0!
0'
#370150000000
1!
0$
b1000 %
1'
0*
b1000 +
#370160000000
0!
0'
#370170000000
1!
b1001 %
1'
b1001 +
#370180000000
0!
0'
#370190000000
1!
b0 %
1'
b0 +
#370200000000
0!
0'
#370210000000
1!
1$
b1 %
1'
1*
b1 +
#370220000000
0!
0'
#370230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#370240000000
0!
0'
#370250000000
1!
b11 %
1'
b11 +
#370260000000
0!
0'
#370270000000
1!
b100 %
1'
b100 +
#370280000000
0!
0'
#370290000000
1!
b101 %
1'
b101 +
#370300000000
0!
0'
#370310000000
1!
0$
b110 %
1'
0*
b110 +
#370320000000
0!
0'
#370330000000
1!
b111 %
1'
b111 +
#370340000000
0!
0'
#370350000000
1!
b1000 %
1'
b1000 +
#370360000000
0!
0'
#370370000000
1!
b1001 %
1'
b1001 +
#370380000000
0!
0'
#370390000000
1!
b0 %
1'
b0 +
#370400000000
0!
0'
#370410000000
1!
1$
b1 %
1'
1*
b1 +
#370420000000
0!
0'
#370430000000
1!
b10 %
1'
b10 +
#370440000000
1"
1(
#370450000000
0!
0"
b100 &
0'
0(
b100 ,
#370460000000
1!
b11 %
1'
b11 +
#370470000000
0!
0'
#370480000000
1!
b100 %
1'
b100 +
#370490000000
0!
0'
#370500000000
1!
b101 %
1'
b101 +
#370510000000
0!
0'
#370520000000
1!
b110 %
1'
b110 +
#370530000000
0!
0'
#370540000000
1!
b111 %
1'
b111 +
#370550000000
0!
0'
#370560000000
1!
0$
b1000 %
1'
0*
b1000 +
#370570000000
0!
0'
#370580000000
1!
b1001 %
1'
b1001 +
#370590000000
0!
0'
#370600000000
1!
b0 %
1'
b0 +
#370610000000
0!
0'
#370620000000
1!
1$
b1 %
1'
1*
b1 +
#370630000000
0!
0'
#370640000000
1!
b10 %
1'
b10 +
#370650000000
0!
0'
#370660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#370670000000
0!
0'
#370680000000
1!
b100 %
1'
b100 +
#370690000000
0!
0'
#370700000000
1!
b101 %
1'
b101 +
#370710000000
0!
0'
#370720000000
1!
0$
b110 %
1'
0*
b110 +
#370730000000
0!
0'
#370740000000
1!
b111 %
1'
b111 +
#370750000000
0!
0'
#370760000000
1!
b1000 %
1'
b1000 +
#370770000000
0!
0'
#370780000000
1!
b1001 %
1'
b1001 +
#370790000000
0!
0'
#370800000000
1!
b0 %
1'
b0 +
#370810000000
0!
0'
#370820000000
1!
1$
b1 %
1'
1*
b1 +
#370830000000
0!
0'
#370840000000
1!
b10 %
1'
b10 +
#370850000000
0!
0'
#370860000000
1!
b11 %
1'
b11 +
#370870000000
1"
1(
#370880000000
0!
0"
b100 &
0'
0(
b100 ,
#370890000000
1!
b100 %
1'
b100 +
#370900000000
0!
0'
#370910000000
1!
b101 %
1'
b101 +
#370920000000
0!
0'
#370930000000
1!
b110 %
1'
b110 +
#370940000000
0!
0'
#370950000000
1!
b111 %
1'
b111 +
#370960000000
0!
0'
#370970000000
1!
0$
b1000 %
1'
0*
b1000 +
#370980000000
0!
0'
#370990000000
1!
b1001 %
1'
b1001 +
#371000000000
0!
0'
#371010000000
1!
b0 %
1'
b0 +
#371020000000
0!
0'
#371030000000
1!
1$
b1 %
1'
1*
b1 +
#371040000000
0!
0'
#371050000000
1!
b10 %
1'
b10 +
#371060000000
0!
0'
#371070000000
1!
b11 %
1'
b11 +
#371080000000
0!
0'
#371090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#371100000000
0!
0'
#371110000000
1!
b101 %
1'
b101 +
#371120000000
0!
0'
#371130000000
1!
0$
b110 %
1'
0*
b110 +
#371140000000
0!
0'
#371150000000
1!
b111 %
1'
b111 +
#371160000000
0!
0'
#371170000000
1!
b1000 %
1'
b1000 +
#371180000000
0!
0'
#371190000000
1!
b1001 %
1'
b1001 +
#371200000000
0!
0'
#371210000000
1!
b0 %
1'
b0 +
#371220000000
0!
0'
#371230000000
1!
1$
b1 %
1'
1*
b1 +
#371240000000
0!
0'
#371250000000
1!
b10 %
1'
b10 +
#371260000000
0!
0'
#371270000000
1!
b11 %
1'
b11 +
#371280000000
0!
0'
#371290000000
1!
b100 %
1'
b100 +
#371300000000
1"
1(
#371310000000
0!
0"
b100 &
0'
0(
b100 ,
#371320000000
1!
b101 %
1'
b101 +
#371330000000
0!
0'
#371340000000
1!
b110 %
1'
b110 +
#371350000000
0!
0'
#371360000000
1!
b111 %
1'
b111 +
#371370000000
0!
0'
#371380000000
1!
0$
b1000 %
1'
0*
b1000 +
#371390000000
0!
0'
#371400000000
1!
b1001 %
1'
b1001 +
#371410000000
0!
0'
#371420000000
1!
b0 %
1'
b0 +
#371430000000
0!
0'
#371440000000
1!
1$
b1 %
1'
1*
b1 +
#371450000000
0!
0'
#371460000000
1!
b10 %
1'
b10 +
#371470000000
0!
0'
#371480000000
1!
b11 %
1'
b11 +
#371490000000
0!
0'
#371500000000
1!
b100 %
1'
b100 +
#371510000000
0!
0'
#371520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#371530000000
0!
0'
#371540000000
1!
0$
b110 %
1'
0*
b110 +
#371550000000
0!
0'
#371560000000
1!
b111 %
1'
b111 +
#371570000000
0!
0'
#371580000000
1!
b1000 %
1'
b1000 +
#371590000000
0!
0'
#371600000000
1!
b1001 %
1'
b1001 +
#371610000000
0!
0'
#371620000000
1!
b0 %
1'
b0 +
#371630000000
0!
0'
#371640000000
1!
1$
b1 %
1'
1*
b1 +
#371650000000
0!
0'
#371660000000
1!
b10 %
1'
b10 +
#371670000000
0!
0'
#371680000000
1!
b11 %
1'
b11 +
#371690000000
0!
0'
#371700000000
1!
b100 %
1'
b100 +
#371710000000
0!
0'
#371720000000
1!
b101 %
1'
b101 +
#371730000000
1"
1(
#371740000000
0!
0"
b100 &
0'
0(
b100 ,
#371750000000
1!
b110 %
1'
b110 +
#371760000000
0!
0'
#371770000000
1!
b111 %
1'
b111 +
#371780000000
0!
0'
#371790000000
1!
0$
b1000 %
1'
0*
b1000 +
#371800000000
0!
0'
#371810000000
1!
b1001 %
1'
b1001 +
#371820000000
0!
0'
#371830000000
1!
b0 %
1'
b0 +
#371840000000
0!
0'
#371850000000
1!
1$
b1 %
1'
1*
b1 +
#371860000000
0!
0'
#371870000000
1!
b10 %
1'
b10 +
#371880000000
0!
0'
#371890000000
1!
b11 %
1'
b11 +
#371900000000
0!
0'
#371910000000
1!
b100 %
1'
b100 +
#371920000000
0!
0'
#371930000000
1!
b101 %
1'
b101 +
#371940000000
0!
0'
#371950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#371960000000
0!
0'
#371970000000
1!
b111 %
1'
b111 +
#371980000000
0!
0'
#371990000000
1!
b1000 %
1'
b1000 +
#372000000000
0!
0'
#372010000000
1!
b1001 %
1'
b1001 +
#372020000000
0!
0'
#372030000000
1!
b0 %
1'
b0 +
#372040000000
0!
0'
#372050000000
1!
1$
b1 %
1'
1*
b1 +
#372060000000
0!
0'
#372070000000
1!
b10 %
1'
b10 +
#372080000000
0!
0'
#372090000000
1!
b11 %
1'
b11 +
#372100000000
0!
0'
#372110000000
1!
b100 %
1'
b100 +
#372120000000
0!
0'
#372130000000
1!
b101 %
1'
b101 +
#372140000000
0!
0'
#372150000000
1!
0$
b110 %
1'
0*
b110 +
#372160000000
1"
1(
#372170000000
0!
0"
b100 &
0'
0(
b100 ,
#372180000000
1!
1$
b111 %
1'
1*
b111 +
#372190000000
0!
0'
#372200000000
1!
0$
b1000 %
1'
0*
b1000 +
#372210000000
0!
0'
#372220000000
1!
b1001 %
1'
b1001 +
#372230000000
0!
0'
#372240000000
1!
b0 %
1'
b0 +
#372250000000
0!
0'
#372260000000
1!
1$
b1 %
1'
1*
b1 +
#372270000000
0!
0'
#372280000000
1!
b10 %
1'
b10 +
#372290000000
0!
0'
#372300000000
1!
b11 %
1'
b11 +
#372310000000
0!
0'
#372320000000
1!
b100 %
1'
b100 +
#372330000000
0!
0'
#372340000000
1!
b101 %
1'
b101 +
#372350000000
0!
0'
#372360000000
1!
b110 %
1'
b110 +
#372370000000
0!
0'
#372380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#372390000000
0!
0'
#372400000000
1!
b1000 %
1'
b1000 +
#372410000000
0!
0'
#372420000000
1!
b1001 %
1'
b1001 +
#372430000000
0!
0'
#372440000000
1!
b0 %
1'
b0 +
#372450000000
0!
0'
#372460000000
1!
1$
b1 %
1'
1*
b1 +
#372470000000
0!
0'
#372480000000
1!
b10 %
1'
b10 +
#372490000000
0!
0'
#372500000000
1!
b11 %
1'
b11 +
#372510000000
0!
0'
#372520000000
1!
b100 %
1'
b100 +
#372530000000
0!
0'
#372540000000
1!
b101 %
1'
b101 +
#372550000000
0!
0'
#372560000000
1!
0$
b110 %
1'
0*
b110 +
#372570000000
0!
0'
#372580000000
1!
b111 %
1'
b111 +
#372590000000
1"
1(
#372600000000
0!
0"
b100 &
0'
0(
b100 ,
#372610000000
1!
b1000 %
1'
b1000 +
#372620000000
0!
0'
#372630000000
1!
b1001 %
1'
b1001 +
#372640000000
0!
0'
#372650000000
1!
b0 %
1'
b0 +
#372660000000
0!
0'
#372670000000
1!
1$
b1 %
1'
1*
b1 +
#372680000000
0!
0'
#372690000000
1!
b10 %
1'
b10 +
#372700000000
0!
0'
#372710000000
1!
b11 %
1'
b11 +
#372720000000
0!
0'
#372730000000
1!
b100 %
1'
b100 +
#372740000000
0!
0'
#372750000000
1!
b101 %
1'
b101 +
#372760000000
0!
0'
#372770000000
1!
b110 %
1'
b110 +
#372780000000
0!
0'
#372790000000
1!
b111 %
1'
b111 +
#372800000000
0!
0'
#372810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#372820000000
0!
0'
#372830000000
1!
b1001 %
1'
b1001 +
#372840000000
0!
0'
#372850000000
1!
b0 %
1'
b0 +
#372860000000
0!
0'
#372870000000
1!
1$
b1 %
1'
1*
b1 +
#372880000000
0!
0'
#372890000000
1!
b10 %
1'
b10 +
#372900000000
0!
0'
#372910000000
1!
b11 %
1'
b11 +
#372920000000
0!
0'
#372930000000
1!
b100 %
1'
b100 +
#372940000000
0!
0'
#372950000000
1!
b101 %
1'
b101 +
#372960000000
0!
0'
#372970000000
1!
0$
b110 %
1'
0*
b110 +
#372980000000
0!
0'
#372990000000
1!
b111 %
1'
b111 +
#373000000000
0!
0'
#373010000000
1!
b1000 %
1'
b1000 +
#373020000000
1"
1(
#373030000000
0!
0"
b100 &
0'
0(
b100 ,
#373040000000
1!
b1001 %
1'
b1001 +
#373050000000
0!
0'
#373060000000
1!
b0 %
1'
b0 +
#373070000000
0!
0'
#373080000000
1!
1$
b1 %
1'
1*
b1 +
#373090000000
0!
0'
#373100000000
1!
b10 %
1'
b10 +
#373110000000
0!
0'
#373120000000
1!
b11 %
1'
b11 +
#373130000000
0!
0'
#373140000000
1!
b100 %
1'
b100 +
#373150000000
0!
0'
#373160000000
1!
b101 %
1'
b101 +
#373170000000
0!
0'
#373180000000
1!
b110 %
1'
b110 +
#373190000000
0!
0'
#373200000000
1!
b111 %
1'
b111 +
#373210000000
0!
0'
#373220000000
1!
0$
b1000 %
1'
0*
b1000 +
#373230000000
0!
0'
#373240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#373250000000
0!
0'
#373260000000
1!
b0 %
1'
b0 +
#373270000000
0!
0'
#373280000000
1!
1$
b1 %
1'
1*
b1 +
#373290000000
0!
0'
#373300000000
1!
b10 %
1'
b10 +
#373310000000
0!
0'
#373320000000
1!
b11 %
1'
b11 +
#373330000000
0!
0'
#373340000000
1!
b100 %
1'
b100 +
#373350000000
0!
0'
#373360000000
1!
b101 %
1'
b101 +
#373370000000
0!
0'
#373380000000
1!
0$
b110 %
1'
0*
b110 +
#373390000000
0!
0'
#373400000000
1!
b111 %
1'
b111 +
#373410000000
0!
0'
#373420000000
1!
b1000 %
1'
b1000 +
#373430000000
0!
0'
#373440000000
1!
b1001 %
1'
b1001 +
#373450000000
1"
1(
#373460000000
0!
0"
b100 &
0'
0(
b100 ,
#373470000000
1!
b0 %
1'
b0 +
#373480000000
0!
0'
#373490000000
1!
1$
b1 %
1'
1*
b1 +
#373500000000
0!
0'
#373510000000
1!
b10 %
1'
b10 +
#373520000000
0!
0'
#373530000000
1!
b11 %
1'
b11 +
#373540000000
0!
0'
#373550000000
1!
b100 %
1'
b100 +
#373560000000
0!
0'
#373570000000
1!
b101 %
1'
b101 +
#373580000000
0!
0'
#373590000000
1!
b110 %
1'
b110 +
#373600000000
0!
0'
#373610000000
1!
b111 %
1'
b111 +
#373620000000
0!
0'
#373630000000
1!
0$
b1000 %
1'
0*
b1000 +
#373640000000
0!
0'
#373650000000
1!
b1001 %
1'
b1001 +
#373660000000
0!
0'
#373670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#373680000000
0!
0'
#373690000000
1!
1$
b1 %
1'
1*
b1 +
#373700000000
0!
0'
#373710000000
1!
b10 %
1'
b10 +
#373720000000
0!
0'
#373730000000
1!
b11 %
1'
b11 +
#373740000000
0!
0'
#373750000000
1!
b100 %
1'
b100 +
#373760000000
0!
0'
#373770000000
1!
b101 %
1'
b101 +
#373780000000
0!
0'
#373790000000
1!
0$
b110 %
1'
0*
b110 +
#373800000000
0!
0'
#373810000000
1!
b111 %
1'
b111 +
#373820000000
0!
0'
#373830000000
1!
b1000 %
1'
b1000 +
#373840000000
0!
0'
#373850000000
1!
b1001 %
1'
b1001 +
#373860000000
0!
0'
#373870000000
1!
b0 %
1'
b0 +
#373880000000
1"
1(
#373890000000
0!
0"
b100 &
0'
0(
b100 ,
#373900000000
1!
1$
b1 %
1'
1*
b1 +
#373910000000
0!
0'
#373920000000
1!
b10 %
1'
b10 +
#373930000000
0!
0'
#373940000000
1!
b11 %
1'
b11 +
#373950000000
0!
0'
#373960000000
1!
b100 %
1'
b100 +
#373970000000
0!
0'
#373980000000
1!
b101 %
1'
b101 +
#373990000000
0!
0'
#374000000000
1!
b110 %
1'
b110 +
#374010000000
0!
0'
#374020000000
1!
b111 %
1'
b111 +
#374030000000
0!
0'
#374040000000
1!
0$
b1000 %
1'
0*
b1000 +
#374050000000
0!
0'
#374060000000
1!
b1001 %
1'
b1001 +
#374070000000
0!
0'
#374080000000
1!
b0 %
1'
b0 +
#374090000000
0!
0'
#374100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#374110000000
0!
0'
#374120000000
1!
b10 %
1'
b10 +
#374130000000
0!
0'
#374140000000
1!
b11 %
1'
b11 +
#374150000000
0!
0'
#374160000000
1!
b100 %
1'
b100 +
#374170000000
0!
0'
#374180000000
1!
b101 %
1'
b101 +
#374190000000
0!
0'
#374200000000
1!
0$
b110 %
1'
0*
b110 +
#374210000000
0!
0'
#374220000000
1!
b111 %
1'
b111 +
#374230000000
0!
0'
#374240000000
1!
b1000 %
1'
b1000 +
#374250000000
0!
0'
#374260000000
1!
b1001 %
1'
b1001 +
#374270000000
0!
0'
#374280000000
1!
b0 %
1'
b0 +
#374290000000
0!
0'
#374300000000
1!
1$
b1 %
1'
1*
b1 +
#374310000000
1"
1(
#374320000000
0!
0"
b100 &
0'
0(
b100 ,
#374330000000
1!
b10 %
1'
b10 +
#374340000000
0!
0'
#374350000000
1!
b11 %
1'
b11 +
#374360000000
0!
0'
#374370000000
1!
b100 %
1'
b100 +
#374380000000
0!
0'
#374390000000
1!
b101 %
1'
b101 +
#374400000000
0!
0'
#374410000000
1!
b110 %
1'
b110 +
#374420000000
0!
0'
#374430000000
1!
b111 %
1'
b111 +
#374440000000
0!
0'
#374450000000
1!
0$
b1000 %
1'
0*
b1000 +
#374460000000
0!
0'
#374470000000
1!
b1001 %
1'
b1001 +
#374480000000
0!
0'
#374490000000
1!
b0 %
1'
b0 +
#374500000000
0!
0'
#374510000000
1!
1$
b1 %
1'
1*
b1 +
#374520000000
0!
0'
#374530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#374540000000
0!
0'
#374550000000
1!
b11 %
1'
b11 +
#374560000000
0!
0'
#374570000000
1!
b100 %
1'
b100 +
#374580000000
0!
0'
#374590000000
1!
b101 %
1'
b101 +
#374600000000
0!
0'
#374610000000
1!
0$
b110 %
1'
0*
b110 +
#374620000000
0!
0'
#374630000000
1!
b111 %
1'
b111 +
#374640000000
0!
0'
#374650000000
1!
b1000 %
1'
b1000 +
#374660000000
0!
0'
#374670000000
1!
b1001 %
1'
b1001 +
#374680000000
0!
0'
#374690000000
1!
b0 %
1'
b0 +
#374700000000
0!
0'
#374710000000
1!
1$
b1 %
1'
1*
b1 +
#374720000000
0!
0'
#374730000000
1!
b10 %
1'
b10 +
#374740000000
1"
1(
#374750000000
0!
0"
b100 &
0'
0(
b100 ,
#374760000000
1!
b11 %
1'
b11 +
#374770000000
0!
0'
#374780000000
1!
b100 %
1'
b100 +
#374790000000
0!
0'
#374800000000
1!
b101 %
1'
b101 +
#374810000000
0!
0'
#374820000000
1!
b110 %
1'
b110 +
#374830000000
0!
0'
#374840000000
1!
b111 %
1'
b111 +
#374850000000
0!
0'
#374860000000
1!
0$
b1000 %
1'
0*
b1000 +
#374870000000
0!
0'
#374880000000
1!
b1001 %
1'
b1001 +
#374890000000
0!
0'
#374900000000
1!
b0 %
1'
b0 +
#374910000000
0!
0'
#374920000000
1!
1$
b1 %
1'
1*
b1 +
#374930000000
0!
0'
#374940000000
1!
b10 %
1'
b10 +
#374950000000
0!
0'
#374960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#374970000000
0!
0'
#374980000000
1!
b100 %
1'
b100 +
#374990000000
0!
0'
#375000000000
1!
b101 %
1'
b101 +
#375010000000
0!
0'
#375020000000
1!
0$
b110 %
1'
0*
b110 +
#375030000000
0!
0'
#375040000000
1!
b111 %
1'
b111 +
#375050000000
0!
0'
#375060000000
1!
b1000 %
1'
b1000 +
#375070000000
0!
0'
#375080000000
1!
b1001 %
1'
b1001 +
#375090000000
0!
0'
#375100000000
1!
b0 %
1'
b0 +
#375110000000
0!
0'
#375120000000
1!
1$
b1 %
1'
1*
b1 +
#375130000000
0!
0'
#375140000000
1!
b10 %
1'
b10 +
#375150000000
0!
0'
#375160000000
1!
b11 %
1'
b11 +
#375170000000
1"
1(
#375180000000
0!
0"
b100 &
0'
0(
b100 ,
#375190000000
1!
b100 %
1'
b100 +
#375200000000
0!
0'
#375210000000
1!
b101 %
1'
b101 +
#375220000000
0!
0'
#375230000000
1!
b110 %
1'
b110 +
#375240000000
0!
0'
#375250000000
1!
b111 %
1'
b111 +
#375260000000
0!
0'
#375270000000
1!
0$
b1000 %
1'
0*
b1000 +
#375280000000
0!
0'
#375290000000
1!
b1001 %
1'
b1001 +
#375300000000
0!
0'
#375310000000
1!
b0 %
1'
b0 +
#375320000000
0!
0'
#375330000000
1!
1$
b1 %
1'
1*
b1 +
#375340000000
0!
0'
#375350000000
1!
b10 %
1'
b10 +
#375360000000
0!
0'
#375370000000
1!
b11 %
1'
b11 +
#375380000000
0!
0'
#375390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#375400000000
0!
0'
#375410000000
1!
b101 %
1'
b101 +
#375420000000
0!
0'
#375430000000
1!
0$
b110 %
1'
0*
b110 +
#375440000000
0!
0'
#375450000000
1!
b111 %
1'
b111 +
#375460000000
0!
0'
#375470000000
1!
b1000 %
1'
b1000 +
#375480000000
0!
0'
#375490000000
1!
b1001 %
1'
b1001 +
#375500000000
0!
0'
#375510000000
1!
b0 %
1'
b0 +
#375520000000
0!
0'
#375530000000
1!
1$
b1 %
1'
1*
b1 +
#375540000000
0!
0'
#375550000000
1!
b10 %
1'
b10 +
#375560000000
0!
0'
#375570000000
1!
b11 %
1'
b11 +
#375580000000
0!
0'
#375590000000
1!
b100 %
1'
b100 +
#375600000000
1"
1(
#375610000000
0!
0"
b100 &
0'
0(
b100 ,
#375620000000
1!
b101 %
1'
b101 +
#375630000000
0!
0'
#375640000000
1!
b110 %
1'
b110 +
#375650000000
0!
0'
#375660000000
1!
b111 %
1'
b111 +
#375670000000
0!
0'
#375680000000
1!
0$
b1000 %
1'
0*
b1000 +
#375690000000
0!
0'
#375700000000
1!
b1001 %
1'
b1001 +
#375710000000
0!
0'
#375720000000
1!
b0 %
1'
b0 +
#375730000000
0!
0'
#375740000000
1!
1$
b1 %
1'
1*
b1 +
#375750000000
0!
0'
#375760000000
1!
b10 %
1'
b10 +
#375770000000
0!
0'
#375780000000
1!
b11 %
1'
b11 +
#375790000000
0!
0'
#375800000000
1!
b100 %
1'
b100 +
#375810000000
0!
0'
#375820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#375830000000
0!
0'
#375840000000
1!
0$
b110 %
1'
0*
b110 +
#375850000000
0!
0'
#375860000000
1!
b111 %
1'
b111 +
#375870000000
0!
0'
#375880000000
1!
b1000 %
1'
b1000 +
#375890000000
0!
0'
#375900000000
1!
b1001 %
1'
b1001 +
#375910000000
0!
0'
#375920000000
1!
b0 %
1'
b0 +
#375930000000
0!
0'
#375940000000
1!
1$
b1 %
1'
1*
b1 +
#375950000000
0!
0'
#375960000000
1!
b10 %
1'
b10 +
#375970000000
0!
0'
#375980000000
1!
b11 %
1'
b11 +
#375990000000
0!
0'
#376000000000
1!
b100 %
1'
b100 +
#376010000000
0!
0'
#376020000000
1!
b101 %
1'
b101 +
#376030000000
1"
1(
#376040000000
0!
0"
b100 &
0'
0(
b100 ,
#376050000000
1!
b110 %
1'
b110 +
#376060000000
0!
0'
#376070000000
1!
b111 %
1'
b111 +
#376080000000
0!
0'
#376090000000
1!
0$
b1000 %
1'
0*
b1000 +
#376100000000
0!
0'
#376110000000
1!
b1001 %
1'
b1001 +
#376120000000
0!
0'
#376130000000
1!
b0 %
1'
b0 +
#376140000000
0!
0'
#376150000000
1!
1$
b1 %
1'
1*
b1 +
#376160000000
0!
0'
#376170000000
1!
b10 %
1'
b10 +
#376180000000
0!
0'
#376190000000
1!
b11 %
1'
b11 +
#376200000000
0!
0'
#376210000000
1!
b100 %
1'
b100 +
#376220000000
0!
0'
#376230000000
1!
b101 %
1'
b101 +
#376240000000
0!
0'
#376250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#376260000000
0!
0'
#376270000000
1!
b111 %
1'
b111 +
#376280000000
0!
0'
#376290000000
1!
b1000 %
1'
b1000 +
#376300000000
0!
0'
#376310000000
1!
b1001 %
1'
b1001 +
#376320000000
0!
0'
#376330000000
1!
b0 %
1'
b0 +
#376340000000
0!
0'
#376350000000
1!
1$
b1 %
1'
1*
b1 +
#376360000000
0!
0'
#376370000000
1!
b10 %
1'
b10 +
#376380000000
0!
0'
#376390000000
1!
b11 %
1'
b11 +
#376400000000
0!
0'
#376410000000
1!
b100 %
1'
b100 +
#376420000000
0!
0'
#376430000000
1!
b101 %
1'
b101 +
#376440000000
0!
0'
#376450000000
1!
0$
b110 %
1'
0*
b110 +
#376460000000
1"
1(
#376470000000
0!
0"
b100 &
0'
0(
b100 ,
#376480000000
1!
1$
b111 %
1'
1*
b111 +
#376490000000
0!
0'
#376500000000
1!
0$
b1000 %
1'
0*
b1000 +
#376510000000
0!
0'
#376520000000
1!
b1001 %
1'
b1001 +
#376530000000
0!
0'
#376540000000
1!
b0 %
1'
b0 +
#376550000000
0!
0'
#376560000000
1!
1$
b1 %
1'
1*
b1 +
#376570000000
0!
0'
#376580000000
1!
b10 %
1'
b10 +
#376590000000
0!
0'
#376600000000
1!
b11 %
1'
b11 +
#376610000000
0!
0'
#376620000000
1!
b100 %
1'
b100 +
#376630000000
0!
0'
#376640000000
1!
b101 %
1'
b101 +
#376650000000
0!
0'
#376660000000
1!
b110 %
1'
b110 +
#376670000000
0!
0'
#376680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#376690000000
0!
0'
#376700000000
1!
b1000 %
1'
b1000 +
#376710000000
0!
0'
#376720000000
1!
b1001 %
1'
b1001 +
#376730000000
0!
0'
#376740000000
1!
b0 %
1'
b0 +
#376750000000
0!
0'
#376760000000
1!
1$
b1 %
1'
1*
b1 +
#376770000000
0!
0'
#376780000000
1!
b10 %
1'
b10 +
#376790000000
0!
0'
#376800000000
1!
b11 %
1'
b11 +
#376810000000
0!
0'
#376820000000
1!
b100 %
1'
b100 +
#376830000000
0!
0'
#376840000000
1!
b101 %
1'
b101 +
#376850000000
0!
0'
#376860000000
1!
0$
b110 %
1'
0*
b110 +
#376870000000
0!
0'
#376880000000
1!
b111 %
1'
b111 +
#376890000000
1"
1(
#376900000000
0!
0"
b100 &
0'
0(
b100 ,
#376910000000
1!
b1000 %
1'
b1000 +
#376920000000
0!
0'
#376930000000
1!
b1001 %
1'
b1001 +
#376940000000
0!
0'
#376950000000
1!
b0 %
1'
b0 +
#376960000000
0!
0'
#376970000000
1!
1$
b1 %
1'
1*
b1 +
#376980000000
0!
0'
#376990000000
1!
b10 %
1'
b10 +
#377000000000
0!
0'
#377010000000
1!
b11 %
1'
b11 +
#377020000000
0!
0'
#377030000000
1!
b100 %
1'
b100 +
#377040000000
0!
0'
#377050000000
1!
b101 %
1'
b101 +
#377060000000
0!
0'
#377070000000
1!
b110 %
1'
b110 +
#377080000000
0!
0'
#377090000000
1!
b111 %
1'
b111 +
#377100000000
0!
0'
#377110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#377120000000
0!
0'
#377130000000
1!
b1001 %
1'
b1001 +
#377140000000
0!
0'
#377150000000
1!
b0 %
1'
b0 +
#377160000000
0!
0'
#377170000000
1!
1$
b1 %
1'
1*
b1 +
#377180000000
0!
0'
#377190000000
1!
b10 %
1'
b10 +
#377200000000
0!
0'
#377210000000
1!
b11 %
1'
b11 +
#377220000000
0!
0'
#377230000000
1!
b100 %
1'
b100 +
#377240000000
0!
0'
#377250000000
1!
b101 %
1'
b101 +
#377260000000
0!
0'
#377270000000
1!
0$
b110 %
1'
0*
b110 +
#377280000000
0!
0'
#377290000000
1!
b111 %
1'
b111 +
#377300000000
0!
0'
#377310000000
1!
b1000 %
1'
b1000 +
#377320000000
1"
1(
#377330000000
0!
0"
b100 &
0'
0(
b100 ,
#377340000000
1!
b1001 %
1'
b1001 +
#377350000000
0!
0'
#377360000000
1!
b0 %
1'
b0 +
#377370000000
0!
0'
#377380000000
1!
1$
b1 %
1'
1*
b1 +
#377390000000
0!
0'
#377400000000
1!
b10 %
1'
b10 +
#377410000000
0!
0'
#377420000000
1!
b11 %
1'
b11 +
#377430000000
0!
0'
#377440000000
1!
b100 %
1'
b100 +
#377450000000
0!
0'
#377460000000
1!
b101 %
1'
b101 +
#377470000000
0!
0'
#377480000000
1!
b110 %
1'
b110 +
#377490000000
0!
0'
#377500000000
1!
b111 %
1'
b111 +
#377510000000
0!
0'
#377520000000
1!
0$
b1000 %
1'
0*
b1000 +
#377530000000
0!
0'
#377540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#377550000000
0!
0'
#377560000000
1!
b0 %
1'
b0 +
#377570000000
0!
0'
#377580000000
1!
1$
b1 %
1'
1*
b1 +
#377590000000
0!
0'
#377600000000
1!
b10 %
1'
b10 +
#377610000000
0!
0'
#377620000000
1!
b11 %
1'
b11 +
#377630000000
0!
0'
#377640000000
1!
b100 %
1'
b100 +
#377650000000
0!
0'
#377660000000
1!
b101 %
1'
b101 +
#377670000000
0!
0'
#377680000000
1!
0$
b110 %
1'
0*
b110 +
#377690000000
0!
0'
#377700000000
1!
b111 %
1'
b111 +
#377710000000
0!
0'
#377720000000
1!
b1000 %
1'
b1000 +
#377730000000
0!
0'
#377740000000
1!
b1001 %
1'
b1001 +
#377750000000
1"
1(
#377760000000
0!
0"
b100 &
0'
0(
b100 ,
#377770000000
1!
b0 %
1'
b0 +
#377780000000
0!
0'
#377790000000
1!
1$
b1 %
1'
1*
b1 +
#377800000000
0!
0'
#377810000000
1!
b10 %
1'
b10 +
#377820000000
0!
0'
#377830000000
1!
b11 %
1'
b11 +
#377840000000
0!
0'
#377850000000
1!
b100 %
1'
b100 +
#377860000000
0!
0'
#377870000000
1!
b101 %
1'
b101 +
#377880000000
0!
0'
#377890000000
1!
b110 %
1'
b110 +
#377900000000
0!
0'
#377910000000
1!
b111 %
1'
b111 +
#377920000000
0!
0'
#377930000000
1!
0$
b1000 %
1'
0*
b1000 +
#377940000000
0!
0'
#377950000000
1!
b1001 %
1'
b1001 +
#377960000000
0!
0'
#377970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#377980000000
0!
0'
#377990000000
1!
1$
b1 %
1'
1*
b1 +
#378000000000
0!
0'
#378010000000
1!
b10 %
1'
b10 +
#378020000000
0!
0'
#378030000000
1!
b11 %
1'
b11 +
#378040000000
0!
0'
#378050000000
1!
b100 %
1'
b100 +
#378060000000
0!
0'
#378070000000
1!
b101 %
1'
b101 +
#378080000000
0!
0'
#378090000000
1!
0$
b110 %
1'
0*
b110 +
#378100000000
0!
0'
#378110000000
1!
b111 %
1'
b111 +
#378120000000
0!
0'
#378130000000
1!
b1000 %
1'
b1000 +
#378140000000
0!
0'
#378150000000
1!
b1001 %
1'
b1001 +
#378160000000
0!
0'
#378170000000
1!
b0 %
1'
b0 +
#378180000000
1"
1(
#378190000000
0!
0"
b100 &
0'
0(
b100 ,
#378200000000
1!
1$
b1 %
1'
1*
b1 +
#378210000000
0!
0'
#378220000000
1!
b10 %
1'
b10 +
#378230000000
0!
0'
#378240000000
1!
b11 %
1'
b11 +
#378250000000
0!
0'
#378260000000
1!
b100 %
1'
b100 +
#378270000000
0!
0'
#378280000000
1!
b101 %
1'
b101 +
#378290000000
0!
0'
#378300000000
1!
b110 %
1'
b110 +
#378310000000
0!
0'
#378320000000
1!
b111 %
1'
b111 +
#378330000000
0!
0'
#378340000000
1!
0$
b1000 %
1'
0*
b1000 +
#378350000000
0!
0'
#378360000000
1!
b1001 %
1'
b1001 +
#378370000000
0!
0'
#378380000000
1!
b0 %
1'
b0 +
#378390000000
0!
0'
#378400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#378410000000
0!
0'
#378420000000
1!
b10 %
1'
b10 +
#378430000000
0!
0'
#378440000000
1!
b11 %
1'
b11 +
#378450000000
0!
0'
#378460000000
1!
b100 %
1'
b100 +
#378470000000
0!
0'
#378480000000
1!
b101 %
1'
b101 +
#378490000000
0!
0'
#378500000000
1!
0$
b110 %
1'
0*
b110 +
#378510000000
0!
0'
#378520000000
1!
b111 %
1'
b111 +
#378530000000
0!
0'
#378540000000
1!
b1000 %
1'
b1000 +
#378550000000
0!
0'
#378560000000
1!
b1001 %
1'
b1001 +
#378570000000
0!
0'
#378580000000
1!
b0 %
1'
b0 +
#378590000000
0!
0'
#378600000000
1!
1$
b1 %
1'
1*
b1 +
#378610000000
1"
1(
#378620000000
0!
0"
b100 &
0'
0(
b100 ,
#378630000000
1!
b10 %
1'
b10 +
#378640000000
0!
0'
#378650000000
1!
b11 %
1'
b11 +
#378660000000
0!
0'
#378670000000
1!
b100 %
1'
b100 +
#378680000000
0!
0'
#378690000000
1!
b101 %
1'
b101 +
#378700000000
0!
0'
#378710000000
1!
b110 %
1'
b110 +
#378720000000
0!
0'
#378730000000
1!
b111 %
1'
b111 +
#378740000000
0!
0'
#378750000000
1!
0$
b1000 %
1'
0*
b1000 +
#378760000000
0!
0'
#378770000000
1!
b1001 %
1'
b1001 +
#378780000000
0!
0'
#378790000000
1!
b0 %
1'
b0 +
#378800000000
0!
0'
#378810000000
1!
1$
b1 %
1'
1*
b1 +
#378820000000
0!
0'
#378830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#378840000000
0!
0'
#378850000000
1!
b11 %
1'
b11 +
#378860000000
0!
0'
#378870000000
1!
b100 %
1'
b100 +
#378880000000
0!
0'
#378890000000
1!
b101 %
1'
b101 +
#378900000000
0!
0'
#378910000000
1!
0$
b110 %
1'
0*
b110 +
#378920000000
0!
0'
#378930000000
1!
b111 %
1'
b111 +
#378940000000
0!
0'
#378950000000
1!
b1000 %
1'
b1000 +
#378960000000
0!
0'
#378970000000
1!
b1001 %
1'
b1001 +
#378980000000
0!
0'
#378990000000
1!
b0 %
1'
b0 +
#379000000000
0!
0'
#379010000000
1!
1$
b1 %
1'
1*
b1 +
#379020000000
0!
0'
#379030000000
1!
b10 %
1'
b10 +
#379040000000
1"
1(
#379050000000
0!
0"
b100 &
0'
0(
b100 ,
#379060000000
1!
b11 %
1'
b11 +
#379070000000
0!
0'
#379080000000
1!
b100 %
1'
b100 +
#379090000000
0!
0'
#379100000000
1!
b101 %
1'
b101 +
#379110000000
0!
0'
#379120000000
1!
b110 %
1'
b110 +
#379130000000
0!
0'
#379140000000
1!
b111 %
1'
b111 +
#379150000000
0!
0'
#379160000000
1!
0$
b1000 %
1'
0*
b1000 +
#379170000000
0!
0'
#379180000000
1!
b1001 %
1'
b1001 +
#379190000000
0!
0'
#379200000000
1!
b0 %
1'
b0 +
#379210000000
0!
0'
#379220000000
1!
1$
b1 %
1'
1*
b1 +
#379230000000
0!
0'
#379240000000
1!
b10 %
1'
b10 +
#379250000000
0!
0'
#379260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#379270000000
0!
0'
#379280000000
1!
b100 %
1'
b100 +
#379290000000
0!
0'
#379300000000
1!
b101 %
1'
b101 +
#379310000000
0!
0'
#379320000000
1!
0$
b110 %
1'
0*
b110 +
#379330000000
0!
0'
#379340000000
1!
b111 %
1'
b111 +
#379350000000
0!
0'
#379360000000
1!
b1000 %
1'
b1000 +
#379370000000
0!
0'
#379380000000
1!
b1001 %
1'
b1001 +
#379390000000
0!
0'
#379400000000
1!
b0 %
1'
b0 +
#379410000000
0!
0'
#379420000000
1!
1$
b1 %
1'
1*
b1 +
#379430000000
0!
0'
#379440000000
1!
b10 %
1'
b10 +
#379450000000
0!
0'
#379460000000
1!
b11 %
1'
b11 +
#379470000000
1"
1(
#379480000000
0!
0"
b100 &
0'
0(
b100 ,
#379490000000
1!
b100 %
1'
b100 +
#379500000000
0!
0'
#379510000000
1!
b101 %
1'
b101 +
#379520000000
0!
0'
#379530000000
1!
b110 %
1'
b110 +
#379540000000
0!
0'
#379550000000
1!
b111 %
1'
b111 +
#379560000000
0!
0'
#379570000000
1!
0$
b1000 %
1'
0*
b1000 +
#379580000000
0!
0'
#379590000000
1!
b1001 %
1'
b1001 +
#379600000000
0!
0'
#379610000000
1!
b0 %
1'
b0 +
#379620000000
0!
0'
#379630000000
1!
1$
b1 %
1'
1*
b1 +
#379640000000
0!
0'
#379650000000
1!
b10 %
1'
b10 +
#379660000000
0!
0'
#379670000000
1!
b11 %
1'
b11 +
#379680000000
0!
0'
#379690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#379700000000
0!
0'
#379710000000
1!
b101 %
1'
b101 +
#379720000000
0!
0'
#379730000000
1!
0$
b110 %
1'
0*
b110 +
#379740000000
0!
0'
#379750000000
1!
b111 %
1'
b111 +
#379760000000
0!
0'
#379770000000
1!
b1000 %
1'
b1000 +
#379780000000
0!
0'
#379790000000
1!
b1001 %
1'
b1001 +
#379800000000
0!
0'
#379810000000
1!
b0 %
1'
b0 +
#379820000000
0!
0'
#379830000000
1!
1$
b1 %
1'
1*
b1 +
#379840000000
0!
0'
#379850000000
1!
b10 %
1'
b10 +
#379860000000
0!
0'
#379870000000
1!
b11 %
1'
b11 +
#379880000000
0!
0'
#379890000000
1!
b100 %
1'
b100 +
#379900000000
1"
1(
#379910000000
0!
0"
b100 &
0'
0(
b100 ,
#379920000000
1!
b101 %
1'
b101 +
#379930000000
0!
0'
#379940000000
1!
b110 %
1'
b110 +
#379950000000
0!
0'
#379960000000
1!
b111 %
1'
b111 +
#379970000000
0!
0'
#379980000000
1!
0$
b1000 %
1'
0*
b1000 +
#379990000000
0!
0'
#380000000000
1!
b1001 %
1'
b1001 +
#380010000000
0!
0'
#380020000000
1!
b0 %
1'
b0 +
#380030000000
0!
0'
#380040000000
1!
1$
b1 %
1'
1*
b1 +
#380050000000
0!
0'
#380060000000
1!
b10 %
1'
b10 +
#380070000000
0!
0'
#380080000000
1!
b11 %
1'
b11 +
#380090000000
0!
0'
#380100000000
1!
b100 %
1'
b100 +
#380110000000
0!
0'
#380120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#380130000000
0!
0'
#380140000000
1!
0$
b110 %
1'
0*
b110 +
#380150000000
0!
0'
#380160000000
1!
b111 %
1'
b111 +
#380170000000
0!
0'
#380180000000
1!
b1000 %
1'
b1000 +
#380190000000
0!
0'
#380200000000
1!
b1001 %
1'
b1001 +
#380210000000
0!
0'
#380220000000
1!
b0 %
1'
b0 +
#380230000000
0!
0'
#380240000000
1!
1$
b1 %
1'
1*
b1 +
#380250000000
0!
0'
#380260000000
1!
b10 %
1'
b10 +
#380270000000
0!
0'
#380280000000
1!
b11 %
1'
b11 +
#380290000000
0!
0'
#380300000000
1!
b100 %
1'
b100 +
#380310000000
0!
0'
#380320000000
1!
b101 %
1'
b101 +
#380330000000
1"
1(
#380340000000
0!
0"
b100 &
0'
0(
b100 ,
#380350000000
1!
b110 %
1'
b110 +
#380360000000
0!
0'
#380370000000
1!
b111 %
1'
b111 +
#380380000000
0!
0'
#380390000000
1!
0$
b1000 %
1'
0*
b1000 +
#380400000000
0!
0'
#380410000000
1!
b1001 %
1'
b1001 +
#380420000000
0!
0'
#380430000000
1!
b0 %
1'
b0 +
#380440000000
0!
0'
#380450000000
1!
1$
b1 %
1'
1*
b1 +
#380460000000
0!
0'
#380470000000
1!
b10 %
1'
b10 +
#380480000000
0!
0'
#380490000000
1!
b11 %
1'
b11 +
#380500000000
0!
0'
#380510000000
1!
b100 %
1'
b100 +
#380520000000
0!
0'
#380530000000
1!
b101 %
1'
b101 +
#380540000000
0!
0'
#380550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#380560000000
0!
0'
#380570000000
1!
b111 %
1'
b111 +
#380580000000
0!
0'
#380590000000
1!
b1000 %
1'
b1000 +
#380600000000
0!
0'
#380610000000
1!
b1001 %
1'
b1001 +
#380620000000
0!
0'
#380630000000
1!
b0 %
1'
b0 +
#380640000000
0!
0'
#380650000000
1!
1$
b1 %
1'
1*
b1 +
#380660000000
0!
0'
#380670000000
1!
b10 %
1'
b10 +
#380680000000
0!
0'
#380690000000
1!
b11 %
1'
b11 +
#380700000000
0!
0'
#380710000000
1!
b100 %
1'
b100 +
#380720000000
0!
0'
#380730000000
1!
b101 %
1'
b101 +
#380740000000
0!
0'
#380750000000
1!
0$
b110 %
1'
0*
b110 +
#380760000000
1"
1(
#380770000000
0!
0"
b100 &
0'
0(
b100 ,
#380780000000
1!
1$
b111 %
1'
1*
b111 +
#380790000000
0!
0'
#380800000000
1!
0$
b1000 %
1'
0*
b1000 +
#380810000000
0!
0'
#380820000000
1!
b1001 %
1'
b1001 +
#380830000000
0!
0'
#380840000000
1!
b0 %
1'
b0 +
#380850000000
0!
0'
#380860000000
1!
1$
b1 %
1'
1*
b1 +
#380870000000
0!
0'
#380880000000
1!
b10 %
1'
b10 +
#380890000000
0!
0'
#380900000000
1!
b11 %
1'
b11 +
#380910000000
0!
0'
#380920000000
1!
b100 %
1'
b100 +
#380930000000
0!
0'
#380940000000
1!
b101 %
1'
b101 +
#380950000000
0!
0'
#380960000000
1!
b110 %
1'
b110 +
#380970000000
0!
0'
#380980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#380990000000
0!
0'
#381000000000
1!
b1000 %
1'
b1000 +
#381010000000
0!
0'
#381020000000
1!
b1001 %
1'
b1001 +
#381030000000
0!
0'
#381040000000
1!
b0 %
1'
b0 +
#381050000000
0!
0'
#381060000000
1!
1$
b1 %
1'
1*
b1 +
#381070000000
0!
0'
#381080000000
1!
b10 %
1'
b10 +
#381090000000
0!
0'
#381100000000
1!
b11 %
1'
b11 +
#381110000000
0!
0'
#381120000000
1!
b100 %
1'
b100 +
#381130000000
0!
0'
#381140000000
1!
b101 %
1'
b101 +
#381150000000
0!
0'
#381160000000
1!
0$
b110 %
1'
0*
b110 +
#381170000000
0!
0'
#381180000000
1!
b111 %
1'
b111 +
#381190000000
1"
1(
#381200000000
0!
0"
b100 &
0'
0(
b100 ,
#381210000000
1!
b1000 %
1'
b1000 +
#381220000000
0!
0'
#381230000000
1!
b1001 %
1'
b1001 +
#381240000000
0!
0'
#381250000000
1!
b0 %
1'
b0 +
#381260000000
0!
0'
#381270000000
1!
1$
b1 %
1'
1*
b1 +
#381280000000
0!
0'
#381290000000
1!
b10 %
1'
b10 +
#381300000000
0!
0'
#381310000000
1!
b11 %
1'
b11 +
#381320000000
0!
0'
#381330000000
1!
b100 %
1'
b100 +
#381340000000
0!
0'
#381350000000
1!
b101 %
1'
b101 +
#381360000000
0!
0'
#381370000000
1!
b110 %
1'
b110 +
#381380000000
0!
0'
#381390000000
1!
b111 %
1'
b111 +
#381400000000
0!
0'
#381410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#381420000000
0!
0'
#381430000000
1!
b1001 %
1'
b1001 +
#381440000000
0!
0'
#381450000000
1!
b0 %
1'
b0 +
#381460000000
0!
0'
#381470000000
1!
1$
b1 %
1'
1*
b1 +
#381480000000
0!
0'
#381490000000
1!
b10 %
1'
b10 +
#381500000000
0!
0'
#381510000000
1!
b11 %
1'
b11 +
#381520000000
0!
0'
#381530000000
1!
b100 %
1'
b100 +
#381540000000
0!
0'
#381550000000
1!
b101 %
1'
b101 +
#381560000000
0!
0'
#381570000000
1!
0$
b110 %
1'
0*
b110 +
#381580000000
0!
0'
#381590000000
1!
b111 %
1'
b111 +
#381600000000
0!
0'
#381610000000
1!
b1000 %
1'
b1000 +
#381620000000
1"
1(
#381630000000
0!
0"
b100 &
0'
0(
b100 ,
#381640000000
1!
b1001 %
1'
b1001 +
#381650000000
0!
0'
#381660000000
1!
b0 %
1'
b0 +
#381670000000
0!
0'
#381680000000
1!
1$
b1 %
1'
1*
b1 +
#381690000000
0!
0'
#381700000000
1!
b10 %
1'
b10 +
#381710000000
0!
0'
#381720000000
1!
b11 %
1'
b11 +
#381730000000
0!
0'
#381740000000
1!
b100 %
1'
b100 +
#381750000000
0!
0'
#381760000000
1!
b101 %
1'
b101 +
#381770000000
0!
0'
#381780000000
1!
b110 %
1'
b110 +
#381790000000
0!
0'
#381800000000
1!
b111 %
1'
b111 +
#381810000000
0!
0'
#381820000000
1!
0$
b1000 %
1'
0*
b1000 +
#381830000000
0!
0'
#381840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#381850000000
0!
0'
#381860000000
1!
b0 %
1'
b0 +
#381870000000
0!
0'
#381880000000
1!
1$
b1 %
1'
1*
b1 +
#381890000000
0!
0'
#381900000000
1!
b10 %
1'
b10 +
#381910000000
0!
0'
#381920000000
1!
b11 %
1'
b11 +
#381930000000
0!
0'
#381940000000
1!
b100 %
1'
b100 +
#381950000000
0!
0'
#381960000000
1!
b101 %
1'
b101 +
#381970000000
0!
0'
#381980000000
1!
0$
b110 %
1'
0*
b110 +
#381990000000
0!
0'
#382000000000
1!
b111 %
1'
b111 +
#382010000000
0!
0'
#382020000000
1!
b1000 %
1'
b1000 +
#382030000000
0!
0'
#382040000000
1!
b1001 %
1'
b1001 +
#382050000000
1"
1(
#382060000000
0!
0"
b100 &
0'
0(
b100 ,
#382070000000
1!
b0 %
1'
b0 +
#382080000000
0!
0'
#382090000000
1!
1$
b1 %
1'
1*
b1 +
#382100000000
0!
0'
#382110000000
1!
b10 %
1'
b10 +
#382120000000
0!
0'
#382130000000
1!
b11 %
1'
b11 +
#382140000000
0!
0'
#382150000000
1!
b100 %
1'
b100 +
#382160000000
0!
0'
#382170000000
1!
b101 %
1'
b101 +
#382180000000
0!
0'
#382190000000
1!
b110 %
1'
b110 +
#382200000000
0!
0'
#382210000000
1!
b111 %
1'
b111 +
#382220000000
0!
0'
#382230000000
1!
0$
b1000 %
1'
0*
b1000 +
#382240000000
0!
0'
#382250000000
1!
b1001 %
1'
b1001 +
#382260000000
0!
0'
#382270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#382280000000
0!
0'
#382290000000
1!
1$
b1 %
1'
1*
b1 +
#382300000000
0!
0'
#382310000000
1!
b10 %
1'
b10 +
#382320000000
0!
0'
#382330000000
1!
b11 %
1'
b11 +
#382340000000
0!
0'
#382350000000
1!
b100 %
1'
b100 +
#382360000000
0!
0'
#382370000000
1!
b101 %
1'
b101 +
#382380000000
0!
0'
#382390000000
1!
0$
b110 %
1'
0*
b110 +
#382400000000
0!
0'
#382410000000
1!
b111 %
1'
b111 +
#382420000000
0!
0'
#382430000000
1!
b1000 %
1'
b1000 +
#382440000000
0!
0'
#382450000000
1!
b1001 %
1'
b1001 +
#382460000000
0!
0'
#382470000000
1!
b0 %
1'
b0 +
#382480000000
1"
1(
#382490000000
0!
0"
b100 &
0'
0(
b100 ,
#382500000000
1!
1$
b1 %
1'
1*
b1 +
#382510000000
0!
0'
#382520000000
1!
b10 %
1'
b10 +
#382530000000
0!
0'
#382540000000
1!
b11 %
1'
b11 +
#382550000000
0!
0'
#382560000000
1!
b100 %
1'
b100 +
#382570000000
0!
0'
#382580000000
1!
b101 %
1'
b101 +
#382590000000
0!
0'
#382600000000
1!
b110 %
1'
b110 +
#382610000000
0!
0'
#382620000000
1!
b111 %
1'
b111 +
#382630000000
0!
0'
#382640000000
1!
0$
b1000 %
1'
0*
b1000 +
#382650000000
0!
0'
#382660000000
1!
b1001 %
1'
b1001 +
#382670000000
0!
0'
#382680000000
1!
b0 %
1'
b0 +
#382690000000
0!
0'
#382700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#382710000000
0!
0'
#382720000000
1!
b10 %
1'
b10 +
#382730000000
0!
0'
#382740000000
1!
b11 %
1'
b11 +
#382750000000
0!
0'
#382760000000
1!
b100 %
1'
b100 +
#382770000000
0!
0'
#382780000000
1!
b101 %
1'
b101 +
#382790000000
0!
0'
#382800000000
1!
0$
b110 %
1'
0*
b110 +
#382810000000
0!
0'
#382820000000
1!
b111 %
1'
b111 +
#382830000000
0!
0'
#382840000000
1!
b1000 %
1'
b1000 +
#382850000000
0!
0'
#382860000000
1!
b1001 %
1'
b1001 +
#382870000000
0!
0'
#382880000000
1!
b0 %
1'
b0 +
#382890000000
0!
0'
#382900000000
1!
1$
b1 %
1'
1*
b1 +
#382910000000
1"
1(
#382920000000
0!
0"
b100 &
0'
0(
b100 ,
#382930000000
1!
b10 %
1'
b10 +
#382940000000
0!
0'
#382950000000
1!
b11 %
1'
b11 +
#382960000000
0!
0'
#382970000000
1!
b100 %
1'
b100 +
#382980000000
0!
0'
#382990000000
1!
b101 %
1'
b101 +
#383000000000
0!
0'
#383010000000
1!
b110 %
1'
b110 +
#383020000000
0!
0'
#383030000000
1!
b111 %
1'
b111 +
#383040000000
0!
0'
#383050000000
1!
0$
b1000 %
1'
0*
b1000 +
#383060000000
0!
0'
#383070000000
1!
b1001 %
1'
b1001 +
#383080000000
0!
0'
#383090000000
1!
b0 %
1'
b0 +
#383100000000
0!
0'
#383110000000
1!
1$
b1 %
1'
1*
b1 +
#383120000000
0!
0'
#383130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#383140000000
0!
0'
#383150000000
1!
b11 %
1'
b11 +
#383160000000
0!
0'
#383170000000
1!
b100 %
1'
b100 +
#383180000000
0!
0'
#383190000000
1!
b101 %
1'
b101 +
#383200000000
0!
0'
#383210000000
1!
0$
b110 %
1'
0*
b110 +
#383220000000
0!
0'
#383230000000
1!
b111 %
1'
b111 +
#383240000000
0!
0'
#383250000000
1!
b1000 %
1'
b1000 +
#383260000000
0!
0'
#383270000000
1!
b1001 %
1'
b1001 +
#383280000000
0!
0'
#383290000000
1!
b0 %
1'
b0 +
#383300000000
0!
0'
#383310000000
1!
1$
b1 %
1'
1*
b1 +
#383320000000
0!
0'
#383330000000
1!
b10 %
1'
b10 +
#383340000000
1"
1(
#383350000000
0!
0"
b100 &
0'
0(
b100 ,
#383360000000
1!
b11 %
1'
b11 +
#383370000000
0!
0'
#383380000000
1!
b100 %
1'
b100 +
#383390000000
0!
0'
#383400000000
1!
b101 %
1'
b101 +
#383410000000
0!
0'
#383420000000
1!
b110 %
1'
b110 +
#383430000000
0!
0'
#383440000000
1!
b111 %
1'
b111 +
#383450000000
0!
0'
#383460000000
1!
0$
b1000 %
1'
0*
b1000 +
#383470000000
0!
0'
#383480000000
1!
b1001 %
1'
b1001 +
#383490000000
0!
0'
#383500000000
1!
b0 %
1'
b0 +
#383510000000
0!
0'
#383520000000
1!
1$
b1 %
1'
1*
b1 +
#383530000000
0!
0'
#383540000000
1!
b10 %
1'
b10 +
#383550000000
0!
0'
#383560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#383570000000
0!
0'
#383580000000
1!
b100 %
1'
b100 +
#383590000000
0!
0'
#383600000000
1!
b101 %
1'
b101 +
#383610000000
0!
0'
#383620000000
1!
0$
b110 %
1'
0*
b110 +
#383630000000
0!
0'
#383640000000
1!
b111 %
1'
b111 +
#383650000000
0!
0'
#383660000000
1!
b1000 %
1'
b1000 +
#383670000000
0!
0'
#383680000000
1!
b1001 %
1'
b1001 +
#383690000000
0!
0'
#383700000000
1!
b0 %
1'
b0 +
#383710000000
0!
0'
#383720000000
1!
1$
b1 %
1'
1*
b1 +
#383730000000
0!
0'
#383740000000
1!
b10 %
1'
b10 +
#383750000000
0!
0'
#383760000000
1!
b11 %
1'
b11 +
#383770000000
1"
1(
#383780000000
0!
0"
b100 &
0'
0(
b100 ,
#383790000000
1!
b100 %
1'
b100 +
#383800000000
0!
0'
#383810000000
1!
b101 %
1'
b101 +
#383820000000
0!
0'
#383830000000
1!
b110 %
1'
b110 +
#383840000000
0!
0'
#383850000000
1!
b111 %
1'
b111 +
#383860000000
0!
0'
#383870000000
1!
0$
b1000 %
1'
0*
b1000 +
#383880000000
0!
0'
#383890000000
1!
b1001 %
1'
b1001 +
#383900000000
0!
0'
#383910000000
1!
b0 %
1'
b0 +
#383920000000
0!
0'
#383930000000
1!
1$
b1 %
1'
1*
b1 +
#383940000000
0!
0'
#383950000000
1!
b10 %
1'
b10 +
#383960000000
0!
0'
#383970000000
1!
b11 %
1'
b11 +
#383980000000
0!
0'
#383990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#384000000000
0!
0'
#384010000000
1!
b101 %
1'
b101 +
#384020000000
0!
0'
#384030000000
1!
0$
b110 %
1'
0*
b110 +
#384040000000
0!
0'
#384050000000
1!
b111 %
1'
b111 +
#384060000000
0!
0'
#384070000000
1!
b1000 %
1'
b1000 +
#384080000000
0!
0'
#384090000000
1!
b1001 %
1'
b1001 +
#384100000000
0!
0'
#384110000000
1!
b0 %
1'
b0 +
#384120000000
0!
0'
#384130000000
1!
1$
b1 %
1'
1*
b1 +
#384140000000
0!
0'
#384150000000
1!
b10 %
1'
b10 +
#384160000000
0!
0'
#384170000000
1!
b11 %
1'
b11 +
#384180000000
0!
0'
#384190000000
1!
b100 %
1'
b100 +
#384200000000
1"
1(
#384210000000
0!
0"
b100 &
0'
0(
b100 ,
#384220000000
1!
b101 %
1'
b101 +
#384230000000
0!
0'
#384240000000
1!
b110 %
1'
b110 +
#384250000000
0!
0'
#384260000000
1!
b111 %
1'
b111 +
#384270000000
0!
0'
#384280000000
1!
0$
b1000 %
1'
0*
b1000 +
#384290000000
0!
0'
#384300000000
1!
b1001 %
1'
b1001 +
#384310000000
0!
0'
#384320000000
1!
b0 %
1'
b0 +
#384330000000
0!
0'
#384340000000
1!
1$
b1 %
1'
1*
b1 +
#384350000000
0!
0'
#384360000000
1!
b10 %
1'
b10 +
#384370000000
0!
0'
#384380000000
1!
b11 %
1'
b11 +
#384390000000
0!
0'
#384400000000
1!
b100 %
1'
b100 +
#384410000000
0!
0'
#384420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#384430000000
0!
0'
#384440000000
1!
0$
b110 %
1'
0*
b110 +
#384450000000
0!
0'
#384460000000
1!
b111 %
1'
b111 +
#384470000000
0!
0'
#384480000000
1!
b1000 %
1'
b1000 +
#384490000000
0!
0'
#384500000000
1!
b1001 %
1'
b1001 +
#384510000000
0!
0'
#384520000000
1!
b0 %
1'
b0 +
#384530000000
0!
0'
#384540000000
1!
1$
b1 %
1'
1*
b1 +
#384550000000
0!
0'
#384560000000
1!
b10 %
1'
b10 +
#384570000000
0!
0'
#384580000000
1!
b11 %
1'
b11 +
#384590000000
0!
0'
#384600000000
1!
b100 %
1'
b100 +
#384610000000
0!
0'
#384620000000
1!
b101 %
1'
b101 +
#384630000000
1"
1(
#384640000000
0!
0"
b100 &
0'
0(
b100 ,
#384650000000
1!
b110 %
1'
b110 +
#384660000000
0!
0'
#384670000000
1!
b111 %
1'
b111 +
#384680000000
0!
0'
#384690000000
1!
0$
b1000 %
1'
0*
b1000 +
#384700000000
0!
0'
#384710000000
1!
b1001 %
1'
b1001 +
#384720000000
0!
0'
#384730000000
1!
b0 %
1'
b0 +
#384740000000
0!
0'
#384750000000
1!
1$
b1 %
1'
1*
b1 +
#384760000000
0!
0'
#384770000000
1!
b10 %
1'
b10 +
#384780000000
0!
0'
#384790000000
1!
b11 %
1'
b11 +
#384800000000
0!
0'
#384810000000
1!
b100 %
1'
b100 +
#384820000000
0!
0'
#384830000000
1!
b101 %
1'
b101 +
#384840000000
0!
0'
#384850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#384860000000
0!
0'
#384870000000
1!
b111 %
1'
b111 +
#384880000000
0!
0'
#384890000000
1!
b1000 %
1'
b1000 +
#384900000000
0!
0'
#384910000000
1!
b1001 %
1'
b1001 +
#384920000000
0!
0'
#384930000000
1!
b0 %
1'
b0 +
#384940000000
0!
0'
#384950000000
1!
1$
b1 %
1'
1*
b1 +
#384960000000
0!
0'
#384970000000
1!
b10 %
1'
b10 +
#384980000000
0!
0'
#384990000000
1!
b11 %
1'
b11 +
#385000000000
0!
0'
#385010000000
1!
b100 %
1'
b100 +
#385020000000
0!
0'
#385030000000
1!
b101 %
1'
b101 +
#385040000000
0!
0'
#385050000000
1!
0$
b110 %
1'
0*
b110 +
#385060000000
1"
1(
#385070000000
0!
0"
b100 &
0'
0(
b100 ,
#385080000000
1!
1$
b111 %
1'
1*
b111 +
#385090000000
0!
0'
#385100000000
1!
0$
b1000 %
1'
0*
b1000 +
#385110000000
0!
0'
#385120000000
1!
b1001 %
1'
b1001 +
#385130000000
0!
0'
#385140000000
1!
b0 %
1'
b0 +
#385150000000
0!
0'
#385160000000
1!
1$
b1 %
1'
1*
b1 +
#385170000000
0!
0'
#385180000000
1!
b10 %
1'
b10 +
#385190000000
0!
0'
#385200000000
1!
b11 %
1'
b11 +
#385210000000
0!
0'
#385220000000
1!
b100 %
1'
b100 +
#385230000000
0!
0'
#385240000000
1!
b101 %
1'
b101 +
#385250000000
0!
0'
#385260000000
1!
b110 %
1'
b110 +
#385270000000
0!
0'
#385280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#385290000000
0!
0'
#385300000000
1!
b1000 %
1'
b1000 +
#385310000000
0!
0'
#385320000000
1!
b1001 %
1'
b1001 +
#385330000000
0!
0'
#385340000000
1!
b0 %
1'
b0 +
#385350000000
0!
0'
#385360000000
1!
1$
b1 %
1'
1*
b1 +
#385370000000
0!
0'
#385380000000
1!
b10 %
1'
b10 +
#385390000000
0!
0'
#385400000000
1!
b11 %
1'
b11 +
#385410000000
0!
0'
#385420000000
1!
b100 %
1'
b100 +
#385430000000
0!
0'
#385440000000
1!
b101 %
1'
b101 +
#385450000000
0!
0'
#385460000000
1!
0$
b110 %
1'
0*
b110 +
#385470000000
0!
0'
#385480000000
1!
b111 %
1'
b111 +
#385490000000
1"
1(
#385500000000
0!
0"
b100 &
0'
0(
b100 ,
#385510000000
1!
b1000 %
1'
b1000 +
#385520000000
0!
0'
#385530000000
1!
b1001 %
1'
b1001 +
#385540000000
0!
0'
#385550000000
1!
b0 %
1'
b0 +
#385560000000
0!
0'
#385570000000
1!
1$
b1 %
1'
1*
b1 +
#385580000000
0!
0'
#385590000000
1!
b10 %
1'
b10 +
#385600000000
0!
0'
#385610000000
1!
b11 %
1'
b11 +
#385620000000
0!
0'
#385630000000
1!
b100 %
1'
b100 +
#385640000000
0!
0'
#385650000000
1!
b101 %
1'
b101 +
#385660000000
0!
0'
#385670000000
1!
b110 %
1'
b110 +
#385680000000
0!
0'
#385690000000
1!
b111 %
1'
b111 +
#385700000000
0!
0'
#385710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#385720000000
0!
0'
#385730000000
1!
b1001 %
1'
b1001 +
#385740000000
0!
0'
#385750000000
1!
b0 %
1'
b0 +
#385760000000
0!
0'
#385770000000
1!
1$
b1 %
1'
1*
b1 +
#385780000000
0!
0'
#385790000000
1!
b10 %
1'
b10 +
#385800000000
0!
0'
#385810000000
1!
b11 %
1'
b11 +
#385820000000
0!
0'
#385830000000
1!
b100 %
1'
b100 +
#385840000000
0!
0'
#385850000000
1!
b101 %
1'
b101 +
#385860000000
0!
0'
#385870000000
1!
0$
b110 %
1'
0*
b110 +
#385880000000
0!
0'
#385890000000
1!
b111 %
1'
b111 +
#385900000000
0!
0'
#385910000000
1!
b1000 %
1'
b1000 +
#385920000000
1"
1(
#385930000000
0!
0"
b100 &
0'
0(
b100 ,
#385940000000
1!
b1001 %
1'
b1001 +
#385950000000
0!
0'
#385960000000
1!
b0 %
1'
b0 +
#385970000000
0!
0'
#385980000000
1!
1$
b1 %
1'
1*
b1 +
#385990000000
0!
0'
#386000000000
1!
b10 %
1'
b10 +
#386010000000
0!
0'
#386020000000
1!
b11 %
1'
b11 +
#386030000000
0!
0'
#386040000000
1!
b100 %
1'
b100 +
#386050000000
0!
0'
#386060000000
1!
b101 %
1'
b101 +
#386070000000
0!
0'
#386080000000
1!
b110 %
1'
b110 +
#386090000000
0!
0'
#386100000000
1!
b111 %
1'
b111 +
#386110000000
0!
0'
#386120000000
1!
0$
b1000 %
1'
0*
b1000 +
#386130000000
0!
0'
#386140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#386150000000
0!
0'
#386160000000
1!
b0 %
1'
b0 +
#386170000000
0!
0'
#386180000000
1!
1$
b1 %
1'
1*
b1 +
#386190000000
0!
0'
#386200000000
1!
b10 %
1'
b10 +
#386210000000
0!
0'
#386220000000
1!
b11 %
1'
b11 +
#386230000000
0!
0'
#386240000000
1!
b100 %
1'
b100 +
#386250000000
0!
0'
#386260000000
1!
b101 %
1'
b101 +
#386270000000
0!
0'
#386280000000
1!
0$
b110 %
1'
0*
b110 +
#386290000000
0!
0'
#386300000000
1!
b111 %
1'
b111 +
#386310000000
0!
0'
#386320000000
1!
b1000 %
1'
b1000 +
#386330000000
0!
0'
#386340000000
1!
b1001 %
1'
b1001 +
#386350000000
1"
1(
#386360000000
0!
0"
b100 &
0'
0(
b100 ,
#386370000000
1!
b0 %
1'
b0 +
#386380000000
0!
0'
#386390000000
1!
1$
b1 %
1'
1*
b1 +
#386400000000
0!
0'
#386410000000
1!
b10 %
1'
b10 +
#386420000000
0!
0'
#386430000000
1!
b11 %
1'
b11 +
#386440000000
0!
0'
#386450000000
1!
b100 %
1'
b100 +
#386460000000
0!
0'
#386470000000
1!
b101 %
1'
b101 +
#386480000000
0!
0'
#386490000000
1!
b110 %
1'
b110 +
#386500000000
0!
0'
#386510000000
1!
b111 %
1'
b111 +
#386520000000
0!
0'
#386530000000
1!
0$
b1000 %
1'
0*
b1000 +
#386540000000
0!
0'
#386550000000
1!
b1001 %
1'
b1001 +
#386560000000
0!
0'
#386570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#386580000000
0!
0'
#386590000000
1!
1$
b1 %
1'
1*
b1 +
#386600000000
0!
0'
#386610000000
1!
b10 %
1'
b10 +
#386620000000
0!
0'
#386630000000
1!
b11 %
1'
b11 +
#386640000000
0!
0'
#386650000000
1!
b100 %
1'
b100 +
#386660000000
0!
0'
#386670000000
1!
b101 %
1'
b101 +
#386680000000
0!
0'
#386690000000
1!
0$
b110 %
1'
0*
b110 +
#386700000000
0!
0'
#386710000000
1!
b111 %
1'
b111 +
#386720000000
0!
0'
#386730000000
1!
b1000 %
1'
b1000 +
#386740000000
0!
0'
#386750000000
1!
b1001 %
1'
b1001 +
#386760000000
0!
0'
#386770000000
1!
b0 %
1'
b0 +
#386780000000
1"
1(
#386790000000
0!
0"
b100 &
0'
0(
b100 ,
#386800000000
1!
1$
b1 %
1'
1*
b1 +
#386810000000
0!
0'
#386820000000
1!
b10 %
1'
b10 +
#386830000000
0!
0'
#386840000000
1!
b11 %
1'
b11 +
#386850000000
0!
0'
#386860000000
1!
b100 %
1'
b100 +
#386870000000
0!
0'
#386880000000
1!
b101 %
1'
b101 +
#386890000000
0!
0'
#386900000000
1!
b110 %
1'
b110 +
#386910000000
0!
0'
#386920000000
1!
b111 %
1'
b111 +
#386930000000
0!
0'
#386940000000
1!
0$
b1000 %
1'
0*
b1000 +
#386950000000
0!
0'
#386960000000
1!
b1001 %
1'
b1001 +
#386970000000
0!
0'
#386980000000
1!
b0 %
1'
b0 +
#386990000000
0!
0'
#387000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#387010000000
0!
0'
#387020000000
1!
b10 %
1'
b10 +
#387030000000
0!
0'
#387040000000
1!
b11 %
1'
b11 +
#387050000000
0!
0'
#387060000000
1!
b100 %
1'
b100 +
#387070000000
0!
0'
#387080000000
1!
b101 %
1'
b101 +
#387090000000
0!
0'
#387100000000
1!
0$
b110 %
1'
0*
b110 +
#387110000000
0!
0'
#387120000000
1!
b111 %
1'
b111 +
#387130000000
0!
0'
#387140000000
1!
b1000 %
1'
b1000 +
#387150000000
0!
0'
#387160000000
1!
b1001 %
1'
b1001 +
#387170000000
0!
0'
#387180000000
1!
b0 %
1'
b0 +
#387190000000
0!
0'
#387200000000
1!
1$
b1 %
1'
1*
b1 +
#387210000000
1"
1(
#387220000000
0!
0"
b100 &
0'
0(
b100 ,
#387230000000
1!
b10 %
1'
b10 +
#387240000000
0!
0'
#387250000000
1!
b11 %
1'
b11 +
#387260000000
0!
0'
#387270000000
1!
b100 %
1'
b100 +
#387280000000
0!
0'
#387290000000
1!
b101 %
1'
b101 +
#387300000000
0!
0'
#387310000000
1!
b110 %
1'
b110 +
#387320000000
0!
0'
#387330000000
1!
b111 %
1'
b111 +
#387340000000
0!
0'
#387350000000
1!
0$
b1000 %
1'
0*
b1000 +
#387360000000
0!
0'
#387370000000
1!
b1001 %
1'
b1001 +
#387380000000
0!
0'
#387390000000
1!
b0 %
1'
b0 +
#387400000000
0!
0'
#387410000000
1!
1$
b1 %
1'
1*
b1 +
#387420000000
0!
0'
#387430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#387440000000
0!
0'
#387450000000
1!
b11 %
1'
b11 +
#387460000000
0!
0'
#387470000000
1!
b100 %
1'
b100 +
#387480000000
0!
0'
#387490000000
1!
b101 %
1'
b101 +
#387500000000
0!
0'
#387510000000
1!
0$
b110 %
1'
0*
b110 +
#387520000000
0!
0'
#387530000000
1!
b111 %
1'
b111 +
#387540000000
0!
0'
#387550000000
1!
b1000 %
1'
b1000 +
#387560000000
0!
0'
#387570000000
1!
b1001 %
1'
b1001 +
#387580000000
0!
0'
#387590000000
1!
b0 %
1'
b0 +
#387600000000
0!
0'
#387610000000
1!
1$
b1 %
1'
1*
b1 +
#387620000000
0!
0'
#387630000000
1!
b10 %
1'
b10 +
#387640000000
1"
1(
#387650000000
0!
0"
b100 &
0'
0(
b100 ,
#387660000000
1!
b11 %
1'
b11 +
#387670000000
0!
0'
#387680000000
1!
b100 %
1'
b100 +
#387690000000
0!
0'
#387700000000
1!
b101 %
1'
b101 +
#387710000000
0!
0'
#387720000000
1!
b110 %
1'
b110 +
#387730000000
0!
0'
#387740000000
1!
b111 %
1'
b111 +
#387750000000
0!
0'
#387760000000
1!
0$
b1000 %
1'
0*
b1000 +
#387770000000
0!
0'
#387780000000
1!
b1001 %
1'
b1001 +
#387790000000
0!
0'
#387800000000
1!
b0 %
1'
b0 +
#387810000000
0!
0'
#387820000000
1!
1$
b1 %
1'
1*
b1 +
#387830000000
0!
0'
#387840000000
1!
b10 %
1'
b10 +
#387850000000
0!
0'
#387860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#387870000000
0!
0'
#387880000000
1!
b100 %
1'
b100 +
#387890000000
0!
0'
#387900000000
1!
b101 %
1'
b101 +
#387910000000
0!
0'
#387920000000
1!
0$
b110 %
1'
0*
b110 +
#387930000000
0!
0'
#387940000000
1!
b111 %
1'
b111 +
#387950000000
0!
0'
#387960000000
1!
b1000 %
1'
b1000 +
#387970000000
0!
0'
#387980000000
1!
b1001 %
1'
b1001 +
#387990000000
0!
0'
#388000000000
1!
b0 %
1'
b0 +
#388010000000
0!
0'
#388020000000
1!
1$
b1 %
1'
1*
b1 +
#388030000000
0!
0'
#388040000000
1!
b10 %
1'
b10 +
#388050000000
0!
0'
#388060000000
1!
b11 %
1'
b11 +
#388070000000
1"
1(
#388080000000
0!
0"
b100 &
0'
0(
b100 ,
#388090000000
1!
b100 %
1'
b100 +
#388100000000
0!
0'
#388110000000
1!
b101 %
1'
b101 +
#388120000000
0!
0'
#388130000000
1!
b110 %
1'
b110 +
#388140000000
0!
0'
#388150000000
1!
b111 %
1'
b111 +
#388160000000
0!
0'
#388170000000
1!
0$
b1000 %
1'
0*
b1000 +
#388180000000
0!
0'
#388190000000
1!
b1001 %
1'
b1001 +
#388200000000
0!
0'
#388210000000
1!
b0 %
1'
b0 +
#388220000000
0!
0'
#388230000000
1!
1$
b1 %
1'
1*
b1 +
#388240000000
0!
0'
#388250000000
1!
b10 %
1'
b10 +
#388260000000
0!
0'
#388270000000
1!
b11 %
1'
b11 +
#388280000000
0!
0'
#388290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#388300000000
0!
0'
#388310000000
1!
b101 %
1'
b101 +
#388320000000
0!
0'
#388330000000
1!
0$
b110 %
1'
0*
b110 +
#388340000000
0!
0'
#388350000000
1!
b111 %
1'
b111 +
#388360000000
0!
0'
#388370000000
1!
b1000 %
1'
b1000 +
#388380000000
0!
0'
#388390000000
1!
b1001 %
1'
b1001 +
#388400000000
0!
0'
#388410000000
1!
b0 %
1'
b0 +
#388420000000
0!
0'
#388430000000
1!
1$
b1 %
1'
1*
b1 +
#388440000000
0!
0'
#388450000000
1!
b10 %
1'
b10 +
#388460000000
0!
0'
#388470000000
1!
b11 %
1'
b11 +
#388480000000
0!
0'
#388490000000
1!
b100 %
1'
b100 +
#388500000000
1"
1(
#388510000000
0!
0"
b100 &
0'
0(
b100 ,
#388520000000
1!
b101 %
1'
b101 +
#388530000000
0!
0'
#388540000000
1!
b110 %
1'
b110 +
#388550000000
0!
0'
#388560000000
1!
b111 %
1'
b111 +
#388570000000
0!
0'
#388580000000
1!
0$
b1000 %
1'
0*
b1000 +
#388590000000
0!
0'
#388600000000
1!
b1001 %
1'
b1001 +
#388610000000
0!
0'
#388620000000
1!
b0 %
1'
b0 +
#388630000000
0!
0'
#388640000000
1!
1$
b1 %
1'
1*
b1 +
#388650000000
0!
0'
#388660000000
1!
b10 %
1'
b10 +
#388670000000
0!
0'
#388680000000
1!
b11 %
1'
b11 +
#388690000000
0!
0'
#388700000000
1!
b100 %
1'
b100 +
#388710000000
0!
0'
#388720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#388730000000
0!
0'
#388740000000
1!
0$
b110 %
1'
0*
b110 +
#388750000000
0!
0'
#388760000000
1!
b111 %
1'
b111 +
#388770000000
0!
0'
#388780000000
1!
b1000 %
1'
b1000 +
#388790000000
0!
0'
#388800000000
1!
b1001 %
1'
b1001 +
#388810000000
0!
0'
#388820000000
1!
b0 %
1'
b0 +
#388830000000
0!
0'
#388840000000
1!
1$
b1 %
1'
1*
b1 +
#388850000000
0!
0'
#388860000000
1!
b10 %
1'
b10 +
#388870000000
0!
0'
#388880000000
1!
b11 %
1'
b11 +
#388890000000
0!
0'
#388900000000
1!
b100 %
1'
b100 +
#388910000000
0!
0'
#388920000000
1!
b101 %
1'
b101 +
#388930000000
1"
1(
#388940000000
0!
0"
b100 &
0'
0(
b100 ,
#388950000000
1!
b110 %
1'
b110 +
#388960000000
0!
0'
#388970000000
1!
b111 %
1'
b111 +
#388980000000
0!
0'
#388990000000
1!
0$
b1000 %
1'
0*
b1000 +
#389000000000
0!
0'
#389010000000
1!
b1001 %
1'
b1001 +
#389020000000
0!
0'
#389030000000
1!
b0 %
1'
b0 +
#389040000000
0!
0'
#389050000000
1!
1$
b1 %
1'
1*
b1 +
#389060000000
0!
0'
#389070000000
1!
b10 %
1'
b10 +
#389080000000
0!
0'
#389090000000
1!
b11 %
1'
b11 +
#389100000000
0!
0'
#389110000000
1!
b100 %
1'
b100 +
#389120000000
0!
0'
#389130000000
1!
b101 %
1'
b101 +
#389140000000
0!
0'
#389150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#389160000000
0!
0'
#389170000000
1!
b111 %
1'
b111 +
#389180000000
0!
0'
#389190000000
1!
b1000 %
1'
b1000 +
#389200000000
0!
0'
#389210000000
1!
b1001 %
1'
b1001 +
#389220000000
0!
0'
#389230000000
1!
b0 %
1'
b0 +
#389240000000
0!
0'
#389250000000
1!
1$
b1 %
1'
1*
b1 +
#389260000000
0!
0'
#389270000000
1!
b10 %
1'
b10 +
#389280000000
0!
0'
#389290000000
1!
b11 %
1'
b11 +
#389300000000
0!
0'
#389310000000
1!
b100 %
1'
b100 +
#389320000000
0!
0'
#389330000000
1!
b101 %
1'
b101 +
#389340000000
0!
0'
#389350000000
1!
0$
b110 %
1'
0*
b110 +
#389360000000
1"
1(
#389370000000
0!
0"
b100 &
0'
0(
b100 ,
#389380000000
1!
1$
b111 %
1'
1*
b111 +
#389390000000
0!
0'
#389400000000
1!
0$
b1000 %
1'
0*
b1000 +
#389410000000
0!
0'
#389420000000
1!
b1001 %
1'
b1001 +
#389430000000
0!
0'
#389440000000
1!
b0 %
1'
b0 +
#389450000000
0!
0'
#389460000000
1!
1$
b1 %
1'
1*
b1 +
#389470000000
0!
0'
#389480000000
1!
b10 %
1'
b10 +
#389490000000
0!
0'
#389500000000
1!
b11 %
1'
b11 +
#389510000000
0!
0'
#389520000000
1!
b100 %
1'
b100 +
#389530000000
0!
0'
#389540000000
1!
b101 %
1'
b101 +
#389550000000
0!
0'
#389560000000
1!
b110 %
1'
b110 +
#389570000000
0!
0'
#389580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#389590000000
0!
0'
#389600000000
1!
b1000 %
1'
b1000 +
#389610000000
0!
0'
#389620000000
1!
b1001 %
1'
b1001 +
#389630000000
0!
0'
#389640000000
1!
b0 %
1'
b0 +
#389650000000
0!
0'
#389660000000
1!
1$
b1 %
1'
1*
b1 +
#389670000000
0!
0'
#389680000000
1!
b10 %
1'
b10 +
#389690000000
0!
0'
#389700000000
1!
b11 %
1'
b11 +
#389710000000
0!
0'
#389720000000
1!
b100 %
1'
b100 +
#389730000000
0!
0'
#389740000000
1!
b101 %
1'
b101 +
#389750000000
0!
0'
#389760000000
1!
0$
b110 %
1'
0*
b110 +
#389770000000
0!
0'
#389780000000
1!
b111 %
1'
b111 +
#389790000000
1"
1(
#389800000000
0!
0"
b100 &
0'
0(
b100 ,
#389810000000
1!
b1000 %
1'
b1000 +
#389820000000
0!
0'
#389830000000
1!
b1001 %
1'
b1001 +
#389840000000
0!
0'
#389850000000
1!
b0 %
1'
b0 +
#389860000000
0!
0'
#389870000000
1!
1$
b1 %
1'
1*
b1 +
#389880000000
0!
0'
#389890000000
1!
b10 %
1'
b10 +
#389900000000
0!
0'
#389910000000
1!
b11 %
1'
b11 +
#389920000000
0!
0'
#389930000000
1!
b100 %
1'
b100 +
#389940000000
0!
0'
#389950000000
1!
b101 %
1'
b101 +
#389960000000
0!
0'
#389970000000
1!
b110 %
1'
b110 +
#389980000000
0!
0'
#389990000000
1!
b111 %
1'
b111 +
#390000000000
0!
0'
#390010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#390020000000
0!
0'
#390030000000
1!
b1001 %
1'
b1001 +
#390040000000
0!
0'
#390050000000
1!
b0 %
1'
b0 +
#390060000000
0!
0'
#390070000000
1!
1$
b1 %
1'
1*
b1 +
#390080000000
0!
0'
#390090000000
1!
b10 %
1'
b10 +
#390100000000
0!
0'
#390110000000
1!
b11 %
1'
b11 +
#390120000000
0!
0'
#390130000000
1!
b100 %
1'
b100 +
#390140000000
0!
0'
#390150000000
1!
b101 %
1'
b101 +
#390160000000
0!
0'
#390170000000
1!
0$
b110 %
1'
0*
b110 +
#390180000000
0!
0'
#390190000000
1!
b111 %
1'
b111 +
#390200000000
0!
0'
#390210000000
1!
b1000 %
1'
b1000 +
#390220000000
1"
1(
#390230000000
0!
0"
b100 &
0'
0(
b100 ,
#390240000000
1!
b1001 %
1'
b1001 +
#390250000000
0!
0'
#390260000000
1!
b0 %
1'
b0 +
#390270000000
0!
0'
#390280000000
1!
1$
b1 %
1'
1*
b1 +
#390290000000
0!
0'
#390300000000
1!
b10 %
1'
b10 +
#390310000000
0!
0'
#390320000000
1!
b11 %
1'
b11 +
#390330000000
0!
0'
#390340000000
1!
b100 %
1'
b100 +
#390350000000
0!
0'
#390360000000
1!
b101 %
1'
b101 +
#390370000000
0!
0'
#390380000000
1!
b110 %
1'
b110 +
#390390000000
0!
0'
#390400000000
1!
b111 %
1'
b111 +
#390410000000
0!
0'
#390420000000
1!
0$
b1000 %
1'
0*
b1000 +
#390430000000
0!
0'
#390440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#390450000000
0!
0'
#390460000000
1!
b0 %
1'
b0 +
#390470000000
0!
0'
#390480000000
1!
1$
b1 %
1'
1*
b1 +
#390490000000
0!
0'
#390500000000
1!
b10 %
1'
b10 +
#390510000000
0!
0'
#390520000000
1!
b11 %
1'
b11 +
#390530000000
0!
0'
#390540000000
1!
b100 %
1'
b100 +
#390550000000
0!
0'
#390560000000
1!
b101 %
1'
b101 +
#390570000000
0!
0'
#390580000000
1!
0$
b110 %
1'
0*
b110 +
#390590000000
0!
0'
#390600000000
1!
b111 %
1'
b111 +
#390610000000
0!
0'
#390620000000
1!
b1000 %
1'
b1000 +
#390630000000
0!
0'
#390640000000
1!
b1001 %
1'
b1001 +
#390650000000
1"
1(
#390660000000
0!
0"
b100 &
0'
0(
b100 ,
#390670000000
1!
b0 %
1'
b0 +
#390680000000
0!
0'
#390690000000
1!
1$
b1 %
1'
1*
b1 +
#390700000000
0!
0'
#390710000000
1!
b10 %
1'
b10 +
#390720000000
0!
0'
#390730000000
1!
b11 %
1'
b11 +
#390740000000
0!
0'
#390750000000
1!
b100 %
1'
b100 +
#390760000000
0!
0'
#390770000000
1!
b101 %
1'
b101 +
#390780000000
0!
0'
#390790000000
1!
b110 %
1'
b110 +
#390800000000
0!
0'
#390810000000
1!
b111 %
1'
b111 +
#390820000000
0!
0'
#390830000000
1!
0$
b1000 %
1'
0*
b1000 +
#390840000000
0!
0'
#390850000000
1!
b1001 %
1'
b1001 +
#390860000000
0!
0'
#390870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#390880000000
0!
0'
#390890000000
1!
1$
b1 %
1'
1*
b1 +
#390900000000
0!
0'
#390910000000
1!
b10 %
1'
b10 +
#390920000000
0!
0'
#390930000000
1!
b11 %
1'
b11 +
#390940000000
0!
0'
#390950000000
1!
b100 %
1'
b100 +
#390960000000
0!
0'
#390970000000
1!
b101 %
1'
b101 +
#390980000000
0!
0'
#390990000000
1!
0$
b110 %
1'
0*
b110 +
#391000000000
0!
0'
#391010000000
1!
b111 %
1'
b111 +
#391020000000
0!
0'
#391030000000
1!
b1000 %
1'
b1000 +
#391040000000
0!
0'
#391050000000
1!
b1001 %
1'
b1001 +
#391060000000
0!
0'
#391070000000
1!
b0 %
1'
b0 +
#391080000000
1"
1(
#391090000000
0!
0"
b100 &
0'
0(
b100 ,
#391100000000
1!
1$
b1 %
1'
1*
b1 +
#391110000000
0!
0'
#391120000000
1!
b10 %
1'
b10 +
#391130000000
0!
0'
#391140000000
1!
b11 %
1'
b11 +
#391150000000
0!
0'
#391160000000
1!
b100 %
1'
b100 +
#391170000000
0!
0'
#391180000000
1!
b101 %
1'
b101 +
#391190000000
0!
0'
#391200000000
1!
b110 %
1'
b110 +
#391210000000
0!
0'
#391220000000
1!
b111 %
1'
b111 +
#391230000000
0!
0'
#391240000000
1!
0$
b1000 %
1'
0*
b1000 +
#391250000000
0!
0'
#391260000000
1!
b1001 %
1'
b1001 +
#391270000000
0!
0'
#391280000000
1!
b0 %
1'
b0 +
#391290000000
0!
0'
#391300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#391310000000
0!
0'
#391320000000
1!
b10 %
1'
b10 +
#391330000000
0!
0'
#391340000000
1!
b11 %
1'
b11 +
#391350000000
0!
0'
#391360000000
1!
b100 %
1'
b100 +
#391370000000
0!
0'
#391380000000
1!
b101 %
1'
b101 +
#391390000000
0!
0'
#391400000000
1!
0$
b110 %
1'
0*
b110 +
#391410000000
0!
0'
#391420000000
1!
b111 %
1'
b111 +
#391430000000
0!
0'
#391440000000
1!
b1000 %
1'
b1000 +
#391450000000
0!
0'
#391460000000
1!
b1001 %
1'
b1001 +
#391470000000
0!
0'
#391480000000
1!
b0 %
1'
b0 +
#391490000000
0!
0'
#391500000000
1!
1$
b1 %
1'
1*
b1 +
#391510000000
1"
1(
#391520000000
0!
0"
b100 &
0'
0(
b100 ,
#391530000000
1!
b10 %
1'
b10 +
#391540000000
0!
0'
#391550000000
1!
b11 %
1'
b11 +
#391560000000
0!
0'
#391570000000
1!
b100 %
1'
b100 +
#391580000000
0!
0'
#391590000000
1!
b101 %
1'
b101 +
#391600000000
0!
0'
#391610000000
1!
b110 %
1'
b110 +
#391620000000
0!
0'
#391630000000
1!
b111 %
1'
b111 +
#391640000000
0!
0'
#391650000000
1!
0$
b1000 %
1'
0*
b1000 +
#391660000000
0!
0'
#391670000000
1!
b1001 %
1'
b1001 +
#391680000000
0!
0'
#391690000000
1!
b0 %
1'
b0 +
#391700000000
0!
0'
#391710000000
1!
1$
b1 %
1'
1*
b1 +
#391720000000
0!
0'
#391730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#391740000000
0!
0'
#391750000000
1!
b11 %
1'
b11 +
#391760000000
0!
0'
#391770000000
1!
b100 %
1'
b100 +
#391780000000
0!
0'
#391790000000
1!
b101 %
1'
b101 +
#391800000000
0!
0'
#391810000000
1!
0$
b110 %
1'
0*
b110 +
#391820000000
0!
0'
#391830000000
1!
b111 %
1'
b111 +
#391840000000
0!
0'
#391850000000
1!
b1000 %
1'
b1000 +
#391860000000
0!
0'
#391870000000
1!
b1001 %
1'
b1001 +
#391880000000
0!
0'
#391890000000
1!
b0 %
1'
b0 +
#391900000000
0!
0'
#391910000000
1!
1$
b1 %
1'
1*
b1 +
#391920000000
0!
0'
#391930000000
1!
b10 %
1'
b10 +
#391940000000
1"
1(
#391950000000
0!
0"
b100 &
0'
0(
b100 ,
#391960000000
1!
b11 %
1'
b11 +
#391970000000
0!
0'
#391980000000
1!
b100 %
1'
b100 +
#391990000000
0!
0'
#392000000000
1!
b101 %
1'
b101 +
#392010000000
0!
0'
#392020000000
1!
b110 %
1'
b110 +
#392030000000
0!
0'
#392040000000
1!
b111 %
1'
b111 +
#392050000000
0!
0'
#392060000000
1!
0$
b1000 %
1'
0*
b1000 +
#392070000000
0!
0'
#392080000000
1!
b1001 %
1'
b1001 +
#392090000000
0!
0'
#392100000000
1!
b0 %
1'
b0 +
#392110000000
0!
0'
#392120000000
1!
1$
b1 %
1'
1*
b1 +
#392130000000
0!
0'
#392140000000
1!
b10 %
1'
b10 +
#392150000000
0!
0'
#392160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#392170000000
0!
0'
#392180000000
1!
b100 %
1'
b100 +
#392190000000
0!
0'
#392200000000
1!
b101 %
1'
b101 +
#392210000000
0!
0'
#392220000000
1!
0$
b110 %
1'
0*
b110 +
#392230000000
0!
0'
#392240000000
1!
b111 %
1'
b111 +
#392250000000
0!
0'
#392260000000
1!
b1000 %
1'
b1000 +
#392270000000
0!
0'
#392280000000
1!
b1001 %
1'
b1001 +
#392290000000
0!
0'
#392300000000
1!
b0 %
1'
b0 +
#392310000000
0!
0'
#392320000000
1!
1$
b1 %
1'
1*
b1 +
#392330000000
0!
0'
#392340000000
1!
b10 %
1'
b10 +
#392350000000
0!
0'
#392360000000
1!
b11 %
1'
b11 +
#392370000000
1"
1(
#392380000000
0!
0"
b100 &
0'
0(
b100 ,
#392390000000
1!
b100 %
1'
b100 +
#392400000000
0!
0'
#392410000000
1!
b101 %
1'
b101 +
#392420000000
0!
0'
#392430000000
1!
b110 %
1'
b110 +
#392440000000
0!
0'
#392450000000
1!
b111 %
1'
b111 +
#392460000000
0!
0'
#392470000000
1!
0$
b1000 %
1'
0*
b1000 +
#392480000000
0!
0'
#392490000000
1!
b1001 %
1'
b1001 +
#392500000000
0!
0'
#392510000000
1!
b0 %
1'
b0 +
#392520000000
0!
0'
#392530000000
1!
1$
b1 %
1'
1*
b1 +
#392540000000
0!
0'
#392550000000
1!
b10 %
1'
b10 +
#392560000000
0!
0'
#392570000000
1!
b11 %
1'
b11 +
#392580000000
0!
0'
#392590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#392600000000
0!
0'
#392610000000
1!
b101 %
1'
b101 +
#392620000000
0!
0'
#392630000000
1!
0$
b110 %
1'
0*
b110 +
#392640000000
0!
0'
#392650000000
1!
b111 %
1'
b111 +
#392660000000
0!
0'
#392670000000
1!
b1000 %
1'
b1000 +
#392680000000
0!
0'
#392690000000
1!
b1001 %
1'
b1001 +
#392700000000
0!
0'
#392710000000
1!
b0 %
1'
b0 +
#392720000000
0!
0'
#392730000000
1!
1$
b1 %
1'
1*
b1 +
#392740000000
0!
0'
#392750000000
1!
b10 %
1'
b10 +
#392760000000
0!
0'
#392770000000
1!
b11 %
1'
b11 +
#392780000000
0!
0'
#392790000000
1!
b100 %
1'
b100 +
#392800000000
1"
1(
#392810000000
0!
0"
b100 &
0'
0(
b100 ,
#392820000000
1!
b101 %
1'
b101 +
#392830000000
0!
0'
#392840000000
1!
b110 %
1'
b110 +
#392850000000
0!
0'
#392860000000
1!
b111 %
1'
b111 +
#392870000000
0!
0'
#392880000000
1!
0$
b1000 %
1'
0*
b1000 +
#392890000000
0!
0'
#392900000000
1!
b1001 %
1'
b1001 +
#392910000000
0!
0'
#392920000000
1!
b0 %
1'
b0 +
#392930000000
0!
0'
#392940000000
1!
1$
b1 %
1'
1*
b1 +
#392950000000
0!
0'
#392960000000
1!
b10 %
1'
b10 +
#392970000000
0!
0'
#392980000000
1!
b11 %
1'
b11 +
#392990000000
0!
0'
#393000000000
1!
b100 %
1'
b100 +
#393010000000
0!
0'
#393020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#393030000000
0!
0'
#393040000000
1!
0$
b110 %
1'
0*
b110 +
#393050000000
0!
0'
#393060000000
1!
b111 %
1'
b111 +
#393070000000
0!
0'
#393080000000
1!
b1000 %
1'
b1000 +
#393090000000
0!
0'
#393100000000
1!
b1001 %
1'
b1001 +
#393110000000
0!
0'
#393120000000
1!
b0 %
1'
b0 +
#393130000000
0!
0'
#393140000000
1!
1$
b1 %
1'
1*
b1 +
#393150000000
0!
0'
#393160000000
1!
b10 %
1'
b10 +
#393170000000
0!
0'
#393180000000
1!
b11 %
1'
b11 +
#393190000000
0!
0'
#393200000000
1!
b100 %
1'
b100 +
#393210000000
0!
0'
#393220000000
1!
b101 %
1'
b101 +
#393230000000
1"
1(
#393240000000
0!
0"
b100 &
0'
0(
b100 ,
#393250000000
1!
b110 %
1'
b110 +
#393260000000
0!
0'
#393270000000
1!
b111 %
1'
b111 +
#393280000000
0!
0'
#393290000000
1!
0$
b1000 %
1'
0*
b1000 +
#393300000000
0!
0'
#393310000000
1!
b1001 %
1'
b1001 +
#393320000000
0!
0'
#393330000000
1!
b0 %
1'
b0 +
#393340000000
0!
0'
#393350000000
1!
1$
b1 %
1'
1*
b1 +
#393360000000
0!
0'
#393370000000
1!
b10 %
1'
b10 +
#393380000000
0!
0'
#393390000000
1!
b11 %
1'
b11 +
#393400000000
0!
0'
#393410000000
1!
b100 %
1'
b100 +
#393420000000
0!
0'
#393430000000
1!
b101 %
1'
b101 +
#393440000000
0!
0'
#393450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#393460000000
0!
0'
#393470000000
1!
b111 %
1'
b111 +
#393480000000
0!
0'
#393490000000
1!
b1000 %
1'
b1000 +
#393500000000
0!
0'
#393510000000
1!
b1001 %
1'
b1001 +
#393520000000
0!
0'
#393530000000
1!
b0 %
1'
b0 +
#393540000000
0!
0'
#393550000000
1!
1$
b1 %
1'
1*
b1 +
#393560000000
0!
0'
#393570000000
1!
b10 %
1'
b10 +
#393580000000
0!
0'
#393590000000
1!
b11 %
1'
b11 +
#393600000000
0!
0'
#393610000000
1!
b100 %
1'
b100 +
#393620000000
0!
0'
#393630000000
1!
b101 %
1'
b101 +
#393640000000
0!
0'
#393650000000
1!
0$
b110 %
1'
0*
b110 +
#393660000000
1"
1(
#393670000000
0!
0"
b100 &
0'
0(
b100 ,
#393680000000
1!
1$
b111 %
1'
1*
b111 +
#393690000000
0!
0'
#393700000000
1!
0$
b1000 %
1'
0*
b1000 +
#393710000000
0!
0'
#393720000000
1!
b1001 %
1'
b1001 +
#393730000000
0!
0'
#393740000000
1!
b0 %
1'
b0 +
#393750000000
0!
0'
#393760000000
1!
1$
b1 %
1'
1*
b1 +
#393770000000
0!
0'
#393780000000
1!
b10 %
1'
b10 +
#393790000000
0!
0'
#393800000000
1!
b11 %
1'
b11 +
#393810000000
0!
0'
#393820000000
1!
b100 %
1'
b100 +
#393830000000
0!
0'
#393840000000
1!
b101 %
1'
b101 +
#393850000000
0!
0'
#393860000000
1!
b110 %
1'
b110 +
#393870000000
0!
0'
#393880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#393890000000
0!
0'
#393900000000
1!
b1000 %
1'
b1000 +
#393910000000
0!
0'
#393920000000
1!
b1001 %
1'
b1001 +
#393930000000
0!
0'
#393940000000
1!
b0 %
1'
b0 +
#393950000000
0!
0'
#393960000000
1!
1$
b1 %
1'
1*
b1 +
#393970000000
0!
0'
#393980000000
1!
b10 %
1'
b10 +
#393990000000
0!
0'
#394000000000
1!
b11 %
1'
b11 +
#394010000000
0!
0'
#394020000000
1!
b100 %
1'
b100 +
#394030000000
0!
0'
#394040000000
1!
b101 %
1'
b101 +
#394050000000
0!
0'
#394060000000
1!
0$
b110 %
1'
0*
b110 +
#394070000000
0!
0'
#394080000000
1!
b111 %
1'
b111 +
#394090000000
1"
1(
#394100000000
0!
0"
b100 &
0'
0(
b100 ,
#394110000000
1!
b1000 %
1'
b1000 +
#394120000000
0!
0'
#394130000000
1!
b1001 %
1'
b1001 +
#394140000000
0!
0'
#394150000000
1!
b0 %
1'
b0 +
#394160000000
0!
0'
#394170000000
1!
1$
b1 %
1'
1*
b1 +
#394180000000
0!
0'
#394190000000
1!
b10 %
1'
b10 +
#394200000000
0!
0'
#394210000000
1!
b11 %
1'
b11 +
#394220000000
0!
0'
#394230000000
1!
b100 %
1'
b100 +
#394240000000
0!
0'
#394250000000
1!
b101 %
1'
b101 +
#394260000000
0!
0'
#394270000000
1!
b110 %
1'
b110 +
#394280000000
0!
0'
#394290000000
1!
b111 %
1'
b111 +
#394300000000
0!
0'
#394310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#394320000000
0!
0'
#394330000000
1!
b1001 %
1'
b1001 +
#394340000000
0!
0'
#394350000000
1!
b0 %
1'
b0 +
#394360000000
0!
0'
#394370000000
1!
1$
b1 %
1'
1*
b1 +
#394380000000
0!
0'
#394390000000
1!
b10 %
1'
b10 +
#394400000000
0!
0'
#394410000000
1!
b11 %
1'
b11 +
#394420000000
0!
0'
#394430000000
1!
b100 %
1'
b100 +
#394440000000
0!
0'
#394450000000
1!
b101 %
1'
b101 +
#394460000000
0!
0'
#394470000000
1!
0$
b110 %
1'
0*
b110 +
#394480000000
0!
0'
#394490000000
1!
b111 %
1'
b111 +
#394500000000
0!
0'
#394510000000
1!
b1000 %
1'
b1000 +
#394520000000
1"
1(
#394530000000
0!
0"
b100 &
0'
0(
b100 ,
#394540000000
1!
b1001 %
1'
b1001 +
#394550000000
0!
0'
#394560000000
1!
b0 %
1'
b0 +
#394570000000
0!
0'
#394580000000
1!
1$
b1 %
1'
1*
b1 +
#394590000000
0!
0'
#394600000000
1!
b10 %
1'
b10 +
#394610000000
0!
0'
#394620000000
1!
b11 %
1'
b11 +
#394630000000
0!
0'
#394640000000
1!
b100 %
1'
b100 +
#394650000000
0!
0'
#394660000000
1!
b101 %
1'
b101 +
#394670000000
0!
0'
#394680000000
1!
b110 %
1'
b110 +
#394690000000
0!
0'
#394700000000
1!
b111 %
1'
b111 +
#394710000000
0!
0'
#394720000000
1!
0$
b1000 %
1'
0*
b1000 +
#394730000000
0!
0'
#394740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#394750000000
0!
0'
#394760000000
1!
b0 %
1'
b0 +
#394770000000
0!
0'
#394780000000
1!
1$
b1 %
1'
1*
b1 +
#394790000000
0!
0'
#394800000000
1!
b10 %
1'
b10 +
#394810000000
0!
0'
#394820000000
1!
b11 %
1'
b11 +
#394830000000
0!
0'
#394840000000
1!
b100 %
1'
b100 +
#394850000000
0!
0'
#394860000000
1!
b101 %
1'
b101 +
#394870000000
0!
0'
#394880000000
1!
0$
b110 %
1'
0*
b110 +
#394890000000
0!
0'
#394900000000
1!
b111 %
1'
b111 +
#394910000000
0!
0'
#394920000000
1!
b1000 %
1'
b1000 +
#394930000000
0!
0'
#394940000000
1!
b1001 %
1'
b1001 +
#394950000000
1"
1(
#394960000000
0!
0"
b100 &
0'
0(
b100 ,
#394970000000
1!
b0 %
1'
b0 +
#394980000000
0!
0'
#394990000000
1!
1$
b1 %
1'
1*
b1 +
#395000000000
0!
0'
#395010000000
1!
b10 %
1'
b10 +
#395020000000
0!
0'
#395030000000
1!
b11 %
1'
b11 +
#395040000000
0!
0'
#395050000000
1!
b100 %
1'
b100 +
#395060000000
0!
0'
#395070000000
1!
b101 %
1'
b101 +
#395080000000
0!
0'
#395090000000
1!
b110 %
1'
b110 +
#395100000000
0!
0'
#395110000000
1!
b111 %
1'
b111 +
#395120000000
0!
0'
#395130000000
1!
0$
b1000 %
1'
0*
b1000 +
#395140000000
0!
0'
#395150000000
1!
b1001 %
1'
b1001 +
#395160000000
0!
0'
#395170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#395180000000
0!
0'
#395190000000
1!
1$
b1 %
1'
1*
b1 +
#395200000000
0!
0'
#395210000000
1!
b10 %
1'
b10 +
#395220000000
0!
0'
#395230000000
1!
b11 %
1'
b11 +
#395240000000
0!
0'
#395250000000
1!
b100 %
1'
b100 +
#395260000000
0!
0'
#395270000000
1!
b101 %
1'
b101 +
#395280000000
0!
0'
#395290000000
1!
0$
b110 %
1'
0*
b110 +
#395300000000
0!
0'
#395310000000
1!
b111 %
1'
b111 +
#395320000000
0!
0'
#395330000000
1!
b1000 %
1'
b1000 +
#395340000000
0!
0'
#395350000000
1!
b1001 %
1'
b1001 +
#395360000000
0!
0'
#395370000000
1!
b0 %
1'
b0 +
#395380000000
1"
1(
#395390000000
0!
0"
b100 &
0'
0(
b100 ,
#395400000000
1!
1$
b1 %
1'
1*
b1 +
#395410000000
0!
0'
#395420000000
1!
b10 %
1'
b10 +
#395430000000
0!
0'
#395440000000
1!
b11 %
1'
b11 +
#395450000000
0!
0'
#395460000000
1!
b100 %
1'
b100 +
#395470000000
0!
0'
#395480000000
1!
b101 %
1'
b101 +
#395490000000
0!
0'
#395500000000
1!
b110 %
1'
b110 +
#395510000000
0!
0'
#395520000000
1!
b111 %
1'
b111 +
#395530000000
0!
0'
#395540000000
1!
0$
b1000 %
1'
0*
b1000 +
#395550000000
0!
0'
#395560000000
1!
b1001 %
1'
b1001 +
#395570000000
0!
0'
#395580000000
1!
b0 %
1'
b0 +
#395590000000
0!
0'
#395600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#395610000000
0!
0'
#395620000000
1!
b10 %
1'
b10 +
#395630000000
0!
0'
#395640000000
1!
b11 %
1'
b11 +
#395650000000
0!
0'
#395660000000
1!
b100 %
1'
b100 +
#395670000000
0!
0'
#395680000000
1!
b101 %
1'
b101 +
#395690000000
0!
0'
#395700000000
1!
0$
b110 %
1'
0*
b110 +
#395710000000
0!
0'
#395720000000
1!
b111 %
1'
b111 +
#395730000000
0!
0'
#395740000000
1!
b1000 %
1'
b1000 +
#395750000000
0!
0'
#395760000000
1!
b1001 %
1'
b1001 +
#395770000000
0!
0'
#395780000000
1!
b0 %
1'
b0 +
#395790000000
0!
0'
#395800000000
1!
1$
b1 %
1'
1*
b1 +
#395810000000
1"
1(
#395820000000
0!
0"
b100 &
0'
0(
b100 ,
#395830000000
1!
b10 %
1'
b10 +
#395840000000
0!
0'
#395850000000
1!
b11 %
1'
b11 +
#395860000000
0!
0'
#395870000000
1!
b100 %
1'
b100 +
#395880000000
0!
0'
#395890000000
1!
b101 %
1'
b101 +
#395900000000
0!
0'
#395910000000
1!
b110 %
1'
b110 +
#395920000000
0!
0'
#395930000000
1!
b111 %
1'
b111 +
#395940000000
0!
0'
#395950000000
1!
0$
b1000 %
1'
0*
b1000 +
#395960000000
0!
0'
#395970000000
1!
b1001 %
1'
b1001 +
#395980000000
0!
0'
#395990000000
1!
b0 %
1'
b0 +
#396000000000
0!
0'
#396010000000
1!
1$
b1 %
1'
1*
b1 +
#396020000000
0!
0'
#396030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#396040000000
0!
0'
#396050000000
1!
b11 %
1'
b11 +
#396060000000
0!
0'
#396070000000
1!
b100 %
1'
b100 +
#396080000000
0!
0'
#396090000000
1!
b101 %
1'
b101 +
#396100000000
0!
0'
#396110000000
1!
0$
b110 %
1'
0*
b110 +
#396120000000
0!
0'
#396130000000
1!
b111 %
1'
b111 +
#396140000000
0!
0'
#396150000000
1!
b1000 %
1'
b1000 +
#396160000000
0!
0'
#396170000000
1!
b1001 %
1'
b1001 +
#396180000000
0!
0'
#396190000000
1!
b0 %
1'
b0 +
#396200000000
0!
0'
#396210000000
1!
1$
b1 %
1'
1*
b1 +
#396220000000
0!
0'
#396230000000
1!
b10 %
1'
b10 +
#396240000000
1"
1(
#396250000000
0!
0"
b100 &
0'
0(
b100 ,
#396260000000
1!
b11 %
1'
b11 +
#396270000000
0!
0'
#396280000000
1!
b100 %
1'
b100 +
#396290000000
0!
0'
#396300000000
1!
b101 %
1'
b101 +
#396310000000
0!
0'
#396320000000
1!
b110 %
1'
b110 +
#396330000000
0!
0'
#396340000000
1!
b111 %
1'
b111 +
#396350000000
0!
0'
#396360000000
1!
0$
b1000 %
1'
0*
b1000 +
#396370000000
0!
0'
#396380000000
1!
b1001 %
1'
b1001 +
#396390000000
0!
0'
#396400000000
1!
b0 %
1'
b0 +
#396410000000
0!
0'
#396420000000
1!
1$
b1 %
1'
1*
b1 +
#396430000000
0!
0'
#396440000000
1!
b10 %
1'
b10 +
#396450000000
0!
0'
#396460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#396470000000
0!
0'
#396480000000
1!
b100 %
1'
b100 +
#396490000000
0!
0'
#396500000000
1!
b101 %
1'
b101 +
#396510000000
0!
0'
#396520000000
1!
0$
b110 %
1'
0*
b110 +
#396530000000
0!
0'
#396540000000
1!
b111 %
1'
b111 +
#396550000000
0!
0'
#396560000000
1!
b1000 %
1'
b1000 +
#396570000000
0!
0'
#396580000000
1!
b1001 %
1'
b1001 +
#396590000000
0!
0'
#396600000000
1!
b0 %
1'
b0 +
#396610000000
0!
0'
#396620000000
1!
1$
b1 %
1'
1*
b1 +
#396630000000
0!
0'
#396640000000
1!
b10 %
1'
b10 +
#396650000000
0!
0'
#396660000000
1!
b11 %
1'
b11 +
#396670000000
1"
1(
#396680000000
0!
0"
b100 &
0'
0(
b100 ,
#396690000000
1!
b100 %
1'
b100 +
#396700000000
0!
0'
#396710000000
1!
b101 %
1'
b101 +
#396720000000
0!
0'
#396730000000
1!
b110 %
1'
b110 +
#396740000000
0!
0'
#396750000000
1!
b111 %
1'
b111 +
#396760000000
0!
0'
#396770000000
1!
0$
b1000 %
1'
0*
b1000 +
#396780000000
0!
0'
#396790000000
1!
b1001 %
1'
b1001 +
#396800000000
0!
0'
#396810000000
1!
b0 %
1'
b0 +
#396820000000
0!
0'
#396830000000
1!
1$
b1 %
1'
1*
b1 +
#396840000000
0!
0'
#396850000000
1!
b10 %
1'
b10 +
#396860000000
0!
0'
#396870000000
1!
b11 %
1'
b11 +
#396880000000
0!
0'
#396890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#396900000000
0!
0'
#396910000000
1!
b101 %
1'
b101 +
#396920000000
0!
0'
#396930000000
1!
0$
b110 %
1'
0*
b110 +
#396940000000
0!
0'
#396950000000
1!
b111 %
1'
b111 +
#396960000000
0!
0'
#396970000000
1!
b1000 %
1'
b1000 +
#396980000000
0!
0'
#396990000000
1!
b1001 %
1'
b1001 +
#397000000000
0!
0'
#397010000000
1!
b0 %
1'
b0 +
#397020000000
0!
0'
#397030000000
1!
1$
b1 %
1'
1*
b1 +
#397040000000
0!
0'
#397050000000
1!
b10 %
1'
b10 +
#397060000000
0!
0'
#397070000000
1!
b11 %
1'
b11 +
#397080000000
0!
0'
#397090000000
1!
b100 %
1'
b100 +
#397100000000
1"
1(
#397110000000
0!
0"
b100 &
0'
0(
b100 ,
#397120000000
1!
b101 %
1'
b101 +
#397130000000
0!
0'
#397140000000
1!
b110 %
1'
b110 +
#397150000000
0!
0'
#397160000000
1!
b111 %
1'
b111 +
#397170000000
0!
0'
#397180000000
1!
0$
b1000 %
1'
0*
b1000 +
#397190000000
0!
0'
#397200000000
1!
b1001 %
1'
b1001 +
#397210000000
0!
0'
#397220000000
1!
b0 %
1'
b0 +
#397230000000
0!
0'
#397240000000
1!
1$
b1 %
1'
1*
b1 +
#397250000000
0!
0'
#397260000000
1!
b10 %
1'
b10 +
#397270000000
0!
0'
#397280000000
1!
b11 %
1'
b11 +
#397290000000
0!
0'
#397300000000
1!
b100 %
1'
b100 +
#397310000000
0!
0'
#397320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#397330000000
0!
0'
#397340000000
1!
0$
b110 %
1'
0*
b110 +
#397350000000
0!
0'
#397360000000
1!
b111 %
1'
b111 +
#397370000000
0!
0'
#397380000000
1!
b1000 %
1'
b1000 +
#397390000000
0!
0'
#397400000000
1!
b1001 %
1'
b1001 +
#397410000000
0!
0'
#397420000000
1!
b0 %
1'
b0 +
#397430000000
0!
0'
#397440000000
1!
1$
b1 %
1'
1*
b1 +
#397450000000
0!
0'
#397460000000
1!
b10 %
1'
b10 +
#397470000000
0!
0'
#397480000000
1!
b11 %
1'
b11 +
#397490000000
0!
0'
#397500000000
1!
b100 %
1'
b100 +
#397510000000
0!
0'
#397520000000
1!
b101 %
1'
b101 +
#397530000000
1"
1(
#397540000000
0!
0"
b100 &
0'
0(
b100 ,
#397550000000
1!
b110 %
1'
b110 +
#397560000000
0!
0'
#397570000000
1!
b111 %
1'
b111 +
#397580000000
0!
0'
#397590000000
1!
0$
b1000 %
1'
0*
b1000 +
#397600000000
0!
0'
#397610000000
1!
b1001 %
1'
b1001 +
#397620000000
0!
0'
#397630000000
1!
b0 %
1'
b0 +
#397640000000
0!
0'
#397650000000
1!
1$
b1 %
1'
1*
b1 +
#397660000000
0!
0'
#397670000000
1!
b10 %
1'
b10 +
#397680000000
0!
0'
#397690000000
1!
b11 %
1'
b11 +
#397700000000
0!
0'
#397710000000
1!
b100 %
1'
b100 +
#397720000000
0!
0'
#397730000000
1!
b101 %
1'
b101 +
#397740000000
0!
0'
#397750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#397760000000
0!
0'
#397770000000
1!
b111 %
1'
b111 +
#397780000000
0!
0'
#397790000000
1!
b1000 %
1'
b1000 +
#397800000000
0!
0'
#397810000000
1!
b1001 %
1'
b1001 +
#397820000000
0!
0'
#397830000000
1!
b0 %
1'
b0 +
#397840000000
0!
0'
#397850000000
1!
1$
b1 %
1'
1*
b1 +
#397860000000
0!
0'
#397870000000
1!
b10 %
1'
b10 +
#397880000000
0!
0'
#397890000000
1!
b11 %
1'
b11 +
#397900000000
0!
0'
#397910000000
1!
b100 %
1'
b100 +
#397920000000
0!
0'
#397930000000
1!
b101 %
1'
b101 +
#397940000000
0!
0'
#397950000000
1!
0$
b110 %
1'
0*
b110 +
#397960000000
1"
1(
#397970000000
0!
0"
b100 &
0'
0(
b100 ,
#397980000000
1!
1$
b111 %
1'
1*
b111 +
#397990000000
0!
0'
#398000000000
1!
0$
b1000 %
1'
0*
b1000 +
#398010000000
0!
0'
#398020000000
1!
b1001 %
1'
b1001 +
#398030000000
0!
0'
#398040000000
1!
b0 %
1'
b0 +
#398050000000
0!
0'
#398060000000
1!
1$
b1 %
1'
1*
b1 +
#398070000000
0!
0'
#398080000000
1!
b10 %
1'
b10 +
#398090000000
0!
0'
#398100000000
1!
b11 %
1'
b11 +
#398110000000
0!
0'
#398120000000
1!
b100 %
1'
b100 +
#398130000000
0!
0'
#398140000000
1!
b101 %
1'
b101 +
#398150000000
0!
0'
#398160000000
1!
b110 %
1'
b110 +
#398170000000
0!
0'
#398180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#398190000000
0!
0'
#398200000000
1!
b1000 %
1'
b1000 +
#398210000000
0!
0'
#398220000000
1!
b1001 %
1'
b1001 +
#398230000000
0!
0'
#398240000000
1!
b0 %
1'
b0 +
#398250000000
0!
0'
#398260000000
1!
1$
b1 %
1'
1*
b1 +
#398270000000
0!
0'
#398280000000
1!
b10 %
1'
b10 +
#398290000000
0!
0'
#398300000000
1!
b11 %
1'
b11 +
#398310000000
0!
0'
#398320000000
1!
b100 %
1'
b100 +
#398330000000
0!
0'
#398340000000
1!
b101 %
1'
b101 +
#398350000000
0!
0'
#398360000000
1!
0$
b110 %
1'
0*
b110 +
#398370000000
0!
0'
#398380000000
1!
b111 %
1'
b111 +
#398390000000
1"
1(
#398400000000
0!
0"
b100 &
0'
0(
b100 ,
#398410000000
1!
b1000 %
1'
b1000 +
#398420000000
0!
0'
#398430000000
1!
b1001 %
1'
b1001 +
#398440000000
0!
0'
#398450000000
1!
b0 %
1'
b0 +
#398460000000
0!
0'
#398470000000
1!
1$
b1 %
1'
1*
b1 +
#398480000000
0!
0'
#398490000000
1!
b10 %
1'
b10 +
#398500000000
0!
0'
#398510000000
1!
b11 %
1'
b11 +
#398520000000
0!
0'
#398530000000
1!
b100 %
1'
b100 +
#398540000000
0!
0'
#398550000000
1!
b101 %
1'
b101 +
#398560000000
0!
0'
#398570000000
1!
b110 %
1'
b110 +
#398580000000
0!
0'
#398590000000
1!
b111 %
1'
b111 +
#398600000000
0!
0'
#398610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#398620000000
0!
0'
#398630000000
1!
b1001 %
1'
b1001 +
#398640000000
0!
0'
#398650000000
1!
b0 %
1'
b0 +
#398660000000
0!
0'
#398670000000
1!
1$
b1 %
1'
1*
b1 +
#398680000000
0!
0'
#398690000000
1!
b10 %
1'
b10 +
#398700000000
0!
0'
#398710000000
1!
b11 %
1'
b11 +
#398720000000
0!
0'
#398730000000
1!
b100 %
1'
b100 +
#398740000000
0!
0'
#398750000000
1!
b101 %
1'
b101 +
#398760000000
0!
0'
#398770000000
1!
0$
b110 %
1'
0*
b110 +
#398780000000
0!
0'
#398790000000
1!
b111 %
1'
b111 +
#398800000000
0!
0'
#398810000000
1!
b1000 %
1'
b1000 +
#398820000000
1"
1(
#398830000000
0!
0"
b100 &
0'
0(
b100 ,
#398840000000
1!
b1001 %
1'
b1001 +
#398850000000
0!
0'
#398860000000
1!
b0 %
1'
b0 +
#398870000000
0!
0'
#398880000000
1!
1$
b1 %
1'
1*
b1 +
#398890000000
0!
0'
#398900000000
1!
b10 %
1'
b10 +
#398910000000
0!
0'
#398920000000
1!
b11 %
1'
b11 +
#398930000000
0!
0'
#398940000000
1!
b100 %
1'
b100 +
#398950000000
0!
0'
#398960000000
1!
b101 %
1'
b101 +
#398970000000
0!
0'
#398980000000
1!
b110 %
1'
b110 +
#398990000000
0!
0'
#399000000000
1!
b111 %
1'
b111 +
#399010000000
0!
0'
#399020000000
1!
0$
b1000 %
1'
0*
b1000 +
#399030000000
0!
0'
#399040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#399050000000
0!
0'
#399060000000
1!
b0 %
1'
b0 +
#399070000000
0!
0'
#399080000000
1!
1$
b1 %
1'
1*
b1 +
#399090000000
0!
0'
#399100000000
1!
b10 %
1'
b10 +
#399110000000
0!
0'
#399120000000
1!
b11 %
1'
b11 +
#399130000000
0!
0'
#399140000000
1!
b100 %
1'
b100 +
#399150000000
0!
0'
#399160000000
1!
b101 %
1'
b101 +
#399170000000
0!
0'
#399180000000
1!
0$
b110 %
1'
0*
b110 +
#399190000000
0!
0'
#399200000000
1!
b111 %
1'
b111 +
#399210000000
0!
0'
#399220000000
1!
b1000 %
1'
b1000 +
#399230000000
0!
0'
#399240000000
1!
b1001 %
1'
b1001 +
#399250000000
1"
1(
#399260000000
0!
0"
b100 &
0'
0(
b100 ,
#399270000000
1!
b0 %
1'
b0 +
#399280000000
0!
0'
#399290000000
1!
1$
b1 %
1'
1*
b1 +
#399300000000
0!
0'
#399310000000
1!
b10 %
1'
b10 +
#399320000000
0!
0'
#399330000000
1!
b11 %
1'
b11 +
#399340000000
0!
0'
#399350000000
1!
b100 %
1'
b100 +
#399360000000
0!
0'
#399370000000
1!
b101 %
1'
b101 +
#399380000000
0!
0'
#399390000000
1!
b110 %
1'
b110 +
#399400000000
0!
0'
#399410000000
1!
b111 %
1'
b111 +
#399420000000
0!
0'
#399430000000
1!
0$
b1000 %
1'
0*
b1000 +
#399440000000
0!
0'
#399450000000
1!
b1001 %
1'
b1001 +
#399460000000
0!
0'
#399470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#399480000000
0!
0'
#399490000000
1!
1$
b1 %
1'
1*
b1 +
#399500000000
0!
0'
#399510000000
1!
b10 %
1'
b10 +
#399520000000
0!
0'
#399530000000
1!
b11 %
1'
b11 +
#399540000000
0!
0'
#399550000000
1!
b100 %
1'
b100 +
#399560000000
0!
0'
#399570000000
1!
b101 %
1'
b101 +
#399580000000
0!
0'
#399590000000
1!
0$
b110 %
1'
0*
b110 +
#399600000000
0!
0'
#399610000000
1!
b111 %
1'
b111 +
#399620000000
0!
0'
#399630000000
1!
b1000 %
1'
b1000 +
#399640000000
0!
0'
#399650000000
1!
b1001 %
1'
b1001 +
#399660000000
0!
0'
#399670000000
1!
b0 %
1'
b0 +
#399680000000
1"
1(
#399690000000
0!
0"
b100 &
0'
0(
b100 ,
#399700000000
1!
1$
b1 %
1'
1*
b1 +
#399710000000
0!
0'
#399720000000
1!
b10 %
1'
b10 +
#399730000000
0!
0'
#399740000000
1!
b11 %
1'
b11 +
#399750000000
0!
0'
#399760000000
1!
b100 %
1'
b100 +
#399770000000
0!
0'
#399780000000
1!
b101 %
1'
b101 +
#399790000000
0!
0'
#399800000000
1!
b110 %
1'
b110 +
#399810000000
0!
0'
#399820000000
1!
b111 %
1'
b111 +
#399830000000
0!
0'
#399840000000
1!
0$
b1000 %
1'
0*
b1000 +
#399850000000
0!
0'
#399860000000
1!
b1001 %
1'
b1001 +
#399870000000
0!
0'
#399880000000
1!
b0 %
1'
b0 +
#399890000000
0!
0'
#399900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#399910000000
0!
0'
#399920000000
1!
b10 %
1'
b10 +
#399930000000
0!
0'
#399940000000
1!
b11 %
1'
b11 +
#399950000000
0!
0'
#399960000000
1!
b100 %
1'
b100 +
#399970000000
0!
0'
#399980000000
1!
b101 %
1'
b101 +
#399990000000
0!
0'
#400000000000
1!
0$
b110 %
1'
0*
b110 +
#400010000000
0!
0'
#400020000000
1!
b111 %
1'
b111 +
#400030000000
0!
0'
#400040000000
1!
b1000 %
1'
b1000 +
#400050000000
0!
0'
#400060000000
1!
b1001 %
1'
b1001 +
#400070000000
0!
0'
#400080000000
1!
b0 %
1'
b0 +
#400090000000
0!
0'
#400100000000
1!
1$
b1 %
1'
1*
b1 +
#400110000000
1"
1(
#400120000000
0!
0"
b100 &
0'
0(
b100 ,
#400130000000
1!
b10 %
1'
b10 +
#400140000000
0!
0'
#400150000000
1!
b11 %
1'
b11 +
#400160000000
0!
0'
#400170000000
1!
b100 %
1'
b100 +
#400180000000
0!
0'
#400190000000
1!
b101 %
1'
b101 +
#400200000000
0!
0'
#400210000000
1!
b110 %
1'
b110 +
#400220000000
0!
0'
#400230000000
1!
b111 %
1'
b111 +
#400240000000
0!
0'
#400250000000
1!
0$
b1000 %
1'
0*
b1000 +
#400260000000
0!
0'
#400270000000
1!
b1001 %
1'
b1001 +
#400280000000
0!
0'
#400290000000
1!
b0 %
1'
b0 +
#400300000000
0!
0'
#400310000000
1!
1$
b1 %
1'
1*
b1 +
#400320000000
0!
0'
#400330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#400340000000
0!
0'
#400350000000
1!
b11 %
1'
b11 +
#400360000000
0!
0'
#400370000000
1!
b100 %
1'
b100 +
#400380000000
0!
0'
#400390000000
1!
b101 %
1'
b101 +
#400400000000
0!
0'
#400410000000
1!
0$
b110 %
1'
0*
b110 +
#400420000000
0!
0'
#400430000000
1!
b111 %
1'
b111 +
#400440000000
0!
0'
#400450000000
1!
b1000 %
1'
b1000 +
#400460000000
0!
0'
#400470000000
1!
b1001 %
1'
b1001 +
#400480000000
0!
0'
#400490000000
1!
b0 %
1'
b0 +
#400500000000
0!
0'
#400510000000
1!
1$
b1 %
1'
1*
b1 +
#400520000000
0!
0'
#400530000000
1!
b10 %
1'
b10 +
#400540000000
1"
1(
#400550000000
0!
0"
b100 &
0'
0(
b100 ,
#400560000000
1!
b11 %
1'
b11 +
#400570000000
0!
0'
#400580000000
1!
b100 %
1'
b100 +
#400590000000
0!
0'
#400600000000
1!
b101 %
1'
b101 +
#400610000000
0!
0'
#400620000000
1!
b110 %
1'
b110 +
#400630000000
0!
0'
#400640000000
1!
b111 %
1'
b111 +
#400650000000
0!
0'
#400660000000
1!
0$
b1000 %
1'
0*
b1000 +
#400670000000
0!
0'
#400680000000
1!
b1001 %
1'
b1001 +
#400690000000
0!
0'
#400700000000
1!
b0 %
1'
b0 +
#400710000000
0!
0'
#400720000000
1!
1$
b1 %
1'
1*
b1 +
#400730000000
0!
0'
#400740000000
1!
b10 %
1'
b10 +
#400750000000
0!
0'
#400760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#400770000000
0!
0'
#400780000000
1!
b100 %
1'
b100 +
#400790000000
0!
0'
#400800000000
1!
b101 %
1'
b101 +
#400810000000
0!
0'
#400820000000
1!
0$
b110 %
1'
0*
b110 +
#400830000000
0!
0'
#400840000000
1!
b111 %
1'
b111 +
#400850000000
0!
0'
#400860000000
1!
b1000 %
1'
b1000 +
#400870000000
0!
0'
#400880000000
1!
b1001 %
1'
b1001 +
#400890000000
0!
0'
#400900000000
1!
b0 %
1'
b0 +
#400910000000
0!
0'
#400920000000
1!
1$
b1 %
1'
1*
b1 +
#400930000000
0!
0'
#400940000000
1!
b10 %
1'
b10 +
#400950000000
0!
0'
#400960000000
1!
b11 %
1'
b11 +
#400970000000
1"
1(
#400980000000
0!
0"
b100 &
0'
0(
b100 ,
#400990000000
1!
b100 %
1'
b100 +
#401000000000
0!
0'
#401010000000
1!
b101 %
1'
b101 +
#401020000000
0!
0'
#401030000000
1!
b110 %
1'
b110 +
#401040000000
0!
0'
#401050000000
1!
b111 %
1'
b111 +
#401060000000
0!
0'
#401070000000
1!
0$
b1000 %
1'
0*
b1000 +
#401080000000
0!
0'
#401090000000
1!
b1001 %
1'
b1001 +
#401100000000
0!
0'
#401110000000
1!
b0 %
1'
b0 +
#401120000000
0!
0'
#401130000000
1!
1$
b1 %
1'
1*
b1 +
#401140000000
0!
0'
#401150000000
1!
b10 %
1'
b10 +
#401160000000
0!
0'
#401170000000
1!
b11 %
1'
b11 +
#401180000000
0!
0'
#401190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#401200000000
0!
0'
#401210000000
1!
b101 %
1'
b101 +
#401220000000
0!
0'
#401230000000
1!
0$
b110 %
1'
0*
b110 +
#401240000000
0!
0'
#401250000000
1!
b111 %
1'
b111 +
#401260000000
0!
0'
#401270000000
1!
b1000 %
1'
b1000 +
#401280000000
0!
0'
#401290000000
1!
b1001 %
1'
b1001 +
#401300000000
0!
0'
#401310000000
1!
b0 %
1'
b0 +
#401320000000
0!
0'
#401330000000
1!
1$
b1 %
1'
1*
b1 +
#401340000000
0!
0'
#401350000000
1!
b10 %
1'
b10 +
#401360000000
0!
0'
#401370000000
1!
b11 %
1'
b11 +
#401380000000
0!
0'
#401390000000
1!
b100 %
1'
b100 +
#401400000000
1"
1(
#401410000000
0!
0"
b100 &
0'
0(
b100 ,
#401420000000
1!
b101 %
1'
b101 +
#401430000000
0!
0'
#401440000000
1!
b110 %
1'
b110 +
#401450000000
0!
0'
#401460000000
1!
b111 %
1'
b111 +
#401470000000
0!
0'
#401480000000
1!
0$
b1000 %
1'
0*
b1000 +
#401490000000
0!
0'
#401500000000
1!
b1001 %
1'
b1001 +
#401510000000
0!
0'
#401520000000
1!
b0 %
1'
b0 +
#401530000000
0!
0'
#401540000000
1!
1$
b1 %
1'
1*
b1 +
#401550000000
0!
0'
#401560000000
1!
b10 %
1'
b10 +
#401570000000
0!
0'
#401580000000
1!
b11 %
1'
b11 +
#401590000000
0!
0'
#401600000000
1!
b100 %
1'
b100 +
#401610000000
0!
0'
#401620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#401630000000
0!
0'
#401640000000
1!
0$
b110 %
1'
0*
b110 +
#401650000000
0!
0'
#401660000000
1!
b111 %
1'
b111 +
#401670000000
0!
0'
#401680000000
1!
b1000 %
1'
b1000 +
#401690000000
0!
0'
#401700000000
1!
b1001 %
1'
b1001 +
#401710000000
0!
0'
#401720000000
1!
b0 %
1'
b0 +
#401730000000
0!
0'
#401740000000
1!
1$
b1 %
1'
1*
b1 +
#401750000000
0!
0'
#401760000000
1!
b10 %
1'
b10 +
#401770000000
0!
0'
#401780000000
1!
b11 %
1'
b11 +
#401790000000
0!
0'
#401800000000
1!
b100 %
1'
b100 +
#401810000000
0!
0'
#401820000000
1!
b101 %
1'
b101 +
#401830000000
1"
1(
#401840000000
0!
0"
b100 &
0'
0(
b100 ,
#401850000000
1!
b110 %
1'
b110 +
#401860000000
0!
0'
#401870000000
1!
b111 %
1'
b111 +
#401880000000
0!
0'
#401890000000
1!
0$
b1000 %
1'
0*
b1000 +
#401900000000
0!
0'
#401910000000
1!
b1001 %
1'
b1001 +
#401920000000
0!
0'
#401930000000
1!
b0 %
1'
b0 +
#401940000000
0!
0'
#401950000000
1!
1$
b1 %
1'
1*
b1 +
#401960000000
0!
0'
#401970000000
1!
b10 %
1'
b10 +
#401980000000
0!
0'
#401990000000
1!
b11 %
1'
b11 +
#402000000000
0!
0'
#402010000000
1!
b100 %
1'
b100 +
#402020000000
0!
0'
#402030000000
1!
b101 %
1'
b101 +
#402040000000
0!
0'
#402050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#402060000000
0!
0'
#402070000000
1!
b111 %
1'
b111 +
#402080000000
0!
0'
#402090000000
1!
b1000 %
1'
b1000 +
#402100000000
0!
0'
#402110000000
1!
b1001 %
1'
b1001 +
#402120000000
0!
0'
#402130000000
1!
b0 %
1'
b0 +
#402140000000
0!
0'
#402150000000
1!
1$
b1 %
1'
1*
b1 +
#402160000000
0!
0'
#402170000000
1!
b10 %
1'
b10 +
#402180000000
0!
0'
#402190000000
1!
b11 %
1'
b11 +
#402200000000
0!
0'
#402210000000
1!
b100 %
1'
b100 +
#402220000000
0!
0'
#402230000000
1!
b101 %
1'
b101 +
#402240000000
0!
0'
#402250000000
1!
0$
b110 %
1'
0*
b110 +
#402260000000
1"
1(
#402270000000
0!
0"
b100 &
0'
0(
b100 ,
#402280000000
1!
1$
b111 %
1'
1*
b111 +
#402290000000
0!
0'
#402300000000
1!
0$
b1000 %
1'
0*
b1000 +
#402310000000
0!
0'
#402320000000
1!
b1001 %
1'
b1001 +
#402330000000
0!
0'
#402340000000
1!
b0 %
1'
b0 +
#402350000000
0!
0'
#402360000000
1!
1$
b1 %
1'
1*
b1 +
#402370000000
0!
0'
#402380000000
1!
b10 %
1'
b10 +
#402390000000
0!
0'
#402400000000
1!
b11 %
1'
b11 +
#402410000000
0!
0'
#402420000000
1!
b100 %
1'
b100 +
#402430000000
0!
0'
#402440000000
1!
b101 %
1'
b101 +
#402450000000
0!
0'
#402460000000
1!
b110 %
1'
b110 +
#402470000000
0!
0'
#402480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#402490000000
0!
0'
#402500000000
1!
b1000 %
1'
b1000 +
#402510000000
0!
0'
#402520000000
1!
b1001 %
1'
b1001 +
#402530000000
0!
0'
#402540000000
1!
b0 %
1'
b0 +
#402550000000
0!
0'
#402560000000
1!
1$
b1 %
1'
1*
b1 +
#402570000000
0!
0'
#402580000000
1!
b10 %
1'
b10 +
#402590000000
0!
0'
#402600000000
1!
b11 %
1'
b11 +
#402610000000
0!
0'
#402620000000
1!
b100 %
1'
b100 +
#402630000000
0!
0'
#402640000000
1!
b101 %
1'
b101 +
#402650000000
0!
0'
#402660000000
1!
0$
b110 %
1'
0*
b110 +
#402670000000
0!
0'
#402680000000
1!
b111 %
1'
b111 +
#402690000000
1"
1(
#402700000000
0!
0"
b100 &
0'
0(
b100 ,
#402710000000
1!
b1000 %
1'
b1000 +
#402720000000
0!
0'
#402730000000
1!
b1001 %
1'
b1001 +
#402740000000
0!
0'
#402750000000
1!
b0 %
1'
b0 +
#402760000000
0!
0'
#402770000000
1!
1$
b1 %
1'
1*
b1 +
#402780000000
0!
0'
#402790000000
1!
b10 %
1'
b10 +
#402800000000
0!
0'
#402810000000
1!
b11 %
1'
b11 +
#402820000000
0!
0'
#402830000000
1!
b100 %
1'
b100 +
#402840000000
0!
0'
#402850000000
1!
b101 %
1'
b101 +
#402860000000
0!
0'
#402870000000
1!
b110 %
1'
b110 +
#402880000000
0!
0'
#402890000000
1!
b111 %
1'
b111 +
#402900000000
0!
0'
#402910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#402920000000
0!
0'
#402930000000
1!
b1001 %
1'
b1001 +
#402940000000
0!
0'
#402950000000
1!
b0 %
1'
b0 +
#402960000000
0!
0'
#402970000000
1!
1$
b1 %
1'
1*
b1 +
#402980000000
0!
0'
#402990000000
1!
b10 %
1'
b10 +
#403000000000
0!
0'
#403010000000
1!
b11 %
1'
b11 +
#403020000000
0!
0'
#403030000000
1!
b100 %
1'
b100 +
#403040000000
0!
0'
#403050000000
1!
b101 %
1'
b101 +
#403060000000
0!
0'
#403070000000
1!
0$
b110 %
1'
0*
b110 +
#403080000000
0!
0'
#403090000000
1!
b111 %
1'
b111 +
#403100000000
0!
0'
#403110000000
1!
b1000 %
1'
b1000 +
#403120000000
1"
1(
#403130000000
0!
0"
b100 &
0'
0(
b100 ,
#403140000000
1!
b1001 %
1'
b1001 +
#403150000000
0!
0'
#403160000000
1!
b0 %
1'
b0 +
#403170000000
0!
0'
#403180000000
1!
1$
b1 %
1'
1*
b1 +
#403190000000
0!
0'
#403200000000
1!
b10 %
1'
b10 +
#403210000000
0!
0'
#403220000000
1!
b11 %
1'
b11 +
#403230000000
0!
0'
#403240000000
1!
b100 %
1'
b100 +
#403250000000
0!
0'
#403260000000
1!
b101 %
1'
b101 +
#403270000000
0!
0'
#403280000000
1!
b110 %
1'
b110 +
#403290000000
0!
0'
#403300000000
1!
b111 %
1'
b111 +
#403310000000
0!
0'
#403320000000
1!
0$
b1000 %
1'
0*
b1000 +
#403330000000
0!
0'
#403340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#403350000000
0!
0'
#403360000000
1!
b0 %
1'
b0 +
#403370000000
0!
0'
#403380000000
1!
1$
b1 %
1'
1*
b1 +
#403390000000
0!
0'
#403400000000
1!
b10 %
1'
b10 +
#403410000000
0!
0'
#403420000000
1!
b11 %
1'
b11 +
#403430000000
0!
0'
#403440000000
1!
b100 %
1'
b100 +
#403450000000
0!
0'
#403460000000
1!
b101 %
1'
b101 +
#403470000000
0!
0'
#403480000000
1!
0$
b110 %
1'
0*
b110 +
#403490000000
0!
0'
#403500000000
1!
b111 %
1'
b111 +
#403510000000
0!
0'
#403520000000
1!
b1000 %
1'
b1000 +
#403530000000
0!
0'
#403540000000
1!
b1001 %
1'
b1001 +
#403550000000
1"
1(
#403560000000
0!
0"
b100 &
0'
0(
b100 ,
#403570000000
1!
b0 %
1'
b0 +
#403580000000
0!
0'
#403590000000
1!
1$
b1 %
1'
1*
b1 +
#403600000000
0!
0'
#403610000000
1!
b10 %
1'
b10 +
#403620000000
0!
0'
#403630000000
1!
b11 %
1'
b11 +
#403640000000
0!
0'
#403650000000
1!
b100 %
1'
b100 +
#403660000000
0!
0'
#403670000000
1!
b101 %
1'
b101 +
#403680000000
0!
0'
#403690000000
1!
b110 %
1'
b110 +
#403700000000
0!
0'
#403710000000
1!
b111 %
1'
b111 +
#403720000000
0!
0'
#403730000000
1!
0$
b1000 %
1'
0*
b1000 +
#403740000000
0!
0'
#403750000000
1!
b1001 %
1'
b1001 +
#403760000000
0!
0'
#403770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#403780000000
0!
0'
#403790000000
1!
1$
b1 %
1'
1*
b1 +
#403800000000
0!
0'
#403810000000
1!
b10 %
1'
b10 +
#403820000000
0!
0'
#403830000000
1!
b11 %
1'
b11 +
#403840000000
0!
0'
#403850000000
1!
b100 %
1'
b100 +
#403860000000
0!
0'
#403870000000
1!
b101 %
1'
b101 +
#403880000000
0!
0'
#403890000000
1!
0$
b110 %
1'
0*
b110 +
#403900000000
0!
0'
#403910000000
1!
b111 %
1'
b111 +
#403920000000
0!
0'
#403930000000
1!
b1000 %
1'
b1000 +
#403940000000
0!
0'
#403950000000
1!
b1001 %
1'
b1001 +
#403960000000
0!
0'
#403970000000
1!
b0 %
1'
b0 +
#403980000000
1"
1(
#403990000000
0!
0"
b100 &
0'
0(
b100 ,
#404000000000
1!
1$
b1 %
1'
1*
b1 +
#404010000000
0!
0'
#404020000000
1!
b10 %
1'
b10 +
#404030000000
0!
0'
#404040000000
1!
b11 %
1'
b11 +
#404050000000
0!
0'
#404060000000
1!
b100 %
1'
b100 +
#404070000000
0!
0'
#404080000000
1!
b101 %
1'
b101 +
#404090000000
0!
0'
#404100000000
1!
b110 %
1'
b110 +
#404110000000
0!
0'
#404120000000
1!
b111 %
1'
b111 +
#404130000000
0!
0'
#404140000000
1!
0$
b1000 %
1'
0*
b1000 +
#404150000000
0!
0'
#404160000000
1!
b1001 %
1'
b1001 +
#404170000000
0!
0'
#404180000000
1!
b0 %
1'
b0 +
#404190000000
0!
0'
#404200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#404210000000
0!
0'
#404220000000
1!
b10 %
1'
b10 +
#404230000000
0!
0'
#404240000000
1!
b11 %
1'
b11 +
#404250000000
0!
0'
#404260000000
1!
b100 %
1'
b100 +
#404270000000
0!
0'
#404280000000
1!
b101 %
1'
b101 +
#404290000000
0!
0'
#404300000000
1!
0$
b110 %
1'
0*
b110 +
#404310000000
0!
0'
#404320000000
1!
b111 %
1'
b111 +
#404330000000
0!
0'
#404340000000
1!
b1000 %
1'
b1000 +
#404350000000
0!
0'
#404360000000
1!
b1001 %
1'
b1001 +
#404370000000
0!
0'
#404380000000
1!
b0 %
1'
b0 +
#404390000000
0!
0'
#404400000000
1!
1$
b1 %
1'
1*
b1 +
#404410000000
1"
1(
#404420000000
0!
0"
b100 &
0'
0(
b100 ,
#404430000000
1!
b10 %
1'
b10 +
#404440000000
0!
0'
#404450000000
1!
b11 %
1'
b11 +
#404460000000
0!
0'
#404470000000
1!
b100 %
1'
b100 +
#404480000000
0!
0'
#404490000000
1!
b101 %
1'
b101 +
#404500000000
0!
0'
#404510000000
1!
b110 %
1'
b110 +
#404520000000
0!
0'
#404530000000
1!
b111 %
1'
b111 +
#404540000000
0!
0'
#404550000000
1!
0$
b1000 %
1'
0*
b1000 +
#404560000000
0!
0'
#404570000000
1!
b1001 %
1'
b1001 +
#404580000000
0!
0'
#404590000000
1!
b0 %
1'
b0 +
#404600000000
0!
0'
#404610000000
1!
1$
b1 %
1'
1*
b1 +
#404620000000
0!
0'
#404630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#404640000000
0!
0'
#404650000000
1!
b11 %
1'
b11 +
#404660000000
0!
0'
#404670000000
1!
b100 %
1'
b100 +
#404680000000
0!
0'
#404690000000
1!
b101 %
1'
b101 +
#404700000000
0!
0'
#404710000000
1!
0$
b110 %
1'
0*
b110 +
#404720000000
0!
0'
#404730000000
1!
b111 %
1'
b111 +
#404740000000
0!
0'
#404750000000
1!
b1000 %
1'
b1000 +
#404760000000
0!
0'
#404770000000
1!
b1001 %
1'
b1001 +
#404780000000
0!
0'
#404790000000
1!
b0 %
1'
b0 +
#404800000000
0!
0'
#404810000000
1!
1$
b1 %
1'
1*
b1 +
#404820000000
0!
0'
#404830000000
1!
b10 %
1'
b10 +
#404840000000
1"
1(
#404850000000
0!
0"
b100 &
0'
0(
b100 ,
#404860000000
1!
b11 %
1'
b11 +
#404870000000
0!
0'
#404880000000
1!
b100 %
1'
b100 +
#404890000000
0!
0'
#404900000000
1!
b101 %
1'
b101 +
#404910000000
0!
0'
#404920000000
1!
b110 %
1'
b110 +
#404930000000
0!
0'
#404940000000
1!
b111 %
1'
b111 +
#404950000000
0!
0'
#404960000000
1!
0$
b1000 %
1'
0*
b1000 +
#404970000000
0!
0'
#404980000000
1!
b1001 %
1'
b1001 +
#404990000000
0!
0'
#405000000000
1!
b0 %
1'
b0 +
#405010000000
0!
0'
#405020000000
1!
1$
b1 %
1'
1*
b1 +
#405030000000
0!
0'
#405040000000
1!
b10 %
1'
b10 +
#405050000000
0!
0'
#405060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#405070000000
0!
0'
#405080000000
1!
b100 %
1'
b100 +
#405090000000
0!
0'
#405100000000
1!
b101 %
1'
b101 +
#405110000000
0!
0'
#405120000000
1!
0$
b110 %
1'
0*
b110 +
#405130000000
0!
0'
#405140000000
1!
b111 %
1'
b111 +
#405150000000
0!
0'
#405160000000
1!
b1000 %
1'
b1000 +
#405170000000
0!
0'
#405180000000
1!
b1001 %
1'
b1001 +
#405190000000
0!
0'
#405200000000
1!
b0 %
1'
b0 +
#405210000000
0!
0'
#405220000000
1!
1$
b1 %
1'
1*
b1 +
#405230000000
0!
0'
#405240000000
1!
b10 %
1'
b10 +
#405250000000
0!
0'
#405260000000
1!
b11 %
1'
b11 +
#405270000000
1"
1(
#405280000000
0!
0"
b100 &
0'
0(
b100 ,
#405290000000
1!
b100 %
1'
b100 +
#405300000000
0!
0'
#405310000000
1!
b101 %
1'
b101 +
#405320000000
0!
0'
#405330000000
1!
b110 %
1'
b110 +
#405340000000
0!
0'
#405350000000
1!
b111 %
1'
b111 +
#405360000000
0!
0'
#405370000000
1!
0$
b1000 %
1'
0*
b1000 +
#405380000000
0!
0'
#405390000000
1!
b1001 %
1'
b1001 +
#405400000000
0!
0'
#405410000000
1!
b0 %
1'
b0 +
#405420000000
0!
0'
#405430000000
1!
1$
b1 %
1'
1*
b1 +
#405440000000
0!
0'
#405450000000
1!
b10 %
1'
b10 +
#405460000000
0!
0'
#405470000000
1!
b11 %
1'
b11 +
#405480000000
0!
0'
#405490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#405500000000
0!
0'
#405510000000
1!
b101 %
1'
b101 +
#405520000000
0!
0'
#405530000000
1!
0$
b110 %
1'
0*
b110 +
#405540000000
0!
0'
#405550000000
1!
b111 %
1'
b111 +
#405560000000
0!
0'
#405570000000
1!
b1000 %
1'
b1000 +
#405580000000
0!
0'
#405590000000
1!
b1001 %
1'
b1001 +
#405600000000
0!
0'
#405610000000
1!
b0 %
1'
b0 +
#405620000000
0!
0'
#405630000000
1!
1$
b1 %
1'
1*
b1 +
#405640000000
0!
0'
#405650000000
1!
b10 %
1'
b10 +
#405660000000
0!
0'
#405670000000
1!
b11 %
1'
b11 +
#405680000000
0!
0'
#405690000000
1!
b100 %
1'
b100 +
#405700000000
1"
1(
#405710000000
0!
0"
b100 &
0'
0(
b100 ,
#405720000000
1!
b101 %
1'
b101 +
#405730000000
0!
0'
#405740000000
1!
b110 %
1'
b110 +
#405750000000
0!
0'
#405760000000
1!
b111 %
1'
b111 +
#405770000000
0!
0'
#405780000000
1!
0$
b1000 %
1'
0*
b1000 +
#405790000000
0!
0'
#405800000000
1!
b1001 %
1'
b1001 +
#405810000000
0!
0'
#405820000000
1!
b0 %
1'
b0 +
#405830000000
0!
0'
#405840000000
1!
1$
b1 %
1'
1*
b1 +
#405850000000
0!
0'
#405860000000
1!
b10 %
1'
b10 +
#405870000000
0!
0'
#405880000000
1!
b11 %
1'
b11 +
#405890000000
0!
0'
#405900000000
1!
b100 %
1'
b100 +
#405910000000
0!
0'
#405920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#405930000000
0!
0'
#405940000000
1!
0$
b110 %
1'
0*
b110 +
#405950000000
0!
0'
#405960000000
1!
b111 %
1'
b111 +
#405970000000
0!
0'
#405980000000
1!
b1000 %
1'
b1000 +
#405990000000
0!
0'
#406000000000
1!
b1001 %
1'
b1001 +
#406010000000
0!
0'
#406020000000
1!
b0 %
1'
b0 +
#406030000000
0!
0'
#406040000000
1!
1$
b1 %
1'
1*
b1 +
#406050000000
0!
0'
#406060000000
1!
b10 %
1'
b10 +
#406070000000
0!
0'
#406080000000
1!
b11 %
1'
b11 +
#406090000000
0!
0'
#406100000000
1!
b100 %
1'
b100 +
#406110000000
0!
0'
#406120000000
1!
b101 %
1'
b101 +
#406130000000
1"
1(
#406140000000
0!
0"
b100 &
0'
0(
b100 ,
#406150000000
1!
b110 %
1'
b110 +
#406160000000
0!
0'
#406170000000
1!
b111 %
1'
b111 +
#406180000000
0!
0'
#406190000000
1!
0$
b1000 %
1'
0*
b1000 +
#406200000000
0!
0'
#406210000000
1!
b1001 %
1'
b1001 +
#406220000000
0!
0'
#406230000000
1!
b0 %
1'
b0 +
#406240000000
0!
0'
#406250000000
1!
1$
b1 %
1'
1*
b1 +
#406260000000
0!
0'
#406270000000
1!
b10 %
1'
b10 +
#406280000000
0!
0'
#406290000000
1!
b11 %
1'
b11 +
#406300000000
0!
0'
#406310000000
1!
b100 %
1'
b100 +
#406320000000
0!
0'
#406330000000
1!
b101 %
1'
b101 +
#406340000000
0!
0'
#406350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#406360000000
0!
0'
#406370000000
1!
b111 %
1'
b111 +
#406380000000
0!
0'
#406390000000
1!
b1000 %
1'
b1000 +
#406400000000
0!
0'
#406410000000
1!
b1001 %
1'
b1001 +
#406420000000
0!
0'
#406430000000
1!
b0 %
1'
b0 +
#406440000000
0!
0'
#406450000000
1!
1$
b1 %
1'
1*
b1 +
#406460000000
0!
0'
#406470000000
1!
b10 %
1'
b10 +
#406480000000
0!
0'
#406490000000
1!
b11 %
1'
b11 +
#406500000000
0!
0'
#406510000000
1!
b100 %
1'
b100 +
#406520000000
0!
0'
#406530000000
1!
b101 %
1'
b101 +
#406540000000
0!
0'
#406550000000
1!
0$
b110 %
1'
0*
b110 +
#406560000000
1"
1(
#406570000000
0!
0"
b100 &
0'
0(
b100 ,
#406580000000
1!
1$
b111 %
1'
1*
b111 +
#406590000000
0!
0'
#406600000000
1!
0$
b1000 %
1'
0*
b1000 +
#406610000000
0!
0'
#406620000000
1!
b1001 %
1'
b1001 +
#406630000000
0!
0'
#406640000000
1!
b0 %
1'
b0 +
#406650000000
0!
0'
#406660000000
1!
1$
b1 %
1'
1*
b1 +
#406670000000
0!
0'
#406680000000
1!
b10 %
1'
b10 +
#406690000000
0!
0'
#406700000000
1!
b11 %
1'
b11 +
#406710000000
0!
0'
#406720000000
1!
b100 %
1'
b100 +
#406730000000
0!
0'
#406740000000
1!
b101 %
1'
b101 +
#406750000000
0!
0'
#406760000000
1!
b110 %
1'
b110 +
#406770000000
0!
0'
#406780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#406790000000
0!
0'
#406800000000
1!
b1000 %
1'
b1000 +
#406810000000
0!
0'
#406820000000
1!
b1001 %
1'
b1001 +
#406830000000
0!
0'
#406840000000
1!
b0 %
1'
b0 +
#406850000000
0!
0'
#406860000000
1!
1$
b1 %
1'
1*
b1 +
#406870000000
0!
0'
#406880000000
1!
b10 %
1'
b10 +
#406890000000
0!
0'
#406900000000
1!
b11 %
1'
b11 +
#406910000000
0!
0'
#406920000000
1!
b100 %
1'
b100 +
#406930000000
0!
0'
#406940000000
1!
b101 %
1'
b101 +
#406950000000
0!
0'
#406960000000
1!
0$
b110 %
1'
0*
b110 +
#406970000000
0!
0'
#406980000000
1!
b111 %
1'
b111 +
#406990000000
1"
1(
#407000000000
0!
0"
b100 &
0'
0(
b100 ,
#407010000000
1!
b1000 %
1'
b1000 +
#407020000000
0!
0'
#407030000000
1!
b1001 %
1'
b1001 +
#407040000000
0!
0'
#407050000000
1!
b0 %
1'
b0 +
#407060000000
0!
0'
#407070000000
1!
1$
b1 %
1'
1*
b1 +
#407080000000
0!
0'
#407090000000
1!
b10 %
1'
b10 +
#407100000000
0!
0'
#407110000000
1!
b11 %
1'
b11 +
#407120000000
0!
0'
#407130000000
1!
b100 %
1'
b100 +
#407140000000
0!
0'
#407150000000
1!
b101 %
1'
b101 +
#407160000000
0!
0'
#407170000000
1!
b110 %
1'
b110 +
#407180000000
0!
0'
#407190000000
1!
b111 %
1'
b111 +
#407200000000
0!
0'
#407210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#407220000000
0!
0'
#407230000000
1!
b1001 %
1'
b1001 +
#407240000000
0!
0'
#407250000000
1!
b0 %
1'
b0 +
#407260000000
0!
0'
#407270000000
1!
1$
b1 %
1'
1*
b1 +
#407280000000
0!
0'
#407290000000
1!
b10 %
1'
b10 +
#407300000000
0!
0'
#407310000000
1!
b11 %
1'
b11 +
#407320000000
0!
0'
#407330000000
1!
b100 %
1'
b100 +
#407340000000
0!
0'
#407350000000
1!
b101 %
1'
b101 +
#407360000000
0!
0'
#407370000000
1!
0$
b110 %
1'
0*
b110 +
#407380000000
0!
0'
#407390000000
1!
b111 %
1'
b111 +
#407400000000
0!
0'
#407410000000
1!
b1000 %
1'
b1000 +
#407420000000
1"
1(
#407430000000
0!
0"
b100 &
0'
0(
b100 ,
#407440000000
1!
b1001 %
1'
b1001 +
#407450000000
0!
0'
#407460000000
1!
b0 %
1'
b0 +
#407470000000
0!
0'
#407480000000
1!
1$
b1 %
1'
1*
b1 +
#407490000000
0!
0'
#407500000000
1!
b10 %
1'
b10 +
#407510000000
0!
0'
#407520000000
1!
b11 %
1'
b11 +
#407530000000
0!
0'
#407540000000
1!
b100 %
1'
b100 +
#407550000000
0!
0'
#407560000000
1!
b101 %
1'
b101 +
#407570000000
0!
0'
#407580000000
1!
b110 %
1'
b110 +
#407590000000
0!
0'
#407600000000
1!
b111 %
1'
b111 +
#407610000000
0!
0'
#407620000000
1!
0$
b1000 %
1'
0*
b1000 +
#407630000000
0!
0'
#407640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#407650000000
0!
0'
#407660000000
1!
b0 %
1'
b0 +
#407670000000
0!
0'
#407680000000
1!
1$
b1 %
1'
1*
b1 +
#407690000000
0!
0'
#407700000000
1!
b10 %
1'
b10 +
#407710000000
0!
0'
#407720000000
1!
b11 %
1'
b11 +
#407730000000
0!
0'
#407740000000
1!
b100 %
1'
b100 +
#407750000000
0!
0'
#407760000000
1!
b101 %
1'
b101 +
#407770000000
0!
0'
#407780000000
1!
0$
b110 %
1'
0*
b110 +
#407790000000
0!
0'
#407800000000
1!
b111 %
1'
b111 +
#407810000000
0!
0'
#407820000000
1!
b1000 %
1'
b1000 +
#407830000000
0!
0'
#407840000000
1!
b1001 %
1'
b1001 +
#407850000000
1"
1(
#407860000000
0!
0"
b100 &
0'
0(
b100 ,
#407870000000
1!
b0 %
1'
b0 +
#407880000000
0!
0'
#407890000000
1!
1$
b1 %
1'
1*
b1 +
#407900000000
0!
0'
#407910000000
1!
b10 %
1'
b10 +
#407920000000
0!
0'
#407930000000
1!
b11 %
1'
b11 +
#407940000000
0!
0'
#407950000000
1!
b100 %
1'
b100 +
#407960000000
0!
0'
#407970000000
1!
b101 %
1'
b101 +
#407980000000
0!
0'
#407990000000
1!
b110 %
1'
b110 +
#408000000000
0!
0'
#408010000000
1!
b111 %
1'
b111 +
#408020000000
0!
0'
#408030000000
1!
0$
b1000 %
1'
0*
b1000 +
#408040000000
0!
0'
#408050000000
1!
b1001 %
1'
b1001 +
#408060000000
0!
0'
#408070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#408080000000
0!
0'
#408090000000
1!
1$
b1 %
1'
1*
b1 +
#408100000000
0!
0'
#408110000000
1!
b10 %
1'
b10 +
#408120000000
0!
0'
#408130000000
1!
b11 %
1'
b11 +
#408140000000
0!
0'
#408150000000
1!
b100 %
1'
b100 +
#408160000000
0!
0'
#408170000000
1!
b101 %
1'
b101 +
#408180000000
0!
0'
#408190000000
1!
0$
b110 %
1'
0*
b110 +
#408200000000
0!
0'
#408210000000
1!
b111 %
1'
b111 +
#408220000000
0!
0'
#408230000000
1!
b1000 %
1'
b1000 +
#408240000000
0!
0'
#408250000000
1!
b1001 %
1'
b1001 +
#408260000000
0!
0'
#408270000000
1!
b0 %
1'
b0 +
#408280000000
1"
1(
#408290000000
0!
0"
b100 &
0'
0(
b100 ,
#408300000000
1!
1$
b1 %
1'
1*
b1 +
#408310000000
0!
0'
#408320000000
1!
b10 %
1'
b10 +
#408330000000
0!
0'
#408340000000
1!
b11 %
1'
b11 +
#408350000000
0!
0'
#408360000000
1!
b100 %
1'
b100 +
#408370000000
0!
0'
#408380000000
1!
b101 %
1'
b101 +
#408390000000
0!
0'
#408400000000
1!
b110 %
1'
b110 +
#408410000000
0!
0'
#408420000000
1!
b111 %
1'
b111 +
#408430000000
0!
0'
#408440000000
1!
0$
b1000 %
1'
0*
b1000 +
#408450000000
0!
0'
#408460000000
1!
b1001 %
1'
b1001 +
#408470000000
0!
0'
#408480000000
1!
b0 %
1'
b0 +
#408490000000
0!
0'
#408500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#408510000000
0!
0'
#408520000000
1!
b10 %
1'
b10 +
#408530000000
0!
0'
#408540000000
1!
b11 %
1'
b11 +
#408550000000
0!
0'
#408560000000
1!
b100 %
1'
b100 +
#408570000000
0!
0'
#408580000000
1!
b101 %
1'
b101 +
#408590000000
0!
0'
#408600000000
1!
0$
b110 %
1'
0*
b110 +
#408610000000
0!
0'
#408620000000
1!
b111 %
1'
b111 +
#408630000000
0!
0'
#408640000000
1!
b1000 %
1'
b1000 +
#408650000000
0!
0'
#408660000000
1!
b1001 %
1'
b1001 +
#408670000000
0!
0'
#408680000000
1!
b0 %
1'
b0 +
#408690000000
0!
0'
#408700000000
1!
1$
b1 %
1'
1*
b1 +
#408710000000
1"
1(
#408720000000
0!
0"
b100 &
0'
0(
b100 ,
#408730000000
1!
b10 %
1'
b10 +
#408740000000
0!
0'
#408750000000
1!
b11 %
1'
b11 +
#408760000000
0!
0'
#408770000000
1!
b100 %
1'
b100 +
#408780000000
0!
0'
#408790000000
1!
b101 %
1'
b101 +
#408800000000
0!
0'
#408810000000
1!
b110 %
1'
b110 +
#408820000000
0!
0'
#408830000000
1!
b111 %
1'
b111 +
#408840000000
0!
0'
#408850000000
1!
0$
b1000 %
1'
0*
b1000 +
#408860000000
0!
0'
#408870000000
1!
b1001 %
1'
b1001 +
#408880000000
0!
0'
#408890000000
1!
b0 %
1'
b0 +
#408900000000
0!
0'
#408910000000
1!
1$
b1 %
1'
1*
b1 +
#408920000000
0!
0'
#408930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#408940000000
0!
0'
#408950000000
1!
b11 %
1'
b11 +
#408960000000
0!
0'
#408970000000
1!
b100 %
1'
b100 +
#408980000000
0!
0'
#408990000000
1!
b101 %
1'
b101 +
#409000000000
0!
0'
#409010000000
1!
0$
b110 %
1'
0*
b110 +
#409020000000
0!
0'
#409030000000
1!
b111 %
1'
b111 +
#409040000000
0!
0'
#409050000000
1!
b1000 %
1'
b1000 +
#409060000000
0!
0'
#409070000000
1!
b1001 %
1'
b1001 +
#409080000000
0!
0'
#409090000000
1!
b0 %
1'
b0 +
#409100000000
0!
0'
#409110000000
1!
1$
b1 %
1'
1*
b1 +
#409120000000
0!
0'
#409130000000
1!
b10 %
1'
b10 +
#409140000000
1"
1(
#409150000000
0!
0"
b100 &
0'
0(
b100 ,
#409160000000
1!
b11 %
1'
b11 +
#409170000000
0!
0'
#409180000000
1!
b100 %
1'
b100 +
#409190000000
0!
0'
#409200000000
1!
b101 %
1'
b101 +
#409210000000
0!
0'
#409220000000
1!
b110 %
1'
b110 +
#409230000000
0!
0'
#409240000000
1!
b111 %
1'
b111 +
#409250000000
0!
0'
#409260000000
1!
0$
b1000 %
1'
0*
b1000 +
#409270000000
0!
0'
#409280000000
1!
b1001 %
1'
b1001 +
#409290000000
0!
0'
#409300000000
1!
b0 %
1'
b0 +
#409310000000
0!
0'
#409320000000
1!
1$
b1 %
1'
1*
b1 +
#409330000000
0!
0'
#409340000000
1!
b10 %
1'
b10 +
#409350000000
0!
0'
#409360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#409370000000
0!
0'
#409380000000
1!
b100 %
1'
b100 +
#409390000000
0!
0'
#409400000000
1!
b101 %
1'
b101 +
#409410000000
0!
0'
#409420000000
1!
0$
b110 %
1'
0*
b110 +
#409430000000
0!
0'
#409440000000
1!
b111 %
1'
b111 +
#409450000000
0!
0'
#409460000000
1!
b1000 %
1'
b1000 +
#409470000000
0!
0'
#409480000000
1!
b1001 %
1'
b1001 +
#409490000000
0!
0'
#409500000000
1!
b0 %
1'
b0 +
#409510000000
0!
0'
#409520000000
1!
1$
b1 %
1'
1*
b1 +
#409530000000
0!
0'
#409540000000
1!
b10 %
1'
b10 +
#409550000000
0!
0'
#409560000000
1!
b11 %
1'
b11 +
#409570000000
1"
1(
#409580000000
0!
0"
b100 &
0'
0(
b100 ,
#409590000000
1!
b100 %
1'
b100 +
#409600000000
0!
0'
#409610000000
1!
b101 %
1'
b101 +
#409620000000
0!
0'
#409630000000
1!
b110 %
1'
b110 +
#409640000000
0!
0'
#409650000000
1!
b111 %
1'
b111 +
#409660000000
0!
0'
#409670000000
1!
0$
b1000 %
1'
0*
b1000 +
#409680000000
0!
0'
#409690000000
1!
b1001 %
1'
b1001 +
#409700000000
0!
0'
#409710000000
1!
b0 %
1'
b0 +
#409720000000
0!
0'
#409730000000
1!
1$
b1 %
1'
1*
b1 +
#409740000000
0!
0'
#409750000000
1!
b10 %
1'
b10 +
#409760000000
0!
0'
#409770000000
1!
b11 %
1'
b11 +
#409780000000
0!
0'
#409790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#409800000000
0!
0'
#409810000000
1!
b101 %
1'
b101 +
#409820000000
0!
0'
#409830000000
1!
0$
b110 %
1'
0*
b110 +
#409840000000
0!
0'
#409850000000
1!
b111 %
1'
b111 +
#409860000000
0!
0'
#409870000000
1!
b1000 %
1'
b1000 +
#409880000000
0!
0'
#409890000000
1!
b1001 %
1'
b1001 +
#409900000000
0!
0'
#409910000000
1!
b0 %
1'
b0 +
#409920000000
0!
0'
#409930000000
1!
1$
b1 %
1'
1*
b1 +
#409940000000
0!
0'
#409950000000
1!
b10 %
1'
b10 +
#409960000000
0!
0'
#409970000000
1!
b11 %
1'
b11 +
#409980000000
0!
0'
#409990000000
1!
b100 %
1'
b100 +
#410000000000
1"
1(
#410010000000
0!
0"
b100 &
0'
0(
b100 ,
#410020000000
1!
b101 %
1'
b101 +
#410030000000
0!
0'
#410040000000
1!
b110 %
1'
b110 +
#410050000000
0!
0'
#410060000000
1!
b111 %
1'
b111 +
#410070000000
0!
0'
#410080000000
1!
0$
b1000 %
1'
0*
b1000 +
#410090000000
0!
0'
#410100000000
1!
b1001 %
1'
b1001 +
#410110000000
0!
0'
#410120000000
1!
b0 %
1'
b0 +
#410130000000
0!
0'
#410140000000
1!
1$
b1 %
1'
1*
b1 +
#410150000000
0!
0'
#410160000000
1!
b10 %
1'
b10 +
#410170000000
0!
0'
#410180000000
1!
b11 %
1'
b11 +
#410190000000
0!
0'
#410200000000
1!
b100 %
1'
b100 +
#410210000000
0!
0'
#410220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#410230000000
0!
0'
#410240000000
1!
0$
b110 %
1'
0*
b110 +
#410250000000
0!
0'
#410260000000
1!
b111 %
1'
b111 +
#410270000000
0!
0'
#410280000000
1!
b1000 %
1'
b1000 +
#410290000000
0!
0'
#410300000000
1!
b1001 %
1'
b1001 +
#410310000000
0!
0'
#410320000000
1!
b0 %
1'
b0 +
#410330000000
0!
0'
#410340000000
1!
1$
b1 %
1'
1*
b1 +
#410350000000
0!
0'
#410360000000
1!
b10 %
1'
b10 +
#410370000000
0!
0'
#410380000000
1!
b11 %
1'
b11 +
#410390000000
0!
0'
#410400000000
1!
b100 %
1'
b100 +
#410410000000
0!
0'
#410420000000
1!
b101 %
1'
b101 +
#410430000000
1"
1(
#410440000000
0!
0"
b100 &
0'
0(
b100 ,
#410450000000
1!
b110 %
1'
b110 +
#410460000000
0!
0'
#410470000000
1!
b111 %
1'
b111 +
#410480000000
0!
0'
#410490000000
1!
0$
b1000 %
1'
0*
b1000 +
#410500000000
0!
0'
#410510000000
1!
b1001 %
1'
b1001 +
#410520000000
0!
0'
#410530000000
1!
b0 %
1'
b0 +
#410540000000
0!
0'
#410550000000
1!
1$
b1 %
1'
1*
b1 +
#410560000000
0!
0'
#410570000000
1!
b10 %
1'
b10 +
#410580000000
0!
0'
#410590000000
1!
b11 %
1'
b11 +
#410600000000
0!
0'
#410610000000
1!
b100 %
1'
b100 +
#410620000000
0!
0'
#410630000000
1!
b101 %
1'
b101 +
#410640000000
0!
0'
#410650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#410660000000
0!
0'
#410670000000
1!
b111 %
1'
b111 +
#410680000000
0!
0'
#410690000000
1!
b1000 %
1'
b1000 +
#410700000000
0!
0'
#410710000000
1!
b1001 %
1'
b1001 +
#410720000000
0!
0'
#410730000000
1!
b0 %
1'
b0 +
#410740000000
0!
0'
#410750000000
1!
1$
b1 %
1'
1*
b1 +
#410760000000
0!
0'
#410770000000
1!
b10 %
1'
b10 +
#410780000000
0!
0'
#410790000000
1!
b11 %
1'
b11 +
#410800000000
0!
0'
#410810000000
1!
b100 %
1'
b100 +
#410820000000
0!
0'
#410830000000
1!
b101 %
1'
b101 +
#410840000000
0!
0'
#410850000000
1!
0$
b110 %
1'
0*
b110 +
#410860000000
1"
1(
#410870000000
0!
0"
b100 &
0'
0(
b100 ,
#410880000000
1!
1$
b111 %
1'
1*
b111 +
#410890000000
0!
0'
#410900000000
1!
0$
b1000 %
1'
0*
b1000 +
#410910000000
0!
0'
#410920000000
1!
b1001 %
1'
b1001 +
#410930000000
0!
0'
#410940000000
1!
b0 %
1'
b0 +
#410950000000
0!
0'
#410960000000
1!
1$
b1 %
1'
1*
b1 +
#410970000000
0!
0'
#410980000000
1!
b10 %
1'
b10 +
#410990000000
0!
0'
#411000000000
1!
b11 %
1'
b11 +
#411010000000
0!
0'
#411020000000
1!
b100 %
1'
b100 +
#411030000000
0!
0'
#411040000000
1!
b101 %
1'
b101 +
#411050000000
0!
0'
#411060000000
1!
b110 %
1'
b110 +
#411070000000
0!
0'
#411080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#411090000000
0!
0'
#411100000000
1!
b1000 %
1'
b1000 +
#411110000000
0!
0'
#411120000000
1!
b1001 %
1'
b1001 +
#411130000000
0!
0'
#411140000000
1!
b0 %
1'
b0 +
#411150000000
0!
0'
#411160000000
1!
1$
b1 %
1'
1*
b1 +
#411170000000
0!
0'
#411180000000
1!
b10 %
1'
b10 +
#411190000000
0!
0'
#411200000000
1!
b11 %
1'
b11 +
#411210000000
0!
0'
#411220000000
1!
b100 %
1'
b100 +
#411230000000
0!
0'
#411240000000
1!
b101 %
1'
b101 +
#411250000000
0!
0'
#411260000000
1!
0$
b110 %
1'
0*
b110 +
#411270000000
0!
0'
#411280000000
1!
b111 %
1'
b111 +
#411290000000
1"
1(
#411300000000
0!
0"
b100 &
0'
0(
b100 ,
#411310000000
1!
b1000 %
1'
b1000 +
#411320000000
0!
0'
#411330000000
1!
b1001 %
1'
b1001 +
#411340000000
0!
0'
#411350000000
1!
b0 %
1'
b0 +
#411360000000
0!
0'
#411370000000
1!
1$
b1 %
1'
1*
b1 +
#411380000000
0!
0'
#411390000000
1!
b10 %
1'
b10 +
#411400000000
0!
0'
#411410000000
1!
b11 %
1'
b11 +
#411420000000
0!
0'
#411430000000
1!
b100 %
1'
b100 +
#411440000000
0!
0'
#411450000000
1!
b101 %
1'
b101 +
#411460000000
0!
0'
#411470000000
1!
b110 %
1'
b110 +
#411480000000
0!
0'
#411490000000
1!
b111 %
1'
b111 +
#411500000000
0!
0'
#411510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#411520000000
0!
0'
#411530000000
1!
b1001 %
1'
b1001 +
#411540000000
0!
0'
#411550000000
1!
b0 %
1'
b0 +
#411560000000
0!
0'
#411570000000
1!
1$
b1 %
1'
1*
b1 +
#411580000000
0!
0'
#411590000000
1!
b10 %
1'
b10 +
#411600000000
0!
0'
#411610000000
1!
b11 %
1'
b11 +
#411620000000
0!
0'
#411630000000
1!
b100 %
1'
b100 +
#411640000000
0!
0'
#411650000000
1!
b101 %
1'
b101 +
#411660000000
0!
0'
#411670000000
1!
0$
b110 %
1'
0*
b110 +
#411680000000
0!
0'
#411690000000
1!
b111 %
1'
b111 +
#411700000000
0!
0'
#411710000000
1!
b1000 %
1'
b1000 +
#411720000000
1"
1(
#411730000000
0!
0"
b100 &
0'
0(
b100 ,
#411740000000
1!
b1001 %
1'
b1001 +
#411750000000
0!
0'
#411760000000
1!
b0 %
1'
b0 +
#411770000000
0!
0'
#411780000000
1!
1$
b1 %
1'
1*
b1 +
#411790000000
0!
0'
#411800000000
1!
b10 %
1'
b10 +
#411810000000
0!
0'
#411820000000
1!
b11 %
1'
b11 +
#411830000000
0!
0'
#411840000000
1!
b100 %
1'
b100 +
#411850000000
0!
0'
#411860000000
1!
b101 %
1'
b101 +
#411870000000
0!
0'
#411880000000
1!
b110 %
1'
b110 +
#411890000000
0!
0'
#411900000000
1!
b111 %
1'
b111 +
#411910000000
0!
0'
#411920000000
1!
0$
b1000 %
1'
0*
b1000 +
#411930000000
0!
0'
#411940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#411950000000
0!
0'
#411960000000
1!
b0 %
1'
b0 +
#411970000000
0!
0'
#411980000000
1!
1$
b1 %
1'
1*
b1 +
#411990000000
0!
0'
#412000000000
1!
b10 %
1'
b10 +
#412010000000
0!
0'
#412020000000
1!
b11 %
1'
b11 +
#412030000000
0!
0'
#412040000000
1!
b100 %
1'
b100 +
#412050000000
0!
0'
#412060000000
1!
b101 %
1'
b101 +
#412070000000
0!
0'
#412080000000
1!
0$
b110 %
1'
0*
b110 +
#412090000000
0!
0'
#412100000000
1!
b111 %
1'
b111 +
#412110000000
0!
0'
#412120000000
1!
b1000 %
1'
b1000 +
#412130000000
0!
0'
#412140000000
1!
b1001 %
1'
b1001 +
#412150000000
1"
1(
#412160000000
0!
0"
b100 &
0'
0(
b100 ,
#412170000000
1!
b0 %
1'
b0 +
#412180000000
0!
0'
#412190000000
1!
1$
b1 %
1'
1*
b1 +
#412200000000
0!
0'
#412210000000
1!
b10 %
1'
b10 +
#412220000000
0!
0'
#412230000000
1!
b11 %
1'
b11 +
#412240000000
0!
0'
#412250000000
1!
b100 %
1'
b100 +
#412260000000
0!
0'
#412270000000
1!
b101 %
1'
b101 +
#412280000000
0!
0'
#412290000000
1!
b110 %
1'
b110 +
#412300000000
0!
0'
#412310000000
1!
b111 %
1'
b111 +
#412320000000
0!
0'
#412330000000
1!
0$
b1000 %
1'
0*
b1000 +
#412340000000
0!
0'
#412350000000
1!
b1001 %
1'
b1001 +
#412360000000
0!
0'
#412370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#412380000000
0!
0'
#412390000000
1!
1$
b1 %
1'
1*
b1 +
#412400000000
0!
0'
#412410000000
1!
b10 %
1'
b10 +
#412420000000
0!
0'
#412430000000
1!
b11 %
1'
b11 +
#412440000000
0!
0'
#412450000000
1!
b100 %
1'
b100 +
#412460000000
0!
0'
#412470000000
1!
b101 %
1'
b101 +
#412480000000
0!
0'
#412490000000
1!
0$
b110 %
1'
0*
b110 +
#412500000000
0!
0'
#412510000000
1!
b111 %
1'
b111 +
#412520000000
0!
0'
#412530000000
1!
b1000 %
1'
b1000 +
#412540000000
0!
0'
#412550000000
1!
b1001 %
1'
b1001 +
#412560000000
0!
0'
#412570000000
1!
b0 %
1'
b0 +
#412580000000
1"
1(
#412590000000
0!
0"
b100 &
0'
0(
b100 ,
#412600000000
1!
1$
b1 %
1'
1*
b1 +
#412610000000
0!
0'
#412620000000
1!
b10 %
1'
b10 +
#412630000000
0!
0'
#412640000000
1!
b11 %
1'
b11 +
#412650000000
0!
0'
#412660000000
1!
b100 %
1'
b100 +
#412670000000
0!
0'
#412680000000
1!
b101 %
1'
b101 +
#412690000000
0!
0'
#412700000000
1!
b110 %
1'
b110 +
#412710000000
0!
0'
#412720000000
1!
b111 %
1'
b111 +
#412730000000
0!
0'
#412740000000
1!
0$
b1000 %
1'
0*
b1000 +
#412750000000
0!
0'
#412760000000
1!
b1001 %
1'
b1001 +
#412770000000
0!
0'
#412780000000
1!
b0 %
1'
b0 +
#412790000000
0!
0'
#412800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#412810000000
0!
0'
#412820000000
1!
b10 %
1'
b10 +
#412830000000
0!
0'
#412840000000
1!
b11 %
1'
b11 +
#412850000000
0!
0'
#412860000000
1!
b100 %
1'
b100 +
#412870000000
0!
0'
#412880000000
1!
b101 %
1'
b101 +
#412890000000
0!
0'
#412900000000
1!
0$
b110 %
1'
0*
b110 +
#412910000000
0!
0'
#412920000000
1!
b111 %
1'
b111 +
#412930000000
0!
0'
#412940000000
1!
b1000 %
1'
b1000 +
#412950000000
0!
0'
#412960000000
1!
b1001 %
1'
b1001 +
#412970000000
0!
0'
#412980000000
1!
b0 %
1'
b0 +
#412990000000
0!
0'
#413000000000
1!
1$
b1 %
1'
1*
b1 +
#413010000000
1"
1(
#413020000000
0!
0"
b100 &
0'
0(
b100 ,
#413030000000
1!
b10 %
1'
b10 +
#413040000000
0!
0'
#413050000000
1!
b11 %
1'
b11 +
#413060000000
0!
0'
#413070000000
1!
b100 %
1'
b100 +
#413080000000
0!
0'
#413090000000
1!
b101 %
1'
b101 +
#413100000000
0!
0'
#413110000000
1!
b110 %
1'
b110 +
#413120000000
0!
0'
#413130000000
1!
b111 %
1'
b111 +
#413140000000
0!
0'
#413150000000
1!
0$
b1000 %
1'
0*
b1000 +
#413160000000
0!
0'
#413170000000
1!
b1001 %
1'
b1001 +
#413180000000
0!
0'
#413190000000
1!
b0 %
1'
b0 +
#413200000000
0!
0'
#413210000000
1!
1$
b1 %
1'
1*
b1 +
#413220000000
0!
0'
#413230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#413240000000
0!
0'
#413250000000
1!
b11 %
1'
b11 +
#413260000000
0!
0'
#413270000000
1!
b100 %
1'
b100 +
#413280000000
0!
0'
#413290000000
1!
b101 %
1'
b101 +
#413300000000
0!
0'
#413310000000
1!
0$
b110 %
1'
0*
b110 +
#413320000000
0!
0'
#413330000000
1!
b111 %
1'
b111 +
#413340000000
0!
0'
#413350000000
1!
b1000 %
1'
b1000 +
#413360000000
0!
0'
#413370000000
1!
b1001 %
1'
b1001 +
#413380000000
0!
0'
#413390000000
1!
b0 %
1'
b0 +
#413400000000
0!
0'
#413410000000
1!
1$
b1 %
1'
1*
b1 +
#413420000000
0!
0'
#413430000000
1!
b10 %
1'
b10 +
#413440000000
1"
1(
#413450000000
0!
0"
b100 &
0'
0(
b100 ,
#413460000000
1!
b11 %
1'
b11 +
#413470000000
0!
0'
#413480000000
1!
b100 %
1'
b100 +
#413490000000
0!
0'
#413500000000
1!
b101 %
1'
b101 +
#413510000000
0!
0'
#413520000000
1!
b110 %
1'
b110 +
#413530000000
0!
0'
#413540000000
1!
b111 %
1'
b111 +
#413550000000
0!
0'
#413560000000
1!
0$
b1000 %
1'
0*
b1000 +
#413570000000
0!
0'
#413580000000
1!
b1001 %
1'
b1001 +
#413590000000
0!
0'
#413600000000
1!
b0 %
1'
b0 +
#413610000000
0!
0'
#413620000000
1!
1$
b1 %
1'
1*
b1 +
#413630000000
0!
0'
#413640000000
1!
b10 %
1'
b10 +
#413650000000
0!
0'
#413660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#413670000000
0!
0'
#413680000000
1!
b100 %
1'
b100 +
#413690000000
0!
0'
#413700000000
1!
b101 %
1'
b101 +
#413710000000
0!
0'
#413720000000
1!
0$
b110 %
1'
0*
b110 +
#413730000000
0!
0'
#413740000000
1!
b111 %
1'
b111 +
#413750000000
0!
0'
#413760000000
1!
b1000 %
1'
b1000 +
#413770000000
0!
0'
#413780000000
1!
b1001 %
1'
b1001 +
#413790000000
0!
0'
#413800000000
1!
b0 %
1'
b0 +
#413810000000
0!
0'
#413820000000
1!
1$
b1 %
1'
1*
b1 +
#413830000000
0!
0'
#413840000000
1!
b10 %
1'
b10 +
#413850000000
0!
0'
#413860000000
1!
b11 %
1'
b11 +
#413870000000
1"
1(
#413880000000
0!
0"
b100 &
0'
0(
b100 ,
#413890000000
1!
b100 %
1'
b100 +
#413900000000
0!
0'
#413910000000
1!
b101 %
1'
b101 +
#413920000000
0!
0'
#413930000000
1!
b110 %
1'
b110 +
#413940000000
0!
0'
#413950000000
1!
b111 %
1'
b111 +
#413960000000
0!
0'
#413970000000
1!
0$
b1000 %
1'
0*
b1000 +
#413980000000
0!
0'
#413990000000
1!
b1001 %
1'
b1001 +
#414000000000
0!
0'
#414010000000
1!
b0 %
1'
b0 +
#414020000000
0!
0'
#414030000000
1!
1$
b1 %
1'
1*
b1 +
#414040000000
0!
0'
#414050000000
1!
b10 %
1'
b10 +
#414060000000
0!
0'
#414070000000
1!
b11 %
1'
b11 +
#414080000000
0!
0'
#414090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#414100000000
0!
0'
#414110000000
1!
b101 %
1'
b101 +
#414120000000
0!
0'
#414130000000
1!
0$
b110 %
1'
0*
b110 +
#414140000000
0!
0'
#414150000000
1!
b111 %
1'
b111 +
#414160000000
0!
0'
#414170000000
1!
b1000 %
1'
b1000 +
#414180000000
0!
0'
#414190000000
1!
b1001 %
1'
b1001 +
#414200000000
0!
0'
#414210000000
1!
b0 %
1'
b0 +
#414220000000
0!
0'
#414230000000
1!
1$
b1 %
1'
1*
b1 +
#414240000000
0!
0'
#414250000000
1!
b10 %
1'
b10 +
#414260000000
0!
0'
#414270000000
1!
b11 %
1'
b11 +
#414280000000
0!
0'
#414290000000
1!
b100 %
1'
b100 +
#414300000000
1"
1(
#414310000000
0!
0"
b100 &
0'
0(
b100 ,
#414320000000
1!
b101 %
1'
b101 +
#414330000000
0!
0'
#414340000000
1!
b110 %
1'
b110 +
#414350000000
0!
0'
#414360000000
1!
b111 %
1'
b111 +
#414370000000
0!
0'
#414380000000
1!
0$
b1000 %
1'
0*
b1000 +
#414390000000
0!
0'
#414400000000
1!
b1001 %
1'
b1001 +
#414410000000
0!
0'
#414420000000
1!
b0 %
1'
b0 +
#414430000000
0!
0'
#414440000000
1!
1$
b1 %
1'
1*
b1 +
#414450000000
0!
0'
#414460000000
1!
b10 %
1'
b10 +
#414470000000
0!
0'
#414480000000
1!
b11 %
1'
b11 +
#414490000000
0!
0'
#414500000000
1!
b100 %
1'
b100 +
#414510000000
0!
0'
#414520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#414530000000
0!
0'
#414540000000
1!
0$
b110 %
1'
0*
b110 +
#414550000000
0!
0'
#414560000000
1!
b111 %
1'
b111 +
#414570000000
0!
0'
#414580000000
1!
b1000 %
1'
b1000 +
#414590000000
0!
0'
#414600000000
1!
b1001 %
1'
b1001 +
#414610000000
0!
0'
#414620000000
1!
b0 %
1'
b0 +
#414630000000
0!
0'
#414640000000
1!
1$
b1 %
1'
1*
b1 +
#414650000000
0!
0'
#414660000000
1!
b10 %
1'
b10 +
#414670000000
0!
0'
#414680000000
1!
b11 %
1'
b11 +
#414690000000
0!
0'
#414700000000
1!
b100 %
1'
b100 +
#414710000000
0!
0'
#414720000000
1!
b101 %
1'
b101 +
#414730000000
1"
1(
#414740000000
0!
0"
b100 &
0'
0(
b100 ,
#414750000000
1!
b110 %
1'
b110 +
#414760000000
0!
0'
#414770000000
1!
b111 %
1'
b111 +
#414780000000
0!
0'
#414790000000
1!
0$
b1000 %
1'
0*
b1000 +
#414800000000
0!
0'
#414810000000
1!
b1001 %
1'
b1001 +
#414820000000
0!
0'
#414830000000
1!
b0 %
1'
b0 +
#414840000000
0!
0'
#414850000000
1!
1$
b1 %
1'
1*
b1 +
#414860000000
0!
0'
#414870000000
1!
b10 %
1'
b10 +
#414880000000
0!
0'
#414890000000
1!
b11 %
1'
b11 +
#414900000000
0!
0'
#414910000000
1!
b100 %
1'
b100 +
#414920000000
0!
0'
#414930000000
1!
b101 %
1'
b101 +
#414940000000
0!
0'
#414950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#414960000000
0!
0'
#414970000000
1!
b111 %
1'
b111 +
#414980000000
0!
0'
#414990000000
1!
b1000 %
1'
b1000 +
#415000000000
0!
0'
#415010000000
1!
b1001 %
1'
b1001 +
#415020000000
0!
0'
#415030000000
1!
b0 %
1'
b0 +
#415040000000
0!
0'
#415050000000
1!
1$
b1 %
1'
1*
b1 +
#415060000000
0!
0'
#415070000000
1!
b10 %
1'
b10 +
#415080000000
0!
0'
#415090000000
1!
b11 %
1'
b11 +
#415100000000
0!
0'
#415110000000
1!
b100 %
1'
b100 +
#415120000000
0!
0'
#415130000000
1!
b101 %
1'
b101 +
#415140000000
0!
0'
#415150000000
1!
0$
b110 %
1'
0*
b110 +
#415160000000
1"
1(
#415170000000
0!
0"
b100 &
0'
0(
b100 ,
#415180000000
1!
1$
b111 %
1'
1*
b111 +
#415190000000
0!
0'
#415200000000
1!
0$
b1000 %
1'
0*
b1000 +
#415210000000
0!
0'
#415220000000
1!
b1001 %
1'
b1001 +
#415230000000
0!
0'
#415240000000
1!
b0 %
1'
b0 +
#415250000000
0!
0'
#415260000000
1!
1$
b1 %
1'
1*
b1 +
#415270000000
0!
0'
#415280000000
1!
b10 %
1'
b10 +
#415290000000
0!
0'
#415300000000
1!
b11 %
1'
b11 +
#415310000000
0!
0'
#415320000000
1!
b100 %
1'
b100 +
#415330000000
0!
0'
#415340000000
1!
b101 %
1'
b101 +
#415350000000
0!
0'
#415360000000
1!
b110 %
1'
b110 +
#415370000000
0!
0'
#415380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#415390000000
0!
0'
#415400000000
1!
b1000 %
1'
b1000 +
#415410000000
0!
0'
#415420000000
1!
b1001 %
1'
b1001 +
#415430000000
0!
0'
#415440000000
1!
b0 %
1'
b0 +
#415450000000
0!
0'
#415460000000
1!
1$
b1 %
1'
1*
b1 +
#415470000000
0!
0'
#415480000000
1!
b10 %
1'
b10 +
#415490000000
0!
0'
#415500000000
1!
b11 %
1'
b11 +
#415510000000
0!
0'
#415520000000
1!
b100 %
1'
b100 +
#415530000000
0!
0'
#415540000000
1!
b101 %
1'
b101 +
#415550000000
0!
0'
#415560000000
1!
0$
b110 %
1'
0*
b110 +
#415570000000
0!
0'
#415580000000
1!
b111 %
1'
b111 +
#415590000000
1"
1(
#415600000000
0!
0"
b100 &
0'
0(
b100 ,
#415610000000
1!
b1000 %
1'
b1000 +
#415620000000
0!
0'
#415630000000
1!
b1001 %
1'
b1001 +
#415640000000
0!
0'
#415650000000
1!
b0 %
1'
b0 +
#415660000000
0!
0'
#415670000000
1!
1$
b1 %
1'
1*
b1 +
#415680000000
0!
0'
#415690000000
1!
b10 %
1'
b10 +
#415700000000
0!
0'
#415710000000
1!
b11 %
1'
b11 +
#415720000000
0!
0'
#415730000000
1!
b100 %
1'
b100 +
#415740000000
0!
0'
#415750000000
1!
b101 %
1'
b101 +
#415760000000
0!
0'
#415770000000
1!
b110 %
1'
b110 +
#415780000000
0!
0'
#415790000000
1!
b111 %
1'
b111 +
#415800000000
0!
0'
#415810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#415820000000
0!
0'
#415830000000
1!
b1001 %
1'
b1001 +
#415840000000
0!
0'
#415850000000
1!
b0 %
1'
b0 +
#415860000000
0!
0'
#415870000000
1!
1$
b1 %
1'
1*
b1 +
#415880000000
0!
0'
#415890000000
1!
b10 %
1'
b10 +
#415900000000
0!
0'
#415910000000
1!
b11 %
1'
b11 +
#415920000000
0!
0'
#415930000000
1!
b100 %
1'
b100 +
#415940000000
0!
0'
#415950000000
1!
b101 %
1'
b101 +
#415960000000
0!
0'
#415970000000
1!
0$
b110 %
1'
0*
b110 +
#415980000000
0!
0'
#415990000000
1!
b111 %
1'
b111 +
#416000000000
0!
0'
#416010000000
1!
b1000 %
1'
b1000 +
#416020000000
1"
1(
#416030000000
0!
0"
b100 &
0'
0(
b100 ,
#416040000000
1!
b1001 %
1'
b1001 +
#416050000000
0!
0'
#416060000000
1!
b0 %
1'
b0 +
#416070000000
0!
0'
#416080000000
1!
1$
b1 %
1'
1*
b1 +
#416090000000
0!
0'
#416100000000
1!
b10 %
1'
b10 +
#416110000000
0!
0'
#416120000000
1!
b11 %
1'
b11 +
#416130000000
0!
0'
#416140000000
1!
b100 %
1'
b100 +
#416150000000
0!
0'
#416160000000
1!
b101 %
1'
b101 +
#416170000000
0!
0'
#416180000000
1!
b110 %
1'
b110 +
#416190000000
0!
0'
#416200000000
1!
b111 %
1'
b111 +
#416210000000
0!
0'
#416220000000
1!
0$
b1000 %
1'
0*
b1000 +
#416230000000
0!
0'
#416240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#416250000000
0!
0'
#416260000000
1!
b0 %
1'
b0 +
#416270000000
0!
0'
#416280000000
1!
1$
b1 %
1'
1*
b1 +
#416290000000
0!
0'
#416300000000
1!
b10 %
1'
b10 +
#416310000000
0!
0'
#416320000000
1!
b11 %
1'
b11 +
#416330000000
0!
0'
#416340000000
1!
b100 %
1'
b100 +
#416350000000
0!
0'
#416360000000
1!
b101 %
1'
b101 +
#416370000000
0!
0'
#416380000000
1!
0$
b110 %
1'
0*
b110 +
#416390000000
0!
0'
#416400000000
1!
b111 %
1'
b111 +
#416410000000
0!
0'
#416420000000
1!
b1000 %
1'
b1000 +
#416430000000
0!
0'
#416440000000
1!
b1001 %
1'
b1001 +
#416450000000
1"
1(
#416460000000
0!
0"
b100 &
0'
0(
b100 ,
#416470000000
1!
b0 %
1'
b0 +
#416480000000
0!
0'
#416490000000
1!
1$
b1 %
1'
1*
b1 +
#416500000000
0!
0'
#416510000000
1!
b10 %
1'
b10 +
#416520000000
0!
0'
#416530000000
1!
b11 %
1'
b11 +
#416540000000
0!
0'
#416550000000
1!
b100 %
1'
b100 +
#416560000000
0!
0'
#416570000000
1!
b101 %
1'
b101 +
#416580000000
0!
0'
#416590000000
1!
b110 %
1'
b110 +
#416600000000
0!
0'
#416610000000
1!
b111 %
1'
b111 +
#416620000000
0!
0'
#416630000000
1!
0$
b1000 %
1'
0*
b1000 +
#416640000000
0!
0'
#416650000000
1!
b1001 %
1'
b1001 +
#416660000000
0!
0'
#416670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#416680000000
0!
0'
#416690000000
1!
1$
b1 %
1'
1*
b1 +
#416700000000
0!
0'
#416710000000
1!
b10 %
1'
b10 +
#416720000000
0!
0'
#416730000000
1!
b11 %
1'
b11 +
#416740000000
0!
0'
#416750000000
1!
b100 %
1'
b100 +
#416760000000
0!
0'
#416770000000
1!
b101 %
1'
b101 +
#416780000000
0!
0'
#416790000000
1!
0$
b110 %
1'
0*
b110 +
#416800000000
0!
0'
#416810000000
1!
b111 %
1'
b111 +
#416820000000
0!
0'
#416830000000
1!
b1000 %
1'
b1000 +
#416840000000
0!
0'
#416850000000
1!
b1001 %
1'
b1001 +
#416860000000
0!
0'
#416870000000
1!
b0 %
1'
b0 +
#416880000000
1"
1(
#416890000000
0!
0"
b100 &
0'
0(
b100 ,
#416900000000
1!
1$
b1 %
1'
1*
b1 +
#416910000000
0!
0'
#416920000000
1!
b10 %
1'
b10 +
#416930000000
0!
0'
#416940000000
1!
b11 %
1'
b11 +
#416950000000
0!
0'
#416960000000
1!
b100 %
1'
b100 +
#416970000000
0!
0'
#416980000000
1!
b101 %
1'
b101 +
#416990000000
0!
0'
#417000000000
1!
b110 %
1'
b110 +
#417010000000
0!
0'
#417020000000
1!
b111 %
1'
b111 +
#417030000000
0!
0'
#417040000000
1!
0$
b1000 %
1'
0*
b1000 +
#417050000000
0!
0'
#417060000000
1!
b1001 %
1'
b1001 +
#417070000000
0!
0'
#417080000000
1!
b0 %
1'
b0 +
#417090000000
0!
0'
#417100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#417110000000
0!
0'
#417120000000
1!
b10 %
1'
b10 +
#417130000000
0!
0'
#417140000000
1!
b11 %
1'
b11 +
#417150000000
0!
0'
#417160000000
1!
b100 %
1'
b100 +
#417170000000
0!
0'
#417180000000
1!
b101 %
1'
b101 +
#417190000000
0!
0'
#417200000000
1!
0$
b110 %
1'
0*
b110 +
#417210000000
0!
0'
#417220000000
1!
b111 %
1'
b111 +
#417230000000
0!
0'
#417240000000
1!
b1000 %
1'
b1000 +
#417250000000
0!
0'
#417260000000
1!
b1001 %
1'
b1001 +
#417270000000
0!
0'
#417280000000
1!
b0 %
1'
b0 +
#417290000000
0!
0'
#417300000000
1!
1$
b1 %
1'
1*
b1 +
#417310000000
1"
1(
#417320000000
0!
0"
b100 &
0'
0(
b100 ,
#417330000000
1!
b10 %
1'
b10 +
#417340000000
0!
0'
#417350000000
1!
b11 %
1'
b11 +
#417360000000
0!
0'
#417370000000
1!
b100 %
1'
b100 +
#417380000000
0!
0'
#417390000000
1!
b101 %
1'
b101 +
#417400000000
0!
0'
#417410000000
1!
b110 %
1'
b110 +
#417420000000
0!
0'
#417430000000
1!
b111 %
1'
b111 +
#417440000000
0!
0'
#417450000000
1!
0$
b1000 %
1'
0*
b1000 +
#417460000000
0!
0'
#417470000000
1!
b1001 %
1'
b1001 +
#417480000000
0!
0'
#417490000000
1!
b0 %
1'
b0 +
#417500000000
0!
0'
#417510000000
1!
1$
b1 %
1'
1*
b1 +
#417520000000
0!
0'
#417530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#417540000000
0!
0'
#417550000000
1!
b11 %
1'
b11 +
#417560000000
0!
0'
#417570000000
1!
b100 %
1'
b100 +
#417580000000
0!
0'
#417590000000
1!
b101 %
1'
b101 +
#417600000000
0!
0'
#417610000000
1!
0$
b110 %
1'
0*
b110 +
#417620000000
0!
0'
#417630000000
1!
b111 %
1'
b111 +
#417640000000
0!
0'
#417650000000
1!
b1000 %
1'
b1000 +
#417660000000
0!
0'
#417670000000
1!
b1001 %
1'
b1001 +
#417680000000
0!
0'
#417690000000
1!
b0 %
1'
b0 +
#417700000000
0!
0'
#417710000000
1!
1$
b1 %
1'
1*
b1 +
#417720000000
0!
0'
#417730000000
1!
b10 %
1'
b10 +
#417740000000
1"
1(
#417750000000
0!
0"
b100 &
0'
0(
b100 ,
#417760000000
1!
b11 %
1'
b11 +
#417770000000
0!
0'
#417780000000
1!
b100 %
1'
b100 +
#417790000000
0!
0'
#417800000000
1!
b101 %
1'
b101 +
#417810000000
0!
0'
#417820000000
1!
b110 %
1'
b110 +
#417830000000
0!
0'
#417840000000
1!
b111 %
1'
b111 +
#417850000000
0!
0'
#417860000000
1!
0$
b1000 %
1'
0*
b1000 +
#417870000000
0!
0'
#417880000000
1!
b1001 %
1'
b1001 +
#417890000000
0!
0'
#417900000000
1!
b0 %
1'
b0 +
#417910000000
0!
0'
#417920000000
1!
1$
b1 %
1'
1*
b1 +
#417930000000
0!
0'
#417940000000
1!
b10 %
1'
b10 +
#417950000000
0!
0'
#417960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#417970000000
0!
0'
#417980000000
1!
b100 %
1'
b100 +
#417990000000
0!
0'
#418000000000
1!
b101 %
1'
b101 +
#418010000000
0!
0'
#418020000000
1!
0$
b110 %
1'
0*
b110 +
#418030000000
0!
0'
#418040000000
1!
b111 %
1'
b111 +
#418050000000
0!
0'
#418060000000
1!
b1000 %
1'
b1000 +
#418070000000
0!
0'
#418080000000
1!
b1001 %
1'
b1001 +
#418090000000
0!
0'
#418100000000
1!
b0 %
1'
b0 +
#418110000000
0!
0'
#418120000000
1!
1$
b1 %
1'
1*
b1 +
#418130000000
0!
0'
#418140000000
1!
b10 %
1'
b10 +
#418150000000
0!
0'
#418160000000
1!
b11 %
1'
b11 +
#418170000000
1"
1(
#418180000000
0!
0"
b100 &
0'
0(
b100 ,
#418190000000
1!
b100 %
1'
b100 +
#418200000000
0!
0'
#418210000000
1!
b101 %
1'
b101 +
#418220000000
0!
0'
#418230000000
1!
b110 %
1'
b110 +
#418240000000
0!
0'
#418250000000
1!
b111 %
1'
b111 +
#418260000000
0!
0'
#418270000000
1!
0$
b1000 %
1'
0*
b1000 +
#418280000000
0!
0'
#418290000000
1!
b1001 %
1'
b1001 +
#418300000000
0!
0'
#418310000000
1!
b0 %
1'
b0 +
#418320000000
0!
0'
#418330000000
1!
1$
b1 %
1'
1*
b1 +
#418340000000
0!
0'
#418350000000
1!
b10 %
1'
b10 +
#418360000000
0!
0'
#418370000000
1!
b11 %
1'
b11 +
#418380000000
0!
0'
#418390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#418400000000
0!
0'
#418410000000
1!
b101 %
1'
b101 +
#418420000000
0!
0'
#418430000000
1!
0$
b110 %
1'
0*
b110 +
#418440000000
0!
0'
#418450000000
1!
b111 %
1'
b111 +
#418460000000
0!
0'
#418470000000
1!
b1000 %
1'
b1000 +
#418480000000
0!
0'
#418490000000
1!
b1001 %
1'
b1001 +
#418500000000
0!
0'
#418510000000
1!
b0 %
1'
b0 +
#418520000000
0!
0'
#418530000000
1!
1$
b1 %
1'
1*
b1 +
#418540000000
0!
0'
#418550000000
1!
b10 %
1'
b10 +
#418560000000
0!
0'
#418570000000
1!
b11 %
1'
b11 +
#418580000000
0!
0'
#418590000000
1!
b100 %
1'
b100 +
#418600000000
1"
1(
#418610000000
0!
0"
b100 &
0'
0(
b100 ,
#418620000000
1!
b101 %
1'
b101 +
#418630000000
0!
0'
#418640000000
1!
b110 %
1'
b110 +
#418650000000
0!
0'
#418660000000
1!
b111 %
1'
b111 +
#418670000000
0!
0'
#418680000000
1!
0$
b1000 %
1'
0*
b1000 +
#418690000000
0!
0'
#418700000000
1!
b1001 %
1'
b1001 +
#418710000000
0!
0'
#418720000000
1!
b0 %
1'
b0 +
#418730000000
0!
0'
#418740000000
1!
1$
b1 %
1'
1*
b1 +
#418750000000
0!
0'
#418760000000
1!
b10 %
1'
b10 +
#418770000000
0!
0'
#418780000000
1!
b11 %
1'
b11 +
#418790000000
0!
0'
#418800000000
1!
b100 %
1'
b100 +
#418810000000
0!
0'
#418820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#418830000000
0!
0'
#418840000000
1!
0$
b110 %
1'
0*
b110 +
#418850000000
0!
0'
#418860000000
1!
b111 %
1'
b111 +
#418870000000
0!
0'
#418880000000
1!
b1000 %
1'
b1000 +
#418890000000
0!
0'
#418900000000
1!
b1001 %
1'
b1001 +
#418910000000
0!
0'
#418920000000
1!
b0 %
1'
b0 +
#418930000000
0!
0'
#418940000000
1!
1$
b1 %
1'
1*
b1 +
#418950000000
0!
0'
#418960000000
1!
b10 %
1'
b10 +
#418970000000
0!
0'
#418980000000
1!
b11 %
1'
b11 +
#418990000000
0!
0'
#419000000000
1!
b100 %
1'
b100 +
#419010000000
0!
0'
#419020000000
1!
b101 %
1'
b101 +
#419030000000
1"
1(
#419040000000
0!
0"
b100 &
0'
0(
b100 ,
#419050000000
1!
b110 %
1'
b110 +
#419060000000
0!
0'
#419070000000
1!
b111 %
1'
b111 +
#419080000000
0!
0'
#419090000000
1!
0$
b1000 %
1'
0*
b1000 +
#419100000000
0!
0'
#419110000000
1!
b1001 %
1'
b1001 +
#419120000000
0!
0'
#419130000000
1!
b0 %
1'
b0 +
#419140000000
0!
0'
#419150000000
1!
1$
b1 %
1'
1*
b1 +
#419160000000
0!
0'
#419170000000
1!
b10 %
1'
b10 +
#419180000000
0!
0'
#419190000000
1!
b11 %
1'
b11 +
#419200000000
0!
0'
#419210000000
1!
b100 %
1'
b100 +
#419220000000
0!
0'
#419230000000
1!
b101 %
1'
b101 +
#419240000000
0!
0'
#419250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#419260000000
0!
0'
#419270000000
1!
b111 %
1'
b111 +
#419280000000
0!
0'
#419290000000
1!
b1000 %
1'
b1000 +
#419300000000
0!
0'
#419310000000
1!
b1001 %
1'
b1001 +
#419320000000
0!
0'
#419330000000
1!
b0 %
1'
b0 +
#419340000000
0!
0'
#419350000000
1!
1$
b1 %
1'
1*
b1 +
#419360000000
0!
0'
#419370000000
1!
b10 %
1'
b10 +
#419380000000
0!
0'
#419390000000
1!
b11 %
1'
b11 +
#419400000000
0!
0'
#419410000000
1!
b100 %
1'
b100 +
#419420000000
0!
0'
#419430000000
1!
b101 %
1'
b101 +
#419440000000
0!
0'
#419450000000
1!
0$
b110 %
1'
0*
b110 +
#419460000000
1"
1(
#419470000000
0!
0"
b100 &
0'
0(
b100 ,
#419480000000
1!
1$
b111 %
1'
1*
b111 +
#419490000000
0!
0'
#419500000000
1!
0$
b1000 %
1'
0*
b1000 +
#419510000000
0!
0'
#419520000000
1!
b1001 %
1'
b1001 +
#419530000000
0!
0'
#419540000000
1!
b0 %
1'
b0 +
#419550000000
0!
0'
#419560000000
1!
1$
b1 %
1'
1*
b1 +
#419570000000
0!
0'
#419580000000
1!
b10 %
1'
b10 +
#419590000000
0!
0'
#419600000000
1!
b11 %
1'
b11 +
#419610000000
0!
0'
#419620000000
1!
b100 %
1'
b100 +
#419630000000
0!
0'
#419640000000
1!
b101 %
1'
b101 +
#419650000000
0!
0'
#419660000000
1!
b110 %
1'
b110 +
#419670000000
0!
0'
#419680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#419690000000
0!
0'
#419700000000
1!
b1000 %
1'
b1000 +
#419710000000
0!
0'
#419720000000
1!
b1001 %
1'
b1001 +
#419730000000
0!
0'
#419740000000
1!
b0 %
1'
b0 +
#419750000000
0!
0'
#419760000000
1!
1$
b1 %
1'
1*
b1 +
#419770000000
0!
0'
#419780000000
1!
b10 %
1'
b10 +
#419790000000
0!
0'
#419800000000
1!
b11 %
1'
b11 +
#419810000000
0!
0'
#419820000000
1!
b100 %
1'
b100 +
#419830000000
0!
0'
#419840000000
1!
b101 %
1'
b101 +
#419850000000
0!
0'
#419860000000
1!
0$
b110 %
1'
0*
b110 +
#419870000000
0!
0'
#419880000000
1!
b111 %
1'
b111 +
#419890000000
1"
1(
#419900000000
0!
0"
b100 &
0'
0(
b100 ,
#419910000000
1!
b1000 %
1'
b1000 +
#419920000000
0!
0'
#419930000000
1!
b1001 %
1'
b1001 +
#419940000000
0!
0'
#419950000000
1!
b0 %
1'
b0 +
#419960000000
0!
0'
#419970000000
1!
1$
b1 %
1'
1*
b1 +
#419980000000
0!
0'
#419990000000
1!
b10 %
1'
b10 +
#420000000000
0!
0'
#420010000000
1!
b11 %
1'
b11 +
#420020000000
0!
0'
#420030000000
1!
b100 %
1'
b100 +
#420040000000
0!
0'
#420050000000
1!
b101 %
1'
b101 +
#420060000000
0!
0'
#420070000000
1!
b110 %
1'
b110 +
#420080000000
0!
0'
#420090000000
1!
b111 %
1'
b111 +
#420100000000
0!
0'
#420110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#420120000000
0!
0'
#420130000000
1!
b1001 %
1'
b1001 +
#420140000000
0!
0'
#420150000000
1!
b0 %
1'
b0 +
#420160000000
0!
0'
#420170000000
1!
1$
b1 %
1'
1*
b1 +
#420180000000
0!
0'
#420190000000
1!
b10 %
1'
b10 +
#420200000000
0!
0'
#420210000000
1!
b11 %
1'
b11 +
#420220000000
0!
0'
#420230000000
1!
b100 %
1'
b100 +
#420240000000
0!
0'
#420250000000
1!
b101 %
1'
b101 +
#420260000000
0!
0'
#420270000000
1!
0$
b110 %
1'
0*
b110 +
#420280000000
0!
0'
#420290000000
1!
b111 %
1'
b111 +
#420300000000
0!
0'
#420310000000
1!
b1000 %
1'
b1000 +
#420320000000
1"
1(
#420330000000
0!
0"
b100 &
0'
0(
b100 ,
#420340000000
1!
b1001 %
1'
b1001 +
#420350000000
0!
0'
#420360000000
1!
b0 %
1'
b0 +
#420370000000
0!
0'
#420380000000
1!
1$
b1 %
1'
1*
b1 +
#420390000000
0!
0'
#420400000000
1!
b10 %
1'
b10 +
#420410000000
0!
0'
#420420000000
1!
b11 %
1'
b11 +
#420430000000
0!
0'
#420440000000
1!
b100 %
1'
b100 +
#420450000000
0!
0'
#420460000000
1!
b101 %
1'
b101 +
#420470000000
0!
0'
#420480000000
1!
b110 %
1'
b110 +
#420490000000
0!
0'
#420500000000
1!
b111 %
1'
b111 +
#420510000000
0!
0'
#420520000000
1!
0$
b1000 %
1'
0*
b1000 +
#420530000000
0!
0'
#420540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#420550000000
0!
0'
#420560000000
1!
b0 %
1'
b0 +
#420570000000
0!
0'
#420580000000
1!
1$
b1 %
1'
1*
b1 +
#420590000000
0!
0'
#420600000000
1!
b10 %
1'
b10 +
#420610000000
0!
0'
#420620000000
1!
b11 %
1'
b11 +
#420630000000
0!
0'
#420640000000
1!
b100 %
1'
b100 +
#420650000000
0!
0'
#420660000000
1!
b101 %
1'
b101 +
#420670000000
0!
0'
#420680000000
1!
0$
b110 %
1'
0*
b110 +
#420690000000
0!
0'
#420700000000
1!
b111 %
1'
b111 +
#420710000000
0!
0'
#420720000000
1!
b1000 %
1'
b1000 +
#420730000000
0!
0'
#420740000000
1!
b1001 %
1'
b1001 +
#420750000000
1"
1(
#420760000000
0!
0"
b100 &
0'
0(
b100 ,
#420770000000
1!
b0 %
1'
b0 +
#420780000000
0!
0'
#420790000000
1!
1$
b1 %
1'
1*
b1 +
#420800000000
0!
0'
#420810000000
1!
b10 %
1'
b10 +
#420820000000
0!
0'
#420830000000
1!
b11 %
1'
b11 +
#420840000000
0!
0'
#420850000000
1!
b100 %
1'
b100 +
#420860000000
0!
0'
#420870000000
1!
b101 %
1'
b101 +
#420880000000
0!
0'
#420890000000
1!
b110 %
1'
b110 +
#420900000000
0!
0'
#420910000000
1!
b111 %
1'
b111 +
#420920000000
0!
0'
#420930000000
1!
0$
b1000 %
1'
0*
b1000 +
#420940000000
0!
0'
#420950000000
1!
b1001 %
1'
b1001 +
#420960000000
0!
0'
#420970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#420980000000
0!
0'
#420990000000
1!
1$
b1 %
1'
1*
b1 +
#421000000000
0!
0'
#421010000000
1!
b10 %
1'
b10 +
#421020000000
0!
0'
#421030000000
1!
b11 %
1'
b11 +
#421040000000
0!
0'
#421050000000
1!
b100 %
1'
b100 +
#421060000000
0!
0'
#421070000000
1!
b101 %
1'
b101 +
#421080000000
0!
0'
#421090000000
1!
0$
b110 %
1'
0*
b110 +
#421100000000
0!
0'
#421110000000
1!
b111 %
1'
b111 +
#421120000000
0!
0'
#421130000000
1!
b1000 %
1'
b1000 +
#421140000000
0!
0'
#421150000000
1!
b1001 %
1'
b1001 +
#421160000000
0!
0'
#421170000000
1!
b0 %
1'
b0 +
#421180000000
1"
1(
#421190000000
0!
0"
b100 &
0'
0(
b100 ,
#421200000000
1!
1$
b1 %
1'
1*
b1 +
#421210000000
0!
0'
#421220000000
1!
b10 %
1'
b10 +
#421230000000
0!
0'
#421240000000
1!
b11 %
1'
b11 +
#421250000000
0!
0'
#421260000000
1!
b100 %
1'
b100 +
#421270000000
0!
0'
#421280000000
1!
b101 %
1'
b101 +
#421290000000
0!
0'
#421300000000
1!
b110 %
1'
b110 +
#421310000000
0!
0'
#421320000000
1!
b111 %
1'
b111 +
#421330000000
0!
0'
#421340000000
1!
0$
b1000 %
1'
0*
b1000 +
#421350000000
0!
0'
#421360000000
1!
b1001 %
1'
b1001 +
#421370000000
0!
0'
#421380000000
1!
b0 %
1'
b0 +
#421390000000
0!
0'
#421400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#421410000000
0!
0'
#421420000000
1!
b10 %
1'
b10 +
#421430000000
0!
0'
#421440000000
1!
b11 %
1'
b11 +
#421450000000
0!
0'
#421460000000
1!
b100 %
1'
b100 +
#421470000000
0!
0'
#421480000000
1!
b101 %
1'
b101 +
#421490000000
0!
0'
#421500000000
1!
0$
b110 %
1'
0*
b110 +
#421510000000
0!
0'
#421520000000
1!
b111 %
1'
b111 +
#421530000000
0!
0'
#421540000000
1!
b1000 %
1'
b1000 +
#421550000000
0!
0'
#421560000000
1!
b1001 %
1'
b1001 +
#421570000000
0!
0'
#421580000000
1!
b0 %
1'
b0 +
#421590000000
0!
0'
#421600000000
1!
1$
b1 %
1'
1*
b1 +
#421610000000
1"
1(
#421620000000
0!
0"
b100 &
0'
0(
b100 ,
#421630000000
1!
b10 %
1'
b10 +
#421640000000
0!
0'
#421650000000
1!
b11 %
1'
b11 +
#421660000000
0!
0'
#421670000000
1!
b100 %
1'
b100 +
#421680000000
0!
0'
#421690000000
1!
b101 %
1'
b101 +
#421700000000
0!
0'
#421710000000
1!
b110 %
1'
b110 +
#421720000000
0!
0'
#421730000000
1!
b111 %
1'
b111 +
#421740000000
0!
0'
#421750000000
1!
0$
b1000 %
1'
0*
b1000 +
#421760000000
0!
0'
#421770000000
1!
b1001 %
1'
b1001 +
#421780000000
0!
0'
#421790000000
1!
b0 %
1'
b0 +
#421800000000
0!
0'
#421810000000
1!
1$
b1 %
1'
1*
b1 +
#421820000000
0!
0'
#421830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#421840000000
0!
0'
#421850000000
1!
b11 %
1'
b11 +
#421860000000
0!
0'
#421870000000
1!
b100 %
1'
b100 +
#421880000000
0!
0'
#421890000000
1!
b101 %
1'
b101 +
#421900000000
0!
0'
#421910000000
1!
0$
b110 %
1'
0*
b110 +
#421920000000
0!
0'
#421930000000
1!
b111 %
1'
b111 +
#421940000000
0!
0'
#421950000000
1!
b1000 %
1'
b1000 +
#421960000000
0!
0'
#421970000000
1!
b1001 %
1'
b1001 +
#421980000000
0!
0'
#421990000000
1!
b0 %
1'
b0 +
#422000000000
0!
0'
#422010000000
1!
1$
b1 %
1'
1*
b1 +
#422020000000
0!
0'
#422030000000
1!
b10 %
1'
b10 +
#422040000000
1"
1(
#422050000000
0!
0"
b100 &
0'
0(
b100 ,
#422060000000
1!
b11 %
1'
b11 +
#422070000000
0!
0'
#422080000000
1!
b100 %
1'
b100 +
#422090000000
0!
0'
#422100000000
1!
b101 %
1'
b101 +
#422110000000
0!
0'
#422120000000
1!
b110 %
1'
b110 +
#422130000000
0!
0'
#422140000000
1!
b111 %
1'
b111 +
#422150000000
0!
0'
#422160000000
1!
0$
b1000 %
1'
0*
b1000 +
#422170000000
0!
0'
#422180000000
1!
b1001 %
1'
b1001 +
#422190000000
0!
0'
#422200000000
1!
b0 %
1'
b0 +
#422210000000
0!
0'
#422220000000
1!
1$
b1 %
1'
1*
b1 +
#422230000000
0!
0'
#422240000000
1!
b10 %
1'
b10 +
#422250000000
0!
0'
#422260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#422270000000
0!
0'
#422280000000
1!
b100 %
1'
b100 +
#422290000000
0!
0'
#422300000000
1!
b101 %
1'
b101 +
#422310000000
0!
0'
#422320000000
1!
0$
b110 %
1'
0*
b110 +
#422330000000
0!
0'
#422340000000
1!
b111 %
1'
b111 +
#422350000000
0!
0'
#422360000000
1!
b1000 %
1'
b1000 +
#422370000000
0!
0'
#422380000000
1!
b1001 %
1'
b1001 +
#422390000000
0!
0'
#422400000000
1!
b0 %
1'
b0 +
#422410000000
0!
0'
#422420000000
1!
1$
b1 %
1'
1*
b1 +
#422430000000
0!
0'
#422440000000
1!
b10 %
1'
b10 +
#422450000000
0!
0'
#422460000000
1!
b11 %
1'
b11 +
#422470000000
1"
1(
#422480000000
0!
0"
b100 &
0'
0(
b100 ,
#422490000000
1!
b100 %
1'
b100 +
#422500000000
0!
0'
#422510000000
1!
b101 %
1'
b101 +
#422520000000
0!
0'
#422530000000
1!
b110 %
1'
b110 +
#422540000000
0!
0'
#422550000000
1!
b111 %
1'
b111 +
#422560000000
0!
0'
#422570000000
1!
0$
b1000 %
1'
0*
b1000 +
#422580000000
0!
0'
#422590000000
1!
b1001 %
1'
b1001 +
#422600000000
0!
0'
#422610000000
1!
b0 %
1'
b0 +
#422620000000
0!
0'
#422630000000
1!
1$
b1 %
1'
1*
b1 +
#422640000000
0!
0'
#422650000000
1!
b10 %
1'
b10 +
#422660000000
0!
0'
#422670000000
1!
b11 %
1'
b11 +
#422680000000
0!
0'
#422690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#422700000000
0!
0'
#422710000000
1!
b101 %
1'
b101 +
#422720000000
0!
0'
#422730000000
1!
0$
b110 %
1'
0*
b110 +
#422740000000
0!
0'
#422750000000
1!
b111 %
1'
b111 +
#422760000000
0!
0'
#422770000000
1!
b1000 %
1'
b1000 +
#422780000000
0!
0'
#422790000000
1!
b1001 %
1'
b1001 +
#422800000000
0!
0'
#422810000000
1!
b0 %
1'
b0 +
#422820000000
0!
0'
#422830000000
1!
1$
b1 %
1'
1*
b1 +
#422840000000
0!
0'
#422850000000
1!
b10 %
1'
b10 +
#422860000000
0!
0'
#422870000000
1!
b11 %
1'
b11 +
#422880000000
0!
0'
#422890000000
1!
b100 %
1'
b100 +
#422900000000
1"
1(
#422910000000
0!
0"
b100 &
0'
0(
b100 ,
#422920000000
1!
b101 %
1'
b101 +
#422930000000
0!
0'
#422940000000
1!
b110 %
1'
b110 +
#422950000000
0!
0'
#422960000000
1!
b111 %
1'
b111 +
#422970000000
0!
0'
#422980000000
1!
0$
b1000 %
1'
0*
b1000 +
#422990000000
0!
0'
#423000000000
1!
b1001 %
1'
b1001 +
#423010000000
0!
0'
#423020000000
1!
b0 %
1'
b0 +
#423030000000
0!
0'
#423040000000
1!
1$
b1 %
1'
1*
b1 +
#423050000000
0!
0'
#423060000000
1!
b10 %
1'
b10 +
#423070000000
0!
0'
#423080000000
1!
b11 %
1'
b11 +
#423090000000
0!
0'
#423100000000
1!
b100 %
1'
b100 +
#423110000000
0!
0'
#423120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#423130000000
0!
0'
#423140000000
1!
0$
b110 %
1'
0*
b110 +
#423150000000
0!
0'
#423160000000
1!
b111 %
1'
b111 +
#423170000000
0!
0'
#423180000000
1!
b1000 %
1'
b1000 +
#423190000000
0!
0'
#423200000000
1!
b1001 %
1'
b1001 +
#423210000000
0!
0'
#423220000000
1!
b0 %
1'
b0 +
#423230000000
0!
0'
#423240000000
1!
1$
b1 %
1'
1*
b1 +
#423250000000
0!
0'
#423260000000
1!
b10 %
1'
b10 +
#423270000000
0!
0'
#423280000000
1!
b11 %
1'
b11 +
#423290000000
0!
0'
#423300000000
1!
b100 %
1'
b100 +
#423310000000
0!
0'
#423320000000
1!
b101 %
1'
b101 +
#423330000000
1"
1(
#423340000000
0!
0"
b100 &
0'
0(
b100 ,
#423350000000
1!
b110 %
1'
b110 +
#423360000000
0!
0'
#423370000000
1!
b111 %
1'
b111 +
#423380000000
0!
0'
#423390000000
1!
0$
b1000 %
1'
0*
b1000 +
#423400000000
0!
0'
#423410000000
1!
b1001 %
1'
b1001 +
#423420000000
0!
0'
#423430000000
1!
b0 %
1'
b0 +
#423440000000
0!
0'
#423450000000
1!
1$
b1 %
1'
1*
b1 +
#423460000000
0!
0'
#423470000000
1!
b10 %
1'
b10 +
#423480000000
0!
0'
#423490000000
1!
b11 %
1'
b11 +
#423500000000
0!
0'
#423510000000
1!
b100 %
1'
b100 +
#423520000000
0!
0'
#423530000000
1!
b101 %
1'
b101 +
#423540000000
0!
0'
#423550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#423560000000
0!
0'
#423570000000
1!
b111 %
1'
b111 +
#423580000000
0!
0'
#423590000000
1!
b1000 %
1'
b1000 +
#423600000000
0!
0'
#423610000000
1!
b1001 %
1'
b1001 +
#423620000000
0!
0'
#423630000000
1!
b0 %
1'
b0 +
#423640000000
0!
0'
#423650000000
1!
1$
b1 %
1'
1*
b1 +
#423660000000
0!
0'
#423670000000
1!
b10 %
1'
b10 +
#423680000000
0!
0'
#423690000000
1!
b11 %
1'
b11 +
#423700000000
0!
0'
#423710000000
1!
b100 %
1'
b100 +
#423720000000
0!
0'
#423730000000
1!
b101 %
1'
b101 +
#423740000000
0!
0'
#423750000000
1!
0$
b110 %
1'
0*
b110 +
#423760000000
1"
1(
#423770000000
0!
0"
b100 &
0'
0(
b100 ,
#423780000000
1!
1$
b111 %
1'
1*
b111 +
#423790000000
0!
0'
#423800000000
1!
0$
b1000 %
1'
0*
b1000 +
#423810000000
0!
0'
#423820000000
1!
b1001 %
1'
b1001 +
#423830000000
0!
0'
#423840000000
1!
b0 %
1'
b0 +
#423850000000
0!
0'
#423860000000
1!
1$
b1 %
1'
1*
b1 +
#423870000000
0!
0'
#423880000000
1!
b10 %
1'
b10 +
#423890000000
0!
0'
#423900000000
1!
b11 %
1'
b11 +
#423910000000
0!
0'
#423920000000
1!
b100 %
1'
b100 +
#423930000000
0!
0'
#423940000000
1!
b101 %
1'
b101 +
#423950000000
0!
0'
#423960000000
1!
b110 %
1'
b110 +
#423970000000
0!
0'
#423980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#423990000000
0!
0'
#424000000000
1!
b1000 %
1'
b1000 +
#424010000000
0!
0'
#424020000000
1!
b1001 %
1'
b1001 +
#424030000000
0!
0'
#424040000000
1!
b0 %
1'
b0 +
#424050000000
0!
0'
#424060000000
1!
1$
b1 %
1'
1*
b1 +
#424070000000
0!
0'
#424080000000
1!
b10 %
1'
b10 +
#424090000000
0!
0'
#424100000000
1!
b11 %
1'
b11 +
#424110000000
0!
0'
#424120000000
1!
b100 %
1'
b100 +
#424130000000
0!
0'
#424140000000
1!
b101 %
1'
b101 +
#424150000000
0!
0'
#424160000000
1!
0$
b110 %
1'
0*
b110 +
#424170000000
0!
0'
#424180000000
1!
b111 %
1'
b111 +
#424190000000
1"
1(
#424200000000
0!
0"
b100 &
0'
0(
b100 ,
#424210000000
1!
b1000 %
1'
b1000 +
#424220000000
0!
0'
#424230000000
1!
b1001 %
1'
b1001 +
#424240000000
0!
0'
#424250000000
1!
b0 %
1'
b0 +
#424260000000
0!
0'
#424270000000
1!
1$
b1 %
1'
1*
b1 +
#424280000000
0!
0'
#424290000000
1!
b10 %
1'
b10 +
#424300000000
0!
0'
#424310000000
1!
b11 %
1'
b11 +
#424320000000
0!
0'
#424330000000
1!
b100 %
1'
b100 +
#424340000000
0!
0'
#424350000000
1!
b101 %
1'
b101 +
#424360000000
0!
0'
#424370000000
1!
b110 %
1'
b110 +
#424380000000
0!
0'
#424390000000
1!
b111 %
1'
b111 +
#424400000000
0!
0'
#424410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#424420000000
0!
0'
#424430000000
1!
b1001 %
1'
b1001 +
#424440000000
0!
0'
#424450000000
1!
b0 %
1'
b0 +
#424460000000
0!
0'
#424470000000
1!
1$
b1 %
1'
1*
b1 +
#424480000000
0!
0'
#424490000000
1!
b10 %
1'
b10 +
#424500000000
0!
0'
#424510000000
1!
b11 %
1'
b11 +
#424520000000
0!
0'
#424530000000
1!
b100 %
1'
b100 +
#424540000000
0!
0'
#424550000000
1!
b101 %
1'
b101 +
#424560000000
0!
0'
#424570000000
1!
0$
b110 %
1'
0*
b110 +
#424580000000
0!
0'
#424590000000
1!
b111 %
1'
b111 +
#424600000000
0!
0'
#424610000000
1!
b1000 %
1'
b1000 +
#424620000000
1"
1(
#424630000000
0!
0"
b100 &
0'
0(
b100 ,
#424640000000
1!
b1001 %
1'
b1001 +
#424650000000
0!
0'
#424660000000
1!
b0 %
1'
b0 +
#424670000000
0!
0'
#424680000000
1!
1$
b1 %
1'
1*
b1 +
#424690000000
0!
0'
#424700000000
1!
b10 %
1'
b10 +
#424710000000
0!
0'
#424720000000
1!
b11 %
1'
b11 +
#424730000000
0!
0'
#424740000000
1!
b100 %
1'
b100 +
#424750000000
0!
0'
#424760000000
1!
b101 %
1'
b101 +
#424770000000
0!
0'
#424780000000
1!
b110 %
1'
b110 +
#424790000000
0!
0'
#424800000000
1!
b111 %
1'
b111 +
#424810000000
0!
0'
#424820000000
1!
0$
b1000 %
1'
0*
b1000 +
#424830000000
0!
0'
#424840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#424850000000
0!
0'
#424860000000
1!
b0 %
1'
b0 +
#424870000000
0!
0'
#424880000000
1!
1$
b1 %
1'
1*
b1 +
#424890000000
0!
0'
#424900000000
1!
b10 %
1'
b10 +
#424910000000
0!
0'
#424920000000
1!
b11 %
1'
b11 +
#424930000000
0!
0'
#424940000000
1!
b100 %
1'
b100 +
#424950000000
0!
0'
#424960000000
1!
b101 %
1'
b101 +
#424970000000
0!
0'
#424980000000
1!
0$
b110 %
1'
0*
b110 +
#424990000000
0!
0'
#425000000000
1!
b111 %
1'
b111 +
#425010000000
0!
0'
#425020000000
1!
b1000 %
1'
b1000 +
#425030000000
0!
0'
#425040000000
1!
b1001 %
1'
b1001 +
#425050000000
1"
1(
#425060000000
0!
0"
b100 &
0'
0(
b100 ,
#425070000000
1!
b0 %
1'
b0 +
#425080000000
0!
0'
#425090000000
1!
1$
b1 %
1'
1*
b1 +
#425100000000
0!
0'
#425110000000
1!
b10 %
1'
b10 +
#425120000000
0!
0'
#425130000000
1!
b11 %
1'
b11 +
#425140000000
0!
0'
#425150000000
1!
b100 %
1'
b100 +
#425160000000
0!
0'
#425170000000
1!
b101 %
1'
b101 +
#425180000000
0!
0'
#425190000000
1!
b110 %
1'
b110 +
#425200000000
0!
0'
#425210000000
1!
b111 %
1'
b111 +
#425220000000
0!
0'
#425230000000
1!
0$
b1000 %
1'
0*
b1000 +
#425240000000
0!
0'
#425250000000
1!
b1001 %
1'
b1001 +
#425260000000
0!
0'
#425270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#425280000000
0!
0'
#425290000000
1!
1$
b1 %
1'
1*
b1 +
#425300000000
0!
0'
#425310000000
1!
b10 %
1'
b10 +
#425320000000
0!
0'
#425330000000
1!
b11 %
1'
b11 +
#425340000000
0!
0'
#425350000000
1!
b100 %
1'
b100 +
#425360000000
0!
0'
#425370000000
1!
b101 %
1'
b101 +
#425380000000
0!
0'
#425390000000
1!
0$
b110 %
1'
0*
b110 +
#425400000000
0!
0'
#425410000000
1!
b111 %
1'
b111 +
#425420000000
0!
0'
#425430000000
1!
b1000 %
1'
b1000 +
#425440000000
0!
0'
#425450000000
1!
b1001 %
1'
b1001 +
#425460000000
0!
0'
#425470000000
1!
b0 %
1'
b0 +
#425480000000
1"
1(
#425490000000
0!
0"
b100 &
0'
0(
b100 ,
#425500000000
1!
1$
b1 %
1'
1*
b1 +
#425510000000
0!
0'
#425520000000
1!
b10 %
1'
b10 +
#425530000000
0!
0'
#425540000000
1!
b11 %
1'
b11 +
#425550000000
0!
0'
#425560000000
1!
b100 %
1'
b100 +
#425570000000
0!
0'
#425580000000
1!
b101 %
1'
b101 +
#425590000000
0!
0'
#425600000000
1!
b110 %
1'
b110 +
#425610000000
0!
0'
#425620000000
1!
b111 %
1'
b111 +
#425630000000
0!
0'
#425640000000
1!
0$
b1000 %
1'
0*
b1000 +
#425650000000
0!
0'
#425660000000
1!
b1001 %
1'
b1001 +
#425670000000
0!
0'
#425680000000
1!
b0 %
1'
b0 +
#425690000000
0!
0'
#425700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#425710000000
0!
0'
#425720000000
1!
b10 %
1'
b10 +
#425730000000
0!
0'
#425740000000
1!
b11 %
1'
b11 +
#425750000000
0!
0'
#425760000000
1!
b100 %
1'
b100 +
#425770000000
0!
0'
#425780000000
1!
b101 %
1'
b101 +
#425790000000
0!
0'
#425800000000
1!
0$
b110 %
1'
0*
b110 +
#425810000000
0!
0'
#425820000000
1!
b111 %
1'
b111 +
#425830000000
0!
0'
#425840000000
1!
b1000 %
1'
b1000 +
#425850000000
0!
0'
#425860000000
1!
b1001 %
1'
b1001 +
#425870000000
0!
0'
#425880000000
1!
b0 %
1'
b0 +
#425890000000
0!
0'
#425900000000
1!
1$
b1 %
1'
1*
b1 +
#425910000000
1"
1(
#425920000000
0!
0"
b100 &
0'
0(
b100 ,
#425930000000
1!
b10 %
1'
b10 +
#425940000000
0!
0'
#425950000000
1!
b11 %
1'
b11 +
#425960000000
0!
0'
#425970000000
1!
b100 %
1'
b100 +
#425980000000
0!
0'
#425990000000
1!
b101 %
1'
b101 +
#426000000000
0!
0'
#426010000000
1!
b110 %
1'
b110 +
#426020000000
0!
0'
#426030000000
1!
b111 %
1'
b111 +
#426040000000
0!
0'
#426050000000
1!
0$
b1000 %
1'
0*
b1000 +
#426060000000
0!
0'
#426070000000
1!
b1001 %
1'
b1001 +
#426080000000
0!
0'
#426090000000
1!
b0 %
1'
b0 +
#426100000000
0!
0'
#426110000000
1!
1$
b1 %
1'
1*
b1 +
#426120000000
0!
0'
#426130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#426140000000
0!
0'
#426150000000
1!
b11 %
1'
b11 +
#426160000000
0!
0'
#426170000000
1!
b100 %
1'
b100 +
#426180000000
0!
0'
#426190000000
1!
b101 %
1'
b101 +
#426200000000
0!
0'
#426210000000
1!
0$
b110 %
1'
0*
b110 +
#426220000000
0!
0'
#426230000000
1!
b111 %
1'
b111 +
#426240000000
0!
0'
#426250000000
1!
b1000 %
1'
b1000 +
#426260000000
0!
0'
#426270000000
1!
b1001 %
1'
b1001 +
#426280000000
0!
0'
#426290000000
1!
b0 %
1'
b0 +
#426300000000
0!
0'
#426310000000
1!
1$
b1 %
1'
1*
b1 +
#426320000000
0!
0'
#426330000000
1!
b10 %
1'
b10 +
#426340000000
1"
1(
#426350000000
0!
0"
b100 &
0'
0(
b100 ,
#426360000000
1!
b11 %
1'
b11 +
#426370000000
0!
0'
#426380000000
1!
b100 %
1'
b100 +
#426390000000
0!
0'
#426400000000
1!
b101 %
1'
b101 +
#426410000000
0!
0'
#426420000000
1!
b110 %
1'
b110 +
#426430000000
0!
0'
#426440000000
1!
b111 %
1'
b111 +
#426450000000
0!
0'
#426460000000
1!
0$
b1000 %
1'
0*
b1000 +
#426470000000
0!
0'
#426480000000
1!
b1001 %
1'
b1001 +
#426490000000
0!
0'
#426500000000
1!
b0 %
1'
b0 +
#426510000000
0!
0'
#426520000000
1!
1$
b1 %
1'
1*
b1 +
#426530000000
0!
0'
#426540000000
1!
b10 %
1'
b10 +
#426550000000
0!
0'
#426560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#426570000000
0!
0'
#426580000000
1!
b100 %
1'
b100 +
#426590000000
0!
0'
#426600000000
1!
b101 %
1'
b101 +
#426610000000
0!
0'
#426620000000
1!
0$
b110 %
1'
0*
b110 +
#426630000000
0!
0'
#426640000000
1!
b111 %
1'
b111 +
#426650000000
0!
0'
#426660000000
1!
b1000 %
1'
b1000 +
#426670000000
0!
0'
#426680000000
1!
b1001 %
1'
b1001 +
#426690000000
0!
0'
#426700000000
1!
b0 %
1'
b0 +
#426710000000
0!
0'
#426720000000
1!
1$
b1 %
1'
1*
b1 +
#426730000000
0!
0'
#426740000000
1!
b10 %
1'
b10 +
#426750000000
0!
0'
#426760000000
1!
b11 %
1'
b11 +
#426770000000
1"
1(
#426780000000
0!
0"
b100 &
0'
0(
b100 ,
#426790000000
1!
b100 %
1'
b100 +
#426800000000
0!
0'
#426810000000
1!
b101 %
1'
b101 +
#426820000000
0!
0'
#426830000000
1!
b110 %
1'
b110 +
#426840000000
0!
0'
#426850000000
1!
b111 %
1'
b111 +
#426860000000
0!
0'
#426870000000
1!
0$
b1000 %
1'
0*
b1000 +
#426880000000
0!
0'
#426890000000
1!
b1001 %
1'
b1001 +
#426900000000
0!
0'
#426910000000
1!
b0 %
1'
b0 +
#426920000000
0!
0'
#426930000000
1!
1$
b1 %
1'
1*
b1 +
#426940000000
0!
0'
#426950000000
1!
b10 %
1'
b10 +
#426960000000
0!
0'
#426970000000
1!
b11 %
1'
b11 +
#426980000000
0!
0'
#426990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#427000000000
0!
0'
#427010000000
1!
b101 %
1'
b101 +
#427020000000
0!
0'
#427030000000
1!
0$
b110 %
1'
0*
b110 +
#427040000000
0!
0'
#427050000000
1!
b111 %
1'
b111 +
#427060000000
0!
0'
#427070000000
1!
b1000 %
1'
b1000 +
#427080000000
0!
0'
#427090000000
1!
b1001 %
1'
b1001 +
#427100000000
0!
0'
#427110000000
1!
b0 %
1'
b0 +
#427120000000
0!
0'
#427130000000
1!
1$
b1 %
1'
1*
b1 +
#427140000000
0!
0'
#427150000000
1!
b10 %
1'
b10 +
#427160000000
0!
0'
#427170000000
1!
b11 %
1'
b11 +
#427180000000
0!
0'
#427190000000
1!
b100 %
1'
b100 +
#427200000000
1"
1(
#427210000000
0!
0"
b100 &
0'
0(
b100 ,
#427220000000
1!
b101 %
1'
b101 +
#427230000000
0!
0'
#427240000000
1!
b110 %
1'
b110 +
#427250000000
0!
0'
#427260000000
1!
b111 %
1'
b111 +
#427270000000
0!
0'
#427280000000
1!
0$
b1000 %
1'
0*
b1000 +
#427290000000
0!
0'
#427300000000
1!
b1001 %
1'
b1001 +
#427310000000
0!
0'
#427320000000
1!
b0 %
1'
b0 +
#427330000000
0!
0'
#427340000000
1!
1$
b1 %
1'
1*
b1 +
#427350000000
0!
0'
#427360000000
1!
b10 %
1'
b10 +
#427370000000
0!
0'
#427380000000
1!
b11 %
1'
b11 +
#427390000000
0!
0'
#427400000000
1!
b100 %
1'
b100 +
#427410000000
0!
0'
#427420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#427430000000
0!
0'
#427440000000
1!
0$
b110 %
1'
0*
b110 +
#427450000000
0!
0'
#427460000000
1!
b111 %
1'
b111 +
#427470000000
0!
0'
#427480000000
1!
b1000 %
1'
b1000 +
#427490000000
0!
0'
#427500000000
1!
b1001 %
1'
b1001 +
#427510000000
0!
0'
#427520000000
1!
b0 %
1'
b0 +
#427530000000
0!
0'
#427540000000
1!
1$
b1 %
1'
1*
b1 +
#427550000000
0!
0'
#427560000000
1!
b10 %
1'
b10 +
#427570000000
0!
0'
#427580000000
1!
b11 %
1'
b11 +
#427590000000
0!
0'
#427600000000
1!
b100 %
1'
b100 +
#427610000000
0!
0'
#427620000000
1!
b101 %
1'
b101 +
#427630000000
1"
1(
#427640000000
0!
0"
b100 &
0'
0(
b100 ,
#427650000000
1!
b110 %
1'
b110 +
#427660000000
0!
0'
#427670000000
1!
b111 %
1'
b111 +
#427680000000
0!
0'
#427690000000
1!
0$
b1000 %
1'
0*
b1000 +
#427700000000
0!
0'
#427710000000
1!
b1001 %
1'
b1001 +
#427720000000
0!
0'
#427730000000
1!
b0 %
1'
b0 +
#427740000000
0!
0'
#427750000000
1!
1$
b1 %
1'
1*
b1 +
#427760000000
0!
0'
#427770000000
1!
b10 %
1'
b10 +
#427780000000
0!
0'
#427790000000
1!
b11 %
1'
b11 +
#427800000000
0!
0'
#427810000000
1!
b100 %
1'
b100 +
#427820000000
0!
0'
#427830000000
1!
b101 %
1'
b101 +
#427840000000
0!
0'
#427850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#427860000000
0!
0'
#427870000000
1!
b111 %
1'
b111 +
#427880000000
0!
0'
#427890000000
1!
b1000 %
1'
b1000 +
#427900000000
0!
0'
#427910000000
1!
b1001 %
1'
b1001 +
#427920000000
0!
0'
#427930000000
1!
b0 %
1'
b0 +
#427940000000
0!
0'
#427950000000
1!
1$
b1 %
1'
1*
b1 +
#427960000000
0!
0'
#427970000000
1!
b10 %
1'
b10 +
#427980000000
0!
0'
#427990000000
1!
b11 %
1'
b11 +
#428000000000
0!
0'
#428010000000
1!
b100 %
1'
b100 +
#428020000000
0!
0'
#428030000000
1!
b101 %
1'
b101 +
#428040000000
0!
0'
#428050000000
1!
0$
b110 %
1'
0*
b110 +
#428060000000
1"
1(
#428070000000
0!
0"
b100 &
0'
0(
b100 ,
#428080000000
1!
1$
b111 %
1'
1*
b111 +
#428090000000
0!
0'
#428100000000
1!
0$
b1000 %
1'
0*
b1000 +
#428110000000
0!
0'
#428120000000
1!
b1001 %
1'
b1001 +
#428130000000
0!
0'
#428140000000
1!
b0 %
1'
b0 +
#428150000000
0!
0'
#428160000000
1!
1$
b1 %
1'
1*
b1 +
#428170000000
0!
0'
#428180000000
1!
b10 %
1'
b10 +
#428190000000
0!
0'
#428200000000
1!
b11 %
1'
b11 +
#428210000000
0!
0'
#428220000000
1!
b100 %
1'
b100 +
#428230000000
0!
0'
#428240000000
1!
b101 %
1'
b101 +
#428250000000
0!
0'
#428260000000
1!
b110 %
1'
b110 +
#428270000000
0!
0'
#428280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#428290000000
0!
0'
#428300000000
1!
b1000 %
1'
b1000 +
#428310000000
0!
0'
#428320000000
1!
b1001 %
1'
b1001 +
#428330000000
0!
0'
#428340000000
1!
b0 %
1'
b0 +
#428350000000
0!
0'
#428360000000
1!
1$
b1 %
1'
1*
b1 +
#428370000000
0!
0'
#428380000000
1!
b10 %
1'
b10 +
#428390000000
0!
0'
#428400000000
1!
b11 %
1'
b11 +
#428410000000
0!
0'
#428420000000
1!
b100 %
1'
b100 +
#428430000000
0!
0'
#428440000000
1!
b101 %
1'
b101 +
#428450000000
0!
0'
#428460000000
1!
0$
b110 %
1'
0*
b110 +
#428470000000
0!
0'
#428480000000
1!
b111 %
1'
b111 +
#428490000000
1"
1(
#428500000000
0!
0"
b100 &
0'
0(
b100 ,
#428510000000
1!
b1000 %
1'
b1000 +
#428520000000
0!
0'
#428530000000
1!
b1001 %
1'
b1001 +
#428540000000
0!
0'
#428550000000
1!
b0 %
1'
b0 +
#428560000000
0!
0'
#428570000000
1!
1$
b1 %
1'
1*
b1 +
#428580000000
0!
0'
#428590000000
1!
b10 %
1'
b10 +
#428600000000
0!
0'
#428610000000
1!
b11 %
1'
b11 +
#428620000000
0!
0'
#428630000000
1!
b100 %
1'
b100 +
#428640000000
0!
0'
#428650000000
1!
b101 %
1'
b101 +
#428660000000
0!
0'
#428670000000
1!
b110 %
1'
b110 +
#428680000000
0!
0'
#428690000000
1!
b111 %
1'
b111 +
#428700000000
0!
0'
#428710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#428720000000
0!
0'
#428730000000
1!
b1001 %
1'
b1001 +
#428740000000
0!
0'
#428750000000
1!
b0 %
1'
b0 +
#428760000000
0!
0'
#428770000000
1!
1$
b1 %
1'
1*
b1 +
#428780000000
0!
0'
#428790000000
1!
b10 %
1'
b10 +
#428800000000
0!
0'
#428810000000
1!
b11 %
1'
b11 +
#428820000000
0!
0'
#428830000000
1!
b100 %
1'
b100 +
#428840000000
0!
0'
#428850000000
1!
b101 %
1'
b101 +
#428860000000
0!
0'
#428870000000
1!
0$
b110 %
1'
0*
b110 +
#428880000000
0!
0'
#428890000000
1!
b111 %
1'
b111 +
#428900000000
0!
0'
#428910000000
1!
b1000 %
1'
b1000 +
#428920000000
1"
1(
#428930000000
0!
0"
b100 &
0'
0(
b100 ,
#428940000000
1!
b1001 %
1'
b1001 +
#428950000000
0!
0'
#428960000000
1!
b0 %
1'
b0 +
#428970000000
0!
0'
#428980000000
1!
1$
b1 %
1'
1*
b1 +
#428990000000
0!
0'
#429000000000
1!
b10 %
1'
b10 +
#429010000000
0!
0'
#429020000000
1!
b11 %
1'
b11 +
#429030000000
0!
0'
#429040000000
1!
b100 %
1'
b100 +
#429050000000
0!
0'
#429060000000
1!
b101 %
1'
b101 +
#429070000000
0!
0'
#429080000000
1!
b110 %
1'
b110 +
#429090000000
0!
0'
#429100000000
1!
b111 %
1'
b111 +
#429110000000
0!
0'
#429120000000
1!
0$
b1000 %
1'
0*
b1000 +
#429130000000
0!
0'
#429140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#429150000000
0!
0'
#429160000000
1!
b0 %
1'
b0 +
#429170000000
0!
0'
#429180000000
1!
1$
b1 %
1'
1*
b1 +
#429190000000
0!
0'
#429200000000
1!
b10 %
1'
b10 +
#429210000000
0!
0'
#429220000000
1!
b11 %
1'
b11 +
#429230000000
0!
0'
#429240000000
1!
b100 %
1'
b100 +
#429250000000
0!
0'
#429260000000
1!
b101 %
1'
b101 +
#429270000000
0!
0'
#429280000000
1!
0$
b110 %
1'
0*
b110 +
#429290000000
0!
0'
#429300000000
1!
b111 %
1'
b111 +
#429310000000
0!
0'
#429320000000
1!
b1000 %
1'
b1000 +
#429330000000
0!
0'
#429340000000
1!
b1001 %
1'
b1001 +
#429350000000
1"
1(
#429360000000
0!
0"
b100 &
0'
0(
b100 ,
#429370000000
1!
b0 %
1'
b0 +
#429380000000
0!
0'
#429390000000
1!
1$
b1 %
1'
1*
b1 +
#429400000000
0!
0'
#429410000000
1!
b10 %
1'
b10 +
#429420000000
0!
0'
#429430000000
1!
b11 %
1'
b11 +
#429440000000
0!
0'
#429450000000
1!
b100 %
1'
b100 +
#429460000000
0!
0'
#429470000000
1!
b101 %
1'
b101 +
#429480000000
0!
0'
#429490000000
1!
b110 %
1'
b110 +
#429500000000
0!
0'
#429510000000
1!
b111 %
1'
b111 +
#429520000000
0!
0'
#429530000000
1!
0$
b1000 %
1'
0*
b1000 +
#429540000000
0!
0'
#429550000000
1!
b1001 %
1'
b1001 +
#429560000000
0!
0'
#429570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#429580000000
0!
0'
#429590000000
1!
1$
b1 %
1'
1*
b1 +
#429600000000
0!
0'
#429610000000
1!
b10 %
1'
b10 +
#429620000000
0!
0'
#429630000000
1!
b11 %
1'
b11 +
#429640000000
0!
0'
#429650000000
1!
b100 %
1'
b100 +
#429660000000
0!
0'
#429670000000
1!
b101 %
1'
b101 +
#429680000000
0!
0'
#429690000000
1!
0$
b110 %
1'
0*
b110 +
#429700000000
0!
0'
#429710000000
1!
b111 %
1'
b111 +
#429720000000
0!
0'
#429730000000
1!
b1000 %
1'
b1000 +
#429740000000
0!
0'
#429750000000
1!
b1001 %
1'
b1001 +
#429760000000
0!
0'
#429770000000
1!
b0 %
1'
b0 +
#429780000000
1"
1(
#429790000000
0!
0"
b100 &
0'
0(
b100 ,
#429800000000
1!
1$
b1 %
1'
1*
b1 +
#429810000000
0!
0'
#429820000000
1!
b10 %
1'
b10 +
#429830000000
0!
0'
#429840000000
1!
b11 %
1'
b11 +
#429850000000
0!
0'
#429860000000
1!
b100 %
1'
b100 +
#429870000000
0!
0'
#429880000000
1!
b101 %
1'
b101 +
#429890000000
0!
0'
#429900000000
1!
b110 %
1'
b110 +
#429910000000
0!
0'
#429920000000
1!
b111 %
1'
b111 +
#429930000000
0!
0'
#429940000000
1!
0$
b1000 %
1'
0*
b1000 +
#429950000000
0!
0'
#429960000000
1!
b1001 %
1'
b1001 +
#429970000000
0!
0'
#429980000000
1!
b0 %
1'
b0 +
#429990000000
0!
0'
#430000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#430010000000
0!
0'
#430020000000
1!
b10 %
1'
b10 +
#430030000000
0!
0'
#430040000000
1!
b11 %
1'
b11 +
#430050000000
0!
0'
#430060000000
1!
b100 %
1'
b100 +
#430070000000
0!
0'
#430080000000
1!
b101 %
1'
b101 +
#430090000000
0!
0'
#430100000000
1!
0$
b110 %
1'
0*
b110 +
#430110000000
0!
0'
#430120000000
1!
b111 %
1'
b111 +
#430130000000
0!
0'
#430140000000
1!
b1000 %
1'
b1000 +
#430150000000
0!
0'
#430160000000
1!
b1001 %
1'
b1001 +
#430170000000
0!
0'
#430180000000
1!
b0 %
1'
b0 +
#430190000000
0!
0'
#430200000000
1!
1$
b1 %
1'
1*
b1 +
#430210000000
1"
1(
#430220000000
0!
0"
b100 &
0'
0(
b100 ,
#430230000000
1!
b10 %
1'
b10 +
#430240000000
0!
0'
#430250000000
1!
b11 %
1'
b11 +
#430260000000
0!
0'
#430270000000
1!
b100 %
1'
b100 +
#430280000000
0!
0'
#430290000000
1!
b101 %
1'
b101 +
#430300000000
0!
0'
#430310000000
1!
b110 %
1'
b110 +
#430320000000
0!
0'
#430330000000
1!
b111 %
1'
b111 +
#430340000000
0!
0'
#430350000000
1!
0$
b1000 %
1'
0*
b1000 +
#430360000000
0!
0'
#430370000000
1!
b1001 %
1'
b1001 +
#430380000000
0!
0'
#430390000000
1!
b0 %
1'
b0 +
#430400000000
0!
0'
#430410000000
1!
1$
b1 %
1'
1*
b1 +
#430420000000
0!
0'
#430430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#430440000000
0!
0'
#430450000000
1!
b11 %
1'
b11 +
#430460000000
0!
0'
#430470000000
1!
b100 %
1'
b100 +
#430480000000
0!
0'
#430490000000
1!
b101 %
1'
b101 +
#430500000000
0!
0'
#430510000000
1!
0$
b110 %
1'
0*
b110 +
#430520000000
0!
0'
#430530000000
1!
b111 %
1'
b111 +
#430540000000
0!
0'
#430550000000
1!
b1000 %
1'
b1000 +
#430560000000
0!
0'
#430570000000
1!
b1001 %
1'
b1001 +
#430580000000
0!
0'
#430590000000
1!
b0 %
1'
b0 +
#430600000000
0!
0'
#430610000000
1!
1$
b1 %
1'
1*
b1 +
#430620000000
0!
0'
#430630000000
1!
b10 %
1'
b10 +
#430640000000
1"
1(
#430650000000
0!
0"
b100 &
0'
0(
b100 ,
#430660000000
1!
b11 %
1'
b11 +
#430670000000
0!
0'
#430680000000
1!
b100 %
1'
b100 +
#430690000000
0!
0'
#430700000000
1!
b101 %
1'
b101 +
#430710000000
0!
0'
#430720000000
1!
b110 %
1'
b110 +
#430730000000
0!
0'
#430740000000
1!
b111 %
1'
b111 +
#430750000000
0!
0'
#430760000000
1!
0$
b1000 %
1'
0*
b1000 +
#430770000000
0!
0'
#430780000000
1!
b1001 %
1'
b1001 +
#430790000000
0!
0'
#430800000000
1!
b0 %
1'
b0 +
#430810000000
0!
0'
#430820000000
1!
1$
b1 %
1'
1*
b1 +
#430830000000
0!
0'
#430840000000
1!
b10 %
1'
b10 +
#430850000000
0!
0'
#430860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#430870000000
0!
0'
#430880000000
1!
b100 %
1'
b100 +
#430890000000
0!
0'
#430900000000
1!
b101 %
1'
b101 +
#430910000000
0!
0'
#430920000000
1!
0$
b110 %
1'
0*
b110 +
#430930000000
0!
0'
#430940000000
1!
b111 %
1'
b111 +
#430950000000
0!
0'
#430960000000
1!
b1000 %
1'
b1000 +
#430970000000
0!
0'
#430980000000
1!
b1001 %
1'
b1001 +
#430990000000
0!
0'
#431000000000
1!
b0 %
1'
b0 +
#431010000000
0!
0'
#431020000000
1!
1$
b1 %
1'
1*
b1 +
#431030000000
0!
0'
#431040000000
1!
b10 %
1'
b10 +
#431050000000
0!
0'
#431060000000
1!
b11 %
1'
b11 +
#431070000000
1"
1(
#431080000000
0!
0"
b100 &
0'
0(
b100 ,
#431090000000
1!
b100 %
1'
b100 +
#431100000000
0!
0'
#431110000000
1!
b101 %
1'
b101 +
#431120000000
0!
0'
#431130000000
1!
b110 %
1'
b110 +
#431140000000
0!
0'
#431150000000
1!
b111 %
1'
b111 +
#431160000000
0!
0'
#431170000000
1!
0$
b1000 %
1'
0*
b1000 +
#431180000000
0!
0'
#431190000000
1!
b1001 %
1'
b1001 +
#431200000000
0!
0'
#431210000000
1!
b0 %
1'
b0 +
#431220000000
0!
0'
#431230000000
1!
1$
b1 %
1'
1*
b1 +
#431240000000
0!
0'
#431250000000
1!
b10 %
1'
b10 +
#431260000000
0!
0'
#431270000000
1!
b11 %
1'
b11 +
#431280000000
0!
0'
#431290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#431300000000
0!
0'
#431310000000
1!
b101 %
1'
b101 +
#431320000000
0!
0'
#431330000000
1!
0$
b110 %
1'
0*
b110 +
#431340000000
0!
0'
#431350000000
1!
b111 %
1'
b111 +
#431360000000
0!
0'
#431370000000
1!
b1000 %
1'
b1000 +
#431380000000
0!
0'
#431390000000
1!
b1001 %
1'
b1001 +
#431400000000
0!
0'
#431410000000
1!
b0 %
1'
b0 +
#431420000000
0!
0'
#431430000000
1!
1$
b1 %
1'
1*
b1 +
#431440000000
0!
0'
#431450000000
1!
b10 %
1'
b10 +
#431460000000
0!
0'
#431470000000
1!
b11 %
1'
b11 +
#431480000000
0!
0'
#431490000000
1!
b100 %
1'
b100 +
#431500000000
1"
1(
#431510000000
0!
0"
b100 &
0'
0(
b100 ,
#431520000000
1!
b101 %
1'
b101 +
#431530000000
0!
0'
#431540000000
1!
b110 %
1'
b110 +
#431550000000
0!
0'
#431560000000
1!
b111 %
1'
b111 +
#431570000000
0!
0'
#431580000000
1!
0$
b1000 %
1'
0*
b1000 +
#431590000000
0!
0'
#431600000000
1!
b1001 %
1'
b1001 +
#431610000000
0!
0'
#431620000000
1!
b0 %
1'
b0 +
#431630000000
0!
0'
#431640000000
1!
1$
b1 %
1'
1*
b1 +
#431650000000
0!
0'
#431660000000
1!
b10 %
1'
b10 +
#431670000000
0!
0'
#431680000000
1!
b11 %
1'
b11 +
#431690000000
0!
0'
#431700000000
1!
b100 %
1'
b100 +
#431710000000
0!
0'
#431720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#431730000000
0!
0'
#431740000000
1!
0$
b110 %
1'
0*
b110 +
#431750000000
0!
0'
#431760000000
1!
b111 %
1'
b111 +
#431770000000
0!
0'
#431780000000
1!
b1000 %
1'
b1000 +
#431790000000
0!
0'
#431800000000
1!
b1001 %
1'
b1001 +
#431810000000
0!
0'
#431820000000
1!
b0 %
1'
b0 +
#431830000000
0!
0'
#431840000000
1!
1$
b1 %
1'
1*
b1 +
#431850000000
0!
0'
#431860000000
1!
b10 %
1'
b10 +
#431870000000
0!
0'
#431880000000
1!
b11 %
1'
b11 +
#431890000000
0!
0'
#431900000000
1!
b100 %
1'
b100 +
#431910000000
0!
0'
#431920000000
1!
b101 %
1'
b101 +
#431930000000
1"
1(
#431940000000
0!
0"
b100 &
0'
0(
b100 ,
#431950000000
1!
b110 %
1'
b110 +
#431960000000
0!
0'
#431970000000
1!
b111 %
1'
b111 +
#431980000000
0!
0'
#431990000000
1!
0$
b1000 %
1'
0*
b1000 +
#432000000000
0!
0'
#432010000000
1!
b1001 %
1'
b1001 +
#432020000000
0!
0'
#432030000000
1!
b0 %
1'
b0 +
#432040000000
0!
0'
#432050000000
1!
1$
b1 %
1'
1*
b1 +
#432060000000
0!
0'
#432070000000
1!
b10 %
1'
b10 +
#432080000000
0!
0'
#432090000000
1!
b11 %
1'
b11 +
#432100000000
0!
0'
#432110000000
1!
b100 %
1'
b100 +
#432120000000
0!
0'
#432130000000
1!
b101 %
1'
b101 +
#432140000000
0!
0'
#432150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#432160000000
0!
0'
#432170000000
1!
b111 %
1'
b111 +
#432180000000
0!
0'
#432190000000
1!
b1000 %
1'
b1000 +
#432200000000
0!
0'
#432210000000
1!
b1001 %
1'
b1001 +
#432220000000
0!
0'
#432230000000
1!
b0 %
1'
b0 +
#432240000000
0!
0'
#432250000000
1!
1$
b1 %
1'
1*
b1 +
#432260000000
0!
0'
#432270000000
1!
b10 %
1'
b10 +
#432280000000
0!
0'
#432290000000
1!
b11 %
1'
b11 +
#432300000000
0!
0'
#432310000000
1!
b100 %
1'
b100 +
#432320000000
0!
0'
#432330000000
1!
b101 %
1'
b101 +
#432340000000
0!
0'
#432350000000
1!
0$
b110 %
1'
0*
b110 +
#432360000000
1"
1(
#432370000000
0!
0"
b100 &
0'
0(
b100 ,
#432380000000
1!
1$
b111 %
1'
1*
b111 +
#432390000000
0!
0'
#432400000000
1!
0$
b1000 %
1'
0*
b1000 +
#432410000000
0!
0'
#432420000000
1!
b1001 %
1'
b1001 +
#432430000000
0!
0'
#432440000000
1!
b0 %
1'
b0 +
#432450000000
0!
0'
#432460000000
1!
1$
b1 %
1'
1*
b1 +
#432470000000
0!
0'
#432480000000
1!
b10 %
1'
b10 +
#432490000000
0!
0'
#432500000000
1!
b11 %
1'
b11 +
#432510000000
0!
0'
#432520000000
1!
b100 %
1'
b100 +
#432530000000
0!
0'
#432540000000
1!
b101 %
1'
b101 +
#432550000000
0!
0'
#432560000000
1!
b110 %
1'
b110 +
#432570000000
0!
0'
#432580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#432590000000
0!
0'
#432600000000
1!
b1000 %
1'
b1000 +
#432610000000
0!
0'
#432620000000
1!
b1001 %
1'
b1001 +
#432630000000
0!
0'
#432640000000
1!
b0 %
1'
b0 +
#432650000000
0!
0'
#432660000000
1!
1$
b1 %
1'
1*
b1 +
#432670000000
0!
0'
#432680000000
1!
b10 %
1'
b10 +
#432690000000
0!
0'
#432700000000
1!
b11 %
1'
b11 +
#432710000000
0!
0'
#432720000000
1!
b100 %
1'
b100 +
#432730000000
0!
0'
#432740000000
1!
b101 %
1'
b101 +
#432750000000
0!
0'
#432760000000
1!
0$
b110 %
1'
0*
b110 +
#432770000000
0!
0'
#432780000000
1!
b111 %
1'
b111 +
#432790000000
1"
1(
#432800000000
0!
0"
b100 &
0'
0(
b100 ,
#432810000000
1!
b1000 %
1'
b1000 +
#432820000000
0!
0'
#432830000000
1!
b1001 %
1'
b1001 +
#432840000000
0!
0'
#432850000000
1!
b0 %
1'
b0 +
#432860000000
0!
0'
#432870000000
1!
1$
b1 %
1'
1*
b1 +
#432880000000
0!
0'
#432890000000
1!
b10 %
1'
b10 +
#432900000000
0!
0'
#432910000000
1!
b11 %
1'
b11 +
#432920000000
0!
0'
#432930000000
1!
b100 %
1'
b100 +
#432940000000
0!
0'
#432950000000
1!
b101 %
1'
b101 +
#432960000000
0!
0'
#432970000000
1!
b110 %
1'
b110 +
#432980000000
0!
0'
#432990000000
1!
b111 %
1'
b111 +
#433000000000
0!
0'
#433010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#433020000000
0!
0'
#433030000000
1!
b1001 %
1'
b1001 +
#433040000000
0!
0'
#433050000000
1!
b0 %
1'
b0 +
#433060000000
0!
0'
#433070000000
1!
1$
b1 %
1'
1*
b1 +
#433080000000
0!
0'
#433090000000
1!
b10 %
1'
b10 +
#433100000000
0!
0'
#433110000000
1!
b11 %
1'
b11 +
#433120000000
0!
0'
#433130000000
1!
b100 %
1'
b100 +
#433140000000
0!
0'
#433150000000
1!
b101 %
1'
b101 +
#433160000000
0!
0'
#433170000000
1!
0$
b110 %
1'
0*
b110 +
#433180000000
0!
0'
#433190000000
1!
b111 %
1'
b111 +
#433200000000
0!
0'
#433210000000
1!
b1000 %
1'
b1000 +
#433220000000
1"
1(
#433230000000
0!
0"
b100 &
0'
0(
b100 ,
#433240000000
1!
b1001 %
1'
b1001 +
#433250000000
0!
0'
#433260000000
1!
b0 %
1'
b0 +
#433270000000
0!
0'
#433280000000
1!
1$
b1 %
1'
1*
b1 +
#433290000000
0!
0'
#433300000000
1!
b10 %
1'
b10 +
#433310000000
0!
0'
#433320000000
1!
b11 %
1'
b11 +
#433330000000
0!
0'
#433340000000
1!
b100 %
1'
b100 +
#433350000000
0!
0'
#433360000000
1!
b101 %
1'
b101 +
#433370000000
0!
0'
#433380000000
1!
b110 %
1'
b110 +
#433390000000
0!
0'
#433400000000
1!
b111 %
1'
b111 +
#433410000000
0!
0'
#433420000000
1!
0$
b1000 %
1'
0*
b1000 +
#433430000000
0!
0'
#433440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#433450000000
0!
0'
#433460000000
1!
b0 %
1'
b0 +
#433470000000
0!
0'
#433480000000
1!
1$
b1 %
1'
1*
b1 +
#433490000000
0!
0'
#433500000000
1!
b10 %
1'
b10 +
#433510000000
0!
0'
#433520000000
1!
b11 %
1'
b11 +
#433530000000
0!
0'
#433540000000
1!
b100 %
1'
b100 +
#433550000000
0!
0'
#433560000000
1!
b101 %
1'
b101 +
#433570000000
0!
0'
#433580000000
1!
0$
b110 %
1'
0*
b110 +
#433590000000
0!
0'
#433600000000
1!
b111 %
1'
b111 +
#433610000000
0!
0'
#433620000000
1!
b1000 %
1'
b1000 +
#433630000000
0!
0'
#433640000000
1!
b1001 %
1'
b1001 +
#433650000000
1"
1(
#433660000000
0!
0"
b100 &
0'
0(
b100 ,
#433670000000
1!
b0 %
1'
b0 +
#433680000000
0!
0'
#433690000000
1!
1$
b1 %
1'
1*
b1 +
#433700000000
0!
0'
#433710000000
1!
b10 %
1'
b10 +
#433720000000
0!
0'
#433730000000
1!
b11 %
1'
b11 +
#433740000000
0!
0'
#433750000000
1!
b100 %
1'
b100 +
#433760000000
0!
0'
#433770000000
1!
b101 %
1'
b101 +
#433780000000
0!
0'
#433790000000
1!
b110 %
1'
b110 +
#433800000000
0!
0'
#433810000000
1!
b111 %
1'
b111 +
#433820000000
0!
0'
#433830000000
1!
0$
b1000 %
1'
0*
b1000 +
#433840000000
0!
0'
#433850000000
1!
b1001 %
1'
b1001 +
#433860000000
0!
0'
#433870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#433880000000
0!
0'
#433890000000
1!
1$
b1 %
1'
1*
b1 +
#433900000000
0!
0'
#433910000000
1!
b10 %
1'
b10 +
#433920000000
0!
0'
#433930000000
1!
b11 %
1'
b11 +
#433940000000
0!
0'
#433950000000
1!
b100 %
1'
b100 +
#433960000000
0!
0'
#433970000000
1!
b101 %
1'
b101 +
#433980000000
0!
0'
#433990000000
1!
0$
b110 %
1'
0*
b110 +
#434000000000
0!
0'
#434010000000
1!
b111 %
1'
b111 +
#434020000000
0!
0'
#434030000000
1!
b1000 %
1'
b1000 +
#434040000000
0!
0'
#434050000000
1!
b1001 %
1'
b1001 +
#434060000000
0!
0'
#434070000000
1!
b0 %
1'
b0 +
#434080000000
1"
1(
#434090000000
0!
0"
b100 &
0'
0(
b100 ,
#434100000000
1!
1$
b1 %
1'
1*
b1 +
#434110000000
0!
0'
#434120000000
1!
b10 %
1'
b10 +
#434130000000
0!
0'
#434140000000
1!
b11 %
1'
b11 +
#434150000000
0!
0'
#434160000000
1!
b100 %
1'
b100 +
#434170000000
0!
0'
#434180000000
1!
b101 %
1'
b101 +
#434190000000
0!
0'
#434200000000
1!
b110 %
1'
b110 +
#434210000000
0!
0'
#434220000000
1!
b111 %
1'
b111 +
#434230000000
0!
0'
#434240000000
1!
0$
b1000 %
1'
0*
b1000 +
#434250000000
0!
0'
#434260000000
1!
b1001 %
1'
b1001 +
#434270000000
0!
0'
#434280000000
1!
b0 %
1'
b0 +
#434290000000
0!
0'
#434300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#434310000000
0!
0'
#434320000000
1!
b10 %
1'
b10 +
#434330000000
0!
0'
#434340000000
1!
b11 %
1'
b11 +
#434350000000
0!
0'
#434360000000
1!
b100 %
1'
b100 +
#434370000000
0!
0'
#434380000000
1!
b101 %
1'
b101 +
#434390000000
0!
0'
#434400000000
1!
0$
b110 %
1'
0*
b110 +
#434410000000
0!
0'
#434420000000
1!
b111 %
1'
b111 +
#434430000000
0!
0'
#434440000000
1!
b1000 %
1'
b1000 +
#434450000000
0!
0'
#434460000000
1!
b1001 %
1'
b1001 +
#434470000000
0!
0'
#434480000000
1!
b0 %
1'
b0 +
#434490000000
0!
0'
#434500000000
1!
1$
b1 %
1'
1*
b1 +
#434510000000
1"
1(
#434520000000
0!
0"
b100 &
0'
0(
b100 ,
#434530000000
1!
b10 %
1'
b10 +
#434540000000
0!
0'
#434550000000
1!
b11 %
1'
b11 +
#434560000000
0!
0'
#434570000000
1!
b100 %
1'
b100 +
#434580000000
0!
0'
#434590000000
1!
b101 %
1'
b101 +
#434600000000
0!
0'
#434610000000
1!
b110 %
1'
b110 +
#434620000000
0!
0'
#434630000000
1!
b111 %
1'
b111 +
#434640000000
0!
0'
#434650000000
1!
0$
b1000 %
1'
0*
b1000 +
#434660000000
0!
0'
#434670000000
1!
b1001 %
1'
b1001 +
#434680000000
0!
0'
#434690000000
1!
b0 %
1'
b0 +
#434700000000
0!
0'
#434710000000
1!
1$
b1 %
1'
1*
b1 +
#434720000000
0!
0'
#434730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#434740000000
0!
0'
#434750000000
1!
b11 %
1'
b11 +
#434760000000
0!
0'
#434770000000
1!
b100 %
1'
b100 +
#434780000000
0!
0'
#434790000000
1!
b101 %
1'
b101 +
#434800000000
0!
0'
#434810000000
1!
0$
b110 %
1'
0*
b110 +
#434820000000
0!
0'
#434830000000
1!
b111 %
1'
b111 +
#434840000000
0!
0'
#434850000000
1!
b1000 %
1'
b1000 +
#434860000000
0!
0'
#434870000000
1!
b1001 %
1'
b1001 +
#434880000000
0!
0'
#434890000000
1!
b0 %
1'
b0 +
#434900000000
0!
0'
#434910000000
1!
1$
b1 %
1'
1*
b1 +
#434920000000
0!
0'
#434930000000
1!
b10 %
1'
b10 +
#434940000000
1"
1(
#434950000000
0!
0"
b100 &
0'
0(
b100 ,
#434960000000
1!
b11 %
1'
b11 +
#434970000000
0!
0'
#434980000000
1!
b100 %
1'
b100 +
#434990000000
0!
0'
#435000000000
1!
b101 %
1'
b101 +
#435010000000
0!
0'
#435020000000
1!
b110 %
1'
b110 +
#435030000000
0!
0'
#435040000000
1!
b111 %
1'
b111 +
#435050000000
0!
0'
#435060000000
1!
0$
b1000 %
1'
0*
b1000 +
#435070000000
0!
0'
#435080000000
1!
b1001 %
1'
b1001 +
#435090000000
0!
0'
#435100000000
1!
b0 %
1'
b0 +
#435110000000
0!
0'
#435120000000
1!
1$
b1 %
1'
1*
b1 +
#435130000000
0!
0'
#435140000000
1!
b10 %
1'
b10 +
#435150000000
0!
0'
#435160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#435170000000
0!
0'
#435180000000
1!
b100 %
1'
b100 +
#435190000000
0!
0'
#435200000000
1!
b101 %
1'
b101 +
#435210000000
0!
0'
#435220000000
1!
0$
b110 %
1'
0*
b110 +
#435230000000
0!
0'
#435240000000
1!
b111 %
1'
b111 +
#435250000000
0!
0'
#435260000000
1!
b1000 %
1'
b1000 +
#435270000000
0!
0'
#435280000000
1!
b1001 %
1'
b1001 +
#435290000000
0!
0'
#435300000000
1!
b0 %
1'
b0 +
#435310000000
0!
0'
#435320000000
1!
1$
b1 %
1'
1*
b1 +
#435330000000
0!
0'
#435340000000
1!
b10 %
1'
b10 +
#435350000000
0!
0'
#435360000000
1!
b11 %
1'
b11 +
#435370000000
1"
1(
#435380000000
0!
0"
b100 &
0'
0(
b100 ,
#435390000000
1!
b100 %
1'
b100 +
#435400000000
0!
0'
#435410000000
1!
b101 %
1'
b101 +
#435420000000
0!
0'
#435430000000
1!
b110 %
1'
b110 +
#435440000000
0!
0'
#435450000000
1!
b111 %
1'
b111 +
#435460000000
0!
0'
#435470000000
1!
0$
b1000 %
1'
0*
b1000 +
#435480000000
0!
0'
#435490000000
1!
b1001 %
1'
b1001 +
#435500000000
0!
0'
#435510000000
1!
b0 %
1'
b0 +
#435520000000
0!
0'
#435530000000
1!
1$
b1 %
1'
1*
b1 +
#435540000000
0!
0'
#435550000000
1!
b10 %
1'
b10 +
#435560000000
0!
0'
#435570000000
1!
b11 %
1'
b11 +
#435580000000
0!
0'
#435590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#435600000000
0!
0'
#435610000000
1!
b101 %
1'
b101 +
#435620000000
0!
0'
#435630000000
1!
0$
b110 %
1'
0*
b110 +
#435640000000
0!
0'
#435650000000
1!
b111 %
1'
b111 +
#435660000000
0!
0'
#435670000000
1!
b1000 %
1'
b1000 +
#435680000000
0!
0'
#435690000000
1!
b1001 %
1'
b1001 +
#435700000000
0!
0'
#435710000000
1!
b0 %
1'
b0 +
#435720000000
0!
0'
#435730000000
1!
1$
b1 %
1'
1*
b1 +
#435740000000
0!
0'
#435750000000
1!
b10 %
1'
b10 +
#435760000000
0!
0'
#435770000000
1!
b11 %
1'
b11 +
#435780000000
0!
0'
#435790000000
1!
b100 %
1'
b100 +
#435800000000
1"
1(
#435810000000
0!
0"
b100 &
0'
0(
b100 ,
#435820000000
1!
b101 %
1'
b101 +
#435830000000
0!
0'
#435840000000
1!
b110 %
1'
b110 +
#435850000000
0!
0'
#435860000000
1!
b111 %
1'
b111 +
#435870000000
0!
0'
#435880000000
1!
0$
b1000 %
1'
0*
b1000 +
#435890000000
0!
0'
#435900000000
1!
b1001 %
1'
b1001 +
#435910000000
0!
0'
#435920000000
1!
b0 %
1'
b0 +
#435930000000
0!
0'
#435940000000
1!
1$
b1 %
1'
1*
b1 +
#435950000000
0!
0'
#435960000000
1!
b10 %
1'
b10 +
#435970000000
0!
0'
#435980000000
1!
b11 %
1'
b11 +
#435990000000
0!
0'
#436000000000
1!
b100 %
1'
b100 +
#436010000000
0!
0'
#436020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#436030000000
0!
0'
#436040000000
1!
0$
b110 %
1'
0*
b110 +
#436050000000
0!
0'
#436060000000
1!
b111 %
1'
b111 +
#436070000000
0!
0'
#436080000000
1!
b1000 %
1'
b1000 +
#436090000000
0!
0'
#436100000000
1!
b1001 %
1'
b1001 +
#436110000000
0!
0'
#436120000000
1!
b0 %
1'
b0 +
#436130000000
0!
0'
#436140000000
1!
1$
b1 %
1'
1*
b1 +
#436150000000
0!
0'
#436160000000
1!
b10 %
1'
b10 +
#436170000000
0!
0'
#436180000000
1!
b11 %
1'
b11 +
#436190000000
0!
0'
#436200000000
1!
b100 %
1'
b100 +
#436210000000
0!
0'
#436220000000
1!
b101 %
1'
b101 +
#436230000000
1"
1(
#436240000000
0!
0"
b100 &
0'
0(
b100 ,
#436250000000
1!
b110 %
1'
b110 +
#436260000000
0!
0'
#436270000000
1!
b111 %
1'
b111 +
#436280000000
0!
0'
#436290000000
1!
0$
b1000 %
1'
0*
b1000 +
#436300000000
0!
0'
#436310000000
1!
b1001 %
1'
b1001 +
#436320000000
0!
0'
#436330000000
1!
b0 %
1'
b0 +
#436340000000
0!
0'
#436350000000
1!
1$
b1 %
1'
1*
b1 +
#436360000000
0!
0'
#436370000000
1!
b10 %
1'
b10 +
#436380000000
0!
0'
#436390000000
1!
b11 %
1'
b11 +
#436400000000
0!
0'
#436410000000
1!
b100 %
1'
b100 +
#436420000000
0!
0'
#436430000000
1!
b101 %
1'
b101 +
#436440000000
0!
0'
#436450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#436460000000
0!
0'
#436470000000
1!
b111 %
1'
b111 +
#436480000000
0!
0'
#436490000000
1!
b1000 %
1'
b1000 +
#436500000000
0!
0'
#436510000000
1!
b1001 %
1'
b1001 +
#436520000000
0!
0'
#436530000000
1!
b0 %
1'
b0 +
#436540000000
0!
0'
#436550000000
1!
1$
b1 %
1'
1*
b1 +
#436560000000
0!
0'
#436570000000
1!
b10 %
1'
b10 +
#436580000000
0!
0'
#436590000000
1!
b11 %
1'
b11 +
#436600000000
0!
0'
#436610000000
1!
b100 %
1'
b100 +
#436620000000
0!
0'
#436630000000
1!
b101 %
1'
b101 +
#436640000000
0!
0'
#436650000000
1!
0$
b110 %
1'
0*
b110 +
#436660000000
1"
1(
#436670000000
0!
0"
b100 &
0'
0(
b100 ,
#436680000000
1!
1$
b111 %
1'
1*
b111 +
#436690000000
0!
0'
#436700000000
1!
0$
b1000 %
1'
0*
b1000 +
#436710000000
0!
0'
#436720000000
1!
b1001 %
1'
b1001 +
#436730000000
0!
0'
#436740000000
1!
b0 %
1'
b0 +
#436750000000
0!
0'
#436760000000
1!
1$
b1 %
1'
1*
b1 +
#436770000000
0!
0'
#436780000000
1!
b10 %
1'
b10 +
#436790000000
0!
0'
#436800000000
1!
b11 %
1'
b11 +
#436810000000
0!
0'
#436820000000
1!
b100 %
1'
b100 +
#436830000000
0!
0'
#436840000000
1!
b101 %
1'
b101 +
#436850000000
0!
0'
#436860000000
1!
b110 %
1'
b110 +
#436870000000
0!
0'
#436880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#436890000000
0!
0'
#436900000000
1!
b1000 %
1'
b1000 +
#436910000000
0!
0'
#436920000000
1!
b1001 %
1'
b1001 +
#436930000000
0!
0'
#436940000000
1!
b0 %
1'
b0 +
#436950000000
0!
0'
#436960000000
1!
1$
b1 %
1'
1*
b1 +
#436970000000
0!
0'
#436980000000
1!
b10 %
1'
b10 +
#436990000000
0!
0'
#437000000000
1!
b11 %
1'
b11 +
#437010000000
0!
0'
#437020000000
1!
b100 %
1'
b100 +
#437030000000
0!
0'
#437040000000
1!
b101 %
1'
b101 +
#437050000000
0!
0'
#437060000000
1!
0$
b110 %
1'
0*
b110 +
#437070000000
0!
0'
#437080000000
1!
b111 %
1'
b111 +
#437090000000
1"
1(
#437100000000
0!
0"
b100 &
0'
0(
b100 ,
#437110000000
1!
b1000 %
1'
b1000 +
#437120000000
0!
0'
#437130000000
1!
b1001 %
1'
b1001 +
#437140000000
0!
0'
#437150000000
1!
b0 %
1'
b0 +
#437160000000
0!
0'
#437170000000
1!
1$
b1 %
1'
1*
b1 +
#437180000000
0!
0'
#437190000000
1!
b10 %
1'
b10 +
#437200000000
0!
0'
#437210000000
1!
b11 %
1'
b11 +
#437220000000
0!
0'
#437230000000
1!
b100 %
1'
b100 +
#437240000000
0!
0'
#437250000000
1!
b101 %
1'
b101 +
#437260000000
0!
0'
#437270000000
1!
b110 %
1'
b110 +
#437280000000
0!
0'
#437290000000
1!
b111 %
1'
b111 +
#437300000000
0!
0'
#437310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#437320000000
0!
0'
#437330000000
1!
b1001 %
1'
b1001 +
#437340000000
0!
0'
#437350000000
1!
b0 %
1'
b0 +
#437360000000
0!
0'
#437370000000
1!
1$
b1 %
1'
1*
b1 +
#437380000000
0!
0'
#437390000000
1!
b10 %
1'
b10 +
#437400000000
0!
0'
#437410000000
1!
b11 %
1'
b11 +
#437420000000
0!
0'
#437430000000
1!
b100 %
1'
b100 +
#437440000000
0!
0'
#437450000000
1!
b101 %
1'
b101 +
#437460000000
0!
0'
#437470000000
1!
0$
b110 %
1'
0*
b110 +
#437480000000
0!
0'
#437490000000
1!
b111 %
1'
b111 +
#437500000000
0!
0'
#437510000000
1!
b1000 %
1'
b1000 +
#437520000000
1"
1(
#437530000000
0!
0"
b100 &
0'
0(
b100 ,
#437540000000
1!
b1001 %
1'
b1001 +
#437550000000
0!
0'
#437560000000
1!
b0 %
1'
b0 +
#437570000000
0!
0'
#437580000000
1!
1$
b1 %
1'
1*
b1 +
#437590000000
0!
0'
#437600000000
1!
b10 %
1'
b10 +
#437610000000
0!
0'
#437620000000
1!
b11 %
1'
b11 +
#437630000000
0!
0'
#437640000000
1!
b100 %
1'
b100 +
#437650000000
0!
0'
#437660000000
1!
b101 %
1'
b101 +
#437670000000
0!
0'
#437680000000
1!
b110 %
1'
b110 +
#437690000000
0!
0'
#437700000000
1!
b111 %
1'
b111 +
#437710000000
0!
0'
#437720000000
1!
0$
b1000 %
1'
0*
b1000 +
#437730000000
0!
0'
#437740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#437750000000
0!
0'
#437760000000
1!
b0 %
1'
b0 +
#437770000000
0!
0'
#437780000000
1!
1$
b1 %
1'
1*
b1 +
#437790000000
0!
0'
#437800000000
1!
b10 %
1'
b10 +
#437810000000
0!
0'
#437820000000
1!
b11 %
1'
b11 +
#437830000000
0!
0'
#437840000000
1!
b100 %
1'
b100 +
#437850000000
0!
0'
#437860000000
1!
b101 %
1'
b101 +
#437870000000
0!
0'
#437880000000
1!
0$
b110 %
1'
0*
b110 +
#437890000000
0!
0'
#437900000000
1!
b111 %
1'
b111 +
#437910000000
0!
0'
#437920000000
1!
b1000 %
1'
b1000 +
#437930000000
0!
0'
#437940000000
1!
b1001 %
1'
b1001 +
#437950000000
1"
1(
#437960000000
0!
0"
b100 &
0'
0(
b100 ,
#437970000000
1!
b0 %
1'
b0 +
#437980000000
0!
0'
#437990000000
1!
1$
b1 %
1'
1*
b1 +
#438000000000
0!
0'
#438010000000
1!
b10 %
1'
b10 +
#438020000000
0!
0'
#438030000000
1!
b11 %
1'
b11 +
#438040000000
0!
0'
#438050000000
1!
b100 %
1'
b100 +
#438060000000
0!
0'
#438070000000
1!
b101 %
1'
b101 +
#438080000000
0!
0'
#438090000000
1!
b110 %
1'
b110 +
#438100000000
0!
0'
#438110000000
1!
b111 %
1'
b111 +
#438120000000
0!
0'
#438130000000
1!
0$
b1000 %
1'
0*
b1000 +
#438140000000
0!
0'
#438150000000
1!
b1001 %
1'
b1001 +
#438160000000
0!
0'
#438170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#438180000000
0!
0'
#438190000000
1!
1$
b1 %
1'
1*
b1 +
#438200000000
0!
0'
#438210000000
1!
b10 %
1'
b10 +
#438220000000
0!
0'
#438230000000
1!
b11 %
1'
b11 +
#438240000000
0!
0'
#438250000000
1!
b100 %
1'
b100 +
#438260000000
0!
0'
#438270000000
1!
b101 %
1'
b101 +
#438280000000
0!
0'
#438290000000
1!
0$
b110 %
1'
0*
b110 +
#438300000000
0!
0'
#438310000000
1!
b111 %
1'
b111 +
#438320000000
0!
0'
#438330000000
1!
b1000 %
1'
b1000 +
#438340000000
0!
0'
#438350000000
1!
b1001 %
1'
b1001 +
#438360000000
0!
0'
#438370000000
1!
b0 %
1'
b0 +
#438380000000
1"
1(
#438390000000
0!
0"
b100 &
0'
0(
b100 ,
#438400000000
1!
1$
b1 %
1'
1*
b1 +
#438410000000
0!
0'
#438420000000
1!
b10 %
1'
b10 +
#438430000000
0!
0'
#438440000000
1!
b11 %
1'
b11 +
#438450000000
0!
0'
#438460000000
1!
b100 %
1'
b100 +
#438470000000
0!
0'
#438480000000
1!
b101 %
1'
b101 +
#438490000000
0!
0'
#438500000000
1!
b110 %
1'
b110 +
#438510000000
0!
0'
#438520000000
1!
b111 %
1'
b111 +
#438530000000
0!
0'
#438540000000
1!
0$
b1000 %
1'
0*
b1000 +
#438550000000
0!
0'
#438560000000
1!
b1001 %
1'
b1001 +
#438570000000
0!
0'
#438580000000
1!
b0 %
1'
b0 +
#438590000000
0!
0'
#438600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#438610000000
0!
0'
#438620000000
1!
b10 %
1'
b10 +
#438630000000
0!
0'
#438640000000
1!
b11 %
1'
b11 +
#438650000000
0!
0'
#438660000000
1!
b100 %
1'
b100 +
#438670000000
0!
0'
#438680000000
1!
b101 %
1'
b101 +
#438690000000
0!
0'
#438700000000
1!
0$
b110 %
1'
0*
b110 +
#438710000000
0!
0'
#438720000000
1!
b111 %
1'
b111 +
#438730000000
0!
0'
#438740000000
1!
b1000 %
1'
b1000 +
#438750000000
0!
0'
#438760000000
1!
b1001 %
1'
b1001 +
#438770000000
0!
0'
#438780000000
1!
b0 %
1'
b0 +
#438790000000
0!
0'
#438800000000
1!
1$
b1 %
1'
1*
b1 +
#438810000000
1"
1(
#438820000000
0!
0"
b100 &
0'
0(
b100 ,
#438830000000
1!
b10 %
1'
b10 +
#438840000000
0!
0'
#438850000000
1!
b11 %
1'
b11 +
#438860000000
0!
0'
#438870000000
1!
b100 %
1'
b100 +
#438880000000
0!
0'
#438890000000
1!
b101 %
1'
b101 +
#438900000000
0!
0'
#438910000000
1!
b110 %
1'
b110 +
#438920000000
0!
0'
#438930000000
1!
b111 %
1'
b111 +
#438940000000
0!
0'
#438950000000
1!
0$
b1000 %
1'
0*
b1000 +
#438960000000
0!
0'
#438970000000
1!
b1001 %
1'
b1001 +
#438980000000
0!
0'
#438990000000
1!
b0 %
1'
b0 +
#439000000000
0!
0'
#439010000000
1!
1$
b1 %
1'
1*
b1 +
#439020000000
0!
0'
#439030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#439040000000
0!
0'
#439050000000
1!
b11 %
1'
b11 +
#439060000000
0!
0'
#439070000000
1!
b100 %
1'
b100 +
#439080000000
0!
0'
#439090000000
1!
b101 %
1'
b101 +
#439100000000
0!
0'
#439110000000
1!
0$
b110 %
1'
0*
b110 +
#439120000000
0!
0'
#439130000000
1!
b111 %
1'
b111 +
#439140000000
0!
0'
#439150000000
1!
b1000 %
1'
b1000 +
#439160000000
0!
0'
#439170000000
1!
b1001 %
1'
b1001 +
#439180000000
0!
0'
#439190000000
1!
b0 %
1'
b0 +
#439200000000
0!
0'
#439210000000
1!
1$
b1 %
1'
1*
b1 +
#439220000000
0!
0'
#439230000000
1!
b10 %
1'
b10 +
#439240000000
1"
1(
#439250000000
0!
0"
b100 &
0'
0(
b100 ,
#439260000000
1!
b11 %
1'
b11 +
#439270000000
0!
0'
#439280000000
1!
b100 %
1'
b100 +
#439290000000
0!
0'
#439300000000
1!
b101 %
1'
b101 +
#439310000000
0!
0'
#439320000000
1!
b110 %
1'
b110 +
#439330000000
0!
0'
#439340000000
1!
b111 %
1'
b111 +
#439350000000
0!
0'
#439360000000
1!
0$
b1000 %
1'
0*
b1000 +
#439370000000
0!
0'
#439380000000
1!
b1001 %
1'
b1001 +
#439390000000
0!
0'
#439400000000
1!
b0 %
1'
b0 +
#439410000000
0!
0'
#439420000000
1!
1$
b1 %
1'
1*
b1 +
#439430000000
0!
0'
#439440000000
1!
b10 %
1'
b10 +
#439450000000
0!
0'
#439460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#439470000000
0!
0'
#439480000000
1!
b100 %
1'
b100 +
#439490000000
0!
0'
#439500000000
1!
b101 %
1'
b101 +
#439510000000
0!
0'
#439520000000
1!
0$
b110 %
1'
0*
b110 +
#439530000000
0!
0'
#439540000000
1!
b111 %
1'
b111 +
#439550000000
0!
0'
#439560000000
1!
b1000 %
1'
b1000 +
#439570000000
0!
0'
#439580000000
1!
b1001 %
1'
b1001 +
#439590000000
0!
0'
#439600000000
1!
b0 %
1'
b0 +
#439610000000
0!
0'
#439620000000
1!
1$
b1 %
1'
1*
b1 +
#439630000000
0!
0'
#439640000000
1!
b10 %
1'
b10 +
#439650000000
0!
0'
#439660000000
1!
b11 %
1'
b11 +
#439670000000
1"
1(
#439680000000
0!
0"
b100 &
0'
0(
b100 ,
#439690000000
1!
b100 %
1'
b100 +
#439700000000
0!
0'
#439710000000
1!
b101 %
1'
b101 +
#439720000000
0!
0'
#439730000000
1!
b110 %
1'
b110 +
#439740000000
0!
0'
#439750000000
1!
b111 %
1'
b111 +
#439760000000
0!
0'
#439770000000
1!
0$
b1000 %
1'
0*
b1000 +
#439780000000
0!
0'
#439790000000
1!
b1001 %
1'
b1001 +
#439800000000
0!
0'
#439810000000
1!
b0 %
1'
b0 +
#439820000000
0!
0'
#439830000000
1!
1$
b1 %
1'
1*
b1 +
#439840000000
0!
0'
#439850000000
1!
b10 %
1'
b10 +
#439860000000
0!
0'
#439870000000
1!
b11 %
1'
b11 +
#439880000000
0!
0'
#439890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#439900000000
0!
0'
#439910000000
1!
b101 %
1'
b101 +
#439920000000
0!
0'
#439930000000
1!
0$
b110 %
1'
0*
b110 +
#439940000000
0!
0'
#439950000000
1!
b111 %
1'
b111 +
#439960000000
0!
0'
#439970000000
1!
b1000 %
1'
b1000 +
#439980000000
0!
0'
#439990000000
1!
b1001 %
1'
b1001 +
#440000000000
0!
0'
#440010000000
1!
b0 %
1'
b0 +
#440020000000
0!
0'
#440030000000
1!
1$
b1 %
1'
1*
b1 +
#440040000000
0!
0'
#440050000000
1!
b10 %
1'
b10 +
#440060000000
0!
0'
#440070000000
1!
b11 %
1'
b11 +
#440080000000
0!
0'
#440090000000
1!
b100 %
1'
b100 +
#440100000000
1"
1(
#440110000000
0!
0"
b100 &
0'
0(
b100 ,
#440120000000
1!
b101 %
1'
b101 +
#440130000000
0!
0'
#440140000000
1!
b110 %
1'
b110 +
#440150000000
0!
0'
#440160000000
1!
b111 %
1'
b111 +
#440170000000
0!
0'
#440180000000
1!
0$
b1000 %
1'
0*
b1000 +
#440190000000
0!
0'
#440200000000
1!
b1001 %
1'
b1001 +
#440210000000
0!
0'
#440220000000
1!
b0 %
1'
b0 +
#440230000000
0!
0'
#440240000000
1!
1$
b1 %
1'
1*
b1 +
#440250000000
0!
0'
#440260000000
1!
b10 %
1'
b10 +
#440270000000
0!
0'
#440280000000
1!
b11 %
1'
b11 +
#440290000000
0!
0'
#440300000000
1!
b100 %
1'
b100 +
#440310000000
0!
0'
#440320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#440330000000
0!
0'
#440340000000
1!
0$
b110 %
1'
0*
b110 +
#440350000000
0!
0'
#440360000000
1!
b111 %
1'
b111 +
#440370000000
0!
0'
#440380000000
1!
b1000 %
1'
b1000 +
#440390000000
0!
0'
#440400000000
1!
b1001 %
1'
b1001 +
#440410000000
0!
0'
#440420000000
1!
b0 %
1'
b0 +
#440430000000
0!
0'
#440440000000
1!
1$
b1 %
1'
1*
b1 +
#440450000000
0!
0'
#440460000000
1!
b10 %
1'
b10 +
#440470000000
0!
0'
#440480000000
1!
b11 %
1'
b11 +
#440490000000
0!
0'
#440500000000
1!
b100 %
1'
b100 +
#440510000000
0!
0'
#440520000000
1!
b101 %
1'
b101 +
#440530000000
1"
1(
#440540000000
0!
0"
b100 &
0'
0(
b100 ,
#440550000000
1!
b110 %
1'
b110 +
#440560000000
0!
0'
#440570000000
1!
b111 %
1'
b111 +
#440580000000
0!
0'
#440590000000
1!
0$
b1000 %
1'
0*
b1000 +
#440600000000
0!
0'
#440610000000
1!
b1001 %
1'
b1001 +
#440620000000
0!
0'
#440630000000
1!
b0 %
1'
b0 +
#440640000000
0!
0'
#440650000000
1!
1$
b1 %
1'
1*
b1 +
#440660000000
0!
0'
#440670000000
1!
b10 %
1'
b10 +
#440680000000
0!
0'
#440690000000
1!
b11 %
1'
b11 +
#440700000000
0!
0'
#440710000000
1!
b100 %
1'
b100 +
#440720000000
0!
0'
#440730000000
1!
b101 %
1'
b101 +
#440740000000
0!
0'
#440750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#440760000000
0!
0'
#440770000000
1!
b111 %
1'
b111 +
#440780000000
0!
0'
#440790000000
1!
b1000 %
1'
b1000 +
#440800000000
0!
0'
#440810000000
1!
b1001 %
1'
b1001 +
#440820000000
0!
0'
#440830000000
1!
b0 %
1'
b0 +
#440840000000
0!
0'
#440850000000
1!
1$
b1 %
1'
1*
b1 +
#440860000000
0!
0'
#440870000000
1!
b10 %
1'
b10 +
#440880000000
0!
0'
#440890000000
1!
b11 %
1'
b11 +
#440900000000
0!
0'
#440910000000
1!
b100 %
1'
b100 +
#440920000000
0!
0'
#440930000000
1!
b101 %
1'
b101 +
#440940000000
0!
0'
#440950000000
1!
0$
b110 %
1'
0*
b110 +
#440960000000
1"
1(
#440970000000
0!
0"
b100 &
0'
0(
b100 ,
#440980000000
1!
1$
b111 %
1'
1*
b111 +
#440990000000
0!
0'
#441000000000
1!
0$
b1000 %
1'
0*
b1000 +
#441010000000
0!
0'
#441020000000
1!
b1001 %
1'
b1001 +
#441030000000
0!
0'
#441040000000
1!
b0 %
1'
b0 +
#441050000000
0!
0'
#441060000000
1!
1$
b1 %
1'
1*
b1 +
#441070000000
0!
0'
#441080000000
1!
b10 %
1'
b10 +
#441090000000
0!
0'
#441100000000
1!
b11 %
1'
b11 +
#441110000000
0!
0'
#441120000000
1!
b100 %
1'
b100 +
#441130000000
0!
0'
#441140000000
1!
b101 %
1'
b101 +
#441150000000
0!
0'
#441160000000
1!
b110 %
1'
b110 +
#441170000000
0!
0'
#441180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#441190000000
0!
0'
#441200000000
1!
b1000 %
1'
b1000 +
#441210000000
0!
0'
#441220000000
1!
b1001 %
1'
b1001 +
#441230000000
0!
0'
#441240000000
1!
b0 %
1'
b0 +
#441250000000
0!
0'
#441260000000
1!
1$
b1 %
1'
1*
b1 +
#441270000000
0!
0'
#441280000000
1!
b10 %
1'
b10 +
#441290000000
0!
0'
#441300000000
1!
b11 %
1'
b11 +
#441310000000
0!
0'
#441320000000
1!
b100 %
1'
b100 +
#441330000000
0!
0'
#441340000000
1!
b101 %
1'
b101 +
#441350000000
0!
0'
#441360000000
1!
0$
b110 %
1'
0*
b110 +
#441370000000
0!
0'
#441380000000
1!
b111 %
1'
b111 +
#441390000000
1"
1(
#441400000000
0!
0"
b100 &
0'
0(
b100 ,
#441410000000
1!
b1000 %
1'
b1000 +
#441420000000
0!
0'
#441430000000
1!
b1001 %
1'
b1001 +
#441440000000
0!
0'
#441450000000
1!
b0 %
1'
b0 +
#441460000000
0!
0'
#441470000000
1!
1$
b1 %
1'
1*
b1 +
#441480000000
0!
0'
#441490000000
1!
b10 %
1'
b10 +
#441500000000
0!
0'
#441510000000
1!
b11 %
1'
b11 +
#441520000000
0!
0'
#441530000000
1!
b100 %
1'
b100 +
#441540000000
0!
0'
#441550000000
1!
b101 %
1'
b101 +
#441560000000
0!
0'
#441570000000
1!
b110 %
1'
b110 +
#441580000000
0!
0'
#441590000000
1!
b111 %
1'
b111 +
#441600000000
0!
0'
#441610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#441620000000
0!
0'
#441630000000
1!
b1001 %
1'
b1001 +
#441640000000
0!
0'
#441650000000
1!
b0 %
1'
b0 +
#441660000000
0!
0'
#441670000000
1!
1$
b1 %
1'
1*
b1 +
#441680000000
0!
0'
#441690000000
1!
b10 %
1'
b10 +
#441700000000
0!
0'
#441710000000
1!
b11 %
1'
b11 +
#441720000000
0!
0'
#441730000000
1!
b100 %
1'
b100 +
#441740000000
0!
0'
#441750000000
1!
b101 %
1'
b101 +
#441760000000
0!
0'
#441770000000
1!
0$
b110 %
1'
0*
b110 +
#441780000000
0!
0'
#441790000000
1!
b111 %
1'
b111 +
#441800000000
0!
0'
#441810000000
1!
b1000 %
1'
b1000 +
#441820000000
1"
1(
#441830000000
0!
0"
b100 &
0'
0(
b100 ,
#441840000000
1!
b1001 %
1'
b1001 +
#441850000000
0!
0'
#441860000000
1!
b0 %
1'
b0 +
#441870000000
0!
0'
#441880000000
1!
1$
b1 %
1'
1*
b1 +
#441890000000
0!
0'
#441900000000
1!
b10 %
1'
b10 +
#441910000000
0!
0'
#441920000000
1!
b11 %
1'
b11 +
#441930000000
0!
0'
#441940000000
1!
b100 %
1'
b100 +
#441950000000
0!
0'
#441960000000
1!
b101 %
1'
b101 +
#441970000000
0!
0'
#441980000000
1!
b110 %
1'
b110 +
#441990000000
0!
0'
#442000000000
1!
b111 %
1'
b111 +
#442010000000
0!
0'
#442020000000
1!
0$
b1000 %
1'
0*
b1000 +
#442030000000
0!
0'
#442040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#442050000000
0!
0'
#442060000000
1!
b0 %
1'
b0 +
#442070000000
0!
0'
#442080000000
1!
1$
b1 %
1'
1*
b1 +
#442090000000
0!
0'
#442100000000
1!
b10 %
1'
b10 +
#442110000000
0!
0'
#442120000000
1!
b11 %
1'
b11 +
#442130000000
0!
0'
#442140000000
1!
b100 %
1'
b100 +
#442150000000
0!
0'
#442160000000
1!
b101 %
1'
b101 +
#442170000000
0!
0'
#442180000000
1!
0$
b110 %
1'
0*
b110 +
#442190000000
0!
0'
#442200000000
1!
b111 %
1'
b111 +
#442210000000
0!
0'
#442220000000
1!
b1000 %
1'
b1000 +
#442230000000
0!
0'
#442240000000
1!
b1001 %
1'
b1001 +
#442250000000
1"
1(
#442260000000
0!
0"
b100 &
0'
0(
b100 ,
#442270000000
1!
b0 %
1'
b0 +
#442280000000
0!
0'
#442290000000
1!
1$
b1 %
1'
1*
b1 +
#442300000000
0!
0'
#442310000000
1!
b10 %
1'
b10 +
#442320000000
0!
0'
#442330000000
1!
b11 %
1'
b11 +
#442340000000
0!
0'
#442350000000
1!
b100 %
1'
b100 +
#442360000000
0!
0'
#442370000000
1!
b101 %
1'
b101 +
#442380000000
0!
0'
#442390000000
1!
b110 %
1'
b110 +
#442400000000
0!
0'
#442410000000
1!
b111 %
1'
b111 +
#442420000000
0!
0'
#442430000000
1!
0$
b1000 %
1'
0*
b1000 +
#442440000000
0!
0'
#442450000000
1!
b1001 %
1'
b1001 +
#442460000000
0!
0'
#442470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#442480000000
0!
0'
#442490000000
1!
1$
b1 %
1'
1*
b1 +
#442500000000
0!
0'
#442510000000
1!
b10 %
1'
b10 +
#442520000000
0!
0'
#442530000000
1!
b11 %
1'
b11 +
#442540000000
0!
0'
#442550000000
1!
b100 %
1'
b100 +
#442560000000
0!
0'
#442570000000
1!
b101 %
1'
b101 +
#442580000000
0!
0'
#442590000000
1!
0$
b110 %
1'
0*
b110 +
#442600000000
0!
0'
#442610000000
1!
b111 %
1'
b111 +
#442620000000
0!
0'
#442630000000
1!
b1000 %
1'
b1000 +
#442640000000
0!
0'
#442650000000
1!
b1001 %
1'
b1001 +
#442660000000
0!
0'
#442670000000
1!
b0 %
1'
b0 +
#442680000000
1"
1(
#442690000000
0!
0"
b100 &
0'
0(
b100 ,
#442700000000
1!
1$
b1 %
1'
1*
b1 +
#442710000000
0!
0'
#442720000000
1!
b10 %
1'
b10 +
#442730000000
0!
0'
#442740000000
1!
b11 %
1'
b11 +
#442750000000
0!
0'
#442760000000
1!
b100 %
1'
b100 +
#442770000000
0!
0'
#442780000000
1!
b101 %
1'
b101 +
#442790000000
0!
0'
#442800000000
1!
b110 %
1'
b110 +
#442810000000
0!
0'
#442820000000
1!
b111 %
1'
b111 +
#442830000000
0!
0'
#442840000000
1!
0$
b1000 %
1'
0*
b1000 +
#442850000000
0!
0'
#442860000000
1!
b1001 %
1'
b1001 +
#442870000000
0!
0'
#442880000000
1!
b0 %
1'
b0 +
#442890000000
0!
0'
#442900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#442910000000
0!
0'
#442920000000
1!
b10 %
1'
b10 +
#442930000000
0!
0'
#442940000000
1!
b11 %
1'
b11 +
#442950000000
0!
0'
#442960000000
1!
b100 %
1'
b100 +
#442970000000
0!
0'
#442980000000
1!
b101 %
1'
b101 +
#442990000000
0!
0'
#443000000000
1!
0$
b110 %
1'
0*
b110 +
#443010000000
0!
0'
#443020000000
1!
b111 %
1'
b111 +
#443030000000
0!
0'
#443040000000
1!
b1000 %
1'
b1000 +
#443050000000
0!
0'
#443060000000
1!
b1001 %
1'
b1001 +
#443070000000
0!
0'
#443080000000
1!
b0 %
1'
b0 +
#443090000000
0!
0'
#443100000000
1!
1$
b1 %
1'
1*
b1 +
#443110000000
1"
1(
#443120000000
0!
0"
b100 &
0'
0(
b100 ,
#443130000000
1!
b10 %
1'
b10 +
#443140000000
0!
0'
#443150000000
1!
b11 %
1'
b11 +
#443160000000
0!
0'
#443170000000
1!
b100 %
1'
b100 +
#443180000000
0!
0'
#443190000000
1!
b101 %
1'
b101 +
#443200000000
0!
0'
#443210000000
1!
b110 %
1'
b110 +
#443220000000
0!
0'
#443230000000
1!
b111 %
1'
b111 +
#443240000000
0!
0'
#443250000000
1!
0$
b1000 %
1'
0*
b1000 +
#443260000000
0!
0'
#443270000000
1!
b1001 %
1'
b1001 +
#443280000000
0!
0'
#443290000000
1!
b0 %
1'
b0 +
#443300000000
0!
0'
#443310000000
1!
1$
b1 %
1'
1*
b1 +
#443320000000
0!
0'
#443330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#443340000000
0!
0'
#443350000000
1!
b11 %
1'
b11 +
#443360000000
0!
0'
#443370000000
1!
b100 %
1'
b100 +
#443380000000
0!
0'
#443390000000
1!
b101 %
1'
b101 +
#443400000000
0!
0'
#443410000000
1!
0$
b110 %
1'
0*
b110 +
#443420000000
0!
0'
#443430000000
1!
b111 %
1'
b111 +
#443440000000
0!
0'
#443450000000
1!
b1000 %
1'
b1000 +
#443460000000
0!
0'
#443470000000
1!
b1001 %
1'
b1001 +
#443480000000
0!
0'
#443490000000
1!
b0 %
1'
b0 +
#443500000000
0!
0'
#443510000000
1!
1$
b1 %
1'
1*
b1 +
#443520000000
0!
0'
#443530000000
1!
b10 %
1'
b10 +
#443540000000
1"
1(
#443550000000
0!
0"
b100 &
0'
0(
b100 ,
#443560000000
1!
b11 %
1'
b11 +
#443570000000
0!
0'
#443580000000
1!
b100 %
1'
b100 +
#443590000000
0!
0'
#443600000000
1!
b101 %
1'
b101 +
#443610000000
0!
0'
#443620000000
1!
b110 %
1'
b110 +
#443630000000
0!
0'
#443640000000
1!
b111 %
1'
b111 +
#443650000000
0!
0'
#443660000000
1!
0$
b1000 %
1'
0*
b1000 +
#443670000000
0!
0'
#443680000000
1!
b1001 %
1'
b1001 +
#443690000000
0!
0'
#443700000000
1!
b0 %
1'
b0 +
#443710000000
0!
0'
#443720000000
1!
1$
b1 %
1'
1*
b1 +
#443730000000
0!
0'
#443740000000
1!
b10 %
1'
b10 +
#443750000000
0!
0'
#443760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#443770000000
0!
0'
#443780000000
1!
b100 %
1'
b100 +
#443790000000
0!
0'
#443800000000
1!
b101 %
1'
b101 +
#443810000000
0!
0'
#443820000000
1!
0$
b110 %
1'
0*
b110 +
#443830000000
0!
0'
#443840000000
1!
b111 %
1'
b111 +
#443850000000
0!
0'
#443860000000
1!
b1000 %
1'
b1000 +
#443870000000
0!
0'
#443880000000
1!
b1001 %
1'
b1001 +
#443890000000
0!
0'
#443900000000
1!
b0 %
1'
b0 +
#443910000000
0!
0'
#443920000000
1!
1$
b1 %
1'
1*
b1 +
#443930000000
0!
0'
#443940000000
1!
b10 %
1'
b10 +
#443950000000
0!
0'
#443960000000
1!
b11 %
1'
b11 +
#443970000000
1"
1(
#443980000000
0!
0"
b100 &
0'
0(
b100 ,
#443990000000
1!
b100 %
1'
b100 +
#444000000000
0!
0'
#444010000000
1!
b101 %
1'
b101 +
#444020000000
0!
0'
#444030000000
1!
b110 %
1'
b110 +
#444040000000
0!
0'
#444050000000
1!
b111 %
1'
b111 +
#444060000000
0!
0'
#444070000000
1!
0$
b1000 %
1'
0*
b1000 +
#444080000000
0!
0'
#444090000000
1!
b1001 %
1'
b1001 +
#444100000000
0!
0'
#444110000000
1!
b0 %
1'
b0 +
#444120000000
0!
0'
#444130000000
1!
1$
b1 %
1'
1*
b1 +
#444140000000
0!
0'
#444150000000
1!
b10 %
1'
b10 +
#444160000000
0!
0'
#444170000000
1!
b11 %
1'
b11 +
#444180000000
0!
0'
#444190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#444200000000
0!
0'
#444210000000
1!
b101 %
1'
b101 +
#444220000000
0!
0'
#444230000000
1!
0$
b110 %
1'
0*
b110 +
#444240000000
0!
0'
#444250000000
1!
b111 %
1'
b111 +
#444260000000
0!
0'
#444270000000
1!
b1000 %
1'
b1000 +
#444280000000
0!
0'
#444290000000
1!
b1001 %
1'
b1001 +
#444300000000
0!
0'
#444310000000
1!
b0 %
1'
b0 +
#444320000000
0!
0'
#444330000000
1!
1$
b1 %
1'
1*
b1 +
#444340000000
0!
0'
#444350000000
1!
b10 %
1'
b10 +
#444360000000
0!
0'
#444370000000
1!
b11 %
1'
b11 +
#444380000000
0!
0'
#444390000000
1!
b100 %
1'
b100 +
#444400000000
1"
1(
#444410000000
0!
0"
b100 &
0'
0(
b100 ,
#444420000000
1!
b101 %
1'
b101 +
#444430000000
0!
0'
#444440000000
1!
b110 %
1'
b110 +
#444450000000
0!
0'
#444460000000
1!
b111 %
1'
b111 +
#444470000000
0!
0'
#444480000000
1!
0$
b1000 %
1'
0*
b1000 +
#444490000000
0!
0'
#444500000000
1!
b1001 %
1'
b1001 +
#444510000000
0!
0'
#444520000000
1!
b0 %
1'
b0 +
#444530000000
0!
0'
#444540000000
1!
1$
b1 %
1'
1*
b1 +
#444550000000
0!
0'
#444560000000
1!
b10 %
1'
b10 +
#444570000000
0!
0'
#444580000000
1!
b11 %
1'
b11 +
#444590000000
0!
0'
#444600000000
1!
b100 %
1'
b100 +
#444610000000
0!
0'
#444620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#444630000000
0!
0'
#444640000000
1!
0$
b110 %
1'
0*
b110 +
#444650000000
0!
0'
#444660000000
1!
b111 %
1'
b111 +
#444670000000
0!
0'
#444680000000
1!
b1000 %
1'
b1000 +
#444690000000
0!
0'
#444700000000
1!
b1001 %
1'
b1001 +
#444710000000
0!
0'
#444720000000
1!
b0 %
1'
b0 +
#444730000000
0!
0'
#444740000000
1!
1$
b1 %
1'
1*
b1 +
#444750000000
0!
0'
#444760000000
1!
b10 %
1'
b10 +
#444770000000
0!
0'
#444780000000
1!
b11 %
1'
b11 +
#444790000000
0!
0'
#444800000000
1!
b100 %
1'
b100 +
#444810000000
0!
0'
#444820000000
1!
b101 %
1'
b101 +
#444830000000
1"
1(
#444840000000
0!
0"
b100 &
0'
0(
b100 ,
#444850000000
1!
b110 %
1'
b110 +
#444860000000
0!
0'
#444870000000
1!
b111 %
1'
b111 +
#444880000000
0!
0'
#444890000000
1!
0$
b1000 %
1'
0*
b1000 +
#444900000000
0!
0'
#444910000000
1!
b1001 %
1'
b1001 +
#444920000000
0!
0'
#444930000000
1!
b0 %
1'
b0 +
#444940000000
0!
0'
#444950000000
1!
1$
b1 %
1'
1*
b1 +
#444960000000
0!
0'
#444970000000
1!
b10 %
1'
b10 +
#444980000000
0!
0'
#444990000000
1!
b11 %
1'
b11 +
#445000000000
0!
0'
#445010000000
1!
b100 %
1'
b100 +
#445020000000
0!
0'
#445030000000
1!
b101 %
1'
b101 +
#445040000000
0!
0'
#445050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#445060000000
0!
0'
#445070000000
1!
b111 %
1'
b111 +
#445080000000
0!
0'
#445090000000
1!
b1000 %
1'
b1000 +
#445100000000
0!
0'
#445110000000
1!
b1001 %
1'
b1001 +
#445120000000
0!
0'
#445130000000
1!
b0 %
1'
b0 +
#445140000000
0!
0'
#445150000000
1!
1$
b1 %
1'
1*
b1 +
#445160000000
0!
0'
#445170000000
1!
b10 %
1'
b10 +
#445180000000
0!
0'
#445190000000
1!
b11 %
1'
b11 +
#445200000000
0!
0'
#445210000000
1!
b100 %
1'
b100 +
#445220000000
0!
0'
#445230000000
1!
b101 %
1'
b101 +
#445240000000
0!
0'
#445250000000
1!
0$
b110 %
1'
0*
b110 +
#445260000000
1"
1(
#445270000000
0!
0"
b100 &
0'
0(
b100 ,
#445280000000
1!
1$
b111 %
1'
1*
b111 +
#445290000000
0!
0'
#445300000000
1!
0$
b1000 %
1'
0*
b1000 +
#445310000000
0!
0'
#445320000000
1!
b1001 %
1'
b1001 +
#445330000000
0!
0'
#445340000000
1!
b0 %
1'
b0 +
#445350000000
0!
0'
#445360000000
1!
1$
b1 %
1'
1*
b1 +
#445370000000
0!
0'
#445380000000
1!
b10 %
1'
b10 +
#445390000000
0!
0'
#445400000000
1!
b11 %
1'
b11 +
#445410000000
0!
0'
#445420000000
1!
b100 %
1'
b100 +
#445430000000
0!
0'
#445440000000
1!
b101 %
1'
b101 +
#445450000000
0!
0'
#445460000000
1!
b110 %
1'
b110 +
#445470000000
0!
0'
#445480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#445490000000
0!
0'
#445500000000
1!
b1000 %
1'
b1000 +
#445510000000
0!
0'
#445520000000
1!
b1001 %
1'
b1001 +
#445530000000
0!
0'
#445540000000
1!
b0 %
1'
b0 +
#445550000000
0!
0'
#445560000000
1!
1$
b1 %
1'
1*
b1 +
#445570000000
0!
0'
#445580000000
1!
b10 %
1'
b10 +
#445590000000
0!
0'
#445600000000
1!
b11 %
1'
b11 +
#445610000000
0!
0'
#445620000000
1!
b100 %
1'
b100 +
#445630000000
0!
0'
#445640000000
1!
b101 %
1'
b101 +
#445650000000
0!
0'
#445660000000
1!
0$
b110 %
1'
0*
b110 +
#445670000000
0!
0'
#445680000000
1!
b111 %
1'
b111 +
#445690000000
1"
1(
#445700000000
0!
0"
b100 &
0'
0(
b100 ,
#445710000000
1!
b1000 %
1'
b1000 +
#445720000000
0!
0'
#445730000000
1!
b1001 %
1'
b1001 +
#445740000000
0!
0'
#445750000000
1!
b0 %
1'
b0 +
#445760000000
0!
0'
#445770000000
1!
1$
b1 %
1'
1*
b1 +
#445780000000
0!
0'
#445790000000
1!
b10 %
1'
b10 +
#445800000000
0!
0'
#445810000000
1!
b11 %
1'
b11 +
#445820000000
0!
0'
#445830000000
1!
b100 %
1'
b100 +
#445840000000
0!
0'
#445850000000
1!
b101 %
1'
b101 +
#445860000000
0!
0'
#445870000000
1!
b110 %
1'
b110 +
#445880000000
0!
0'
#445890000000
1!
b111 %
1'
b111 +
#445900000000
0!
0'
#445910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#445920000000
0!
0'
#445930000000
1!
b1001 %
1'
b1001 +
#445940000000
0!
0'
#445950000000
1!
b0 %
1'
b0 +
#445960000000
0!
0'
#445970000000
1!
1$
b1 %
1'
1*
b1 +
#445980000000
0!
0'
#445990000000
1!
b10 %
1'
b10 +
#446000000000
0!
0'
#446010000000
1!
b11 %
1'
b11 +
#446020000000
0!
0'
#446030000000
1!
b100 %
1'
b100 +
#446040000000
0!
0'
#446050000000
1!
b101 %
1'
b101 +
#446060000000
0!
0'
#446070000000
1!
0$
b110 %
1'
0*
b110 +
#446080000000
0!
0'
#446090000000
1!
b111 %
1'
b111 +
#446100000000
0!
0'
#446110000000
1!
b1000 %
1'
b1000 +
#446120000000
1"
1(
#446130000000
0!
0"
b100 &
0'
0(
b100 ,
#446140000000
1!
b1001 %
1'
b1001 +
#446150000000
0!
0'
#446160000000
1!
b0 %
1'
b0 +
#446170000000
0!
0'
#446180000000
1!
1$
b1 %
1'
1*
b1 +
#446190000000
0!
0'
#446200000000
1!
b10 %
1'
b10 +
#446210000000
0!
0'
#446220000000
1!
b11 %
1'
b11 +
#446230000000
0!
0'
#446240000000
1!
b100 %
1'
b100 +
#446250000000
0!
0'
#446260000000
1!
b101 %
1'
b101 +
#446270000000
0!
0'
#446280000000
1!
b110 %
1'
b110 +
#446290000000
0!
0'
#446300000000
1!
b111 %
1'
b111 +
#446310000000
0!
0'
#446320000000
1!
0$
b1000 %
1'
0*
b1000 +
#446330000000
0!
0'
#446340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#446350000000
0!
0'
#446360000000
1!
b0 %
1'
b0 +
#446370000000
0!
0'
#446380000000
1!
1$
b1 %
1'
1*
b1 +
#446390000000
0!
0'
#446400000000
1!
b10 %
1'
b10 +
#446410000000
0!
0'
#446420000000
1!
b11 %
1'
b11 +
#446430000000
0!
0'
#446440000000
1!
b100 %
1'
b100 +
#446450000000
0!
0'
#446460000000
1!
b101 %
1'
b101 +
#446470000000
0!
0'
#446480000000
1!
0$
b110 %
1'
0*
b110 +
#446490000000
0!
0'
#446500000000
1!
b111 %
1'
b111 +
#446510000000
0!
0'
#446520000000
1!
b1000 %
1'
b1000 +
#446530000000
0!
0'
#446540000000
1!
b1001 %
1'
b1001 +
#446550000000
1"
1(
#446560000000
0!
0"
b100 &
0'
0(
b100 ,
#446570000000
1!
b0 %
1'
b0 +
#446580000000
0!
0'
#446590000000
1!
1$
b1 %
1'
1*
b1 +
#446600000000
0!
0'
#446610000000
1!
b10 %
1'
b10 +
#446620000000
0!
0'
#446630000000
1!
b11 %
1'
b11 +
#446640000000
0!
0'
#446650000000
1!
b100 %
1'
b100 +
#446660000000
0!
0'
#446670000000
1!
b101 %
1'
b101 +
#446680000000
0!
0'
#446690000000
1!
b110 %
1'
b110 +
#446700000000
0!
0'
#446710000000
1!
b111 %
1'
b111 +
#446720000000
0!
0'
#446730000000
1!
0$
b1000 %
1'
0*
b1000 +
#446740000000
0!
0'
#446750000000
1!
b1001 %
1'
b1001 +
#446760000000
0!
0'
#446770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#446780000000
0!
0'
#446790000000
1!
1$
b1 %
1'
1*
b1 +
#446800000000
0!
0'
#446810000000
1!
b10 %
1'
b10 +
#446820000000
0!
0'
#446830000000
1!
b11 %
1'
b11 +
#446840000000
0!
0'
#446850000000
1!
b100 %
1'
b100 +
#446860000000
0!
0'
#446870000000
1!
b101 %
1'
b101 +
#446880000000
0!
0'
#446890000000
1!
0$
b110 %
1'
0*
b110 +
#446900000000
0!
0'
#446910000000
1!
b111 %
1'
b111 +
#446920000000
0!
0'
#446930000000
1!
b1000 %
1'
b1000 +
#446940000000
0!
0'
#446950000000
1!
b1001 %
1'
b1001 +
#446960000000
0!
0'
#446970000000
1!
b0 %
1'
b0 +
#446980000000
1"
1(
#446990000000
0!
0"
b100 &
0'
0(
b100 ,
#447000000000
1!
1$
b1 %
1'
1*
b1 +
#447010000000
0!
0'
#447020000000
1!
b10 %
1'
b10 +
#447030000000
0!
0'
#447040000000
1!
b11 %
1'
b11 +
#447050000000
0!
0'
#447060000000
1!
b100 %
1'
b100 +
#447070000000
0!
0'
#447080000000
1!
b101 %
1'
b101 +
#447090000000
0!
0'
#447100000000
1!
b110 %
1'
b110 +
#447110000000
0!
0'
#447120000000
1!
b111 %
1'
b111 +
#447130000000
0!
0'
#447140000000
1!
0$
b1000 %
1'
0*
b1000 +
#447150000000
0!
0'
#447160000000
1!
b1001 %
1'
b1001 +
#447170000000
0!
0'
#447180000000
1!
b0 %
1'
b0 +
#447190000000
0!
0'
#447200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#447210000000
0!
0'
#447220000000
1!
b10 %
1'
b10 +
#447230000000
0!
0'
#447240000000
1!
b11 %
1'
b11 +
#447250000000
0!
0'
#447260000000
1!
b100 %
1'
b100 +
#447270000000
0!
0'
#447280000000
1!
b101 %
1'
b101 +
#447290000000
0!
0'
#447300000000
1!
0$
b110 %
1'
0*
b110 +
#447310000000
0!
0'
#447320000000
1!
b111 %
1'
b111 +
#447330000000
0!
0'
#447340000000
1!
b1000 %
1'
b1000 +
#447350000000
0!
0'
#447360000000
1!
b1001 %
1'
b1001 +
#447370000000
0!
0'
#447380000000
1!
b0 %
1'
b0 +
#447390000000
0!
0'
#447400000000
1!
1$
b1 %
1'
1*
b1 +
#447410000000
1"
1(
#447420000000
0!
0"
b100 &
0'
0(
b100 ,
#447430000000
1!
b10 %
1'
b10 +
#447440000000
0!
0'
#447450000000
1!
b11 %
1'
b11 +
#447460000000
0!
0'
#447470000000
1!
b100 %
1'
b100 +
#447480000000
0!
0'
#447490000000
1!
b101 %
1'
b101 +
#447500000000
0!
0'
#447510000000
1!
b110 %
1'
b110 +
#447520000000
0!
0'
#447530000000
1!
b111 %
1'
b111 +
#447540000000
0!
0'
#447550000000
1!
0$
b1000 %
1'
0*
b1000 +
#447560000000
0!
0'
#447570000000
1!
b1001 %
1'
b1001 +
#447580000000
0!
0'
#447590000000
1!
b0 %
1'
b0 +
#447600000000
0!
0'
#447610000000
1!
1$
b1 %
1'
1*
b1 +
#447620000000
0!
0'
#447630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#447640000000
0!
0'
#447650000000
1!
b11 %
1'
b11 +
#447660000000
0!
0'
#447670000000
1!
b100 %
1'
b100 +
#447680000000
0!
0'
#447690000000
1!
b101 %
1'
b101 +
#447700000000
0!
0'
#447710000000
1!
0$
b110 %
1'
0*
b110 +
#447720000000
0!
0'
#447730000000
1!
b111 %
1'
b111 +
#447740000000
0!
0'
#447750000000
1!
b1000 %
1'
b1000 +
#447760000000
0!
0'
#447770000000
1!
b1001 %
1'
b1001 +
#447780000000
0!
0'
#447790000000
1!
b0 %
1'
b0 +
#447800000000
0!
0'
#447810000000
1!
1$
b1 %
1'
1*
b1 +
#447820000000
0!
0'
#447830000000
1!
b10 %
1'
b10 +
#447840000000
1"
1(
#447850000000
0!
0"
b100 &
0'
0(
b100 ,
#447860000000
1!
b11 %
1'
b11 +
#447870000000
0!
0'
#447880000000
1!
b100 %
1'
b100 +
#447890000000
0!
0'
#447900000000
1!
b101 %
1'
b101 +
#447910000000
0!
0'
#447920000000
1!
b110 %
1'
b110 +
#447930000000
0!
0'
#447940000000
1!
b111 %
1'
b111 +
#447950000000
0!
0'
#447960000000
1!
0$
b1000 %
1'
0*
b1000 +
#447970000000
0!
0'
#447980000000
1!
b1001 %
1'
b1001 +
#447990000000
0!
0'
#448000000000
1!
b0 %
1'
b0 +
#448010000000
0!
0'
#448020000000
1!
1$
b1 %
1'
1*
b1 +
#448030000000
0!
0'
#448040000000
1!
b10 %
1'
b10 +
#448050000000
0!
0'
#448060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#448070000000
0!
0'
#448080000000
1!
b100 %
1'
b100 +
#448090000000
0!
0'
#448100000000
1!
b101 %
1'
b101 +
#448110000000
0!
0'
#448120000000
1!
0$
b110 %
1'
0*
b110 +
#448130000000
0!
0'
#448140000000
1!
b111 %
1'
b111 +
#448150000000
0!
0'
#448160000000
1!
b1000 %
1'
b1000 +
#448170000000
0!
0'
#448180000000
1!
b1001 %
1'
b1001 +
#448190000000
0!
0'
#448200000000
1!
b0 %
1'
b0 +
#448210000000
0!
0'
#448220000000
1!
1$
b1 %
1'
1*
b1 +
#448230000000
0!
0'
#448240000000
1!
b10 %
1'
b10 +
#448250000000
0!
0'
#448260000000
1!
b11 %
1'
b11 +
#448270000000
1"
1(
#448280000000
0!
0"
b100 &
0'
0(
b100 ,
#448290000000
1!
b100 %
1'
b100 +
#448300000000
0!
0'
#448310000000
1!
b101 %
1'
b101 +
#448320000000
0!
0'
#448330000000
1!
b110 %
1'
b110 +
#448340000000
0!
0'
#448350000000
1!
b111 %
1'
b111 +
#448360000000
0!
0'
#448370000000
1!
0$
b1000 %
1'
0*
b1000 +
#448380000000
0!
0'
#448390000000
1!
b1001 %
1'
b1001 +
#448400000000
0!
0'
#448410000000
1!
b0 %
1'
b0 +
#448420000000
0!
0'
#448430000000
1!
1$
b1 %
1'
1*
b1 +
#448440000000
0!
0'
#448450000000
1!
b10 %
1'
b10 +
#448460000000
0!
0'
#448470000000
1!
b11 %
1'
b11 +
#448480000000
0!
0'
#448490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#448500000000
0!
0'
#448510000000
1!
b101 %
1'
b101 +
#448520000000
0!
0'
#448530000000
1!
0$
b110 %
1'
0*
b110 +
#448540000000
0!
0'
#448550000000
1!
b111 %
1'
b111 +
#448560000000
0!
0'
#448570000000
1!
b1000 %
1'
b1000 +
#448580000000
0!
0'
#448590000000
1!
b1001 %
1'
b1001 +
#448600000000
0!
0'
#448610000000
1!
b0 %
1'
b0 +
#448620000000
0!
0'
#448630000000
1!
1$
b1 %
1'
1*
b1 +
#448640000000
0!
0'
#448650000000
1!
b10 %
1'
b10 +
#448660000000
0!
0'
#448670000000
1!
b11 %
1'
b11 +
#448680000000
0!
0'
#448690000000
1!
b100 %
1'
b100 +
#448700000000
1"
1(
#448710000000
0!
0"
b100 &
0'
0(
b100 ,
#448720000000
1!
b101 %
1'
b101 +
#448730000000
0!
0'
#448740000000
1!
b110 %
1'
b110 +
#448750000000
0!
0'
#448760000000
1!
b111 %
1'
b111 +
#448770000000
0!
0'
#448780000000
1!
0$
b1000 %
1'
0*
b1000 +
#448790000000
0!
0'
#448800000000
1!
b1001 %
1'
b1001 +
#448810000000
0!
0'
#448820000000
1!
b0 %
1'
b0 +
#448830000000
0!
0'
#448840000000
1!
1$
b1 %
1'
1*
b1 +
#448850000000
0!
0'
#448860000000
1!
b10 %
1'
b10 +
#448870000000
0!
0'
#448880000000
1!
b11 %
1'
b11 +
#448890000000
0!
0'
#448900000000
1!
b100 %
1'
b100 +
#448910000000
0!
0'
#448920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#448930000000
0!
0'
#448940000000
1!
0$
b110 %
1'
0*
b110 +
#448950000000
0!
0'
#448960000000
1!
b111 %
1'
b111 +
#448970000000
0!
0'
#448980000000
1!
b1000 %
1'
b1000 +
#448990000000
0!
0'
#449000000000
1!
b1001 %
1'
b1001 +
#449010000000
0!
0'
#449020000000
1!
b0 %
1'
b0 +
#449030000000
0!
0'
#449040000000
1!
1$
b1 %
1'
1*
b1 +
#449050000000
0!
0'
#449060000000
1!
b10 %
1'
b10 +
#449070000000
0!
0'
#449080000000
1!
b11 %
1'
b11 +
#449090000000
0!
0'
#449100000000
1!
b100 %
1'
b100 +
#449110000000
0!
0'
#449120000000
1!
b101 %
1'
b101 +
#449130000000
1"
1(
#449140000000
0!
0"
b100 &
0'
0(
b100 ,
#449150000000
1!
b110 %
1'
b110 +
#449160000000
0!
0'
#449170000000
1!
b111 %
1'
b111 +
#449180000000
0!
0'
#449190000000
1!
0$
b1000 %
1'
0*
b1000 +
#449200000000
0!
0'
#449210000000
1!
b1001 %
1'
b1001 +
#449220000000
0!
0'
#449230000000
1!
b0 %
1'
b0 +
#449240000000
0!
0'
#449250000000
1!
1$
b1 %
1'
1*
b1 +
#449260000000
0!
0'
#449270000000
1!
b10 %
1'
b10 +
#449280000000
0!
0'
#449290000000
1!
b11 %
1'
b11 +
#449300000000
0!
0'
#449310000000
1!
b100 %
1'
b100 +
#449320000000
0!
0'
#449330000000
1!
b101 %
1'
b101 +
#449340000000
0!
0'
#449350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#449360000000
0!
0'
#449370000000
1!
b111 %
1'
b111 +
#449380000000
0!
0'
#449390000000
1!
b1000 %
1'
b1000 +
#449400000000
0!
0'
#449410000000
1!
b1001 %
1'
b1001 +
#449420000000
0!
0'
#449430000000
1!
b0 %
1'
b0 +
#449440000000
0!
0'
#449450000000
1!
1$
b1 %
1'
1*
b1 +
#449460000000
0!
0'
#449470000000
1!
b10 %
1'
b10 +
#449480000000
0!
0'
#449490000000
1!
b11 %
1'
b11 +
#449500000000
0!
0'
#449510000000
1!
b100 %
1'
b100 +
#449520000000
0!
0'
#449530000000
1!
b101 %
1'
b101 +
#449540000000
0!
0'
#449550000000
1!
0$
b110 %
1'
0*
b110 +
#449560000000
1"
1(
#449570000000
0!
0"
b100 &
0'
0(
b100 ,
#449580000000
1!
1$
b111 %
1'
1*
b111 +
#449590000000
0!
0'
#449600000000
1!
0$
b1000 %
1'
0*
b1000 +
#449610000000
0!
0'
#449620000000
1!
b1001 %
1'
b1001 +
#449630000000
0!
0'
#449640000000
1!
b0 %
1'
b0 +
#449650000000
0!
0'
#449660000000
1!
1$
b1 %
1'
1*
b1 +
#449670000000
0!
0'
#449680000000
1!
b10 %
1'
b10 +
#449690000000
0!
0'
#449700000000
1!
b11 %
1'
b11 +
#449710000000
0!
0'
#449720000000
1!
b100 %
1'
b100 +
#449730000000
0!
0'
#449740000000
1!
b101 %
1'
b101 +
#449750000000
0!
0'
#449760000000
1!
b110 %
1'
b110 +
#449770000000
0!
0'
#449780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#449790000000
0!
0'
#449800000000
1!
b1000 %
1'
b1000 +
#449810000000
0!
0'
#449820000000
1!
b1001 %
1'
b1001 +
#449830000000
0!
0'
#449840000000
1!
b0 %
1'
b0 +
#449850000000
0!
0'
#449860000000
1!
1$
b1 %
1'
1*
b1 +
#449870000000
0!
0'
#449880000000
1!
b10 %
1'
b10 +
#449890000000
0!
0'
#449900000000
1!
b11 %
1'
b11 +
#449910000000
0!
0'
#449920000000
1!
b100 %
1'
b100 +
#449930000000
0!
0'
#449940000000
1!
b101 %
1'
b101 +
#449950000000
0!
0'
#449960000000
1!
0$
b110 %
1'
0*
b110 +
#449970000000
0!
0'
#449980000000
1!
b111 %
1'
b111 +
#449990000000
1"
1(
#450000000000
0!
0"
b100 &
0'
0(
b100 ,
#450010000000
1!
b1000 %
1'
b1000 +
#450020000000
0!
0'
#450030000000
1!
b1001 %
1'
b1001 +
#450040000000
0!
0'
#450050000000
1!
b0 %
1'
b0 +
#450060000000
0!
0'
#450070000000
1!
1$
b1 %
1'
1*
b1 +
#450080000000
0!
0'
#450090000000
1!
b10 %
1'
b10 +
#450100000000
0!
0'
#450110000000
1!
b11 %
1'
b11 +
#450120000000
0!
0'
#450130000000
1!
b100 %
1'
b100 +
#450140000000
0!
0'
#450150000000
1!
b101 %
1'
b101 +
#450160000000
0!
0'
#450170000000
1!
b110 %
1'
b110 +
#450180000000
0!
0'
#450190000000
1!
b111 %
1'
b111 +
#450200000000
0!
0'
#450210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#450220000000
0!
0'
#450230000000
1!
b1001 %
1'
b1001 +
#450240000000
0!
0'
#450250000000
1!
b0 %
1'
b0 +
#450260000000
0!
0'
#450270000000
1!
1$
b1 %
1'
1*
b1 +
#450280000000
0!
0'
#450290000000
1!
b10 %
1'
b10 +
#450300000000
0!
0'
#450310000000
1!
b11 %
1'
b11 +
#450320000000
0!
0'
#450330000000
1!
b100 %
1'
b100 +
#450340000000
0!
0'
#450350000000
1!
b101 %
1'
b101 +
#450360000000
0!
0'
#450370000000
1!
0$
b110 %
1'
0*
b110 +
#450380000000
0!
0'
#450390000000
1!
b111 %
1'
b111 +
#450400000000
0!
0'
#450410000000
1!
b1000 %
1'
b1000 +
#450420000000
1"
1(
#450430000000
0!
0"
b100 &
0'
0(
b100 ,
#450440000000
1!
b1001 %
1'
b1001 +
#450450000000
0!
0'
#450460000000
1!
b0 %
1'
b0 +
#450470000000
0!
0'
#450480000000
1!
1$
b1 %
1'
1*
b1 +
#450490000000
0!
0'
#450500000000
1!
b10 %
1'
b10 +
#450510000000
0!
0'
#450520000000
1!
b11 %
1'
b11 +
#450530000000
0!
0'
#450540000000
1!
b100 %
1'
b100 +
#450550000000
0!
0'
#450560000000
1!
b101 %
1'
b101 +
#450570000000
0!
0'
#450580000000
1!
b110 %
1'
b110 +
#450590000000
0!
0'
#450600000000
1!
b111 %
1'
b111 +
#450610000000
0!
0'
#450620000000
1!
0$
b1000 %
1'
0*
b1000 +
#450630000000
0!
0'
#450640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#450650000000
0!
0'
#450660000000
1!
b0 %
1'
b0 +
#450670000000
0!
0'
#450680000000
1!
1$
b1 %
1'
1*
b1 +
#450690000000
0!
0'
#450700000000
1!
b10 %
1'
b10 +
#450710000000
0!
0'
#450720000000
1!
b11 %
1'
b11 +
#450730000000
0!
0'
#450740000000
1!
b100 %
1'
b100 +
#450750000000
0!
0'
#450760000000
1!
b101 %
1'
b101 +
#450770000000
0!
0'
#450780000000
1!
0$
b110 %
1'
0*
b110 +
#450790000000
0!
0'
#450800000000
1!
b111 %
1'
b111 +
#450810000000
0!
0'
#450820000000
1!
b1000 %
1'
b1000 +
#450830000000
0!
0'
#450840000000
1!
b1001 %
1'
b1001 +
#450850000000
1"
1(
#450860000000
0!
0"
b100 &
0'
0(
b100 ,
#450870000000
1!
b0 %
1'
b0 +
#450880000000
0!
0'
#450890000000
1!
1$
b1 %
1'
1*
b1 +
#450900000000
0!
0'
#450910000000
1!
b10 %
1'
b10 +
#450920000000
0!
0'
#450930000000
1!
b11 %
1'
b11 +
#450940000000
0!
0'
#450950000000
1!
b100 %
1'
b100 +
#450960000000
0!
0'
#450970000000
1!
b101 %
1'
b101 +
#450980000000
0!
0'
#450990000000
1!
b110 %
1'
b110 +
#451000000000
0!
0'
#451010000000
1!
b111 %
1'
b111 +
#451020000000
0!
0'
#451030000000
1!
0$
b1000 %
1'
0*
b1000 +
#451040000000
0!
0'
#451050000000
1!
b1001 %
1'
b1001 +
#451060000000
0!
0'
#451070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#451080000000
0!
0'
#451090000000
1!
1$
b1 %
1'
1*
b1 +
#451100000000
0!
0'
#451110000000
1!
b10 %
1'
b10 +
#451120000000
0!
0'
#451130000000
1!
b11 %
1'
b11 +
#451140000000
0!
0'
#451150000000
1!
b100 %
1'
b100 +
#451160000000
0!
0'
#451170000000
1!
b101 %
1'
b101 +
#451180000000
0!
0'
#451190000000
1!
0$
b110 %
1'
0*
b110 +
#451200000000
0!
0'
#451210000000
1!
b111 %
1'
b111 +
#451220000000
0!
0'
#451230000000
1!
b1000 %
1'
b1000 +
#451240000000
0!
0'
#451250000000
1!
b1001 %
1'
b1001 +
#451260000000
0!
0'
#451270000000
1!
b0 %
1'
b0 +
#451280000000
1"
1(
#451290000000
0!
0"
b100 &
0'
0(
b100 ,
#451300000000
1!
1$
b1 %
1'
1*
b1 +
#451310000000
0!
0'
#451320000000
1!
b10 %
1'
b10 +
#451330000000
0!
0'
#451340000000
1!
b11 %
1'
b11 +
#451350000000
0!
0'
#451360000000
1!
b100 %
1'
b100 +
#451370000000
0!
0'
#451380000000
1!
b101 %
1'
b101 +
#451390000000
0!
0'
#451400000000
1!
b110 %
1'
b110 +
#451410000000
0!
0'
#451420000000
1!
b111 %
1'
b111 +
#451430000000
0!
0'
#451440000000
1!
0$
b1000 %
1'
0*
b1000 +
#451450000000
0!
0'
#451460000000
1!
b1001 %
1'
b1001 +
#451470000000
0!
0'
#451480000000
1!
b0 %
1'
b0 +
#451490000000
0!
0'
#451500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#451510000000
0!
0'
#451520000000
1!
b10 %
1'
b10 +
#451530000000
0!
0'
#451540000000
1!
b11 %
1'
b11 +
#451550000000
0!
0'
#451560000000
1!
b100 %
1'
b100 +
#451570000000
0!
0'
#451580000000
1!
b101 %
1'
b101 +
#451590000000
0!
0'
#451600000000
1!
0$
b110 %
1'
0*
b110 +
#451610000000
0!
0'
#451620000000
1!
b111 %
1'
b111 +
#451630000000
0!
0'
#451640000000
1!
b1000 %
1'
b1000 +
#451650000000
0!
0'
#451660000000
1!
b1001 %
1'
b1001 +
#451670000000
0!
0'
#451680000000
1!
b0 %
1'
b0 +
#451690000000
0!
0'
#451700000000
1!
1$
b1 %
1'
1*
b1 +
#451710000000
1"
1(
#451720000000
0!
0"
b100 &
0'
0(
b100 ,
#451730000000
1!
b10 %
1'
b10 +
#451740000000
0!
0'
#451750000000
1!
b11 %
1'
b11 +
#451760000000
0!
0'
#451770000000
1!
b100 %
1'
b100 +
#451780000000
0!
0'
#451790000000
1!
b101 %
1'
b101 +
#451800000000
0!
0'
#451810000000
1!
b110 %
1'
b110 +
#451820000000
0!
0'
#451830000000
1!
b111 %
1'
b111 +
#451840000000
0!
0'
#451850000000
1!
0$
b1000 %
1'
0*
b1000 +
#451860000000
0!
0'
#451870000000
1!
b1001 %
1'
b1001 +
#451880000000
0!
0'
#451890000000
1!
b0 %
1'
b0 +
#451900000000
0!
0'
#451910000000
1!
1$
b1 %
1'
1*
b1 +
#451920000000
0!
0'
#451930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#451940000000
0!
0'
#451950000000
1!
b11 %
1'
b11 +
#451960000000
0!
0'
#451970000000
1!
b100 %
1'
b100 +
#451980000000
0!
0'
#451990000000
1!
b101 %
1'
b101 +
#452000000000
0!
0'
#452010000000
1!
0$
b110 %
1'
0*
b110 +
#452020000000
0!
0'
#452030000000
1!
b111 %
1'
b111 +
#452040000000
0!
0'
#452050000000
1!
b1000 %
1'
b1000 +
#452060000000
0!
0'
#452070000000
1!
b1001 %
1'
b1001 +
#452080000000
0!
0'
#452090000000
1!
b0 %
1'
b0 +
#452100000000
0!
0'
#452110000000
1!
1$
b1 %
1'
1*
b1 +
#452120000000
0!
0'
#452130000000
1!
b10 %
1'
b10 +
#452140000000
1"
1(
#452150000000
0!
0"
b100 &
0'
0(
b100 ,
#452160000000
1!
b11 %
1'
b11 +
#452170000000
0!
0'
#452180000000
1!
b100 %
1'
b100 +
#452190000000
0!
0'
#452200000000
1!
b101 %
1'
b101 +
#452210000000
0!
0'
#452220000000
1!
b110 %
1'
b110 +
#452230000000
0!
0'
#452240000000
1!
b111 %
1'
b111 +
#452250000000
0!
0'
#452260000000
1!
0$
b1000 %
1'
0*
b1000 +
#452270000000
0!
0'
#452280000000
1!
b1001 %
1'
b1001 +
#452290000000
0!
0'
#452300000000
1!
b0 %
1'
b0 +
#452310000000
0!
0'
#452320000000
1!
1$
b1 %
1'
1*
b1 +
#452330000000
0!
0'
#452340000000
1!
b10 %
1'
b10 +
#452350000000
0!
0'
#452360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#452370000000
0!
0'
#452380000000
1!
b100 %
1'
b100 +
#452390000000
0!
0'
#452400000000
1!
b101 %
1'
b101 +
#452410000000
0!
0'
#452420000000
1!
0$
b110 %
1'
0*
b110 +
#452430000000
0!
0'
#452440000000
1!
b111 %
1'
b111 +
#452450000000
0!
0'
#452460000000
1!
b1000 %
1'
b1000 +
#452470000000
0!
0'
#452480000000
1!
b1001 %
1'
b1001 +
#452490000000
0!
0'
#452500000000
1!
b0 %
1'
b0 +
#452510000000
0!
0'
#452520000000
1!
1$
b1 %
1'
1*
b1 +
#452530000000
0!
0'
#452540000000
1!
b10 %
1'
b10 +
#452550000000
0!
0'
#452560000000
1!
b11 %
1'
b11 +
#452570000000
1"
1(
#452580000000
0!
0"
b100 &
0'
0(
b100 ,
#452590000000
1!
b100 %
1'
b100 +
#452600000000
0!
0'
#452610000000
1!
b101 %
1'
b101 +
#452620000000
0!
0'
#452630000000
1!
b110 %
1'
b110 +
#452640000000
0!
0'
#452650000000
1!
b111 %
1'
b111 +
#452660000000
0!
0'
#452670000000
1!
0$
b1000 %
1'
0*
b1000 +
#452680000000
0!
0'
#452690000000
1!
b1001 %
1'
b1001 +
#452700000000
0!
0'
#452710000000
1!
b0 %
1'
b0 +
#452720000000
0!
0'
#452730000000
1!
1$
b1 %
1'
1*
b1 +
#452740000000
0!
0'
#452750000000
1!
b10 %
1'
b10 +
#452760000000
0!
0'
#452770000000
1!
b11 %
1'
b11 +
#452780000000
0!
0'
#452790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#452800000000
0!
0'
#452810000000
1!
b101 %
1'
b101 +
#452820000000
0!
0'
#452830000000
1!
0$
b110 %
1'
0*
b110 +
#452840000000
0!
0'
#452850000000
1!
b111 %
1'
b111 +
#452860000000
0!
0'
#452870000000
1!
b1000 %
1'
b1000 +
#452880000000
0!
0'
#452890000000
1!
b1001 %
1'
b1001 +
#452900000000
0!
0'
#452910000000
1!
b0 %
1'
b0 +
#452920000000
0!
0'
#452930000000
1!
1$
b1 %
1'
1*
b1 +
#452940000000
0!
0'
#452950000000
1!
b10 %
1'
b10 +
#452960000000
0!
0'
#452970000000
1!
b11 %
1'
b11 +
#452980000000
0!
0'
#452990000000
1!
b100 %
1'
b100 +
#453000000000
1"
1(
#453010000000
0!
0"
b100 &
0'
0(
b100 ,
#453020000000
1!
b101 %
1'
b101 +
#453030000000
0!
0'
#453040000000
1!
b110 %
1'
b110 +
#453050000000
0!
0'
#453060000000
1!
b111 %
1'
b111 +
#453070000000
0!
0'
#453080000000
1!
0$
b1000 %
1'
0*
b1000 +
#453090000000
0!
0'
#453100000000
1!
b1001 %
1'
b1001 +
#453110000000
0!
0'
#453120000000
1!
b0 %
1'
b0 +
#453130000000
0!
0'
#453140000000
1!
1$
b1 %
1'
1*
b1 +
#453150000000
0!
0'
#453160000000
1!
b10 %
1'
b10 +
#453170000000
0!
0'
#453180000000
1!
b11 %
1'
b11 +
#453190000000
0!
0'
#453200000000
1!
b100 %
1'
b100 +
#453210000000
0!
0'
#453220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#453230000000
0!
0'
#453240000000
1!
0$
b110 %
1'
0*
b110 +
#453250000000
0!
0'
#453260000000
1!
b111 %
1'
b111 +
#453270000000
0!
0'
#453280000000
1!
b1000 %
1'
b1000 +
#453290000000
0!
0'
#453300000000
1!
b1001 %
1'
b1001 +
#453310000000
0!
0'
#453320000000
1!
b0 %
1'
b0 +
#453330000000
0!
0'
#453340000000
1!
1$
b1 %
1'
1*
b1 +
#453350000000
0!
0'
#453360000000
1!
b10 %
1'
b10 +
#453370000000
0!
0'
#453380000000
1!
b11 %
1'
b11 +
#453390000000
0!
0'
#453400000000
1!
b100 %
1'
b100 +
#453410000000
0!
0'
#453420000000
1!
b101 %
1'
b101 +
#453430000000
1"
1(
#453440000000
0!
0"
b100 &
0'
0(
b100 ,
#453450000000
1!
b110 %
1'
b110 +
#453460000000
0!
0'
#453470000000
1!
b111 %
1'
b111 +
#453480000000
0!
0'
#453490000000
1!
0$
b1000 %
1'
0*
b1000 +
#453500000000
0!
0'
#453510000000
1!
b1001 %
1'
b1001 +
#453520000000
0!
0'
#453530000000
1!
b0 %
1'
b0 +
#453540000000
0!
0'
#453550000000
1!
1$
b1 %
1'
1*
b1 +
#453560000000
0!
0'
#453570000000
1!
b10 %
1'
b10 +
#453580000000
0!
0'
#453590000000
1!
b11 %
1'
b11 +
#453600000000
0!
0'
#453610000000
1!
b100 %
1'
b100 +
#453620000000
0!
0'
#453630000000
1!
b101 %
1'
b101 +
#453640000000
0!
0'
#453650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#453660000000
0!
0'
#453670000000
1!
b111 %
1'
b111 +
#453680000000
0!
0'
#453690000000
1!
b1000 %
1'
b1000 +
#453700000000
0!
0'
#453710000000
1!
b1001 %
1'
b1001 +
#453720000000
0!
0'
#453730000000
1!
b0 %
1'
b0 +
#453740000000
0!
0'
#453750000000
1!
1$
b1 %
1'
1*
b1 +
#453760000000
0!
0'
#453770000000
1!
b10 %
1'
b10 +
#453780000000
0!
0'
#453790000000
1!
b11 %
1'
b11 +
#453800000000
0!
0'
#453810000000
1!
b100 %
1'
b100 +
#453820000000
0!
0'
#453830000000
1!
b101 %
1'
b101 +
#453840000000
0!
0'
#453850000000
1!
0$
b110 %
1'
0*
b110 +
#453860000000
1"
1(
#453870000000
0!
0"
b100 &
0'
0(
b100 ,
#453880000000
1!
1$
b111 %
1'
1*
b111 +
#453890000000
0!
0'
#453900000000
1!
0$
b1000 %
1'
0*
b1000 +
#453910000000
0!
0'
#453920000000
1!
b1001 %
1'
b1001 +
#453930000000
0!
0'
#453940000000
1!
b0 %
1'
b0 +
#453950000000
0!
0'
#453960000000
1!
1$
b1 %
1'
1*
b1 +
#453970000000
0!
0'
#453980000000
1!
b10 %
1'
b10 +
#453990000000
0!
0'
#454000000000
1!
b11 %
1'
b11 +
#454010000000
0!
0'
#454020000000
1!
b100 %
1'
b100 +
#454030000000
0!
0'
#454040000000
1!
b101 %
1'
b101 +
#454050000000
0!
0'
#454060000000
1!
b110 %
1'
b110 +
#454070000000
0!
0'
#454080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#454090000000
0!
0'
#454100000000
1!
b1000 %
1'
b1000 +
#454110000000
0!
0'
#454120000000
1!
b1001 %
1'
b1001 +
#454130000000
0!
0'
#454140000000
1!
b0 %
1'
b0 +
#454150000000
0!
0'
#454160000000
1!
1$
b1 %
1'
1*
b1 +
#454170000000
0!
0'
#454180000000
1!
b10 %
1'
b10 +
#454190000000
0!
0'
#454200000000
1!
b11 %
1'
b11 +
#454210000000
0!
0'
#454220000000
1!
b100 %
1'
b100 +
#454230000000
0!
0'
#454240000000
1!
b101 %
1'
b101 +
#454250000000
0!
0'
#454260000000
1!
0$
b110 %
1'
0*
b110 +
#454270000000
0!
0'
#454280000000
1!
b111 %
1'
b111 +
#454290000000
1"
1(
#454300000000
0!
0"
b100 &
0'
0(
b100 ,
#454310000000
1!
b1000 %
1'
b1000 +
#454320000000
0!
0'
#454330000000
1!
b1001 %
1'
b1001 +
#454340000000
0!
0'
#454350000000
1!
b0 %
1'
b0 +
#454360000000
0!
0'
#454370000000
1!
1$
b1 %
1'
1*
b1 +
#454380000000
0!
0'
#454390000000
1!
b10 %
1'
b10 +
#454400000000
0!
0'
#454410000000
1!
b11 %
1'
b11 +
#454420000000
0!
0'
#454430000000
1!
b100 %
1'
b100 +
#454440000000
0!
0'
#454450000000
1!
b101 %
1'
b101 +
#454460000000
0!
0'
#454470000000
1!
b110 %
1'
b110 +
#454480000000
0!
0'
#454490000000
1!
b111 %
1'
b111 +
#454500000000
0!
0'
#454510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#454520000000
0!
0'
#454530000000
1!
b1001 %
1'
b1001 +
#454540000000
0!
0'
#454550000000
1!
b0 %
1'
b0 +
#454560000000
0!
0'
#454570000000
1!
1$
b1 %
1'
1*
b1 +
#454580000000
0!
0'
#454590000000
1!
b10 %
1'
b10 +
#454600000000
0!
0'
#454610000000
1!
b11 %
1'
b11 +
#454620000000
0!
0'
#454630000000
1!
b100 %
1'
b100 +
#454640000000
0!
0'
#454650000000
1!
b101 %
1'
b101 +
#454660000000
0!
0'
#454670000000
1!
0$
b110 %
1'
0*
b110 +
#454680000000
0!
0'
#454690000000
1!
b111 %
1'
b111 +
#454700000000
0!
0'
#454710000000
1!
b1000 %
1'
b1000 +
#454720000000
1"
1(
#454730000000
0!
0"
b100 &
0'
0(
b100 ,
#454740000000
1!
b1001 %
1'
b1001 +
#454750000000
0!
0'
#454760000000
1!
b0 %
1'
b0 +
#454770000000
0!
0'
#454780000000
1!
1$
b1 %
1'
1*
b1 +
#454790000000
0!
0'
#454800000000
1!
b10 %
1'
b10 +
#454810000000
0!
0'
#454820000000
1!
b11 %
1'
b11 +
#454830000000
0!
0'
#454840000000
1!
b100 %
1'
b100 +
#454850000000
0!
0'
#454860000000
1!
b101 %
1'
b101 +
#454870000000
0!
0'
#454880000000
1!
b110 %
1'
b110 +
#454890000000
0!
0'
#454900000000
1!
b111 %
1'
b111 +
#454910000000
0!
0'
#454920000000
1!
0$
b1000 %
1'
0*
b1000 +
#454930000000
0!
0'
#454940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#454950000000
0!
0'
#454960000000
1!
b0 %
1'
b0 +
#454970000000
0!
0'
#454980000000
1!
1$
b1 %
1'
1*
b1 +
#454990000000
0!
0'
#455000000000
1!
b10 %
1'
b10 +
#455010000000
0!
0'
#455020000000
1!
b11 %
1'
b11 +
#455030000000
0!
0'
#455040000000
1!
b100 %
1'
b100 +
#455050000000
0!
0'
#455060000000
1!
b101 %
1'
b101 +
#455070000000
0!
0'
#455080000000
1!
0$
b110 %
1'
0*
b110 +
#455090000000
0!
0'
#455100000000
1!
b111 %
1'
b111 +
#455110000000
0!
0'
#455120000000
1!
b1000 %
1'
b1000 +
#455130000000
0!
0'
#455140000000
1!
b1001 %
1'
b1001 +
#455150000000
1"
1(
#455160000000
0!
0"
b100 &
0'
0(
b100 ,
#455170000000
1!
b0 %
1'
b0 +
#455180000000
0!
0'
#455190000000
1!
1$
b1 %
1'
1*
b1 +
#455200000000
0!
0'
#455210000000
1!
b10 %
1'
b10 +
#455220000000
0!
0'
#455230000000
1!
b11 %
1'
b11 +
#455240000000
0!
0'
#455250000000
1!
b100 %
1'
b100 +
#455260000000
0!
0'
#455270000000
1!
b101 %
1'
b101 +
#455280000000
0!
0'
#455290000000
1!
b110 %
1'
b110 +
#455300000000
0!
0'
#455310000000
1!
b111 %
1'
b111 +
#455320000000
0!
0'
#455330000000
1!
0$
b1000 %
1'
0*
b1000 +
#455340000000
0!
0'
#455350000000
1!
b1001 %
1'
b1001 +
#455360000000
0!
0'
#455370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#455380000000
0!
0'
#455390000000
1!
1$
b1 %
1'
1*
b1 +
#455400000000
0!
0'
#455410000000
1!
b10 %
1'
b10 +
#455420000000
0!
0'
#455430000000
1!
b11 %
1'
b11 +
#455440000000
0!
0'
#455450000000
1!
b100 %
1'
b100 +
#455460000000
0!
0'
#455470000000
1!
b101 %
1'
b101 +
#455480000000
0!
0'
#455490000000
1!
0$
b110 %
1'
0*
b110 +
#455500000000
0!
0'
#455510000000
1!
b111 %
1'
b111 +
#455520000000
0!
0'
#455530000000
1!
b1000 %
1'
b1000 +
#455540000000
0!
0'
#455550000000
1!
b1001 %
1'
b1001 +
#455560000000
0!
0'
#455570000000
1!
b0 %
1'
b0 +
#455580000000
1"
1(
#455590000000
0!
0"
b100 &
0'
0(
b100 ,
#455600000000
1!
1$
b1 %
1'
1*
b1 +
#455610000000
0!
0'
#455620000000
1!
b10 %
1'
b10 +
#455630000000
0!
0'
#455640000000
1!
b11 %
1'
b11 +
#455650000000
0!
0'
#455660000000
1!
b100 %
1'
b100 +
#455670000000
0!
0'
#455680000000
1!
b101 %
1'
b101 +
#455690000000
0!
0'
#455700000000
1!
b110 %
1'
b110 +
#455710000000
0!
0'
#455720000000
1!
b111 %
1'
b111 +
#455730000000
0!
0'
#455740000000
1!
0$
b1000 %
1'
0*
b1000 +
#455750000000
0!
0'
#455760000000
1!
b1001 %
1'
b1001 +
#455770000000
0!
0'
#455780000000
1!
b0 %
1'
b0 +
#455790000000
0!
0'
#455800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#455810000000
0!
0'
#455820000000
1!
b10 %
1'
b10 +
#455830000000
0!
0'
#455840000000
1!
b11 %
1'
b11 +
#455850000000
0!
0'
#455860000000
1!
b100 %
1'
b100 +
#455870000000
0!
0'
#455880000000
1!
b101 %
1'
b101 +
#455890000000
0!
0'
#455900000000
1!
0$
b110 %
1'
0*
b110 +
#455910000000
0!
0'
#455920000000
1!
b111 %
1'
b111 +
#455930000000
0!
0'
#455940000000
1!
b1000 %
1'
b1000 +
#455950000000
0!
0'
#455960000000
1!
b1001 %
1'
b1001 +
#455970000000
0!
0'
#455980000000
1!
b0 %
1'
b0 +
#455990000000
0!
0'
#456000000000
1!
1$
b1 %
1'
1*
b1 +
#456010000000
1"
1(
#456020000000
0!
0"
b100 &
0'
0(
b100 ,
#456030000000
1!
b10 %
1'
b10 +
#456040000000
0!
0'
#456050000000
1!
b11 %
1'
b11 +
#456060000000
0!
0'
#456070000000
1!
b100 %
1'
b100 +
#456080000000
0!
0'
#456090000000
1!
b101 %
1'
b101 +
#456100000000
0!
0'
#456110000000
1!
b110 %
1'
b110 +
#456120000000
0!
0'
#456130000000
1!
b111 %
1'
b111 +
#456140000000
0!
0'
#456150000000
1!
0$
b1000 %
1'
0*
b1000 +
#456160000000
0!
0'
#456170000000
1!
b1001 %
1'
b1001 +
#456180000000
0!
0'
#456190000000
1!
b0 %
1'
b0 +
#456200000000
0!
0'
#456210000000
1!
1$
b1 %
1'
1*
b1 +
#456220000000
0!
0'
#456230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#456240000000
0!
0'
#456250000000
1!
b11 %
1'
b11 +
#456260000000
0!
0'
#456270000000
1!
b100 %
1'
b100 +
#456280000000
0!
0'
#456290000000
1!
b101 %
1'
b101 +
#456300000000
0!
0'
#456310000000
1!
0$
b110 %
1'
0*
b110 +
#456320000000
0!
0'
#456330000000
1!
b111 %
1'
b111 +
#456340000000
0!
0'
#456350000000
1!
b1000 %
1'
b1000 +
#456360000000
0!
0'
#456370000000
1!
b1001 %
1'
b1001 +
#456380000000
0!
0'
#456390000000
1!
b0 %
1'
b0 +
#456400000000
0!
0'
#456410000000
1!
1$
b1 %
1'
1*
b1 +
#456420000000
0!
0'
#456430000000
1!
b10 %
1'
b10 +
#456440000000
1"
1(
#456450000000
0!
0"
b100 &
0'
0(
b100 ,
#456460000000
1!
b11 %
1'
b11 +
#456470000000
0!
0'
#456480000000
1!
b100 %
1'
b100 +
#456490000000
0!
0'
#456500000000
1!
b101 %
1'
b101 +
#456510000000
0!
0'
#456520000000
1!
b110 %
1'
b110 +
#456530000000
0!
0'
#456540000000
1!
b111 %
1'
b111 +
#456550000000
0!
0'
#456560000000
1!
0$
b1000 %
1'
0*
b1000 +
#456570000000
0!
0'
#456580000000
1!
b1001 %
1'
b1001 +
#456590000000
0!
0'
#456600000000
1!
b0 %
1'
b0 +
#456610000000
0!
0'
#456620000000
1!
1$
b1 %
1'
1*
b1 +
#456630000000
0!
0'
#456640000000
1!
b10 %
1'
b10 +
#456650000000
0!
0'
#456660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#456670000000
0!
0'
#456680000000
1!
b100 %
1'
b100 +
#456690000000
0!
0'
#456700000000
1!
b101 %
1'
b101 +
#456710000000
0!
0'
#456720000000
1!
0$
b110 %
1'
0*
b110 +
#456730000000
0!
0'
#456740000000
1!
b111 %
1'
b111 +
#456750000000
0!
0'
#456760000000
1!
b1000 %
1'
b1000 +
#456770000000
0!
0'
#456780000000
1!
b1001 %
1'
b1001 +
#456790000000
0!
0'
#456800000000
1!
b0 %
1'
b0 +
#456810000000
0!
0'
#456820000000
1!
1$
b1 %
1'
1*
b1 +
#456830000000
0!
0'
#456840000000
1!
b10 %
1'
b10 +
#456850000000
0!
0'
#456860000000
1!
b11 %
1'
b11 +
#456870000000
1"
1(
#456880000000
0!
0"
b100 &
0'
0(
b100 ,
#456890000000
1!
b100 %
1'
b100 +
#456900000000
0!
0'
#456910000000
1!
b101 %
1'
b101 +
#456920000000
0!
0'
#456930000000
1!
b110 %
1'
b110 +
#456940000000
0!
0'
#456950000000
1!
b111 %
1'
b111 +
#456960000000
0!
0'
#456970000000
1!
0$
b1000 %
1'
0*
b1000 +
#456980000000
0!
0'
#456990000000
1!
b1001 %
1'
b1001 +
#457000000000
0!
0'
#457010000000
1!
b0 %
1'
b0 +
#457020000000
0!
0'
#457030000000
1!
1$
b1 %
1'
1*
b1 +
#457040000000
0!
0'
#457050000000
1!
b10 %
1'
b10 +
#457060000000
0!
0'
#457070000000
1!
b11 %
1'
b11 +
#457080000000
0!
0'
#457090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#457100000000
0!
0'
#457110000000
1!
b101 %
1'
b101 +
#457120000000
0!
0'
#457130000000
1!
0$
b110 %
1'
0*
b110 +
#457140000000
0!
0'
#457150000000
1!
b111 %
1'
b111 +
#457160000000
0!
0'
#457170000000
1!
b1000 %
1'
b1000 +
#457180000000
0!
0'
#457190000000
1!
b1001 %
1'
b1001 +
#457200000000
0!
0'
#457210000000
1!
b0 %
1'
b0 +
#457220000000
0!
0'
#457230000000
1!
1$
b1 %
1'
1*
b1 +
#457240000000
0!
0'
#457250000000
1!
b10 %
1'
b10 +
#457260000000
0!
0'
#457270000000
1!
b11 %
1'
b11 +
#457280000000
0!
0'
#457290000000
1!
b100 %
1'
b100 +
#457300000000
1"
1(
#457310000000
0!
0"
b100 &
0'
0(
b100 ,
#457320000000
1!
b101 %
1'
b101 +
#457330000000
0!
0'
#457340000000
1!
b110 %
1'
b110 +
#457350000000
0!
0'
#457360000000
1!
b111 %
1'
b111 +
#457370000000
0!
0'
#457380000000
1!
0$
b1000 %
1'
0*
b1000 +
#457390000000
0!
0'
#457400000000
1!
b1001 %
1'
b1001 +
#457410000000
0!
0'
#457420000000
1!
b0 %
1'
b0 +
#457430000000
0!
0'
#457440000000
1!
1$
b1 %
1'
1*
b1 +
#457450000000
0!
0'
#457460000000
1!
b10 %
1'
b10 +
#457470000000
0!
0'
#457480000000
1!
b11 %
1'
b11 +
#457490000000
0!
0'
#457500000000
1!
b100 %
1'
b100 +
#457510000000
0!
0'
#457520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#457530000000
0!
0'
#457540000000
1!
0$
b110 %
1'
0*
b110 +
#457550000000
0!
0'
#457560000000
1!
b111 %
1'
b111 +
#457570000000
0!
0'
#457580000000
1!
b1000 %
1'
b1000 +
#457590000000
0!
0'
#457600000000
1!
b1001 %
1'
b1001 +
#457610000000
0!
0'
#457620000000
1!
b0 %
1'
b0 +
#457630000000
0!
0'
#457640000000
1!
1$
b1 %
1'
1*
b1 +
#457650000000
0!
0'
#457660000000
1!
b10 %
1'
b10 +
#457670000000
0!
0'
#457680000000
1!
b11 %
1'
b11 +
#457690000000
0!
0'
#457700000000
1!
b100 %
1'
b100 +
#457710000000
0!
0'
#457720000000
1!
b101 %
1'
b101 +
#457730000000
1"
1(
#457740000000
0!
0"
b100 &
0'
0(
b100 ,
#457750000000
1!
b110 %
1'
b110 +
#457760000000
0!
0'
#457770000000
1!
b111 %
1'
b111 +
#457780000000
0!
0'
#457790000000
1!
0$
b1000 %
1'
0*
b1000 +
#457800000000
0!
0'
#457810000000
1!
b1001 %
1'
b1001 +
#457820000000
0!
0'
#457830000000
1!
b0 %
1'
b0 +
#457840000000
0!
0'
#457850000000
1!
1$
b1 %
1'
1*
b1 +
#457860000000
0!
0'
#457870000000
1!
b10 %
1'
b10 +
#457880000000
0!
0'
#457890000000
1!
b11 %
1'
b11 +
#457900000000
0!
0'
#457910000000
1!
b100 %
1'
b100 +
#457920000000
0!
0'
#457930000000
1!
b101 %
1'
b101 +
#457940000000
0!
0'
#457950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#457960000000
0!
0'
#457970000000
1!
b111 %
1'
b111 +
#457980000000
0!
0'
#457990000000
1!
b1000 %
1'
b1000 +
#458000000000
0!
0'
#458010000000
1!
b1001 %
1'
b1001 +
#458020000000
0!
0'
#458030000000
1!
b0 %
1'
b0 +
#458040000000
0!
0'
#458050000000
1!
1$
b1 %
1'
1*
b1 +
#458060000000
0!
0'
#458070000000
1!
b10 %
1'
b10 +
#458080000000
0!
0'
#458090000000
1!
b11 %
1'
b11 +
#458100000000
0!
0'
#458110000000
1!
b100 %
1'
b100 +
#458120000000
0!
0'
#458130000000
1!
b101 %
1'
b101 +
#458140000000
0!
0'
#458150000000
1!
0$
b110 %
1'
0*
b110 +
#458160000000
1"
1(
#458170000000
0!
0"
b100 &
0'
0(
b100 ,
#458180000000
1!
1$
b111 %
1'
1*
b111 +
#458190000000
0!
0'
#458200000000
1!
0$
b1000 %
1'
0*
b1000 +
#458210000000
0!
0'
#458220000000
1!
b1001 %
1'
b1001 +
#458230000000
0!
0'
#458240000000
1!
b0 %
1'
b0 +
#458250000000
0!
0'
#458260000000
1!
1$
b1 %
1'
1*
b1 +
#458270000000
0!
0'
#458280000000
1!
b10 %
1'
b10 +
#458290000000
0!
0'
#458300000000
1!
b11 %
1'
b11 +
#458310000000
0!
0'
#458320000000
1!
b100 %
1'
b100 +
#458330000000
0!
0'
#458340000000
1!
b101 %
1'
b101 +
#458350000000
0!
0'
#458360000000
1!
b110 %
1'
b110 +
#458370000000
0!
0'
#458380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#458390000000
0!
0'
#458400000000
1!
b1000 %
1'
b1000 +
#458410000000
0!
0'
#458420000000
1!
b1001 %
1'
b1001 +
#458430000000
0!
0'
#458440000000
1!
b0 %
1'
b0 +
#458450000000
0!
0'
#458460000000
1!
1$
b1 %
1'
1*
b1 +
#458470000000
0!
0'
#458480000000
1!
b10 %
1'
b10 +
#458490000000
0!
0'
#458500000000
1!
b11 %
1'
b11 +
#458510000000
0!
0'
#458520000000
1!
b100 %
1'
b100 +
#458530000000
0!
0'
#458540000000
1!
b101 %
1'
b101 +
#458550000000
0!
0'
#458560000000
1!
0$
b110 %
1'
0*
b110 +
#458570000000
0!
0'
#458580000000
1!
b111 %
1'
b111 +
#458590000000
1"
1(
#458600000000
0!
0"
b100 &
0'
0(
b100 ,
#458610000000
1!
b1000 %
1'
b1000 +
#458620000000
0!
0'
#458630000000
1!
b1001 %
1'
b1001 +
#458640000000
0!
0'
#458650000000
1!
b0 %
1'
b0 +
#458660000000
0!
0'
#458670000000
1!
1$
b1 %
1'
1*
b1 +
#458680000000
0!
0'
#458690000000
1!
b10 %
1'
b10 +
#458700000000
0!
0'
#458710000000
1!
b11 %
1'
b11 +
#458720000000
0!
0'
#458730000000
1!
b100 %
1'
b100 +
#458740000000
0!
0'
#458750000000
1!
b101 %
1'
b101 +
#458760000000
0!
0'
#458770000000
1!
b110 %
1'
b110 +
#458780000000
0!
0'
#458790000000
1!
b111 %
1'
b111 +
#458800000000
0!
0'
#458810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#458820000000
0!
0'
#458830000000
1!
b1001 %
1'
b1001 +
#458840000000
0!
0'
#458850000000
1!
b0 %
1'
b0 +
#458860000000
0!
0'
#458870000000
1!
1$
b1 %
1'
1*
b1 +
#458880000000
0!
0'
#458890000000
1!
b10 %
1'
b10 +
#458900000000
0!
0'
#458910000000
1!
b11 %
1'
b11 +
#458920000000
0!
0'
#458930000000
1!
b100 %
1'
b100 +
#458940000000
0!
0'
#458950000000
1!
b101 %
1'
b101 +
#458960000000
0!
0'
#458970000000
1!
0$
b110 %
1'
0*
b110 +
#458980000000
0!
0'
#458990000000
1!
b111 %
1'
b111 +
#459000000000
0!
0'
#459010000000
1!
b1000 %
1'
b1000 +
#459020000000
1"
1(
#459030000000
0!
0"
b100 &
0'
0(
b100 ,
#459040000000
1!
b1001 %
1'
b1001 +
#459050000000
0!
0'
#459060000000
1!
b0 %
1'
b0 +
#459070000000
0!
0'
#459080000000
1!
1$
b1 %
1'
1*
b1 +
#459090000000
0!
0'
#459100000000
1!
b10 %
1'
b10 +
#459110000000
0!
0'
#459120000000
1!
b11 %
1'
b11 +
#459130000000
0!
0'
#459140000000
1!
b100 %
1'
b100 +
#459150000000
0!
0'
#459160000000
1!
b101 %
1'
b101 +
#459170000000
0!
0'
#459180000000
1!
b110 %
1'
b110 +
#459190000000
0!
0'
#459200000000
1!
b111 %
1'
b111 +
#459210000000
0!
0'
#459220000000
1!
0$
b1000 %
1'
0*
b1000 +
#459230000000
0!
0'
#459240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#459250000000
0!
0'
#459260000000
1!
b0 %
1'
b0 +
#459270000000
0!
0'
#459280000000
1!
1$
b1 %
1'
1*
b1 +
#459290000000
0!
0'
#459300000000
1!
b10 %
1'
b10 +
#459310000000
0!
0'
#459320000000
1!
b11 %
1'
b11 +
#459330000000
0!
0'
#459340000000
1!
b100 %
1'
b100 +
#459350000000
0!
0'
#459360000000
1!
b101 %
1'
b101 +
#459370000000
0!
0'
#459380000000
1!
0$
b110 %
1'
0*
b110 +
#459390000000
0!
0'
#459400000000
1!
b111 %
1'
b111 +
#459410000000
0!
0'
#459420000000
1!
b1000 %
1'
b1000 +
#459430000000
0!
0'
#459440000000
1!
b1001 %
1'
b1001 +
#459450000000
1"
1(
#459460000000
0!
0"
b100 &
0'
0(
b100 ,
#459470000000
1!
b0 %
1'
b0 +
#459480000000
0!
0'
#459490000000
1!
1$
b1 %
1'
1*
b1 +
#459500000000
0!
0'
#459510000000
1!
b10 %
1'
b10 +
#459520000000
0!
0'
#459530000000
1!
b11 %
1'
b11 +
#459540000000
0!
0'
#459550000000
1!
b100 %
1'
b100 +
#459560000000
0!
0'
#459570000000
1!
b101 %
1'
b101 +
#459580000000
0!
0'
#459590000000
1!
b110 %
1'
b110 +
#459600000000
0!
0'
#459610000000
1!
b111 %
1'
b111 +
#459620000000
0!
0'
#459630000000
1!
0$
b1000 %
1'
0*
b1000 +
#459640000000
0!
0'
#459650000000
1!
b1001 %
1'
b1001 +
#459660000000
0!
0'
#459670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#459680000000
0!
0'
#459690000000
1!
1$
b1 %
1'
1*
b1 +
#459700000000
0!
0'
#459710000000
1!
b10 %
1'
b10 +
#459720000000
0!
0'
#459730000000
1!
b11 %
1'
b11 +
#459740000000
0!
0'
#459750000000
1!
b100 %
1'
b100 +
#459760000000
0!
0'
#459770000000
1!
b101 %
1'
b101 +
#459780000000
0!
0'
#459790000000
1!
0$
b110 %
1'
0*
b110 +
#459800000000
0!
0'
#459810000000
1!
b111 %
1'
b111 +
#459820000000
0!
0'
#459830000000
1!
b1000 %
1'
b1000 +
#459840000000
0!
0'
#459850000000
1!
b1001 %
1'
b1001 +
#459860000000
0!
0'
#459870000000
1!
b0 %
1'
b0 +
#459880000000
1"
1(
#459890000000
0!
0"
b100 &
0'
0(
b100 ,
#459900000000
1!
1$
b1 %
1'
1*
b1 +
#459910000000
0!
0'
#459920000000
1!
b10 %
1'
b10 +
#459930000000
0!
0'
#459940000000
1!
b11 %
1'
b11 +
#459950000000
0!
0'
#459960000000
1!
b100 %
1'
b100 +
#459970000000
0!
0'
#459980000000
1!
b101 %
1'
b101 +
#459990000000
0!
0'
#460000000000
1!
b110 %
1'
b110 +
#460010000000
0!
0'
#460020000000
1!
b111 %
1'
b111 +
#460030000000
0!
0'
#460040000000
1!
0$
b1000 %
1'
0*
b1000 +
#460050000000
0!
0'
#460060000000
1!
b1001 %
1'
b1001 +
#460070000000
0!
0'
#460080000000
1!
b0 %
1'
b0 +
#460090000000
0!
0'
#460100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#460110000000
0!
0'
#460120000000
1!
b10 %
1'
b10 +
#460130000000
0!
0'
#460140000000
1!
b11 %
1'
b11 +
#460150000000
0!
0'
#460160000000
1!
b100 %
1'
b100 +
#460170000000
0!
0'
#460180000000
1!
b101 %
1'
b101 +
#460190000000
0!
0'
#460200000000
1!
0$
b110 %
1'
0*
b110 +
#460210000000
0!
0'
#460220000000
1!
b111 %
1'
b111 +
#460230000000
0!
0'
#460240000000
1!
b1000 %
1'
b1000 +
#460250000000
0!
0'
#460260000000
1!
b1001 %
1'
b1001 +
#460270000000
0!
0'
#460280000000
1!
b0 %
1'
b0 +
#460290000000
0!
0'
#460300000000
1!
1$
b1 %
1'
1*
b1 +
#460310000000
1"
1(
#460320000000
0!
0"
b100 &
0'
0(
b100 ,
#460330000000
1!
b10 %
1'
b10 +
#460340000000
0!
0'
#460350000000
1!
b11 %
1'
b11 +
#460360000000
0!
0'
#460370000000
1!
b100 %
1'
b100 +
#460380000000
0!
0'
#460390000000
1!
b101 %
1'
b101 +
#460400000000
0!
0'
#460410000000
1!
b110 %
1'
b110 +
#460420000000
0!
0'
#460430000000
1!
b111 %
1'
b111 +
#460440000000
0!
0'
#460450000000
1!
0$
b1000 %
1'
0*
b1000 +
#460460000000
0!
0'
#460470000000
1!
b1001 %
1'
b1001 +
#460480000000
0!
0'
#460490000000
1!
b0 %
1'
b0 +
#460500000000
0!
0'
#460510000000
1!
1$
b1 %
1'
1*
b1 +
#460520000000
0!
0'
#460530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#460540000000
0!
0'
#460550000000
1!
b11 %
1'
b11 +
#460560000000
0!
0'
#460570000000
1!
b100 %
1'
b100 +
#460580000000
0!
0'
#460590000000
1!
b101 %
1'
b101 +
#460600000000
0!
0'
#460610000000
1!
0$
b110 %
1'
0*
b110 +
#460620000000
0!
0'
#460630000000
1!
b111 %
1'
b111 +
#460640000000
0!
0'
#460650000000
1!
b1000 %
1'
b1000 +
#460660000000
0!
0'
#460670000000
1!
b1001 %
1'
b1001 +
#460680000000
0!
0'
#460690000000
1!
b0 %
1'
b0 +
#460700000000
0!
0'
#460710000000
1!
1$
b1 %
1'
1*
b1 +
#460720000000
0!
0'
#460730000000
1!
b10 %
1'
b10 +
#460740000000
1"
1(
#460750000000
0!
0"
b100 &
0'
0(
b100 ,
#460760000000
1!
b11 %
1'
b11 +
#460770000000
0!
0'
#460780000000
1!
b100 %
1'
b100 +
#460790000000
0!
0'
#460800000000
1!
b101 %
1'
b101 +
#460810000000
0!
0'
#460820000000
1!
b110 %
1'
b110 +
#460830000000
0!
0'
#460840000000
1!
b111 %
1'
b111 +
#460850000000
0!
0'
#460860000000
1!
0$
b1000 %
1'
0*
b1000 +
#460870000000
0!
0'
#460880000000
1!
b1001 %
1'
b1001 +
#460890000000
0!
0'
#460900000000
1!
b0 %
1'
b0 +
#460910000000
0!
0'
#460920000000
1!
1$
b1 %
1'
1*
b1 +
#460930000000
0!
0'
#460940000000
1!
b10 %
1'
b10 +
#460950000000
0!
0'
#460960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#460970000000
0!
0'
#460980000000
1!
b100 %
1'
b100 +
#460990000000
0!
0'
#461000000000
1!
b101 %
1'
b101 +
#461010000000
0!
0'
#461020000000
1!
0$
b110 %
1'
0*
b110 +
#461030000000
0!
0'
#461040000000
1!
b111 %
1'
b111 +
#461050000000
0!
0'
#461060000000
1!
b1000 %
1'
b1000 +
#461070000000
0!
0'
#461080000000
1!
b1001 %
1'
b1001 +
#461090000000
0!
0'
#461100000000
1!
b0 %
1'
b0 +
#461110000000
0!
0'
#461120000000
1!
1$
b1 %
1'
1*
b1 +
#461130000000
0!
0'
#461140000000
1!
b10 %
1'
b10 +
#461150000000
0!
0'
#461160000000
1!
b11 %
1'
b11 +
#461170000000
1"
1(
#461180000000
0!
0"
b100 &
0'
0(
b100 ,
#461190000000
1!
b100 %
1'
b100 +
#461200000000
0!
0'
#461210000000
1!
b101 %
1'
b101 +
#461220000000
0!
0'
#461230000000
1!
b110 %
1'
b110 +
#461240000000
0!
0'
#461250000000
1!
b111 %
1'
b111 +
#461260000000
0!
0'
#461270000000
1!
0$
b1000 %
1'
0*
b1000 +
#461280000000
0!
0'
#461290000000
1!
b1001 %
1'
b1001 +
#461300000000
0!
0'
#461310000000
1!
b0 %
1'
b0 +
#461320000000
0!
0'
#461330000000
1!
1$
b1 %
1'
1*
b1 +
#461340000000
0!
0'
#461350000000
1!
b10 %
1'
b10 +
#461360000000
0!
0'
#461370000000
1!
b11 %
1'
b11 +
#461380000000
0!
0'
#461390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#461400000000
0!
0'
#461410000000
1!
b101 %
1'
b101 +
#461420000000
0!
0'
#461430000000
1!
0$
b110 %
1'
0*
b110 +
#461440000000
0!
0'
#461450000000
1!
b111 %
1'
b111 +
#461460000000
0!
0'
#461470000000
1!
b1000 %
1'
b1000 +
#461480000000
0!
0'
#461490000000
1!
b1001 %
1'
b1001 +
#461500000000
0!
0'
#461510000000
1!
b0 %
1'
b0 +
#461520000000
0!
0'
#461530000000
1!
1$
b1 %
1'
1*
b1 +
#461540000000
0!
0'
#461550000000
1!
b10 %
1'
b10 +
#461560000000
0!
0'
#461570000000
1!
b11 %
1'
b11 +
#461580000000
0!
0'
#461590000000
1!
b100 %
1'
b100 +
#461600000000
1"
1(
#461610000000
0!
0"
b100 &
0'
0(
b100 ,
#461620000000
1!
b101 %
1'
b101 +
#461630000000
0!
0'
#461640000000
1!
b110 %
1'
b110 +
#461650000000
0!
0'
#461660000000
1!
b111 %
1'
b111 +
#461670000000
0!
0'
#461680000000
1!
0$
b1000 %
1'
0*
b1000 +
#461690000000
0!
0'
#461700000000
1!
b1001 %
1'
b1001 +
#461710000000
0!
0'
#461720000000
1!
b0 %
1'
b0 +
#461730000000
0!
0'
#461740000000
1!
1$
b1 %
1'
1*
b1 +
#461750000000
0!
0'
#461760000000
1!
b10 %
1'
b10 +
#461770000000
0!
0'
#461780000000
1!
b11 %
1'
b11 +
#461790000000
0!
0'
#461800000000
1!
b100 %
1'
b100 +
#461810000000
0!
0'
#461820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#461830000000
0!
0'
#461840000000
1!
0$
b110 %
1'
0*
b110 +
#461850000000
0!
0'
#461860000000
1!
b111 %
1'
b111 +
#461870000000
0!
0'
#461880000000
1!
b1000 %
1'
b1000 +
#461890000000
0!
0'
#461900000000
1!
b1001 %
1'
b1001 +
#461910000000
0!
0'
#461920000000
1!
b0 %
1'
b0 +
#461930000000
0!
0'
#461940000000
1!
1$
b1 %
1'
1*
b1 +
#461950000000
0!
0'
#461960000000
1!
b10 %
1'
b10 +
#461970000000
0!
0'
#461980000000
1!
b11 %
1'
b11 +
#461990000000
0!
0'
#462000000000
1!
b100 %
1'
b100 +
#462010000000
0!
0'
#462020000000
1!
b101 %
1'
b101 +
#462030000000
1"
1(
#462040000000
0!
0"
b100 &
0'
0(
b100 ,
#462050000000
1!
b110 %
1'
b110 +
#462060000000
0!
0'
#462070000000
1!
b111 %
1'
b111 +
#462080000000
0!
0'
#462090000000
1!
0$
b1000 %
1'
0*
b1000 +
#462100000000
0!
0'
#462110000000
1!
b1001 %
1'
b1001 +
#462120000000
0!
0'
#462130000000
1!
b0 %
1'
b0 +
#462140000000
0!
0'
#462150000000
1!
1$
b1 %
1'
1*
b1 +
#462160000000
0!
0'
#462170000000
1!
b10 %
1'
b10 +
#462180000000
0!
0'
#462190000000
1!
b11 %
1'
b11 +
#462200000000
0!
0'
#462210000000
1!
b100 %
1'
b100 +
#462220000000
0!
0'
#462230000000
1!
b101 %
1'
b101 +
#462240000000
0!
0'
#462250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#462260000000
0!
0'
#462270000000
1!
b111 %
1'
b111 +
#462280000000
0!
0'
#462290000000
1!
b1000 %
1'
b1000 +
#462300000000
0!
0'
#462310000000
1!
b1001 %
1'
b1001 +
#462320000000
0!
0'
#462330000000
1!
b0 %
1'
b0 +
#462340000000
0!
0'
#462350000000
1!
1$
b1 %
1'
1*
b1 +
#462360000000
0!
0'
#462370000000
1!
b10 %
1'
b10 +
#462380000000
0!
0'
#462390000000
1!
b11 %
1'
b11 +
#462400000000
0!
0'
#462410000000
1!
b100 %
1'
b100 +
#462420000000
0!
0'
#462430000000
1!
b101 %
1'
b101 +
#462440000000
0!
0'
#462450000000
1!
0$
b110 %
1'
0*
b110 +
#462460000000
1"
1(
#462470000000
0!
0"
b100 &
0'
0(
b100 ,
#462480000000
1!
1$
b111 %
1'
1*
b111 +
#462490000000
0!
0'
#462500000000
1!
0$
b1000 %
1'
0*
b1000 +
#462510000000
0!
0'
#462520000000
1!
b1001 %
1'
b1001 +
#462530000000
0!
0'
#462540000000
1!
b0 %
1'
b0 +
#462550000000
0!
0'
#462560000000
1!
1$
b1 %
1'
1*
b1 +
#462570000000
0!
0'
#462580000000
1!
b10 %
1'
b10 +
#462590000000
0!
0'
#462600000000
1!
b11 %
1'
b11 +
#462610000000
0!
0'
#462620000000
1!
b100 %
1'
b100 +
#462630000000
0!
0'
#462640000000
1!
b101 %
1'
b101 +
#462650000000
0!
0'
#462660000000
1!
b110 %
1'
b110 +
#462670000000
0!
0'
#462680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#462690000000
0!
0'
#462700000000
1!
b1000 %
1'
b1000 +
#462710000000
0!
0'
#462720000000
1!
b1001 %
1'
b1001 +
#462730000000
0!
0'
#462740000000
1!
b0 %
1'
b0 +
#462750000000
0!
0'
#462760000000
1!
1$
b1 %
1'
1*
b1 +
#462770000000
0!
0'
#462780000000
1!
b10 %
1'
b10 +
#462790000000
0!
0'
#462800000000
1!
b11 %
1'
b11 +
#462810000000
0!
0'
#462820000000
1!
b100 %
1'
b100 +
#462830000000
0!
0'
#462840000000
1!
b101 %
1'
b101 +
#462850000000
0!
0'
#462860000000
1!
0$
b110 %
1'
0*
b110 +
#462870000000
0!
0'
#462880000000
1!
b111 %
1'
b111 +
#462890000000
1"
1(
#462900000000
0!
0"
b100 &
0'
0(
b100 ,
#462910000000
1!
b1000 %
1'
b1000 +
#462920000000
0!
0'
#462930000000
1!
b1001 %
1'
b1001 +
#462940000000
0!
0'
#462950000000
1!
b0 %
1'
b0 +
#462960000000
0!
0'
#462970000000
1!
1$
b1 %
1'
1*
b1 +
#462980000000
0!
0'
#462990000000
1!
b10 %
1'
b10 +
#463000000000
0!
0'
#463010000000
1!
b11 %
1'
b11 +
#463020000000
0!
0'
#463030000000
1!
b100 %
1'
b100 +
#463040000000
0!
0'
#463050000000
1!
b101 %
1'
b101 +
#463060000000
0!
0'
#463070000000
1!
b110 %
1'
b110 +
#463080000000
0!
0'
#463090000000
1!
b111 %
1'
b111 +
#463100000000
0!
0'
#463110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#463120000000
0!
0'
#463130000000
1!
b1001 %
1'
b1001 +
#463140000000
0!
0'
#463150000000
1!
b0 %
1'
b0 +
#463160000000
0!
0'
#463170000000
1!
1$
b1 %
1'
1*
b1 +
#463180000000
0!
0'
#463190000000
1!
b10 %
1'
b10 +
#463200000000
0!
0'
#463210000000
1!
b11 %
1'
b11 +
#463220000000
0!
0'
#463230000000
1!
b100 %
1'
b100 +
#463240000000
0!
0'
#463250000000
1!
b101 %
1'
b101 +
#463260000000
0!
0'
#463270000000
1!
0$
b110 %
1'
0*
b110 +
#463280000000
0!
0'
#463290000000
1!
b111 %
1'
b111 +
#463300000000
0!
0'
#463310000000
1!
b1000 %
1'
b1000 +
#463320000000
1"
1(
#463330000000
0!
0"
b100 &
0'
0(
b100 ,
#463340000000
1!
b1001 %
1'
b1001 +
#463350000000
0!
0'
#463360000000
1!
b0 %
1'
b0 +
#463370000000
0!
0'
#463380000000
1!
1$
b1 %
1'
1*
b1 +
#463390000000
0!
0'
#463400000000
1!
b10 %
1'
b10 +
#463410000000
0!
0'
#463420000000
1!
b11 %
1'
b11 +
#463430000000
0!
0'
#463440000000
1!
b100 %
1'
b100 +
#463450000000
0!
0'
#463460000000
1!
b101 %
1'
b101 +
#463470000000
0!
0'
#463480000000
1!
b110 %
1'
b110 +
#463490000000
0!
0'
#463500000000
1!
b111 %
1'
b111 +
#463510000000
0!
0'
#463520000000
1!
0$
b1000 %
1'
0*
b1000 +
#463530000000
0!
0'
#463540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#463550000000
0!
0'
#463560000000
1!
b0 %
1'
b0 +
#463570000000
0!
0'
#463580000000
1!
1$
b1 %
1'
1*
b1 +
#463590000000
0!
0'
#463600000000
1!
b10 %
1'
b10 +
#463610000000
0!
0'
#463620000000
1!
b11 %
1'
b11 +
#463630000000
0!
0'
#463640000000
1!
b100 %
1'
b100 +
#463650000000
0!
0'
#463660000000
1!
b101 %
1'
b101 +
#463670000000
0!
0'
#463680000000
1!
0$
b110 %
1'
0*
b110 +
#463690000000
0!
0'
#463700000000
1!
b111 %
1'
b111 +
#463710000000
0!
0'
#463720000000
1!
b1000 %
1'
b1000 +
#463730000000
0!
0'
#463740000000
1!
b1001 %
1'
b1001 +
#463750000000
1"
1(
#463760000000
0!
0"
b100 &
0'
0(
b100 ,
#463770000000
1!
b0 %
1'
b0 +
#463780000000
0!
0'
#463790000000
1!
1$
b1 %
1'
1*
b1 +
#463800000000
0!
0'
#463810000000
1!
b10 %
1'
b10 +
#463820000000
0!
0'
#463830000000
1!
b11 %
1'
b11 +
#463840000000
0!
0'
#463850000000
1!
b100 %
1'
b100 +
#463860000000
0!
0'
#463870000000
1!
b101 %
1'
b101 +
#463880000000
0!
0'
#463890000000
1!
b110 %
1'
b110 +
#463900000000
0!
0'
#463910000000
1!
b111 %
1'
b111 +
#463920000000
0!
0'
#463930000000
1!
0$
b1000 %
1'
0*
b1000 +
#463940000000
0!
0'
#463950000000
1!
b1001 %
1'
b1001 +
#463960000000
0!
0'
#463970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#463980000000
0!
0'
#463990000000
1!
1$
b1 %
1'
1*
b1 +
#464000000000
0!
0'
#464010000000
1!
b10 %
1'
b10 +
#464020000000
0!
0'
#464030000000
1!
b11 %
1'
b11 +
#464040000000
0!
0'
#464050000000
1!
b100 %
1'
b100 +
#464060000000
0!
0'
#464070000000
1!
b101 %
1'
b101 +
#464080000000
0!
0'
#464090000000
1!
0$
b110 %
1'
0*
b110 +
#464100000000
0!
0'
#464110000000
1!
b111 %
1'
b111 +
#464120000000
0!
0'
#464130000000
1!
b1000 %
1'
b1000 +
#464140000000
0!
0'
#464150000000
1!
b1001 %
1'
b1001 +
#464160000000
0!
0'
#464170000000
1!
b0 %
1'
b0 +
#464180000000
1"
1(
#464190000000
0!
0"
b100 &
0'
0(
b100 ,
#464200000000
1!
1$
b1 %
1'
1*
b1 +
#464210000000
0!
0'
#464220000000
1!
b10 %
1'
b10 +
#464230000000
0!
0'
#464240000000
1!
b11 %
1'
b11 +
#464250000000
0!
0'
#464260000000
1!
b100 %
1'
b100 +
#464270000000
0!
0'
#464280000000
1!
b101 %
1'
b101 +
#464290000000
0!
0'
#464300000000
1!
b110 %
1'
b110 +
#464310000000
0!
0'
#464320000000
1!
b111 %
1'
b111 +
#464330000000
0!
0'
#464340000000
1!
0$
b1000 %
1'
0*
b1000 +
#464350000000
0!
0'
#464360000000
1!
b1001 %
1'
b1001 +
#464370000000
0!
0'
#464380000000
1!
b0 %
1'
b0 +
#464390000000
0!
0'
#464400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#464410000000
0!
0'
#464420000000
1!
b10 %
1'
b10 +
#464430000000
0!
0'
#464440000000
1!
b11 %
1'
b11 +
#464450000000
0!
0'
#464460000000
1!
b100 %
1'
b100 +
#464470000000
0!
0'
#464480000000
1!
b101 %
1'
b101 +
#464490000000
0!
0'
#464500000000
1!
0$
b110 %
1'
0*
b110 +
#464510000000
0!
0'
#464520000000
1!
b111 %
1'
b111 +
#464530000000
0!
0'
#464540000000
1!
b1000 %
1'
b1000 +
#464550000000
0!
0'
#464560000000
1!
b1001 %
1'
b1001 +
#464570000000
0!
0'
#464580000000
1!
b0 %
1'
b0 +
#464590000000
0!
0'
#464600000000
1!
1$
b1 %
1'
1*
b1 +
#464610000000
1"
1(
#464620000000
0!
0"
b100 &
0'
0(
b100 ,
#464630000000
1!
b10 %
1'
b10 +
#464640000000
0!
0'
#464650000000
1!
b11 %
1'
b11 +
#464660000000
0!
0'
#464670000000
1!
b100 %
1'
b100 +
#464680000000
0!
0'
#464690000000
1!
b101 %
1'
b101 +
#464700000000
0!
0'
#464710000000
1!
b110 %
1'
b110 +
#464720000000
0!
0'
#464730000000
1!
b111 %
1'
b111 +
#464740000000
0!
0'
#464750000000
1!
0$
b1000 %
1'
0*
b1000 +
#464760000000
0!
0'
#464770000000
1!
b1001 %
1'
b1001 +
#464780000000
0!
0'
#464790000000
1!
b0 %
1'
b0 +
#464800000000
0!
0'
#464810000000
1!
1$
b1 %
1'
1*
b1 +
#464820000000
0!
0'
#464830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#464840000000
0!
0'
#464850000000
1!
b11 %
1'
b11 +
#464860000000
0!
0'
#464870000000
1!
b100 %
1'
b100 +
#464880000000
0!
0'
#464890000000
1!
b101 %
1'
b101 +
#464900000000
0!
0'
#464910000000
1!
0$
b110 %
1'
0*
b110 +
#464920000000
0!
0'
#464930000000
1!
b111 %
1'
b111 +
#464940000000
0!
0'
#464950000000
1!
b1000 %
1'
b1000 +
#464960000000
0!
0'
#464970000000
1!
b1001 %
1'
b1001 +
#464980000000
0!
0'
#464990000000
1!
b0 %
1'
b0 +
#465000000000
0!
0'
#465010000000
1!
1$
b1 %
1'
1*
b1 +
#465020000000
0!
0'
#465030000000
1!
b10 %
1'
b10 +
#465040000000
1"
1(
#465050000000
0!
0"
b100 &
0'
0(
b100 ,
#465060000000
1!
b11 %
1'
b11 +
#465070000000
0!
0'
#465080000000
1!
b100 %
1'
b100 +
#465090000000
0!
0'
#465100000000
1!
b101 %
1'
b101 +
#465110000000
0!
0'
#465120000000
1!
b110 %
1'
b110 +
#465130000000
0!
0'
#465140000000
1!
b111 %
1'
b111 +
#465150000000
0!
0'
#465160000000
1!
0$
b1000 %
1'
0*
b1000 +
#465170000000
0!
0'
#465180000000
1!
b1001 %
1'
b1001 +
#465190000000
0!
0'
#465200000000
1!
b0 %
1'
b0 +
#465210000000
0!
0'
#465220000000
1!
1$
b1 %
1'
1*
b1 +
#465230000000
0!
0'
#465240000000
1!
b10 %
1'
b10 +
#465250000000
0!
0'
#465260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#465270000000
0!
0'
#465280000000
1!
b100 %
1'
b100 +
#465290000000
0!
0'
#465300000000
1!
b101 %
1'
b101 +
#465310000000
0!
0'
#465320000000
1!
0$
b110 %
1'
0*
b110 +
#465330000000
0!
0'
#465340000000
1!
b111 %
1'
b111 +
#465350000000
0!
0'
#465360000000
1!
b1000 %
1'
b1000 +
#465370000000
0!
0'
#465380000000
1!
b1001 %
1'
b1001 +
#465390000000
0!
0'
#465400000000
1!
b0 %
1'
b0 +
#465410000000
0!
0'
#465420000000
1!
1$
b1 %
1'
1*
b1 +
#465430000000
0!
0'
#465440000000
1!
b10 %
1'
b10 +
#465450000000
0!
0'
#465460000000
1!
b11 %
1'
b11 +
#465470000000
1"
1(
#465480000000
0!
0"
b100 &
0'
0(
b100 ,
#465490000000
1!
b100 %
1'
b100 +
#465500000000
0!
0'
#465510000000
1!
b101 %
1'
b101 +
#465520000000
0!
0'
#465530000000
1!
b110 %
1'
b110 +
#465540000000
0!
0'
#465550000000
1!
b111 %
1'
b111 +
#465560000000
0!
0'
#465570000000
1!
0$
b1000 %
1'
0*
b1000 +
#465580000000
0!
0'
#465590000000
1!
b1001 %
1'
b1001 +
#465600000000
0!
0'
#465610000000
1!
b0 %
1'
b0 +
#465620000000
0!
0'
#465630000000
1!
1$
b1 %
1'
1*
b1 +
#465640000000
0!
0'
#465650000000
1!
b10 %
1'
b10 +
#465660000000
0!
0'
#465670000000
1!
b11 %
1'
b11 +
#465680000000
0!
0'
#465690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#465700000000
0!
0'
#465710000000
1!
b101 %
1'
b101 +
#465720000000
0!
0'
#465730000000
1!
0$
b110 %
1'
0*
b110 +
#465740000000
0!
0'
#465750000000
1!
b111 %
1'
b111 +
#465760000000
0!
0'
#465770000000
1!
b1000 %
1'
b1000 +
#465780000000
0!
0'
#465790000000
1!
b1001 %
1'
b1001 +
#465800000000
0!
0'
#465810000000
1!
b0 %
1'
b0 +
#465820000000
0!
0'
#465830000000
1!
1$
b1 %
1'
1*
b1 +
#465840000000
0!
0'
#465850000000
1!
b10 %
1'
b10 +
#465860000000
0!
0'
#465870000000
1!
b11 %
1'
b11 +
#465880000000
0!
0'
#465890000000
1!
b100 %
1'
b100 +
#465900000000
1"
1(
#465910000000
0!
0"
b100 &
0'
0(
b100 ,
#465920000000
1!
b101 %
1'
b101 +
#465930000000
0!
0'
#465940000000
1!
b110 %
1'
b110 +
#465950000000
0!
0'
#465960000000
1!
b111 %
1'
b111 +
#465970000000
0!
0'
#465980000000
1!
0$
b1000 %
1'
0*
b1000 +
#465990000000
0!
0'
#466000000000
1!
b1001 %
1'
b1001 +
#466010000000
0!
0'
#466020000000
1!
b0 %
1'
b0 +
#466030000000
0!
0'
#466040000000
1!
1$
b1 %
1'
1*
b1 +
#466050000000
0!
0'
#466060000000
1!
b10 %
1'
b10 +
#466070000000
0!
0'
#466080000000
1!
b11 %
1'
b11 +
#466090000000
0!
0'
#466100000000
1!
b100 %
1'
b100 +
#466110000000
0!
0'
#466120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#466130000000
0!
0'
#466140000000
1!
0$
b110 %
1'
0*
b110 +
#466150000000
0!
0'
#466160000000
1!
b111 %
1'
b111 +
#466170000000
0!
0'
#466180000000
1!
b1000 %
1'
b1000 +
#466190000000
0!
0'
#466200000000
1!
b1001 %
1'
b1001 +
#466210000000
0!
0'
#466220000000
1!
b0 %
1'
b0 +
#466230000000
0!
0'
#466240000000
1!
1$
b1 %
1'
1*
b1 +
#466250000000
0!
0'
#466260000000
1!
b10 %
1'
b10 +
#466270000000
0!
0'
#466280000000
1!
b11 %
1'
b11 +
#466290000000
0!
0'
#466300000000
1!
b100 %
1'
b100 +
#466310000000
0!
0'
#466320000000
1!
b101 %
1'
b101 +
#466330000000
1"
1(
#466340000000
0!
0"
b100 &
0'
0(
b100 ,
#466350000000
1!
b110 %
1'
b110 +
#466360000000
0!
0'
#466370000000
1!
b111 %
1'
b111 +
#466380000000
0!
0'
#466390000000
1!
0$
b1000 %
1'
0*
b1000 +
#466400000000
0!
0'
#466410000000
1!
b1001 %
1'
b1001 +
#466420000000
0!
0'
#466430000000
1!
b0 %
1'
b0 +
#466440000000
0!
0'
#466450000000
1!
1$
b1 %
1'
1*
b1 +
#466460000000
0!
0'
#466470000000
1!
b10 %
1'
b10 +
#466480000000
0!
0'
#466490000000
1!
b11 %
1'
b11 +
#466500000000
0!
0'
#466510000000
1!
b100 %
1'
b100 +
#466520000000
0!
0'
#466530000000
1!
b101 %
1'
b101 +
#466540000000
0!
0'
#466550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#466560000000
0!
0'
#466570000000
1!
b111 %
1'
b111 +
#466580000000
0!
0'
#466590000000
1!
b1000 %
1'
b1000 +
#466600000000
0!
0'
#466610000000
1!
b1001 %
1'
b1001 +
#466620000000
0!
0'
#466630000000
1!
b0 %
1'
b0 +
#466640000000
0!
0'
#466650000000
1!
1$
b1 %
1'
1*
b1 +
#466660000000
0!
0'
#466670000000
1!
b10 %
1'
b10 +
#466680000000
0!
0'
#466690000000
1!
b11 %
1'
b11 +
#466700000000
0!
0'
#466710000000
1!
b100 %
1'
b100 +
#466720000000
0!
0'
#466730000000
1!
b101 %
1'
b101 +
#466740000000
0!
0'
#466750000000
1!
0$
b110 %
1'
0*
b110 +
#466760000000
1"
1(
#466770000000
0!
0"
b100 &
0'
0(
b100 ,
#466780000000
1!
1$
b111 %
1'
1*
b111 +
#466790000000
0!
0'
#466800000000
1!
0$
b1000 %
1'
0*
b1000 +
#466810000000
0!
0'
#466820000000
1!
b1001 %
1'
b1001 +
#466830000000
0!
0'
#466840000000
1!
b0 %
1'
b0 +
#466850000000
0!
0'
#466860000000
1!
1$
b1 %
1'
1*
b1 +
#466870000000
0!
0'
#466880000000
1!
b10 %
1'
b10 +
#466890000000
0!
0'
#466900000000
1!
b11 %
1'
b11 +
#466910000000
0!
0'
#466920000000
1!
b100 %
1'
b100 +
#466930000000
0!
0'
#466940000000
1!
b101 %
1'
b101 +
#466950000000
0!
0'
#466960000000
1!
b110 %
1'
b110 +
#466970000000
0!
0'
#466980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#466990000000
0!
0'
#467000000000
1!
b1000 %
1'
b1000 +
#467010000000
0!
0'
#467020000000
1!
b1001 %
1'
b1001 +
#467030000000
0!
0'
#467040000000
1!
b0 %
1'
b0 +
#467050000000
0!
0'
#467060000000
1!
1$
b1 %
1'
1*
b1 +
#467070000000
0!
0'
#467080000000
1!
b10 %
1'
b10 +
#467090000000
0!
0'
#467100000000
1!
b11 %
1'
b11 +
#467110000000
0!
0'
#467120000000
1!
b100 %
1'
b100 +
#467130000000
0!
0'
#467140000000
1!
b101 %
1'
b101 +
#467150000000
0!
0'
#467160000000
1!
0$
b110 %
1'
0*
b110 +
#467170000000
0!
0'
#467180000000
1!
b111 %
1'
b111 +
#467190000000
1"
1(
#467200000000
0!
0"
b100 &
0'
0(
b100 ,
#467210000000
1!
b1000 %
1'
b1000 +
#467220000000
0!
0'
#467230000000
1!
b1001 %
1'
b1001 +
#467240000000
0!
0'
#467250000000
1!
b0 %
1'
b0 +
#467260000000
0!
0'
#467270000000
1!
1$
b1 %
1'
1*
b1 +
#467280000000
0!
0'
#467290000000
1!
b10 %
1'
b10 +
#467300000000
0!
0'
#467310000000
1!
b11 %
1'
b11 +
#467320000000
0!
0'
#467330000000
1!
b100 %
1'
b100 +
#467340000000
0!
0'
#467350000000
1!
b101 %
1'
b101 +
#467360000000
0!
0'
#467370000000
1!
b110 %
1'
b110 +
#467380000000
0!
0'
#467390000000
1!
b111 %
1'
b111 +
#467400000000
0!
0'
#467410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#467420000000
0!
0'
#467430000000
1!
b1001 %
1'
b1001 +
#467440000000
0!
0'
#467450000000
1!
b0 %
1'
b0 +
#467460000000
0!
0'
#467470000000
1!
1$
b1 %
1'
1*
b1 +
#467480000000
0!
0'
#467490000000
1!
b10 %
1'
b10 +
#467500000000
0!
0'
#467510000000
1!
b11 %
1'
b11 +
#467520000000
0!
0'
#467530000000
1!
b100 %
1'
b100 +
#467540000000
0!
0'
#467550000000
1!
b101 %
1'
b101 +
#467560000000
0!
0'
#467570000000
1!
0$
b110 %
1'
0*
b110 +
#467580000000
0!
0'
#467590000000
1!
b111 %
1'
b111 +
#467600000000
0!
0'
#467610000000
1!
b1000 %
1'
b1000 +
#467620000000
1"
1(
#467630000000
0!
0"
b100 &
0'
0(
b100 ,
#467640000000
1!
b1001 %
1'
b1001 +
#467650000000
0!
0'
#467660000000
1!
b0 %
1'
b0 +
#467670000000
0!
0'
#467680000000
1!
1$
b1 %
1'
1*
b1 +
#467690000000
0!
0'
#467700000000
1!
b10 %
1'
b10 +
#467710000000
0!
0'
#467720000000
1!
b11 %
1'
b11 +
#467730000000
0!
0'
#467740000000
1!
b100 %
1'
b100 +
#467750000000
0!
0'
#467760000000
1!
b101 %
1'
b101 +
#467770000000
0!
0'
#467780000000
1!
b110 %
1'
b110 +
#467790000000
0!
0'
#467800000000
1!
b111 %
1'
b111 +
#467810000000
0!
0'
#467820000000
1!
0$
b1000 %
1'
0*
b1000 +
#467830000000
0!
0'
#467840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#467850000000
0!
0'
#467860000000
1!
b0 %
1'
b0 +
#467870000000
0!
0'
#467880000000
1!
1$
b1 %
1'
1*
b1 +
#467890000000
0!
0'
#467900000000
1!
b10 %
1'
b10 +
#467910000000
0!
0'
#467920000000
1!
b11 %
1'
b11 +
#467930000000
0!
0'
#467940000000
1!
b100 %
1'
b100 +
#467950000000
0!
0'
#467960000000
1!
b101 %
1'
b101 +
#467970000000
0!
0'
#467980000000
1!
0$
b110 %
1'
0*
b110 +
#467990000000
0!
0'
#468000000000
1!
b111 %
1'
b111 +
#468010000000
0!
0'
#468020000000
1!
b1000 %
1'
b1000 +
#468030000000
0!
0'
#468040000000
1!
b1001 %
1'
b1001 +
#468050000000
1"
1(
#468060000000
0!
0"
b100 &
0'
0(
b100 ,
#468070000000
1!
b0 %
1'
b0 +
#468080000000
0!
0'
#468090000000
1!
1$
b1 %
1'
1*
b1 +
#468100000000
0!
0'
#468110000000
1!
b10 %
1'
b10 +
#468120000000
0!
0'
#468130000000
1!
b11 %
1'
b11 +
#468140000000
0!
0'
#468150000000
1!
b100 %
1'
b100 +
#468160000000
0!
0'
#468170000000
1!
b101 %
1'
b101 +
#468180000000
0!
0'
#468190000000
1!
b110 %
1'
b110 +
#468200000000
0!
0'
#468210000000
1!
b111 %
1'
b111 +
#468220000000
0!
0'
#468230000000
1!
0$
b1000 %
1'
0*
b1000 +
#468240000000
0!
0'
#468250000000
1!
b1001 %
1'
b1001 +
#468260000000
0!
0'
#468270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#468280000000
0!
0'
#468290000000
1!
1$
b1 %
1'
1*
b1 +
#468300000000
0!
0'
#468310000000
1!
b10 %
1'
b10 +
#468320000000
0!
0'
#468330000000
1!
b11 %
1'
b11 +
#468340000000
0!
0'
#468350000000
1!
b100 %
1'
b100 +
#468360000000
0!
0'
#468370000000
1!
b101 %
1'
b101 +
#468380000000
0!
0'
#468390000000
1!
0$
b110 %
1'
0*
b110 +
#468400000000
0!
0'
#468410000000
1!
b111 %
1'
b111 +
#468420000000
0!
0'
#468430000000
1!
b1000 %
1'
b1000 +
#468440000000
0!
0'
#468450000000
1!
b1001 %
1'
b1001 +
#468460000000
0!
0'
#468470000000
1!
b0 %
1'
b0 +
#468480000000
1"
1(
#468490000000
0!
0"
b100 &
0'
0(
b100 ,
#468500000000
1!
1$
b1 %
1'
1*
b1 +
#468510000000
0!
0'
#468520000000
1!
b10 %
1'
b10 +
#468530000000
0!
0'
#468540000000
1!
b11 %
1'
b11 +
#468550000000
0!
0'
#468560000000
1!
b100 %
1'
b100 +
#468570000000
0!
0'
#468580000000
1!
b101 %
1'
b101 +
#468590000000
0!
0'
#468600000000
1!
b110 %
1'
b110 +
#468610000000
0!
0'
#468620000000
1!
b111 %
1'
b111 +
#468630000000
0!
0'
#468640000000
1!
0$
b1000 %
1'
0*
b1000 +
#468650000000
0!
0'
#468660000000
1!
b1001 %
1'
b1001 +
#468670000000
0!
0'
#468680000000
1!
b0 %
1'
b0 +
#468690000000
0!
0'
#468700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#468710000000
0!
0'
#468720000000
1!
b10 %
1'
b10 +
#468730000000
0!
0'
#468740000000
1!
b11 %
1'
b11 +
#468750000000
0!
0'
#468760000000
1!
b100 %
1'
b100 +
#468770000000
0!
0'
#468780000000
1!
b101 %
1'
b101 +
#468790000000
0!
0'
#468800000000
1!
0$
b110 %
1'
0*
b110 +
#468810000000
0!
0'
#468820000000
1!
b111 %
1'
b111 +
#468830000000
0!
0'
#468840000000
1!
b1000 %
1'
b1000 +
#468850000000
0!
0'
#468860000000
1!
b1001 %
1'
b1001 +
#468870000000
0!
0'
#468880000000
1!
b0 %
1'
b0 +
#468890000000
0!
0'
#468900000000
1!
1$
b1 %
1'
1*
b1 +
#468910000000
1"
1(
#468920000000
0!
0"
b100 &
0'
0(
b100 ,
#468930000000
1!
b10 %
1'
b10 +
#468940000000
0!
0'
#468950000000
1!
b11 %
1'
b11 +
#468960000000
0!
0'
#468970000000
1!
b100 %
1'
b100 +
#468980000000
0!
0'
#468990000000
1!
b101 %
1'
b101 +
#469000000000
0!
0'
#469010000000
1!
b110 %
1'
b110 +
#469020000000
0!
0'
#469030000000
1!
b111 %
1'
b111 +
#469040000000
0!
0'
#469050000000
1!
0$
b1000 %
1'
0*
b1000 +
#469060000000
0!
0'
#469070000000
1!
b1001 %
1'
b1001 +
#469080000000
0!
0'
#469090000000
1!
b0 %
1'
b0 +
#469100000000
0!
0'
#469110000000
1!
1$
b1 %
1'
1*
b1 +
#469120000000
0!
0'
#469130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#469140000000
0!
0'
#469150000000
1!
b11 %
1'
b11 +
#469160000000
0!
0'
#469170000000
1!
b100 %
1'
b100 +
#469180000000
0!
0'
#469190000000
1!
b101 %
1'
b101 +
#469200000000
0!
0'
#469210000000
1!
0$
b110 %
1'
0*
b110 +
#469220000000
0!
0'
#469230000000
1!
b111 %
1'
b111 +
#469240000000
0!
0'
#469250000000
1!
b1000 %
1'
b1000 +
#469260000000
0!
0'
#469270000000
1!
b1001 %
1'
b1001 +
#469280000000
0!
0'
#469290000000
1!
b0 %
1'
b0 +
#469300000000
0!
0'
#469310000000
1!
1$
b1 %
1'
1*
b1 +
#469320000000
0!
0'
#469330000000
1!
b10 %
1'
b10 +
#469340000000
1"
1(
#469350000000
0!
0"
b100 &
0'
0(
b100 ,
#469360000000
1!
b11 %
1'
b11 +
#469370000000
0!
0'
#469380000000
1!
b100 %
1'
b100 +
#469390000000
0!
0'
#469400000000
1!
b101 %
1'
b101 +
#469410000000
0!
0'
#469420000000
1!
b110 %
1'
b110 +
#469430000000
0!
0'
#469440000000
1!
b111 %
1'
b111 +
#469450000000
0!
0'
#469460000000
1!
0$
b1000 %
1'
0*
b1000 +
#469470000000
0!
0'
#469480000000
1!
b1001 %
1'
b1001 +
#469490000000
0!
0'
#469500000000
1!
b0 %
1'
b0 +
#469510000000
0!
0'
#469520000000
1!
1$
b1 %
1'
1*
b1 +
#469530000000
0!
0'
#469540000000
1!
b10 %
1'
b10 +
#469550000000
0!
0'
#469560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#469570000000
0!
0'
#469580000000
1!
b100 %
1'
b100 +
#469590000000
0!
0'
#469600000000
1!
b101 %
1'
b101 +
#469610000000
0!
0'
#469620000000
1!
0$
b110 %
1'
0*
b110 +
#469630000000
0!
0'
#469640000000
1!
b111 %
1'
b111 +
#469650000000
0!
0'
#469660000000
1!
b1000 %
1'
b1000 +
#469670000000
0!
0'
#469680000000
1!
b1001 %
1'
b1001 +
#469690000000
0!
0'
#469700000000
1!
b0 %
1'
b0 +
#469710000000
0!
0'
#469720000000
1!
1$
b1 %
1'
1*
b1 +
#469730000000
0!
0'
#469740000000
1!
b10 %
1'
b10 +
#469750000000
0!
0'
#469760000000
1!
b11 %
1'
b11 +
#469770000000
1"
1(
#469780000000
0!
0"
b100 &
0'
0(
b100 ,
#469790000000
1!
b100 %
1'
b100 +
#469800000000
0!
0'
#469810000000
1!
b101 %
1'
b101 +
#469820000000
0!
0'
#469830000000
1!
b110 %
1'
b110 +
#469840000000
0!
0'
#469850000000
1!
b111 %
1'
b111 +
#469860000000
0!
0'
#469870000000
1!
0$
b1000 %
1'
0*
b1000 +
#469880000000
0!
0'
#469890000000
1!
b1001 %
1'
b1001 +
#469900000000
0!
0'
#469910000000
1!
b0 %
1'
b0 +
#469920000000
0!
0'
#469930000000
1!
1$
b1 %
1'
1*
b1 +
#469940000000
0!
0'
#469950000000
1!
b10 %
1'
b10 +
#469960000000
0!
0'
#469970000000
1!
b11 %
1'
b11 +
#469980000000
0!
0'
#469990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#470000000000
0!
0'
#470010000000
1!
b101 %
1'
b101 +
#470020000000
0!
0'
#470030000000
1!
0$
b110 %
1'
0*
b110 +
#470040000000
0!
0'
#470050000000
1!
b111 %
1'
b111 +
#470060000000
0!
0'
#470070000000
1!
b1000 %
1'
b1000 +
#470080000000
0!
0'
#470090000000
1!
b1001 %
1'
b1001 +
#470100000000
0!
0'
#470110000000
1!
b0 %
1'
b0 +
#470120000000
0!
0'
#470130000000
1!
1$
b1 %
1'
1*
b1 +
#470140000000
0!
0'
#470150000000
1!
b10 %
1'
b10 +
#470160000000
0!
0'
#470170000000
1!
b11 %
1'
b11 +
#470180000000
0!
0'
#470190000000
1!
b100 %
1'
b100 +
#470200000000
1"
1(
#470210000000
0!
0"
b100 &
0'
0(
b100 ,
#470220000000
1!
b101 %
1'
b101 +
#470230000000
0!
0'
#470240000000
1!
b110 %
1'
b110 +
#470250000000
0!
0'
#470260000000
1!
b111 %
1'
b111 +
#470270000000
0!
0'
#470280000000
1!
0$
b1000 %
1'
0*
b1000 +
#470290000000
0!
0'
#470300000000
1!
b1001 %
1'
b1001 +
#470310000000
0!
0'
#470320000000
1!
b0 %
1'
b0 +
#470330000000
0!
0'
#470340000000
1!
1$
b1 %
1'
1*
b1 +
#470350000000
0!
0'
#470360000000
1!
b10 %
1'
b10 +
#470370000000
0!
0'
#470380000000
1!
b11 %
1'
b11 +
#470390000000
0!
0'
#470400000000
1!
b100 %
1'
b100 +
#470410000000
0!
0'
#470420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#470430000000
0!
0'
#470440000000
1!
0$
b110 %
1'
0*
b110 +
#470450000000
0!
0'
#470460000000
1!
b111 %
1'
b111 +
#470470000000
0!
0'
#470480000000
1!
b1000 %
1'
b1000 +
#470490000000
0!
0'
#470500000000
1!
b1001 %
1'
b1001 +
#470510000000
0!
0'
#470520000000
1!
b0 %
1'
b0 +
#470530000000
0!
0'
#470540000000
1!
1$
b1 %
1'
1*
b1 +
#470550000000
0!
0'
#470560000000
1!
b10 %
1'
b10 +
#470570000000
0!
0'
#470580000000
1!
b11 %
1'
b11 +
#470590000000
0!
0'
#470600000000
1!
b100 %
1'
b100 +
#470610000000
0!
0'
#470620000000
1!
b101 %
1'
b101 +
#470630000000
1"
1(
#470640000000
0!
0"
b100 &
0'
0(
b100 ,
#470650000000
1!
b110 %
1'
b110 +
#470660000000
0!
0'
#470670000000
1!
b111 %
1'
b111 +
#470680000000
0!
0'
#470690000000
1!
0$
b1000 %
1'
0*
b1000 +
#470700000000
0!
0'
#470710000000
1!
b1001 %
1'
b1001 +
#470720000000
0!
0'
#470730000000
1!
b0 %
1'
b0 +
#470740000000
0!
0'
#470750000000
1!
1$
b1 %
1'
1*
b1 +
#470760000000
0!
0'
#470770000000
1!
b10 %
1'
b10 +
#470780000000
0!
0'
#470790000000
1!
b11 %
1'
b11 +
#470800000000
0!
0'
#470810000000
1!
b100 %
1'
b100 +
#470820000000
0!
0'
#470830000000
1!
b101 %
1'
b101 +
#470840000000
0!
0'
#470850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#470860000000
0!
0'
#470870000000
1!
b111 %
1'
b111 +
#470880000000
0!
0'
#470890000000
1!
b1000 %
1'
b1000 +
#470900000000
0!
0'
#470910000000
1!
b1001 %
1'
b1001 +
#470920000000
0!
0'
#470930000000
1!
b0 %
1'
b0 +
#470940000000
0!
0'
#470950000000
1!
1$
b1 %
1'
1*
b1 +
#470960000000
0!
0'
#470970000000
1!
b10 %
1'
b10 +
#470980000000
0!
0'
#470990000000
1!
b11 %
1'
b11 +
#471000000000
0!
0'
#471010000000
1!
b100 %
1'
b100 +
#471020000000
0!
0'
#471030000000
1!
b101 %
1'
b101 +
#471040000000
0!
0'
#471050000000
1!
0$
b110 %
1'
0*
b110 +
#471060000000
1"
1(
#471070000000
0!
0"
b100 &
0'
0(
b100 ,
#471080000000
1!
1$
b111 %
1'
1*
b111 +
#471090000000
0!
0'
#471100000000
1!
0$
b1000 %
1'
0*
b1000 +
#471110000000
0!
0'
#471120000000
1!
b1001 %
1'
b1001 +
#471130000000
0!
0'
#471140000000
1!
b0 %
1'
b0 +
#471150000000
0!
0'
#471160000000
1!
1$
b1 %
1'
1*
b1 +
#471170000000
0!
0'
#471180000000
1!
b10 %
1'
b10 +
#471190000000
0!
0'
#471200000000
1!
b11 %
1'
b11 +
#471210000000
0!
0'
#471220000000
1!
b100 %
1'
b100 +
#471230000000
0!
0'
#471240000000
1!
b101 %
1'
b101 +
#471250000000
0!
0'
#471260000000
1!
b110 %
1'
b110 +
#471270000000
0!
0'
#471280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#471290000000
0!
0'
#471300000000
1!
b1000 %
1'
b1000 +
#471310000000
0!
0'
#471320000000
1!
b1001 %
1'
b1001 +
#471330000000
0!
0'
#471340000000
1!
b0 %
1'
b0 +
#471350000000
0!
0'
#471360000000
1!
1$
b1 %
1'
1*
b1 +
#471370000000
0!
0'
#471380000000
1!
b10 %
1'
b10 +
#471390000000
0!
0'
#471400000000
1!
b11 %
1'
b11 +
#471410000000
0!
0'
#471420000000
1!
b100 %
1'
b100 +
#471430000000
0!
0'
#471440000000
1!
b101 %
1'
b101 +
#471450000000
0!
0'
#471460000000
1!
0$
b110 %
1'
0*
b110 +
#471470000000
0!
0'
#471480000000
1!
b111 %
1'
b111 +
#471490000000
1"
1(
#471500000000
0!
0"
b100 &
0'
0(
b100 ,
#471510000000
1!
b1000 %
1'
b1000 +
#471520000000
0!
0'
#471530000000
1!
b1001 %
1'
b1001 +
#471540000000
0!
0'
#471550000000
1!
b0 %
1'
b0 +
#471560000000
0!
0'
#471570000000
1!
1$
b1 %
1'
1*
b1 +
#471580000000
0!
0'
#471590000000
1!
b10 %
1'
b10 +
#471600000000
0!
0'
#471610000000
1!
b11 %
1'
b11 +
#471620000000
0!
0'
#471630000000
1!
b100 %
1'
b100 +
#471640000000
0!
0'
#471650000000
1!
b101 %
1'
b101 +
#471660000000
0!
0'
#471670000000
1!
b110 %
1'
b110 +
#471680000000
0!
0'
#471690000000
1!
b111 %
1'
b111 +
#471700000000
0!
0'
#471710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#471720000000
0!
0'
#471730000000
1!
b1001 %
1'
b1001 +
#471740000000
0!
0'
#471750000000
1!
b0 %
1'
b0 +
#471760000000
0!
0'
#471770000000
1!
1$
b1 %
1'
1*
b1 +
#471780000000
0!
0'
#471790000000
1!
b10 %
1'
b10 +
#471800000000
0!
0'
#471810000000
1!
b11 %
1'
b11 +
#471820000000
0!
0'
#471830000000
1!
b100 %
1'
b100 +
#471840000000
0!
0'
#471850000000
1!
b101 %
1'
b101 +
#471860000000
0!
0'
#471870000000
1!
0$
b110 %
1'
0*
b110 +
#471880000000
0!
0'
#471890000000
1!
b111 %
1'
b111 +
#471900000000
0!
0'
#471910000000
1!
b1000 %
1'
b1000 +
#471920000000
1"
1(
#471930000000
0!
0"
b100 &
0'
0(
b100 ,
#471940000000
1!
b1001 %
1'
b1001 +
#471950000000
0!
0'
#471960000000
1!
b0 %
1'
b0 +
#471970000000
0!
0'
#471980000000
1!
1$
b1 %
1'
1*
b1 +
#471990000000
0!
0'
#472000000000
1!
b10 %
1'
b10 +
#472010000000
0!
0'
#472020000000
1!
b11 %
1'
b11 +
#472030000000
0!
0'
#472040000000
1!
b100 %
1'
b100 +
#472050000000
0!
0'
#472060000000
1!
b101 %
1'
b101 +
#472070000000
0!
0'
#472080000000
1!
b110 %
1'
b110 +
#472090000000
0!
0'
#472100000000
1!
b111 %
1'
b111 +
#472110000000
0!
0'
#472120000000
1!
0$
b1000 %
1'
0*
b1000 +
#472130000000
0!
0'
#472140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#472150000000
0!
0'
#472160000000
1!
b0 %
1'
b0 +
#472170000000
0!
0'
#472180000000
1!
1$
b1 %
1'
1*
b1 +
#472190000000
0!
0'
#472200000000
1!
b10 %
1'
b10 +
#472210000000
0!
0'
#472220000000
1!
b11 %
1'
b11 +
#472230000000
0!
0'
#472240000000
1!
b100 %
1'
b100 +
#472250000000
0!
0'
#472260000000
1!
b101 %
1'
b101 +
#472270000000
0!
0'
#472280000000
1!
0$
b110 %
1'
0*
b110 +
#472290000000
0!
0'
#472300000000
1!
b111 %
1'
b111 +
#472310000000
0!
0'
#472320000000
1!
b1000 %
1'
b1000 +
#472330000000
0!
0'
#472340000000
1!
b1001 %
1'
b1001 +
#472350000000
1"
1(
#472360000000
0!
0"
b100 &
0'
0(
b100 ,
#472370000000
1!
b0 %
1'
b0 +
#472380000000
0!
0'
#472390000000
1!
1$
b1 %
1'
1*
b1 +
#472400000000
0!
0'
#472410000000
1!
b10 %
1'
b10 +
#472420000000
0!
0'
#472430000000
1!
b11 %
1'
b11 +
#472440000000
0!
0'
#472450000000
1!
b100 %
1'
b100 +
#472460000000
0!
0'
#472470000000
1!
b101 %
1'
b101 +
#472480000000
0!
0'
#472490000000
1!
b110 %
1'
b110 +
#472500000000
0!
0'
#472510000000
1!
b111 %
1'
b111 +
#472520000000
0!
0'
#472530000000
1!
0$
b1000 %
1'
0*
b1000 +
#472540000000
0!
0'
#472550000000
1!
b1001 %
1'
b1001 +
#472560000000
0!
0'
#472570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#472580000000
0!
0'
#472590000000
1!
1$
b1 %
1'
1*
b1 +
#472600000000
0!
0'
#472610000000
1!
b10 %
1'
b10 +
#472620000000
0!
0'
#472630000000
1!
b11 %
1'
b11 +
#472640000000
0!
0'
#472650000000
1!
b100 %
1'
b100 +
#472660000000
0!
0'
#472670000000
1!
b101 %
1'
b101 +
#472680000000
0!
0'
#472690000000
1!
0$
b110 %
1'
0*
b110 +
#472700000000
0!
0'
#472710000000
1!
b111 %
1'
b111 +
#472720000000
0!
0'
#472730000000
1!
b1000 %
1'
b1000 +
#472740000000
0!
0'
#472750000000
1!
b1001 %
1'
b1001 +
#472760000000
0!
0'
#472770000000
1!
b0 %
1'
b0 +
#472780000000
1"
1(
#472790000000
0!
0"
b100 &
0'
0(
b100 ,
#472800000000
1!
1$
b1 %
1'
1*
b1 +
#472810000000
0!
0'
#472820000000
1!
b10 %
1'
b10 +
#472830000000
0!
0'
#472840000000
1!
b11 %
1'
b11 +
#472850000000
0!
0'
#472860000000
1!
b100 %
1'
b100 +
#472870000000
0!
0'
#472880000000
1!
b101 %
1'
b101 +
#472890000000
0!
0'
#472900000000
1!
b110 %
1'
b110 +
#472910000000
0!
0'
#472920000000
1!
b111 %
1'
b111 +
#472930000000
0!
0'
#472940000000
1!
0$
b1000 %
1'
0*
b1000 +
#472950000000
0!
0'
#472960000000
1!
b1001 %
1'
b1001 +
#472970000000
0!
0'
#472980000000
1!
b0 %
1'
b0 +
#472990000000
0!
0'
#473000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#473010000000
0!
0'
#473020000000
1!
b10 %
1'
b10 +
#473030000000
0!
0'
#473040000000
1!
b11 %
1'
b11 +
#473050000000
0!
0'
#473060000000
1!
b100 %
1'
b100 +
#473070000000
0!
0'
#473080000000
1!
b101 %
1'
b101 +
#473090000000
0!
0'
#473100000000
1!
0$
b110 %
1'
0*
b110 +
#473110000000
0!
0'
#473120000000
1!
b111 %
1'
b111 +
#473130000000
0!
0'
#473140000000
1!
b1000 %
1'
b1000 +
#473150000000
0!
0'
#473160000000
1!
b1001 %
1'
b1001 +
#473170000000
0!
0'
#473180000000
1!
b0 %
1'
b0 +
#473190000000
0!
0'
#473200000000
1!
1$
b1 %
1'
1*
b1 +
#473210000000
1"
1(
#473220000000
0!
0"
b100 &
0'
0(
b100 ,
#473230000000
1!
b10 %
1'
b10 +
#473240000000
0!
0'
#473250000000
1!
b11 %
1'
b11 +
#473260000000
0!
0'
#473270000000
1!
b100 %
1'
b100 +
#473280000000
0!
0'
#473290000000
1!
b101 %
1'
b101 +
#473300000000
0!
0'
#473310000000
1!
b110 %
1'
b110 +
#473320000000
0!
0'
#473330000000
1!
b111 %
1'
b111 +
#473340000000
0!
0'
#473350000000
1!
0$
b1000 %
1'
0*
b1000 +
#473360000000
0!
0'
#473370000000
1!
b1001 %
1'
b1001 +
#473380000000
0!
0'
#473390000000
1!
b0 %
1'
b0 +
#473400000000
0!
0'
#473410000000
1!
1$
b1 %
1'
1*
b1 +
#473420000000
0!
0'
#473430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#473440000000
0!
0'
#473450000000
1!
b11 %
1'
b11 +
#473460000000
0!
0'
#473470000000
1!
b100 %
1'
b100 +
#473480000000
0!
0'
#473490000000
1!
b101 %
1'
b101 +
#473500000000
0!
0'
#473510000000
1!
0$
b110 %
1'
0*
b110 +
#473520000000
0!
0'
#473530000000
1!
b111 %
1'
b111 +
#473540000000
0!
0'
#473550000000
1!
b1000 %
1'
b1000 +
#473560000000
0!
0'
#473570000000
1!
b1001 %
1'
b1001 +
#473580000000
0!
0'
#473590000000
1!
b0 %
1'
b0 +
#473600000000
0!
0'
#473610000000
1!
1$
b1 %
1'
1*
b1 +
#473620000000
0!
0'
#473630000000
1!
b10 %
1'
b10 +
#473640000000
1"
1(
#473650000000
0!
0"
b100 &
0'
0(
b100 ,
#473660000000
1!
b11 %
1'
b11 +
#473670000000
0!
0'
#473680000000
1!
b100 %
1'
b100 +
#473690000000
0!
0'
#473700000000
1!
b101 %
1'
b101 +
#473710000000
0!
0'
#473720000000
1!
b110 %
1'
b110 +
#473730000000
0!
0'
#473740000000
1!
b111 %
1'
b111 +
#473750000000
0!
0'
#473760000000
1!
0$
b1000 %
1'
0*
b1000 +
#473770000000
0!
0'
#473780000000
1!
b1001 %
1'
b1001 +
#473790000000
0!
0'
#473800000000
1!
b0 %
1'
b0 +
#473810000000
0!
0'
#473820000000
1!
1$
b1 %
1'
1*
b1 +
#473830000000
0!
0'
#473840000000
1!
b10 %
1'
b10 +
#473850000000
0!
0'
#473860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#473870000000
0!
0'
#473880000000
1!
b100 %
1'
b100 +
#473890000000
0!
0'
#473900000000
1!
b101 %
1'
b101 +
#473910000000
0!
0'
#473920000000
1!
0$
b110 %
1'
0*
b110 +
#473930000000
0!
0'
#473940000000
1!
b111 %
1'
b111 +
#473950000000
0!
0'
#473960000000
1!
b1000 %
1'
b1000 +
#473970000000
0!
0'
#473980000000
1!
b1001 %
1'
b1001 +
#473990000000
0!
0'
#474000000000
1!
b0 %
1'
b0 +
#474010000000
0!
0'
#474020000000
1!
1$
b1 %
1'
1*
b1 +
#474030000000
0!
0'
#474040000000
1!
b10 %
1'
b10 +
#474050000000
0!
0'
#474060000000
1!
b11 %
1'
b11 +
#474070000000
1"
1(
#474080000000
0!
0"
b100 &
0'
0(
b100 ,
#474090000000
1!
b100 %
1'
b100 +
#474100000000
0!
0'
#474110000000
1!
b101 %
1'
b101 +
#474120000000
0!
0'
#474130000000
1!
b110 %
1'
b110 +
#474140000000
0!
0'
#474150000000
1!
b111 %
1'
b111 +
#474160000000
0!
0'
#474170000000
1!
0$
b1000 %
1'
0*
b1000 +
#474180000000
0!
0'
#474190000000
1!
b1001 %
1'
b1001 +
#474200000000
0!
0'
#474210000000
1!
b0 %
1'
b0 +
#474220000000
0!
0'
#474230000000
1!
1$
b1 %
1'
1*
b1 +
#474240000000
0!
0'
#474250000000
1!
b10 %
1'
b10 +
#474260000000
0!
0'
#474270000000
1!
b11 %
1'
b11 +
#474280000000
0!
0'
#474290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#474300000000
0!
0'
#474310000000
1!
b101 %
1'
b101 +
#474320000000
0!
0'
#474330000000
1!
0$
b110 %
1'
0*
b110 +
#474340000000
0!
0'
#474350000000
1!
b111 %
1'
b111 +
#474360000000
0!
0'
#474370000000
1!
b1000 %
1'
b1000 +
#474380000000
0!
0'
#474390000000
1!
b1001 %
1'
b1001 +
#474400000000
0!
0'
#474410000000
1!
b0 %
1'
b0 +
#474420000000
0!
0'
#474430000000
1!
1$
b1 %
1'
1*
b1 +
#474440000000
0!
0'
#474450000000
1!
b10 %
1'
b10 +
#474460000000
0!
0'
#474470000000
1!
b11 %
1'
b11 +
#474480000000
0!
0'
#474490000000
1!
b100 %
1'
b100 +
#474500000000
1"
1(
#474510000000
0!
0"
b100 &
0'
0(
b100 ,
#474520000000
1!
b101 %
1'
b101 +
#474530000000
0!
0'
#474540000000
1!
b110 %
1'
b110 +
#474550000000
0!
0'
#474560000000
1!
b111 %
1'
b111 +
#474570000000
0!
0'
#474580000000
1!
0$
b1000 %
1'
0*
b1000 +
#474590000000
0!
0'
#474600000000
1!
b1001 %
1'
b1001 +
#474610000000
0!
0'
#474620000000
1!
b0 %
1'
b0 +
#474630000000
0!
0'
#474640000000
1!
1$
b1 %
1'
1*
b1 +
#474650000000
0!
0'
#474660000000
1!
b10 %
1'
b10 +
#474670000000
0!
0'
#474680000000
1!
b11 %
1'
b11 +
#474690000000
0!
0'
#474700000000
1!
b100 %
1'
b100 +
#474710000000
0!
0'
#474720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#474730000000
0!
0'
#474740000000
1!
0$
b110 %
1'
0*
b110 +
#474750000000
0!
0'
#474760000000
1!
b111 %
1'
b111 +
#474770000000
0!
0'
#474780000000
1!
b1000 %
1'
b1000 +
#474790000000
0!
0'
#474800000000
1!
b1001 %
1'
b1001 +
#474810000000
0!
0'
#474820000000
1!
b0 %
1'
b0 +
#474830000000
0!
0'
#474840000000
1!
1$
b1 %
1'
1*
b1 +
#474850000000
0!
0'
#474860000000
1!
b10 %
1'
b10 +
#474870000000
0!
0'
#474880000000
1!
b11 %
1'
b11 +
#474890000000
0!
0'
#474900000000
1!
b100 %
1'
b100 +
#474910000000
0!
0'
#474920000000
1!
b101 %
1'
b101 +
#474930000000
1"
1(
#474940000000
0!
0"
b100 &
0'
0(
b100 ,
#474950000000
1!
b110 %
1'
b110 +
#474960000000
0!
0'
#474970000000
1!
b111 %
1'
b111 +
#474980000000
0!
0'
#474990000000
1!
0$
b1000 %
1'
0*
b1000 +
#475000000000
0!
0'
#475010000000
1!
b1001 %
1'
b1001 +
#475020000000
0!
0'
#475030000000
1!
b0 %
1'
b0 +
#475040000000
0!
0'
#475050000000
1!
1$
b1 %
1'
1*
b1 +
#475060000000
0!
0'
#475070000000
1!
b10 %
1'
b10 +
#475080000000
0!
0'
#475090000000
1!
b11 %
1'
b11 +
#475100000000
0!
0'
#475110000000
1!
b100 %
1'
b100 +
#475120000000
0!
0'
#475130000000
1!
b101 %
1'
b101 +
#475140000000
0!
0'
#475150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#475160000000
0!
0'
#475170000000
1!
b111 %
1'
b111 +
#475180000000
0!
0'
#475190000000
1!
b1000 %
1'
b1000 +
#475200000000
0!
0'
#475210000000
1!
b1001 %
1'
b1001 +
#475220000000
0!
0'
#475230000000
1!
b0 %
1'
b0 +
#475240000000
0!
0'
#475250000000
1!
1$
b1 %
1'
1*
b1 +
#475260000000
0!
0'
#475270000000
1!
b10 %
1'
b10 +
#475280000000
0!
0'
#475290000000
1!
b11 %
1'
b11 +
#475300000000
0!
0'
#475310000000
1!
b100 %
1'
b100 +
#475320000000
0!
0'
#475330000000
1!
b101 %
1'
b101 +
#475340000000
0!
0'
#475350000000
1!
0$
b110 %
1'
0*
b110 +
#475360000000
1"
1(
#475370000000
0!
0"
b100 &
0'
0(
b100 ,
#475380000000
1!
1$
b111 %
1'
1*
b111 +
#475390000000
0!
0'
#475400000000
1!
0$
b1000 %
1'
0*
b1000 +
#475410000000
0!
0'
#475420000000
1!
b1001 %
1'
b1001 +
#475430000000
0!
0'
#475440000000
1!
b0 %
1'
b0 +
#475450000000
0!
0'
#475460000000
1!
1$
b1 %
1'
1*
b1 +
#475470000000
0!
0'
#475480000000
1!
b10 %
1'
b10 +
#475490000000
0!
0'
#475500000000
1!
b11 %
1'
b11 +
#475510000000
0!
0'
#475520000000
1!
b100 %
1'
b100 +
#475530000000
0!
0'
#475540000000
1!
b101 %
1'
b101 +
#475550000000
0!
0'
#475560000000
1!
b110 %
1'
b110 +
#475570000000
0!
0'
#475580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#475590000000
0!
0'
#475600000000
1!
b1000 %
1'
b1000 +
#475610000000
0!
0'
#475620000000
1!
b1001 %
1'
b1001 +
#475630000000
0!
0'
#475640000000
1!
b0 %
1'
b0 +
#475650000000
0!
0'
#475660000000
1!
1$
b1 %
1'
1*
b1 +
#475670000000
0!
0'
#475680000000
1!
b10 %
1'
b10 +
#475690000000
0!
0'
#475700000000
1!
b11 %
1'
b11 +
#475710000000
0!
0'
#475720000000
1!
b100 %
1'
b100 +
#475730000000
0!
0'
#475740000000
1!
b101 %
1'
b101 +
#475750000000
0!
0'
#475760000000
1!
0$
b110 %
1'
0*
b110 +
#475770000000
0!
0'
#475780000000
1!
b111 %
1'
b111 +
#475790000000
1"
1(
#475800000000
0!
0"
b100 &
0'
0(
b100 ,
#475810000000
1!
b1000 %
1'
b1000 +
#475820000000
0!
0'
#475830000000
1!
b1001 %
1'
b1001 +
#475840000000
0!
0'
#475850000000
1!
b0 %
1'
b0 +
#475860000000
0!
0'
#475870000000
1!
1$
b1 %
1'
1*
b1 +
#475880000000
0!
0'
#475890000000
1!
b10 %
1'
b10 +
#475900000000
0!
0'
#475910000000
1!
b11 %
1'
b11 +
#475920000000
0!
0'
#475930000000
1!
b100 %
1'
b100 +
#475940000000
0!
0'
#475950000000
1!
b101 %
1'
b101 +
#475960000000
0!
0'
#475970000000
1!
b110 %
1'
b110 +
#475980000000
0!
0'
#475990000000
1!
b111 %
1'
b111 +
#476000000000
0!
0'
#476010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#476020000000
0!
0'
#476030000000
1!
b1001 %
1'
b1001 +
#476040000000
0!
0'
#476050000000
1!
b0 %
1'
b0 +
#476060000000
0!
0'
#476070000000
1!
1$
b1 %
1'
1*
b1 +
#476080000000
0!
0'
#476090000000
1!
b10 %
1'
b10 +
#476100000000
0!
0'
#476110000000
1!
b11 %
1'
b11 +
#476120000000
0!
0'
#476130000000
1!
b100 %
1'
b100 +
#476140000000
0!
0'
#476150000000
1!
b101 %
1'
b101 +
#476160000000
0!
0'
#476170000000
1!
0$
b110 %
1'
0*
b110 +
#476180000000
0!
0'
#476190000000
1!
b111 %
1'
b111 +
#476200000000
0!
0'
#476210000000
1!
b1000 %
1'
b1000 +
#476220000000
1"
1(
#476230000000
0!
0"
b100 &
0'
0(
b100 ,
#476240000000
1!
b1001 %
1'
b1001 +
#476250000000
0!
0'
#476260000000
1!
b0 %
1'
b0 +
#476270000000
0!
0'
#476280000000
1!
1$
b1 %
1'
1*
b1 +
#476290000000
0!
0'
#476300000000
1!
b10 %
1'
b10 +
#476310000000
0!
0'
#476320000000
1!
b11 %
1'
b11 +
#476330000000
0!
0'
#476340000000
1!
b100 %
1'
b100 +
#476350000000
0!
0'
#476360000000
1!
b101 %
1'
b101 +
#476370000000
0!
0'
#476380000000
1!
b110 %
1'
b110 +
#476390000000
0!
0'
#476400000000
1!
b111 %
1'
b111 +
#476410000000
0!
0'
#476420000000
1!
0$
b1000 %
1'
0*
b1000 +
#476430000000
0!
0'
#476440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#476450000000
0!
0'
#476460000000
1!
b0 %
1'
b0 +
#476470000000
0!
0'
#476480000000
1!
1$
b1 %
1'
1*
b1 +
#476490000000
0!
0'
#476500000000
1!
b10 %
1'
b10 +
#476510000000
0!
0'
#476520000000
1!
b11 %
1'
b11 +
#476530000000
0!
0'
#476540000000
1!
b100 %
1'
b100 +
#476550000000
0!
0'
#476560000000
1!
b101 %
1'
b101 +
#476570000000
0!
0'
#476580000000
1!
0$
b110 %
1'
0*
b110 +
#476590000000
0!
0'
#476600000000
1!
b111 %
1'
b111 +
#476610000000
0!
0'
#476620000000
1!
b1000 %
1'
b1000 +
#476630000000
0!
0'
#476640000000
1!
b1001 %
1'
b1001 +
#476650000000
1"
1(
#476660000000
0!
0"
b100 &
0'
0(
b100 ,
#476670000000
1!
b0 %
1'
b0 +
#476680000000
0!
0'
#476690000000
1!
1$
b1 %
1'
1*
b1 +
#476700000000
0!
0'
#476710000000
1!
b10 %
1'
b10 +
#476720000000
0!
0'
#476730000000
1!
b11 %
1'
b11 +
#476740000000
0!
0'
#476750000000
1!
b100 %
1'
b100 +
#476760000000
0!
0'
#476770000000
1!
b101 %
1'
b101 +
#476780000000
0!
0'
#476790000000
1!
b110 %
1'
b110 +
#476800000000
0!
0'
#476810000000
1!
b111 %
1'
b111 +
#476820000000
0!
0'
#476830000000
1!
0$
b1000 %
1'
0*
b1000 +
#476840000000
0!
0'
#476850000000
1!
b1001 %
1'
b1001 +
#476860000000
0!
0'
#476870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#476880000000
0!
0'
#476890000000
1!
1$
b1 %
1'
1*
b1 +
#476900000000
0!
0'
#476910000000
1!
b10 %
1'
b10 +
#476920000000
0!
0'
#476930000000
1!
b11 %
1'
b11 +
#476940000000
0!
0'
#476950000000
1!
b100 %
1'
b100 +
#476960000000
0!
0'
#476970000000
1!
b101 %
1'
b101 +
#476980000000
0!
0'
#476990000000
1!
0$
b110 %
1'
0*
b110 +
#477000000000
0!
0'
#477010000000
1!
b111 %
1'
b111 +
#477020000000
0!
0'
#477030000000
1!
b1000 %
1'
b1000 +
#477040000000
0!
0'
#477050000000
1!
b1001 %
1'
b1001 +
#477060000000
0!
0'
#477070000000
1!
b0 %
1'
b0 +
#477080000000
1"
1(
#477090000000
0!
0"
b100 &
0'
0(
b100 ,
#477100000000
1!
1$
b1 %
1'
1*
b1 +
#477110000000
0!
0'
#477120000000
1!
b10 %
1'
b10 +
#477130000000
0!
0'
#477140000000
1!
b11 %
1'
b11 +
#477150000000
0!
0'
#477160000000
1!
b100 %
1'
b100 +
#477170000000
0!
0'
#477180000000
1!
b101 %
1'
b101 +
#477190000000
0!
0'
#477200000000
1!
b110 %
1'
b110 +
#477210000000
0!
0'
#477220000000
1!
b111 %
1'
b111 +
#477230000000
0!
0'
#477240000000
1!
0$
b1000 %
1'
0*
b1000 +
#477250000000
0!
0'
#477260000000
1!
b1001 %
1'
b1001 +
#477270000000
0!
0'
#477280000000
1!
b0 %
1'
b0 +
#477290000000
0!
0'
#477300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#477310000000
0!
0'
#477320000000
1!
b10 %
1'
b10 +
#477330000000
0!
0'
#477340000000
1!
b11 %
1'
b11 +
#477350000000
0!
0'
#477360000000
1!
b100 %
1'
b100 +
#477370000000
0!
0'
#477380000000
1!
b101 %
1'
b101 +
#477390000000
0!
0'
#477400000000
1!
0$
b110 %
1'
0*
b110 +
#477410000000
0!
0'
#477420000000
1!
b111 %
1'
b111 +
#477430000000
0!
0'
#477440000000
1!
b1000 %
1'
b1000 +
#477450000000
0!
0'
#477460000000
1!
b1001 %
1'
b1001 +
#477470000000
0!
0'
#477480000000
1!
b0 %
1'
b0 +
#477490000000
0!
0'
#477500000000
1!
1$
b1 %
1'
1*
b1 +
#477510000000
1"
1(
#477520000000
0!
0"
b100 &
0'
0(
b100 ,
#477530000000
1!
b10 %
1'
b10 +
#477540000000
0!
0'
#477550000000
1!
b11 %
1'
b11 +
#477560000000
0!
0'
#477570000000
1!
b100 %
1'
b100 +
#477580000000
0!
0'
#477590000000
1!
b101 %
1'
b101 +
#477600000000
0!
0'
#477610000000
1!
b110 %
1'
b110 +
#477620000000
0!
0'
#477630000000
1!
b111 %
1'
b111 +
#477640000000
0!
0'
#477650000000
1!
0$
b1000 %
1'
0*
b1000 +
#477660000000
0!
0'
#477670000000
1!
b1001 %
1'
b1001 +
#477680000000
0!
0'
#477690000000
1!
b0 %
1'
b0 +
#477700000000
0!
0'
#477710000000
1!
1$
b1 %
1'
1*
b1 +
#477720000000
0!
0'
#477730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#477740000000
0!
0'
#477750000000
1!
b11 %
1'
b11 +
#477760000000
0!
0'
#477770000000
1!
b100 %
1'
b100 +
#477780000000
0!
0'
#477790000000
1!
b101 %
1'
b101 +
#477800000000
0!
0'
#477810000000
1!
0$
b110 %
1'
0*
b110 +
#477820000000
0!
0'
#477830000000
1!
b111 %
1'
b111 +
#477840000000
0!
0'
#477850000000
1!
b1000 %
1'
b1000 +
#477860000000
0!
0'
#477870000000
1!
b1001 %
1'
b1001 +
#477880000000
0!
0'
#477890000000
1!
b0 %
1'
b0 +
#477900000000
0!
0'
#477910000000
1!
1$
b1 %
1'
1*
b1 +
#477920000000
0!
0'
#477930000000
1!
b10 %
1'
b10 +
#477940000000
1"
1(
#477950000000
0!
0"
b100 &
0'
0(
b100 ,
#477960000000
1!
b11 %
1'
b11 +
#477970000000
0!
0'
#477980000000
1!
b100 %
1'
b100 +
#477990000000
0!
0'
#478000000000
1!
b101 %
1'
b101 +
#478010000000
0!
0'
#478020000000
1!
b110 %
1'
b110 +
#478030000000
0!
0'
#478040000000
1!
b111 %
1'
b111 +
#478050000000
0!
0'
#478060000000
1!
0$
b1000 %
1'
0*
b1000 +
#478070000000
0!
0'
#478080000000
1!
b1001 %
1'
b1001 +
#478090000000
0!
0'
#478100000000
1!
b0 %
1'
b0 +
#478110000000
0!
0'
#478120000000
1!
1$
b1 %
1'
1*
b1 +
#478130000000
0!
0'
#478140000000
1!
b10 %
1'
b10 +
#478150000000
0!
0'
#478160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#478170000000
0!
0'
#478180000000
1!
b100 %
1'
b100 +
#478190000000
0!
0'
#478200000000
1!
b101 %
1'
b101 +
#478210000000
0!
0'
#478220000000
1!
0$
b110 %
1'
0*
b110 +
#478230000000
0!
0'
#478240000000
1!
b111 %
1'
b111 +
#478250000000
0!
0'
#478260000000
1!
b1000 %
1'
b1000 +
#478270000000
0!
0'
#478280000000
1!
b1001 %
1'
b1001 +
#478290000000
0!
0'
#478300000000
1!
b0 %
1'
b0 +
#478310000000
0!
0'
#478320000000
1!
1$
b1 %
1'
1*
b1 +
#478330000000
0!
0'
#478340000000
1!
b10 %
1'
b10 +
#478350000000
0!
0'
#478360000000
1!
b11 %
1'
b11 +
#478370000000
1"
1(
#478380000000
0!
0"
b100 &
0'
0(
b100 ,
#478390000000
1!
b100 %
1'
b100 +
#478400000000
0!
0'
#478410000000
1!
b101 %
1'
b101 +
#478420000000
0!
0'
#478430000000
1!
b110 %
1'
b110 +
#478440000000
0!
0'
#478450000000
1!
b111 %
1'
b111 +
#478460000000
0!
0'
#478470000000
1!
0$
b1000 %
1'
0*
b1000 +
#478480000000
0!
0'
#478490000000
1!
b1001 %
1'
b1001 +
#478500000000
0!
0'
#478510000000
1!
b0 %
1'
b0 +
#478520000000
0!
0'
#478530000000
1!
1$
b1 %
1'
1*
b1 +
#478540000000
0!
0'
#478550000000
1!
b10 %
1'
b10 +
#478560000000
0!
0'
#478570000000
1!
b11 %
1'
b11 +
#478580000000
0!
0'
#478590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#478600000000
0!
0'
#478610000000
1!
b101 %
1'
b101 +
#478620000000
0!
0'
#478630000000
1!
0$
b110 %
1'
0*
b110 +
#478640000000
0!
0'
#478650000000
1!
b111 %
1'
b111 +
#478660000000
0!
0'
#478670000000
1!
b1000 %
1'
b1000 +
#478680000000
0!
0'
#478690000000
1!
b1001 %
1'
b1001 +
#478700000000
0!
0'
#478710000000
1!
b0 %
1'
b0 +
#478720000000
0!
0'
#478730000000
1!
1$
b1 %
1'
1*
b1 +
#478740000000
0!
0'
#478750000000
1!
b10 %
1'
b10 +
#478760000000
0!
0'
#478770000000
1!
b11 %
1'
b11 +
#478780000000
0!
0'
#478790000000
1!
b100 %
1'
b100 +
#478800000000
1"
1(
#478810000000
0!
0"
b100 &
0'
0(
b100 ,
#478820000000
1!
b101 %
1'
b101 +
#478830000000
0!
0'
#478840000000
1!
b110 %
1'
b110 +
#478850000000
0!
0'
#478860000000
1!
b111 %
1'
b111 +
#478870000000
0!
0'
#478880000000
1!
0$
b1000 %
1'
0*
b1000 +
#478890000000
0!
0'
#478900000000
1!
b1001 %
1'
b1001 +
#478910000000
0!
0'
#478920000000
1!
b0 %
1'
b0 +
#478930000000
0!
0'
#478940000000
1!
1$
b1 %
1'
1*
b1 +
#478950000000
0!
0'
#478960000000
1!
b10 %
1'
b10 +
#478970000000
0!
0'
#478980000000
1!
b11 %
1'
b11 +
#478990000000
0!
0'
#479000000000
1!
b100 %
1'
b100 +
#479010000000
0!
0'
#479020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#479030000000
0!
0'
#479040000000
1!
0$
b110 %
1'
0*
b110 +
#479050000000
0!
0'
#479060000000
1!
b111 %
1'
b111 +
#479070000000
0!
0'
#479080000000
1!
b1000 %
1'
b1000 +
#479090000000
0!
0'
#479100000000
1!
b1001 %
1'
b1001 +
#479110000000
0!
0'
#479120000000
1!
b0 %
1'
b0 +
#479130000000
0!
0'
#479140000000
1!
1$
b1 %
1'
1*
b1 +
#479150000000
0!
0'
#479160000000
1!
b10 %
1'
b10 +
#479170000000
0!
0'
#479180000000
1!
b11 %
1'
b11 +
#479190000000
0!
0'
#479200000000
1!
b100 %
1'
b100 +
#479210000000
0!
0'
#479220000000
1!
b101 %
1'
b101 +
#479230000000
1"
1(
#479240000000
0!
0"
b100 &
0'
0(
b100 ,
#479250000000
1!
b110 %
1'
b110 +
#479260000000
0!
0'
#479270000000
1!
b111 %
1'
b111 +
#479280000000
0!
0'
#479290000000
1!
0$
b1000 %
1'
0*
b1000 +
#479300000000
0!
0'
#479310000000
1!
b1001 %
1'
b1001 +
#479320000000
0!
0'
#479330000000
1!
b0 %
1'
b0 +
#479340000000
0!
0'
#479350000000
1!
1$
b1 %
1'
1*
b1 +
#479360000000
0!
0'
#479370000000
1!
b10 %
1'
b10 +
#479380000000
0!
0'
#479390000000
1!
b11 %
1'
b11 +
#479400000000
0!
0'
#479410000000
1!
b100 %
1'
b100 +
#479420000000
0!
0'
#479430000000
1!
b101 %
1'
b101 +
#479440000000
0!
0'
#479450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#479460000000
0!
0'
#479470000000
1!
b111 %
1'
b111 +
#479480000000
0!
0'
#479490000000
1!
b1000 %
1'
b1000 +
#479500000000
0!
0'
#479510000000
1!
b1001 %
1'
b1001 +
#479520000000
0!
0'
#479530000000
1!
b0 %
1'
b0 +
#479540000000
0!
0'
#479550000000
1!
1$
b1 %
1'
1*
b1 +
#479560000000
0!
0'
#479570000000
1!
b10 %
1'
b10 +
#479580000000
0!
0'
#479590000000
1!
b11 %
1'
b11 +
#479600000000
0!
0'
#479610000000
1!
b100 %
1'
b100 +
#479620000000
0!
0'
#479630000000
1!
b101 %
1'
b101 +
#479640000000
0!
0'
#479650000000
1!
0$
b110 %
1'
0*
b110 +
#479660000000
1"
1(
#479670000000
0!
0"
b100 &
0'
0(
b100 ,
#479680000000
1!
1$
b111 %
1'
1*
b111 +
#479690000000
0!
0'
#479700000000
1!
0$
b1000 %
1'
0*
b1000 +
#479710000000
0!
0'
#479720000000
1!
b1001 %
1'
b1001 +
#479730000000
0!
0'
#479740000000
1!
b0 %
1'
b0 +
#479750000000
0!
0'
#479760000000
1!
1$
b1 %
1'
1*
b1 +
#479770000000
0!
0'
#479780000000
1!
b10 %
1'
b10 +
#479790000000
0!
0'
#479800000000
1!
b11 %
1'
b11 +
#479810000000
0!
0'
#479820000000
1!
b100 %
1'
b100 +
#479830000000
0!
0'
#479840000000
1!
b101 %
1'
b101 +
#479850000000
0!
0'
#479860000000
1!
b110 %
1'
b110 +
#479870000000
0!
0'
#479880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#479890000000
0!
0'
#479900000000
1!
b1000 %
1'
b1000 +
#479910000000
0!
0'
#479920000000
1!
b1001 %
1'
b1001 +
#479930000000
0!
0'
#479940000000
1!
b0 %
1'
b0 +
#479950000000
0!
0'
#479960000000
1!
1$
b1 %
1'
1*
b1 +
#479970000000
0!
0'
#479980000000
1!
b10 %
1'
b10 +
#479990000000
0!
0'
#480000000000
1!
b11 %
1'
b11 +
#480010000000
0!
0'
#480020000000
1!
b100 %
1'
b100 +
#480030000000
0!
0'
#480040000000
1!
b101 %
1'
b101 +
#480050000000
0!
0'
#480060000000
1!
0$
b110 %
1'
0*
b110 +
#480070000000
0!
0'
#480080000000
1!
b111 %
1'
b111 +
#480090000000
1"
1(
#480100000000
0!
0"
b100 &
0'
0(
b100 ,
#480110000000
1!
b1000 %
1'
b1000 +
#480120000000
0!
0'
#480130000000
1!
b1001 %
1'
b1001 +
#480140000000
0!
0'
#480150000000
1!
b0 %
1'
b0 +
#480160000000
0!
0'
#480170000000
1!
1$
b1 %
1'
1*
b1 +
#480180000000
0!
0'
#480190000000
1!
b10 %
1'
b10 +
#480200000000
0!
0'
#480210000000
1!
b11 %
1'
b11 +
#480220000000
0!
0'
#480230000000
1!
b100 %
1'
b100 +
#480240000000
0!
0'
#480250000000
1!
b101 %
1'
b101 +
#480260000000
0!
0'
#480270000000
1!
b110 %
1'
b110 +
#480280000000
0!
0'
#480290000000
1!
b111 %
1'
b111 +
#480300000000
0!
0'
#480310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#480320000000
0!
0'
#480330000000
1!
b1001 %
1'
b1001 +
#480340000000
0!
0'
#480350000000
1!
b0 %
1'
b0 +
#480360000000
0!
0'
#480370000000
1!
1$
b1 %
1'
1*
b1 +
#480380000000
0!
0'
#480390000000
1!
b10 %
1'
b10 +
#480400000000
0!
0'
#480410000000
1!
b11 %
1'
b11 +
#480420000000
0!
0'
#480430000000
1!
b100 %
1'
b100 +
#480440000000
0!
0'
#480450000000
1!
b101 %
1'
b101 +
#480460000000
0!
0'
#480470000000
1!
0$
b110 %
1'
0*
b110 +
#480480000000
0!
0'
#480490000000
1!
b111 %
1'
b111 +
#480500000000
0!
0'
#480510000000
1!
b1000 %
1'
b1000 +
#480520000000
1"
1(
#480530000000
0!
0"
b100 &
0'
0(
b100 ,
#480540000000
1!
b1001 %
1'
b1001 +
#480550000000
0!
0'
#480560000000
1!
b0 %
1'
b0 +
#480570000000
0!
0'
#480580000000
1!
1$
b1 %
1'
1*
b1 +
#480590000000
0!
0'
#480600000000
1!
b10 %
1'
b10 +
#480610000000
0!
0'
#480620000000
1!
b11 %
1'
b11 +
#480630000000
0!
0'
#480640000000
1!
b100 %
1'
b100 +
#480650000000
0!
0'
#480660000000
1!
b101 %
1'
b101 +
#480670000000
0!
0'
#480680000000
1!
b110 %
1'
b110 +
#480690000000
0!
0'
#480700000000
1!
b111 %
1'
b111 +
#480710000000
0!
0'
#480720000000
1!
0$
b1000 %
1'
0*
b1000 +
#480730000000
0!
0'
#480740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#480750000000
0!
0'
#480760000000
1!
b0 %
1'
b0 +
#480770000000
0!
0'
#480780000000
1!
1$
b1 %
1'
1*
b1 +
#480790000000
0!
0'
#480800000000
1!
b10 %
1'
b10 +
#480810000000
0!
0'
#480820000000
1!
b11 %
1'
b11 +
#480830000000
0!
0'
#480840000000
1!
b100 %
1'
b100 +
#480850000000
0!
0'
#480860000000
1!
b101 %
1'
b101 +
#480870000000
0!
0'
#480880000000
1!
0$
b110 %
1'
0*
b110 +
#480890000000
0!
0'
#480900000000
1!
b111 %
1'
b111 +
#480910000000
0!
0'
#480920000000
1!
b1000 %
1'
b1000 +
#480930000000
0!
0'
#480940000000
1!
b1001 %
1'
b1001 +
#480950000000
1"
1(
#480960000000
0!
0"
b100 &
0'
0(
b100 ,
#480970000000
1!
b0 %
1'
b0 +
#480980000000
0!
0'
#480990000000
1!
1$
b1 %
1'
1*
b1 +
#481000000000
0!
0'
#481010000000
1!
b10 %
1'
b10 +
#481020000000
0!
0'
#481030000000
1!
b11 %
1'
b11 +
#481040000000
0!
0'
#481050000000
1!
b100 %
1'
b100 +
#481060000000
0!
0'
#481070000000
1!
b101 %
1'
b101 +
#481080000000
0!
0'
#481090000000
1!
b110 %
1'
b110 +
#481100000000
0!
0'
#481110000000
1!
b111 %
1'
b111 +
#481120000000
0!
0'
#481130000000
1!
0$
b1000 %
1'
0*
b1000 +
#481140000000
0!
0'
#481150000000
1!
b1001 %
1'
b1001 +
#481160000000
0!
0'
#481170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#481180000000
0!
0'
#481190000000
1!
1$
b1 %
1'
1*
b1 +
#481200000000
0!
0'
#481210000000
1!
b10 %
1'
b10 +
#481220000000
0!
0'
#481230000000
1!
b11 %
1'
b11 +
#481240000000
0!
0'
#481250000000
1!
b100 %
1'
b100 +
#481260000000
0!
0'
#481270000000
1!
b101 %
1'
b101 +
#481280000000
0!
0'
#481290000000
1!
0$
b110 %
1'
0*
b110 +
#481300000000
0!
0'
#481310000000
1!
b111 %
1'
b111 +
#481320000000
0!
0'
#481330000000
1!
b1000 %
1'
b1000 +
#481340000000
0!
0'
#481350000000
1!
b1001 %
1'
b1001 +
#481360000000
0!
0'
#481370000000
1!
b0 %
1'
b0 +
#481380000000
1"
1(
#481390000000
0!
0"
b100 &
0'
0(
b100 ,
#481400000000
1!
1$
b1 %
1'
1*
b1 +
#481410000000
0!
0'
#481420000000
1!
b10 %
1'
b10 +
#481430000000
0!
0'
#481440000000
1!
b11 %
1'
b11 +
#481450000000
0!
0'
#481460000000
1!
b100 %
1'
b100 +
#481470000000
0!
0'
#481480000000
1!
b101 %
1'
b101 +
#481490000000
0!
0'
#481500000000
1!
b110 %
1'
b110 +
#481510000000
0!
0'
#481520000000
1!
b111 %
1'
b111 +
#481530000000
0!
0'
#481540000000
1!
0$
b1000 %
1'
0*
b1000 +
#481550000000
0!
0'
#481560000000
1!
b1001 %
1'
b1001 +
#481570000000
0!
0'
#481580000000
1!
b0 %
1'
b0 +
#481590000000
0!
0'
#481600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#481610000000
0!
0'
#481620000000
1!
b10 %
1'
b10 +
#481630000000
0!
0'
#481640000000
1!
b11 %
1'
b11 +
#481650000000
0!
0'
#481660000000
1!
b100 %
1'
b100 +
#481670000000
0!
0'
#481680000000
1!
b101 %
1'
b101 +
#481690000000
0!
0'
#481700000000
1!
0$
b110 %
1'
0*
b110 +
#481710000000
0!
0'
#481720000000
1!
b111 %
1'
b111 +
#481730000000
0!
0'
#481740000000
1!
b1000 %
1'
b1000 +
#481750000000
0!
0'
#481760000000
1!
b1001 %
1'
b1001 +
#481770000000
0!
0'
#481780000000
1!
b0 %
1'
b0 +
#481790000000
0!
0'
#481800000000
1!
1$
b1 %
1'
1*
b1 +
#481810000000
1"
1(
#481820000000
0!
0"
b100 &
0'
0(
b100 ,
#481830000000
1!
b10 %
1'
b10 +
#481840000000
0!
0'
#481850000000
1!
b11 %
1'
b11 +
#481860000000
0!
0'
#481870000000
1!
b100 %
1'
b100 +
#481880000000
0!
0'
#481890000000
1!
b101 %
1'
b101 +
#481900000000
0!
0'
#481910000000
1!
b110 %
1'
b110 +
#481920000000
0!
0'
#481930000000
1!
b111 %
1'
b111 +
#481940000000
0!
0'
#481950000000
1!
0$
b1000 %
1'
0*
b1000 +
#481960000000
0!
0'
#481970000000
1!
b1001 %
1'
b1001 +
#481980000000
0!
0'
#481990000000
1!
b0 %
1'
b0 +
#482000000000
0!
0'
#482010000000
1!
1$
b1 %
1'
1*
b1 +
#482020000000
0!
0'
#482030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#482040000000
0!
0'
#482050000000
1!
b11 %
1'
b11 +
#482060000000
0!
0'
#482070000000
1!
b100 %
1'
b100 +
#482080000000
0!
0'
#482090000000
1!
b101 %
1'
b101 +
#482100000000
0!
0'
#482110000000
1!
0$
b110 %
1'
0*
b110 +
#482120000000
0!
0'
#482130000000
1!
b111 %
1'
b111 +
#482140000000
0!
0'
#482150000000
1!
b1000 %
1'
b1000 +
#482160000000
0!
0'
#482170000000
1!
b1001 %
1'
b1001 +
#482180000000
0!
0'
#482190000000
1!
b0 %
1'
b0 +
#482200000000
0!
0'
#482210000000
1!
1$
b1 %
1'
1*
b1 +
#482220000000
0!
0'
#482230000000
1!
b10 %
1'
b10 +
#482240000000
1"
1(
#482250000000
0!
0"
b100 &
0'
0(
b100 ,
#482260000000
1!
b11 %
1'
b11 +
#482270000000
0!
0'
#482280000000
1!
b100 %
1'
b100 +
#482290000000
0!
0'
#482300000000
1!
b101 %
1'
b101 +
#482310000000
0!
0'
#482320000000
1!
b110 %
1'
b110 +
#482330000000
0!
0'
#482340000000
1!
b111 %
1'
b111 +
#482350000000
0!
0'
#482360000000
1!
0$
b1000 %
1'
0*
b1000 +
#482370000000
0!
0'
#482380000000
1!
b1001 %
1'
b1001 +
#482390000000
0!
0'
#482400000000
1!
b0 %
1'
b0 +
#482410000000
0!
0'
#482420000000
1!
1$
b1 %
1'
1*
b1 +
#482430000000
0!
0'
#482440000000
1!
b10 %
1'
b10 +
#482450000000
0!
0'
#482460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#482470000000
0!
0'
#482480000000
1!
b100 %
1'
b100 +
#482490000000
0!
0'
#482500000000
1!
b101 %
1'
b101 +
#482510000000
0!
0'
#482520000000
1!
0$
b110 %
1'
0*
b110 +
#482530000000
0!
0'
#482540000000
1!
b111 %
1'
b111 +
#482550000000
0!
0'
#482560000000
1!
b1000 %
1'
b1000 +
#482570000000
0!
0'
#482580000000
1!
b1001 %
1'
b1001 +
#482590000000
0!
0'
#482600000000
1!
b0 %
1'
b0 +
#482610000000
0!
0'
#482620000000
1!
1$
b1 %
1'
1*
b1 +
#482630000000
0!
0'
#482640000000
1!
b10 %
1'
b10 +
#482650000000
0!
0'
#482660000000
1!
b11 %
1'
b11 +
#482670000000
1"
1(
#482680000000
0!
0"
b100 &
0'
0(
b100 ,
#482690000000
1!
b100 %
1'
b100 +
#482700000000
0!
0'
#482710000000
1!
b101 %
1'
b101 +
#482720000000
0!
0'
#482730000000
1!
b110 %
1'
b110 +
#482740000000
0!
0'
#482750000000
1!
b111 %
1'
b111 +
#482760000000
0!
0'
#482770000000
1!
0$
b1000 %
1'
0*
b1000 +
#482780000000
0!
0'
#482790000000
1!
b1001 %
1'
b1001 +
#482800000000
0!
0'
#482810000000
1!
b0 %
1'
b0 +
#482820000000
0!
0'
#482830000000
1!
1$
b1 %
1'
1*
b1 +
#482840000000
0!
0'
#482850000000
1!
b10 %
1'
b10 +
#482860000000
0!
0'
#482870000000
1!
b11 %
1'
b11 +
#482880000000
0!
0'
#482890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#482900000000
0!
0'
#482910000000
1!
b101 %
1'
b101 +
#482920000000
0!
0'
#482930000000
1!
0$
b110 %
1'
0*
b110 +
#482940000000
0!
0'
#482950000000
1!
b111 %
1'
b111 +
#482960000000
0!
0'
#482970000000
1!
b1000 %
1'
b1000 +
#482980000000
0!
0'
#482990000000
1!
b1001 %
1'
b1001 +
#483000000000
0!
0'
#483010000000
1!
b0 %
1'
b0 +
#483020000000
0!
0'
#483030000000
1!
1$
b1 %
1'
1*
b1 +
#483040000000
0!
0'
#483050000000
1!
b10 %
1'
b10 +
#483060000000
0!
0'
#483070000000
1!
b11 %
1'
b11 +
#483080000000
0!
0'
#483090000000
1!
b100 %
1'
b100 +
#483100000000
1"
1(
#483110000000
0!
0"
b100 &
0'
0(
b100 ,
#483120000000
1!
b101 %
1'
b101 +
#483130000000
0!
0'
#483140000000
1!
b110 %
1'
b110 +
#483150000000
0!
0'
#483160000000
1!
b111 %
1'
b111 +
#483170000000
0!
0'
#483180000000
1!
0$
b1000 %
1'
0*
b1000 +
#483190000000
0!
0'
#483200000000
1!
b1001 %
1'
b1001 +
#483210000000
0!
0'
#483220000000
1!
b0 %
1'
b0 +
#483230000000
0!
0'
#483240000000
1!
1$
b1 %
1'
1*
b1 +
#483250000000
0!
0'
#483260000000
1!
b10 %
1'
b10 +
#483270000000
0!
0'
#483280000000
1!
b11 %
1'
b11 +
#483290000000
0!
0'
#483300000000
1!
b100 %
1'
b100 +
#483310000000
0!
0'
#483320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#483330000000
0!
0'
#483340000000
1!
0$
b110 %
1'
0*
b110 +
#483350000000
0!
0'
#483360000000
1!
b111 %
1'
b111 +
#483370000000
0!
0'
#483380000000
1!
b1000 %
1'
b1000 +
#483390000000
0!
0'
#483400000000
1!
b1001 %
1'
b1001 +
#483410000000
0!
0'
#483420000000
1!
b0 %
1'
b0 +
#483430000000
0!
0'
#483440000000
1!
1$
b1 %
1'
1*
b1 +
#483450000000
0!
0'
#483460000000
1!
b10 %
1'
b10 +
#483470000000
0!
0'
#483480000000
1!
b11 %
1'
b11 +
#483490000000
0!
0'
#483500000000
1!
b100 %
1'
b100 +
#483510000000
0!
0'
#483520000000
1!
b101 %
1'
b101 +
#483530000000
1"
1(
#483540000000
0!
0"
b100 &
0'
0(
b100 ,
#483550000000
1!
b110 %
1'
b110 +
#483560000000
0!
0'
#483570000000
1!
b111 %
1'
b111 +
#483580000000
0!
0'
#483590000000
1!
0$
b1000 %
1'
0*
b1000 +
#483600000000
0!
0'
#483610000000
1!
b1001 %
1'
b1001 +
#483620000000
0!
0'
#483630000000
1!
b0 %
1'
b0 +
#483640000000
0!
0'
#483650000000
1!
1$
b1 %
1'
1*
b1 +
#483660000000
0!
0'
#483670000000
1!
b10 %
1'
b10 +
#483680000000
0!
0'
#483690000000
1!
b11 %
1'
b11 +
#483700000000
0!
0'
#483710000000
1!
b100 %
1'
b100 +
#483720000000
0!
0'
#483730000000
1!
b101 %
1'
b101 +
#483740000000
0!
0'
#483750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#483760000000
0!
0'
#483770000000
1!
b111 %
1'
b111 +
#483780000000
0!
0'
#483790000000
1!
b1000 %
1'
b1000 +
#483800000000
0!
0'
#483810000000
1!
b1001 %
1'
b1001 +
#483820000000
0!
0'
#483830000000
1!
b0 %
1'
b0 +
#483840000000
0!
0'
#483850000000
1!
1$
b1 %
1'
1*
b1 +
#483860000000
0!
0'
#483870000000
1!
b10 %
1'
b10 +
#483880000000
0!
0'
#483890000000
1!
b11 %
1'
b11 +
#483900000000
0!
0'
#483910000000
1!
b100 %
1'
b100 +
#483920000000
0!
0'
#483930000000
1!
b101 %
1'
b101 +
#483940000000
0!
0'
#483950000000
1!
0$
b110 %
1'
0*
b110 +
#483960000000
1"
1(
#483970000000
0!
0"
b100 &
0'
0(
b100 ,
#483980000000
1!
1$
b111 %
1'
1*
b111 +
#483990000000
0!
0'
#484000000000
1!
0$
b1000 %
1'
0*
b1000 +
#484010000000
0!
0'
#484020000000
1!
b1001 %
1'
b1001 +
#484030000000
0!
0'
#484040000000
1!
b0 %
1'
b0 +
#484050000000
0!
0'
#484060000000
1!
1$
b1 %
1'
1*
b1 +
#484070000000
0!
0'
#484080000000
1!
b10 %
1'
b10 +
#484090000000
0!
0'
#484100000000
1!
b11 %
1'
b11 +
#484110000000
0!
0'
#484120000000
1!
b100 %
1'
b100 +
#484130000000
0!
0'
#484140000000
1!
b101 %
1'
b101 +
#484150000000
0!
0'
#484160000000
1!
b110 %
1'
b110 +
#484170000000
0!
0'
#484180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#484190000000
0!
0'
#484200000000
1!
b1000 %
1'
b1000 +
#484210000000
0!
0'
#484220000000
1!
b1001 %
1'
b1001 +
#484230000000
0!
0'
#484240000000
1!
b0 %
1'
b0 +
#484250000000
0!
0'
#484260000000
1!
1$
b1 %
1'
1*
b1 +
#484270000000
0!
0'
#484280000000
1!
b10 %
1'
b10 +
#484290000000
0!
0'
#484300000000
1!
b11 %
1'
b11 +
#484310000000
0!
0'
#484320000000
1!
b100 %
1'
b100 +
#484330000000
0!
0'
#484340000000
1!
b101 %
1'
b101 +
#484350000000
0!
0'
#484360000000
1!
0$
b110 %
1'
0*
b110 +
#484370000000
0!
0'
#484380000000
1!
b111 %
1'
b111 +
#484390000000
1"
1(
#484400000000
0!
0"
b100 &
0'
0(
b100 ,
#484410000000
1!
b1000 %
1'
b1000 +
#484420000000
0!
0'
#484430000000
1!
b1001 %
1'
b1001 +
#484440000000
0!
0'
#484450000000
1!
b0 %
1'
b0 +
#484460000000
0!
0'
#484470000000
1!
1$
b1 %
1'
1*
b1 +
#484480000000
0!
0'
#484490000000
1!
b10 %
1'
b10 +
#484500000000
0!
0'
#484510000000
1!
b11 %
1'
b11 +
#484520000000
0!
0'
#484530000000
1!
b100 %
1'
b100 +
#484540000000
0!
0'
#484550000000
1!
b101 %
1'
b101 +
#484560000000
0!
0'
#484570000000
1!
b110 %
1'
b110 +
#484580000000
0!
0'
#484590000000
1!
b111 %
1'
b111 +
#484600000000
0!
0'
#484610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#484620000000
0!
0'
#484630000000
1!
b1001 %
1'
b1001 +
#484640000000
0!
0'
#484650000000
1!
b0 %
1'
b0 +
#484660000000
0!
0'
#484670000000
1!
1$
b1 %
1'
1*
b1 +
#484680000000
0!
0'
#484690000000
1!
b10 %
1'
b10 +
#484700000000
0!
0'
#484710000000
1!
b11 %
1'
b11 +
#484720000000
0!
0'
#484730000000
1!
b100 %
1'
b100 +
#484740000000
0!
0'
#484750000000
1!
b101 %
1'
b101 +
#484760000000
0!
0'
#484770000000
1!
0$
b110 %
1'
0*
b110 +
#484780000000
0!
0'
#484790000000
1!
b111 %
1'
b111 +
#484800000000
0!
0'
#484810000000
1!
b1000 %
1'
b1000 +
#484820000000
1"
1(
#484830000000
0!
0"
b100 &
0'
0(
b100 ,
#484840000000
1!
b1001 %
1'
b1001 +
#484850000000
0!
0'
#484860000000
1!
b0 %
1'
b0 +
#484870000000
0!
0'
#484880000000
1!
1$
b1 %
1'
1*
b1 +
#484890000000
0!
0'
#484900000000
1!
b10 %
1'
b10 +
#484910000000
0!
0'
#484920000000
1!
b11 %
1'
b11 +
#484930000000
0!
0'
#484940000000
1!
b100 %
1'
b100 +
#484950000000
0!
0'
#484960000000
1!
b101 %
1'
b101 +
#484970000000
0!
0'
#484980000000
1!
b110 %
1'
b110 +
#484990000000
0!
0'
#485000000000
1!
b111 %
1'
b111 +
#485010000000
0!
0'
#485020000000
1!
0$
b1000 %
1'
0*
b1000 +
#485030000000
0!
0'
#485040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#485050000000
0!
0'
#485060000000
1!
b0 %
1'
b0 +
#485070000000
0!
0'
#485080000000
1!
1$
b1 %
1'
1*
b1 +
#485090000000
0!
0'
#485100000000
1!
b10 %
1'
b10 +
#485110000000
0!
0'
#485120000000
1!
b11 %
1'
b11 +
#485130000000
0!
0'
#485140000000
1!
b100 %
1'
b100 +
#485150000000
0!
0'
#485160000000
1!
b101 %
1'
b101 +
#485170000000
0!
0'
#485180000000
1!
0$
b110 %
1'
0*
b110 +
#485190000000
0!
0'
#485200000000
1!
b111 %
1'
b111 +
#485210000000
0!
0'
#485220000000
1!
b1000 %
1'
b1000 +
#485230000000
0!
0'
#485240000000
1!
b1001 %
1'
b1001 +
#485250000000
1"
1(
#485260000000
0!
0"
b100 &
0'
0(
b100 ,
#485270000000
1!
b0 %
1'
b0 +
#485280000000
0!
0'
#485290000000
1!
1$
b1 %
1'
1*
b1 +
#485300000000
0!
0'
#485310000000
1!
b10 %
1'
b10 +
#485320000000
0!
0'
#485330000000
1!
b11 %
1'
b11 +
#485340000000
0!
0'
#485350000000
1!
b100 %
1'
b100 +
#485360000000
0!
0'
#485370000000
1!
b101 %
1'
b101 +
#485380000000
0!
0'
#485390000000
1!
b110 %
1'
b110 +
#485400000000
0!
0'
#485410000000
1!
b111 %
1'
b111 +
#485420000000
0!
0'
#485430000000
1!
0$
b1000 %
1'
0*
b1000 +
#485440000000
0!
0'
#485450000000
1!
b1001 %
1'
b1001 +
#485460000000
0!
0'
#485470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#485480000000
0!
0'
#485490000000
1!
1$
b1 %
1'
1*
b1 +
#485500000000
0!
0'
#485510000000
1!
b10 %
1'
b10 +
#485520000000
0!
0'
#485530000000
1!
b11 %
1'
b11 +
#485540000000
0!
0'
#485550000000
1!
b100 %
1'
b100 +
#485560000000
0!
0'
#485570000000
1!
b101 %
1'
b101 +
#485580000000
0!
0'
#485590000000
1!
0$
b110 %
1'
0*
b110 +
#485600000000
0!
0'
#485610000000
1!
b111 %
1'
b111 +
#485620000000
0!
0'
#485630000000
1!
b1000 %
1'
b1000 +
#485640000000
0!
0'
#485650000000
1!
b1001 %
1'
b1001 +
#485660000000
0!
0'
#485670000000
1!
b0 %
1'
b0 +
#485680000000
1"
1(
#485690000000
0!
0"
b100 &
0'
0(
b100 ,
#485700000000
1!
1$
b1 %
1'
1*
b1 +
#485710000000
0!
0'
#485720000000
1!
b10 %
1'
b10 +
#485730000000
0!
0'
#485740000000
1!
b11 %
1'
b11 +
#485750000000
0!
0'
#485760000000
1!
b100 %
1'
b100 +
#485770000000
0!
0'
#485780000000
1!
b101 %
1'
b101 +
#485790000000
0!
0'
#485800000000
1!
b110 %
1'
b110 +
#485810000000
0!
0'
#485820000000
1!
b111 %
1'
b111 +
#485830000000
0!
0'
#485840000000
1!
0$
b1000 %
1'
0*
b1000 +
#485850000000
0!
0'
#485860000000
1!
b1001 %
1'
b1001 +
#485870000000
0!
0'
#485880000000
1!
b0 %
1'
b0 +
#485890000000
0!
0'
#485900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#485910000000
0!
0'
#485920000000
1!
b10 %
1'
b10 +
#485930000000
0!
0'
#485940000000
1!
b11 %
1'
b11 +
#485950000000
0!
0'
#485960000000
1!
b100 %
1'
b100 +
#485970000000
0!
0'
#485980000000
1!
b101 %
1'
b101 +
#485990000000
0!
0'
#486000000000
1!
0$
b110 %
1'
0*
b110 +
#486010000000
0!
0'
#486020000000
1!
b111 %
1'
b111 +
#486030000000
0!
0'
#486040000000
1!
b1000 %
1'
b1000 +
#486050000000
0!
0'
#486060000000
1!
b1001 %
1'
b1001 +
#486070000000
0!
0'
#486080000000
1!
b0 %
1'
b0 +
#486090000000
0!
0'
#486100000000
1!
1$
b1 %
1'
1*
b1 +
#486110000000
1"
1(
#486120000000
0!
0"
b100 &
0'
0(
b100 ,
#486130000000
1!
b10 %
1'
b10 +
#486140000000
0!
0'
#486150000000
1!
b11 %
1'
b11 +
#486160000000
0!
0'
#486170000000
1!
b100 %
1'
b100 +
#486180000000
0!
0'
#486190000000
1!
b101 %
1'
b101 +
#486200000000
0!
0'
#486210000000
1!
b110 %
1'
b110 +
#486220000000
0!
0'
#486230000000
1!
b111 %
1'
b111 +
#486240000000
0!
0'
#486250000000
1!
0$
b1000 %
1'
0*
b1000 +
#486260000000
0!
0'
#486270000000
1!
b1001 %
1'
b1001 +
#486280000000
0!
0'
#486290000000
1!
b0 %
1'
b0 +
#486300000000
0!
0'
#486310000000
1!
1$
b1 %
1'
1*
b1 +
#486320000000
0!
0'
#486330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#486340000000
0!
0'
#486350000000
1!
b11 %
1'
b11 +
#486360000000
0!
0'
#486370000000
1!
b100 %
1'
b100 +
#486380000000
0!
0'
#486390000000
1!
b101 %
1'
b101 +
#486400000000
0!
0'
#486410000000
1!
0$
b110 %
1'
0*
b110 +
#486420000000
0!
0'
#486430000000
1!
b111 %
1'
b111 +
#486440000000
0!
0'
#486450000000
1!
b1000 %
1'
b1000 +
#486460000000
0!
0'
#486470000000
1!
b1001 %
1'
b1001 +
#486480000000
0!
0'
#486490000000
1!
b0 %
1'
b0 +
#486500000000
0!
0'
#486510000000
1!
1$
b1 %
1'
1*
b1 +
#486520000000
0!
0'
#486530000000
1!
b10 %
1'
b10 +
#486540000000
1"
1(
#486550000000
0!
0"
b100 &
0'
0(
b100 ,
#486560000000
1!
b11 %
1'
b11 +
#486570000000
0!
0'
#486580000000
1!
b100 %
1'
b100 +
#486590000000
0!
0'
#486600000000
1!
b101 %
1'
b101 +
#486610000000
0!
0'
#486620000000
1!
b110 %
1'
b110 +
#486630000000
0!
0'
#486640000000
1!
b111 %
1'
b111 +
#486650000000
0!
0'
#486660000000
1!
0$
b1000 %
1'
0*
b1000 +
#486670000000
0!
0'
#486680000000
1!
b1001 %
1'
b1001 +
#486690000000
0!
0'
#486700000000
1!
b0 %
1'
b0 +
#486710000000
0!
0'
#486720000000
1!
1$
b1 %
1'
1*
b1 +
#486730000000
0!
0'
#486740000000
1!
b10 %
1'
b10 +
#486750000000
0!
0'
#486760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#486770000000
0!
0'
#486780000000
1!
b100 %
1'
b100 +
#486790000000
0!
0'
#486800000000
1!
b101 %
1'
b101 +
#486810000000
0!
0'
#486820000000
1!
0$
b110 %
1'
0*
b110 +
#486830000000
0!
0'
#486840000000
1!
b111 %
1'
b111 +
#486850000000
0!
0'
#486860000000
1!
b1000 %
1'
b1000 +
#486870000000
0!
0'
#486880000000
1!
b1001 %
1'
b1001 +
#486890000000
0!
0'
#486900000000
1!
b0 %
1'
b0 +
#486910000000
0!
0'
#486920000000
1!
1$
b1 %
1'
1*
b1 +
#486930000000
0!
0'
#486940000000
1!
b10 %
1'
b10 +
#486950000000
0!
0'
#486960000000
1!
b11 %
1'
b11 +
#486970000000
1"
1(
#486980000000
0!
0"
b100 &
0'
0(
b100 ,
#486990000000
1!
b100 %
1'
b100 +
#487000000000
0!
0'
#487010000000
1!
b101 %
1'
b101 +
#487020000000
0!
0'
#487030000000
1!
b110 %
1'
b110 +
#487040000000
0!
0'
#487050000000
1!
b111 %
1'
b111 +
#487060000000
0!
0'
#487070000000
1!
0$
b1000 %
1'
0*
b1000 +
#487080000000
0!
0'
#487090000000
1!
b1001 %
1'
b1001 +
#487100000000
0!
0'
#487110000000
1!
b0 %
1'
b0 +
#487120000000
0!
0'
#487130000000
1!
1$
b1 %
1'
1*
b1 +
#487140000000
0!
0'
#487150000000
1!
b10 %
1'
b10 +
#487160000000
0!
0'
#487170000000
1!
b11 %
1'
b11 +
#487180000000
0!
0'
#487190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#487200000000
0!
0'
#487210000000
1!
b101 %
1'
b101 +
#487220000000
0!
0'
#487230000000
1!
0$
b110 %
1'
0*
b110 +
#487240000000
0!
0'
#487250000000
1!
b111 %
1'
b111 +
#487260000000
0!
0'
#487270000000
1!
b1000 %
1'
b1000 +
#487280000000
0!
0'
#487290000000
1!
b1001 %
1'
b1001 +
#487300000000
0!
0'
#487310000000
1!
b0 %
1'
b0 +
#487320000000
0!
0'
#487330000000
1!
1$
b1 %
1'
1*
b1 +
#487340000000
0!
0'
#487350000000
1!
b10 %
1'
b10 +
#487360000000
0!
0'
#487370000000
1!
b11 %
1'
b11 +
#487380000000
0!
0'
#487390000000
1!
b100 %
1'
b100 +
#487400000000
1"
1(
#487410000000
0!
0"
b100 &
0'
0(
b100 ,
#487420000000
1!
b101 %
1'
b101 +
#487430000000
0!
0'
#487440000000
1!
b110 %
1'
b110 +
#487450000000
0!
0'
#487460000000
1!
b111 %
1'
b111 +
#487470000000
0!
0'
#487480000000
1!
0$
b1000 %
1'
0*
b1000 +
#487490000000
0!
0'
#487500000000
1!
b1001 %
1'
b1001 +
#487510000000
0!
0'
#487520000000
1!
b0 %
1'
b0 +
#487530000000
0!
0'
#487540000000
1!
1$
b1 %
1'
1*
b1 +
#487550000000
0!
0'
#487560000000
1!
b10 %
1'
b10 +
#487570000000
0!
0'
#487580000000
1!
b11 %
1'
b11 +
#487590000000
0!
0'
#487600000000
1!
b100 %
1'
b100 +
#487610000000
0!
0'
#487620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#487630000000
0!
0'
#487640000000
1!
0$
b110 %
1'
0*
b110 +
#487650000000
0!
0'
#487660000000
1!
b111 %
1'
b111 +
#487670000000
0!
0'
#487680000000
1!
b1000 %
1'
b1000 +
#487690000000
0!
0'
#487700000000
1!
b1001 %
1'
b1001 +
#487710000000
0!
0'
#487720000000
1!
b0 %
1'
b0 +
#487730000000
0!
0'
#487740000000
1!
1$
b1 %
1'
1*
b1 +
#487750000000
0!
0'
#487760000000
1!
b10 %
1'
b10 +
#487770000000
0!
0'
#487780000000
1!
b11 %
1'
b11 +
#487790000000
0!
0'
#487800000000
1!
b100 %
1'
b100 +
#487810000000
0!
0'
#487820000000
1!
b101 %
1'
b101 +
#487830000000
1"
1(
#487840000000
0!
0"
b100 &
0'
0(
b100 ,
#487850000000
1!
b110 %
1'
b110 +
#487860000000
0!
0'
#487870000000
1!
b111 %
1'
b111 +
#487880000000
0!
0'
#487890000000
1!
0$
b1000 %
1'
0*
b1000 +
#487900000000
0!
0'
#487910000000
1!
b1001 %
1'
b1001 +
#487920000000
0!
0'
#487930000000
1!
b0 %
1'
b0 +
#487940000000
0!
0'
#487950000000
1!
1$
b1 %
1'
1*
b1 +
#487960000000
0!
0'
#487970000000
1!
b10 %
1'
b10 +
#487980000000
0!
0'
#487990000000
1!
b11 %
1'
b11 +
#488000000000
0!
0'
#488010000000
1!
b100 %
1'
b100 +
#488020000000
0!
0'
#488030000000
1!
b101 %
1'
b101 +
#488040000000
0!
0'
#488050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#488060000000
0!
0'
#488070000000
1!
b111 %
1'
b111 +
#488080000000
0!
0'
#488090000000
1!
b1000 %
1'
b1000 +
#488100000000
0!
0'
#488110000000
1!
b1001 %
1'
b1001 +
#488120000000
0!
0'
#488130000000
1!
b0 %
1'
b0 +
#488140000000
0!
0'
#488150000000
1!
1$
b1 %
1'
1*
b1 +
#488160000000
0!
0'
#488170000000
1!
b10 %
1'
b10 +
#488180000000
0!
0'
#488190000000
1!
b11 %
1'
b11 +
#488200000000
0!
0'
#488210000000
1!
b100 %
1'
b100 +
#488220000000
0!
0'
#488230000000
1!
b101 %
1'
b101 +
#488240000000
0!
0'
#488250000000
1!
0$
b110 %
1'
0*
b110 +
#488260000000
1"
1(
#488270000000
0!
0"
b100 &
0'
0(
b100 ,
#488280000000
1!
1$
b111 %
1'
1*
b111 +
#488290000000
0!
0'
#488300000000
1!
0$
b1000 %
1'
0*
b1000 +
#488310000000
0!
0'
#488320000000
1!
b1001 %
1'
b1001 +
#488330000000
0!
0'
#488340000000
1!
b0 %
1'
b0 +
#488350000000
0!
0'
#488360000000
1!
1$
b1 %
1'
1*
b1 +
#488370000000
0!
0'
#488380000000
1!
b10 %
1'
b10 +
#488390000000
0!
0'
#488400000000
1!
b11 %
1'
b11 +
#488410000000
0!
0'
#488420000000
1!
b100 %
1'
b100 +
#488430000000
0!
0'
#488440000000
1!
b101 %
1'
b101 +
#488450000000
0!
0'
#488460000000
1!
b110 %
1'
b110 +
#488470000000
0!
0'
#488480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#488490000000
0!
0'
#488500000000
1!
b1000 %
1'
b1000 +
#488510000000
0!
0'
#488520000000
1!
b1001 %
1'
b1001 +
#488530000000
0!
0'
#488540000000
1!
b0 %
1'
b0 +
#488550000000
0!
0'
#488560000000
1!
1$
b1 %
1'
1*
b1 +
#488570000000
0!
0'
#488580000000
1!
b10 %
1'
b10 +
#488590000000
0!
0'
#488600000000
1!
b11 %
1'
b11 +
#488610000000
0!
0'
#488620000000
1!
b100 %
1'
b100 +
#488630000000
0!
0'
#488640000000
1!
b101 %
1'
b101 +
#488650000000
0!
0'
#488660000000
1!
0$
b110 %
1'
0*
b110 +
#488670000000
0!
0'
#488680000000
1!
b111 %
1'
b111 +
#488690000000
1"
1(
#488700000000
0!
0"
b100 &
0'
0(
b100 ,
#488710000000
1!
b1000 %
1'
b1000 +
#488720000000
0!
0'
#488730000000
1!
b1001 %
1'
b1001 +
#488740000000
0!
0'
#488750000000
1!
b0 %
1'
b0 +
#488760000000
0!
0'
#488770000000
1!
1$
b1 %
1'
1*
b1 +
#488780000000
0!
0'
#488790000000
1!
b10 %
1'
b10 +
#488800000000
0!
0'
#488810000000
1!
b11 %
1'
b11 +
#488820000000
0!
0'
#488830000000
1!
b100 %
1'
b100 +
#488840000000
0!
0'
#488850000000
1!
b101 %
1'
b101 +
#488860000000
0!
0'
#488870000000
1!
b110 %
1'
b110 +
#488880000000
0!
0'
#488890000000
1!
b111 %
1'
b111 +
#488900000000
0!
0'
#488910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#488920000000
0!
0'
#488930000000
1!
b1001 %
1'
b1001 +
#488940000000
0!
0'
#488950000000
1!
b0 %
1'
b0 +
#488960000000
0!
0'
#488970000000
1!
1$
b1 %
1'
1*
b1 +
#488980000000
0!
0'
#488990000000
1!
b10 %
1'
b10 +
#489000000000
0!
0'
#489010000000
1!
b11 %
1'
b11 +
#489020000000
0!
0'
#489030000000
1!
b100 %
1'
b100 +
#489040000000
0!
0'
#489050000000
1!
b101 %
1'
b101 +
#489060000000
0!
0'
#489070000000
1!
0$
b110 %
1'
0*
b110 +
#489080000000
0!
0'
#489090000000
1!
b111 %
1'
b111 +
#489100000000
0!
0'
#489110000000
1!
b1000 %
1'
b1000 +
#489120000000
1"
1(
#489130000000
0!
0"
b100 &
0'
0(
b100 ,
#489140000000
1!
b1001 %
1'
b1001 +
#489150000000
0!
0'
#489160000000
1!
b0 %
1'
b0 +
#489170000000
0!
0'
#489180000000
1!
1$
b1 %
1'
1*
b1 +
#489190000000
0!
0'
#489200000000
1!
b10 %
1'
b10 +
#489210000000
0!
0'
#489220000000
1!
b11 %
1'
b11 +
#489230000000
0!
0'
#489240000000
1!
b100 %
1'
b100 +
#489250000000
0!
0'
#489260000000
1!
b101 %
1'
b101 +
#489270000000
0!
0'
#489280000000
1!
b110 %
1'
b110 +
#489290000000
0!
0'
#489300000000
1!
b111 %
1'
b111 +
#489310000000
0!
0'
#489320000000
1!
0$
b1000 %
1'
0*
b1000 +
#489330000000
0!
0'
#489340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#489350000000
0!
0'
#489360000000
1!
b0 %
1'
b0 +
#489370000000
0!
0'
#489380000000
1!
1$
b1 %
1'
1*
b1 +
#489390000000
0!
0'
#489400000000
1!
b10 %
1'
b10 +
#489410000000
0!
0'
#489420000000
1!
b11 %
1'
b11 +
#489430000000
0!
0'
#489440000000
1!
b100 %
1'
b100 +
#489450000000
0!
0'
#489460000000
1!
b101 %
1'
b101 +
#489470000000
0!
0'
#489480000000
1!
0$
b110 %
1'
0*
b110 +
#489490000000
0!
0'
#489500000000
1!
b111 %
1'
b111 +
#489510000000
0!
0'
#489520000000
1!
b1000 %
1'
b1000 +
#489530000000
0!
0'
#489540000000
1!
b1001 %
1'
b1001 +
#489550000000
1"
1(
#489560000000
0!
0"
b100 &
0'
0(
b100 ,
#489570000000
1!
b0 %
1'
b0 +
#489580000000
0!
0'
#489590000000
1!
1$
b1 %
1'
1*
b1 +
#489600000000
0!
0'
#489610000000
1!
b10 %
1'
b10 +
#489620000000
0!
0'
#489630000000
1!
b11 %
1'
b11 +
#489640000000
0!
0'
#489650000000
1!
b100 %
1'
b100 +
#489660000000
0!
0'
#489670000000
1!
b101 %
1'
b101 +
#489680000000
0!
0'
#489690000000
1!
b110 %
1'
b110 +
#489700000000
0!
0'
#489710000000
1!
b111 %
1'
b111 +
#489720000000
0!
0'
#489730000000
1!
0$
b1000 %
1'
0*
b1000 +
#489740000000
0!
0'
#489750000000
1!
b1001 %
1'
b1001 +
#489760000000
0!
0'
#489770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#489780000000
0!
0'
#489790000000
1!
1$
b1 %
1'
1*
b1 +
#489800000000
0!
0'
#489810000000
1!
b10 %
1'
b10 +
#489820000000
0!
0'
#489830000000
1!
b11 %
1'
b11 +
#489840000000
0!
0'
#489850000000
1!
b100 %
1'
b100 +
#489860000000
0!
0'
#489870000000
1!
b101 %
1'
b101 +
#489880000000
0!
0'
#489890000000
1!
0$
b110 %
1'
0*
b110 +
#489900000000
0!
0'
#489910000000
1!
b111 %
1'
b111 +
#489920000000
0!
0'
#489930000000
1!
b1000 %
1'
b1000 +
#489940000000
0!
0'
#489950000000
1!
b1001 %
1'
b1001 +
#489960000000
0!
0'
#489970000000
1!
b0 %
1'
b0 +
#489980000000
1"
1(
#489990000000
0!
0"
b100 &
0'
0(
b100 ,
#490000000000
1!
1$
b1 %
1'
1*
b1 +
#490010000000
0!
0'
#490020000000
1!
b10 %
1'
b10 +
#490030000000
0!
0'
#490040000000
1!
b11 %
1'
b11 +
#490050000000
0!
0'
#490060000000
1!
b100 %
1'
b100 +
#490070000000
0!
0'
#490080000000
1!
b101 %
1'
b101 +
#490090000000
0!
0'
#490100000000
1!
b110 %
1'
b110 +
#490110000000
0!
0'
#490120000000
1!
b111 %
1'
b111 +
#490130000000
0!
0'
#490140000000
1!
0$
b1000 %
1'
0*
b1000 +
#490150000000
0!
0'
#490160000000
1!
b1001 %
1'
b1001 +
#490170000000
0!
0'
#490180000000
1!
b0 %
1'
b0 +
#490190000000
0!
0'
#490200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#490210000000
0!
0'
#490220000000
1!
b10 %
1'
b10 +
#490230000000
0!
0'
#490240000000
1!
b11 %
1'
b11 +
#490250000000
0!
0'
#490260000000
1!
b100 %
1'
b100 +
#490270000000
0!
0'
#490280000000
1!
b101 %
1'
b101 +
#490290000000
0!
0'
#490300000000
1!
0$
b110 %
1'
0*
b110 +
#490310000000
0!
0'
#490320000000
1!
b111 %
1'
b111 +
#490330000000
0!
0'
#490340000000
1!
b1000 %
1'
b1000 +
#490350000000
0!
0'
#490360000000
1!
b1001 %
1'
b1001 +
#490370000000
0!
0'
#490380000000
1!
b0 %
1'
b0 +
#490390000000
0!
0'
#490400000000
1!
1$
b1 %
1'
1*
b1 +
#490410000000
1"
1(
#490420000000
0!
0"
b100 &
0'
0(
b100 ,
#490430000000
1!
b10 %
1'
b10 +
#490440000000
0!
0'
#490450000000
1!
b11 %
1'
b11 +
#490460000000
0!
0'
#490470000000
1!
b100 %
1'
b100 +
#490480000000
0!
0'
#490490000000
1!
b101 %
1'
b101 +
#490500000000
0!
0'
#490510000000
1!
b110 %
1'
b110 +
#490520000000
0!
0'
#490530000000
1!
b111 %
1'
b111 +
#490540000000
0!
0'
#490550000000
1!
0$
b1000 %
1'
0*
b1000 +
#490560000000
0!
0'
#490570000000
1!
b1001 %
1'
b1001 +
#490580000000
0!
0'
#490590000000
1!
b0 %
1'
b0 +
#490600000000
0!
0'
#490610000000
1!
1$
b1 %
1'
1*
b1 +
#490620000000
0!
0'
#490630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#490640000000
0!
0'
#490650000000
1!
b11 %
1'
b11 +
#490660000000
0!
0'
#490670000000
1!
b100 %
1'
b100 +
#490680000000
0!
0'
#490690000000
1!
b101 %
1'
b101 +
#490700000000
0!
0'
#490710000000
1!
0$
b110 %
1'
0*
b110 +
#490720000000
0!
0'
#490730000000
1!
b111 %
1'
b111 +
#490740000000
0!
0'
#490750000000
1!
b1000 %
1'
b1000 +
#490760000000
0!
0'
#490770000000
1!
b1001 %
1'
b1001 +
#490780000000
0!
0'
#490790000000
1!
b0 %
1'
b0 +
#490800000000
0!
0'
#490810000000
1!
1$
b1 %
1'
1*
b1 +
#490820000000
0!
0'
#490830000000
1!
b10 %
1'
b10 +
#490840000000
1"
1(
#490850000000
0!
0"
b100 &
0'
0(
b100 ,
#490860000000
1!
b11 %
1'
b11 +
#490870000000
0!
0'
#490880000000
1!
b100 %
1'
b100 +
#490890000000
0!
0'
#490900000000
1!
b101 %
1'
b101 +
#490910000000
0!
0'
#490920000000
1!
b110 %
1'
b110 +
#490930000000
0!
0'
#490940000000
1!
b111 %
1'
b111 +
#490950000000
0!
0'
#490960000000
1!
0$
b1000 %
1'
0*
b1000 +
#490970000000
0!
0'
#490980000000
1!
b1001 %
1'
b1001 +
#490990000000
0!
0'
#491000000000
1!
b0 %
1'
b0 +
#491010000000
0!
0'
#491020000000
1!
1$
b1 %
1'
1*
b1 +
#491030000000
0!
0'
#491040000000
1!
b10 %
1'
b10 +
#491050000000
0!
0'
#491060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#491070000000
0!
0'
#491080000000
1!
b100 %
1'
b100 +
#491090000000
0!
0'
#491100000000
1!
b101 %
1'
b101 +
#491110000000
0!
0'
#491120000000
1!
0$
b110 %
1'
0*
b110 +
#491130000000
0!
0'
#491140000000
1!
b111 %
1'
b111 +
#491150000000
0!
0'
#491160000000
1!
b1000 %
1'
b1000 +
#491170000000
0!
0'
#491180000000
1!
b1001 %
1'
b1001 +
#491190000000
0!
0'
#491200000000
1!
b0 %
1'
b0 +
#491210000000
0!
0'
#491220000000
1!
1$
b1 %
1'
1*
b1 +
#491230000000
0!
0'
#491240000000
1!
b10 %
1'
b10 +
#491250000000
0!
0'
#491260000000
1!
b11 %
1'
b11 +
#491270000000
1"
1(
#491280000000
0!
0"
b100 &
0'
0(
b100 ,
#491290000000
1!
b100 %
1'
b100 +
#491300000000
0!
0'
#491310000000
1!
b101 %
1'
b101 +
#491320000000
0!
0'
#491330000000
1!
b110 %
1'
b110 +
#491340000000
0!
0'
#491350000000
1!
b111 %
1'
b111 +
#491360000000
0!
0'
#491370000000
1!
0$
b1000 %
1'
0*
b1000 +
#491380000000
0!
0'
#491390000000
1!
b1001 %
1'
b1001 +
#491400000000
0!
0'
#491410000000
1!
b0 %
1'
b0 +
#491420000000
0!
0'
#491430000000
1!
1$
b1 %
1'
1*
b1 +
#491440000000
0!
0'
#491450000000
1!
b10 %
1'
b10 +
#491460000000
0!
0'
#491470000000
1!
b11 %
1'
b11 +
#491480000000
0!
0'
#491490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#491500000000
0!
0'
#491510000000
1!
b101 %
1'
b101 +
#491520000000
0!
0'
#491530000000
1!
0$
b110 %
1'
0*
b110 +
#491540000000
0!
0'
#491550000000
1!
b111 %
1'
b111 +
#491560000000
0!
0'
#491570000000
1!
b1000 %
1'
b1000 +
#491580000000
0!
0'
#491590000000
1!
b1001 %
1'
b1001 +
#491600000000
0!
0'
#491610000000
1!
b0 %
1'
b0 +
#491620000000
0!
0'
#491630000000
1!
1$
b1 %
1'
1*
b1 +
#491640000000
0!
0'
#491650000000
1!
b10 %
1'
b10 +
#491660000000
0!
0'
#491670000000
1!
b11 %
1'
b11 +
#491680000000
0!
0'
#491690000000
1!
b100 %
1'
b100 +
#491700000000
1"
1(
#491710000000
0!
0"
b100 &
0'
0(
b100 ,
#491720000000
1!
b101 %
1'
b101 +
#491730000000
0!
0'
#491740000000
1!
b110 %
1'
b110 +
#491750000000
0!
0'
#491760000000
1!
b111 %
1'
b111 +
#491770000000
0!
0'
#491780000000
1!
0$
b1000 %
1'
0*
b1000 +
#491790000000
0!
0'
#491800000000
1!
b1001 %
1'
b1001 +
#491810000000
0!
0'
#491820000000
1!
b0 %
1'
b0 +
#491830000000
0!
0'
#491840000000
1!
1$
b1 %
1'
1*
b1 +
#491850000000
0!
0'
#491860000000
1!
b10 %
1'
b10 +
#491870000000
0!
0'
#491880000000
1!
b11 %
1'
b11 +
#491890000000
0!
0'
#491900000000
1!
b100 %
1'
b100 +
#491910000000
0!
0'
#491920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#491930000000
0!
0'
#491940000000
1!
0$
b110 %
1'
0*
b110 +
#491950000000
0!
0'
#491960000000
1!
b111 %
1'
b111 +
#491970000000
0!
0'
#491980000000
1!
b1000 %
1'
b1000 +
#491990000000
0!
0'
#492000000000
1!
b1001 %
1'
b1001 +
#492010000000
0!
0'
#492020000000
1!
b0 %
1'
b0 +
#492030000000
0!
0'
#492040000000
1!
1$
b1 %
1'
1*
b1 +
#492050000000
0!
0'
#492060000000
1!
b10 %
1'
b10 +
#492070000000
0!
0'
#492080000000
1!
b11 %
1'
b11 +
#492090000000
0!
0'
#492100000000
1!
b100 %
1'
b100 +
#492110000000
0!
0'
#492120000000
1!
b101 %
1'
b101 +
#492130000000
1"
1(
#492140000000
0!
0"
b100 &
0'
0(
b100 ,
#492150000000
1!
b110 %
1'
b110 +
#492160000000
0!
0'
#492170000000
1!
b111 %
1'
b111 +
#492180000000
0!
0'
#492190000000
1!
0$
b1000 %
1'
0*
b1000 +
#492200000000
0!
0'
#492210000000
1!
b1001 %
1'
b1001 +
#492220000000
0!
0'
#492230000000
1!
b0 %
1'
b0 +
#492240000000
0!
0'
#492250000000
1!
1$
b1 %
1'
1*
b1 +
#492260000000
0!
0'
#492270000000
1!
b10 %
1'
b10 +
#492280000000
0!
0'
#492290000000
1!
b11 %
1'
b11 +
#492300000000
0!
0'
#492310000000
1!
b100 %
1'
b100 +
#492320000000
0!
0'
#492330000000
1!
b101 %
1'
b101 +
#492340000000
0!
0'
#492350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#492360000000
0!
0'
#492370000000
1!
b111 %
1'
b111 +
#492380000000
0!
0'
#492390000000
1!
b1000 %
1'
b1000 +
#492400000000
0!
0'
#492410000000
1!
b1001 %
1'
b1001 +
#492420000000
0!
0'
#492430000000
1!
b0 %
1'
b0 +
#492440000000
0!
0'
#492450000000
1!
1$
b1 %
1'
1*
b1 +
#492460000000
0!
0'
#492470000000
1!
b10 %
1'
b10 +
#492480000000
0!
0'
#492490000000
1!
b11 %
1'
b11 +
#492500000000
0!
0'
#492510000000
1!
b100 %
1'
b100 +
#492520000000
0!
0'
#492530000000
1!
b101 %
1'
b101 +
#492540000000
0!
0'
#492550000000
1!
0$
b110 %
1'
0*
b110 +
#492560000000
1"
1(
#492570000000
0!
0"
b100 &
0'
0(
b100 ,
#492580000000
1!
1$
b111 %
1'
1*
b111 +
#492590000000
0!
0'
#492600000000
1!
0$
b1000 %
1'
0*
b1000 +
#492610000000
0!
0'
#492620000000
1!
b1001 %
1'
b1001 +
#492630000000
0!
0'
#492640000000
1!
b0 %
1'
b0 +
#492650000000
0!
0'
#492660000000
1!
1$
b1 %
1'
1*
b1 +
#492670000000
0!
0'
#492680000000
1!
b10 %
1'
b10 +
#492690000000
0!
0'
#492700000000
1!
b11 %
1'
b11 +
#492710000000
0!
0'
#492720000000
1!
b100 %
1'
b100 +
#492730000000
0!
0'
#492740000000
1!
b101 %
1'
b101 +
#492750000000
0!
0'
#492760000000
1!
b110 %
1'
b110 +
#492770000000
0!
0'
#492780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#492790000000
0!
0'
#492800000000
1!
b1000 %
1'
b1000 +
#492810000000
0!
0'
#492820000000
1!
b1001 %
1'
b1001 +
#492830000000
0!
0'
#492840000000
1!
b0 %
1'
b0 +
#492850000000
0!
0'
#492860000000
1!
1$
b1 %
1'
1*
b1 +
#492870000000
0!
0'
#492880000000
1!
b10 %
1'
b10 +
#492890000000
0!
0'
#492900000000
1!
b11 %
1'
b11 +
#492910000000
0!
0'
#492920000000
1!
b100 %
1'
b100 +
#492930000000
0!
0'
#492940000000
1!
b101 %
1'
b101 +
#492950000000
0!
0'
#492960000000
1!
0$
b110 %
1'
0*
b110 +
#492970000000
0!
0'
#492980000000
1!
b111 %
1'
b111 +
#492990000000
1"
1(
#493000000000
0!
0"
b100 &
0'
0(
b100 ,
#493010000000
1!
b1000 %
1'
b1000 +
#493020000000
0!
0'
#493030000000
1!
b1001 %
1'
b1001 +
#493040000000
0!
0'
#493050000000
1!
b0 %
1'
b0 +
#493060000000
0!
0'
#493070000000
1!
1$
b1 %
1'
1*
b1 +
#493080000000
0!
0'
#493090000000
1!
b10 %
1'
b10 +
#493100000000
0!
0'
#493110000000
1!
b11 %
1'
b11 +
#493120000000
0!
0'
#493130000000
1!
b100 %
1'
b100 +
#493140000000
0!
0'
#493150000000
1!
b101 %
1'
b101 +
#493160000000
0!
0'
#493170000000
1!
b110 %
1'
b110 +
#493180000000
0!
0'
#493190000000
1!
b111 %
1'
b111 +
#493200000000
0!
0'
#493210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#493220000000
0!
0'
#493230000000
1!
b1001 %
1'
b1001 +
#493240000000
0!
0'
#493250000000
1!
b0 %
1'
b0 +
#493260000000
0!
0'
#493270000000
1!
1$
b1 %
1'
1*
b1 +
#493280000000
0!
0'
#493290000000
1!
b10 %
1'
b10 +
#493300000000
0!
0'
#493310000000
1!
b11 %
1'
b11 +
#493320000000
0!
0'
#493330000000
1!
b100 %
1'
b100 +
#493340000000
0!
0'
#493350000000
1!
b101 %
1'
b101 +
#493360000000
0!
0'
#493370000000
1!
0$
b110 %
1'
0*
b110 +
#493380000000
0!
0'
#493390000000
1!
b111 %
1'
b111 +
#493400000000
0!
0'
#493410000000
1!
b1000 %
1'
b1000 +
#493420000000
1"
1(
#493430000000
0!
0"
b100 &
0'
0(
b100 ,
#493440000000
1!
b1001 %
1'
b1001 +
#493450000000
0!
0'
#493460000000
1!
b0 %
1'
b0 +
#493470000000
0!
0'
#493480000000
1!
1$
b1 %
1'
1*
b1 +
#493490000000
0!
0'
#493500000000
1!
b10 %
1'
b10 +
#493510000000
0!
0'
#493520000000
1!
b11 %
1'
b11 +
#493530000000
0!
0'
#493540000000
1!
b100 %
1'
b100 +
#493550000000
0!
0'
#493560000000
1!
b101 %
1'
b101 +
#493570000000
0!
0'
#493580000000
1!
b110 %
1'
b110 +
#493590000000
0!
0'
#493600000000
1!
b111 %
1'
b111 +
#493610000000
0!
0'
#493620000000
1!
0$
b1000 %
1'
0*
b1000 +
#493630000000
0!
0'
#493640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#493650000000
0!
0'
#493660000000
1!
b0 %
1'
b0 +
#493670000000
0!
0'
#493680000000
1!
1$
b1 %
1'
1*
b1 +
#493690000000
0!
0'
#493700000000
1!
b10 %
1'
b10 +
#493710000000
0!
0'
#493720000000
1!
b11 %
1'
b11 +
#493730000000
0!
0'
#493740000000
1!
b100 %
1'
b100 +
#493750000000
0!
0'
#493760000000
1!
b101 %
1'
b101 +
#493770000000
0!
0'
#493780000000
1!
0$
b110 %
1'
0*
b110 +
#493790000000
0!
0'
#493800000000
1!
b111 %
1'
b111 +
#493810000000
0!
0'
#493820000000
1!
b1000 %
1'
b1000 +
#493830000000
0!
0'
#493840000000
1!
b1001 %
1'
b1001 +
#493850000000
1"
1(
#493860000000
0!
0"
b100 &
0'
0(
b100 ,
#493870000000
1!
b0 %
1'
b0 +
#493880000000
0!
0'
#493890000000
1!
1$
b1 %
1'
1*
b1 +
#493900000000
0!
0'
#493910000000
1!
b10 %
1'
b10 +
#493920000000
0!
0'
#493930000000
1!
b11 %
1'
b11 +
#493940000000
0!
0'
#493950000000
1!
b100 %
1'
b100 +
#493960000000
0!
0'
#493970000000
1!
b101 %
1'
b101 +
#493980000000
0!
0'
#493990000000
1!
b110 %
1'
b110 +
#494000000000
0!
0'
#494010000000
1!
b111 %
1'
b111 +
#494020000000
0!
0'
#494030000000
1!
0$
b1000 %
1'
0*
b1000 +
#494040000000
0!
0'
#494050000000
1!
b1001 %
1'
b1001 +
#494060000000
0!
0'
#494070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#494080000000
0!
0'
#494090000000
1!
1$
b1 %
1'
1*
b1 +
#494100000000
0!
0'
#494110000000
1!
b10 %
1'
b10 +
#494120000000
0!
0'
#494130000000
1!
b11 %
1'
b11 +
#494140000000
0!
0'
#494150000000
1!
b100 %
1'
b100 +
#494160000000
0!
0'
#494170000000
1!
b101 %
1'
b101 +
#494180000000
0!
0'
#494190000000
1!
0$
b110 %
1'
0*
b110 +
#494200000000
0!
0'
#494210000000
1!
b111 %
1'
b111 +
#494220000000
0!
0'
#494230000000
1!
b1000 %
1'
b1000 +
#494240000000
0!
0'
#494250000000
1!
b1001 %
1'
b1001 +
#494260000000
0!
0'
#494270000000
1!
b0 %
1'
b0 +
#494280000000
1"
1(
#494290000000
0!
0"
b100 &
0'
0(
b100 ,
#494300000000
1!
1$
b1 %
1'
1*
b1 +
#494310000000
0!
0'
#494320000000
1!
b10 %
1'
b10 +
#494330000000
0!
0'
#494340000000
1!
b11 %
1'
b11 +
#494350000000
0!
0'
#494360000000
1!
b100 %
1'
b100 +
#494370000000
0!
0'
#494380000000
1!
b101 %
1'
b101 +
#494390000000
0!
0'
#494400000000
1!
b110 %
1'
b110 +
#494410000000
0!
0'
#494420000000
1!
b111 %
1'
b111 +
#494430000000
0!
0'
#494440000000
1!
0$
b1000 %
1'
0*
b1000 +
#494450000000
0!
0'
#494460000000
1!
b1001 %
1'
b1001 +
#494470000000
0!
0'
#494480000000
1!
b0 %
1'
b0 +
#494490000000
0!
0'
#494500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#494510000000
0!
0'
#494520000000
1!
b10 %
1'
b10 +
#494530000000
0!
0'
#494540000000
1!
b11 %
1'
b11 +
#494550000000
0!
0'
#494560000000
1!
b100 %
1'
b100 +
#494570000000
0!
0'
#494580000000
1!
b101 %
1'
b101 +
#494590000000
0!
0'
#494600000000
1!
0$
b110 %
1'
0*
b110 +
#494610000000
0!
0'
#494620000000
1!
b111 %
1'
b111 +
#494630000000
0!
0'
#494640000000
1!
b1000 %
1'
b1000 +
#494650000000
0!
0'
#494660000000
1!
b1001 %
1'
b1001 +
#494670000000
0!
0'
#494680000000
1!
b0 %
1'
b0 +
#494690000000
0!
0'
#494700000000
1!
1$
b1 %
1'
1*
b1 +
#494710000000
1"
1(
#494720000000
0!
0"
b100 &
0'
0(
b100 ,
#494730000000
1!
b10 %
1'
b10 +
#494740000000
0!
0'
#494750000000
1!
b11 %
1'
b11 +
#494760000000
0!
0'
#494770000000
1!
b100 %
1'
b100 +
#494780000000
0!
0'
#494790000000
1!
b101 %
1'
b101 +
#494800000000
0!
0'
#494810000000
1!
b110 %
1'
b110 +
#494820000000
0!
0'
#494830000000
1!
b111 %
1'
b111 +
#494840000000
0!
0'
#494850000000
1!
0$
b1000 %
1'
0*
b1000 +
#494860000000
0!
0'
#494870000000
1!
b1001 %
1'
b1001 +
#494880000000
0!
0'
#494890000000
1!
b0 %
1'
b0 +
#494900000000
0!
0'
#494910000000
1!
1$
b1 %
1'
1*
b1 +
#494920000000
0!
0'
#494930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#494940000000
0!
0'
#494950000000
1!
b11 %
1'
b11 +
#494960000000
0!
0'
#494970000000
1!
b100 %
1'
b100 +
#494980000000
0!
0'
#494990000000
1!
b101 %
1'
b101 +
#495000000000
0!
0'
#495010000000
1!
0$
b110 %
1'
0*
b110 +
#495020000000
0!
0'
#495030000000
1!
b111 %
1'
b111 +
#495040000000
0!
0'
#495050000000
1!
b1000 %
1'
b1000 +
#495060000000
0!
0'
#495070000000
1!
b1001 %
1'
b1001 +
#495080000000
0!
0'
#495090000000
1!
b0 %
1'
b0 +
#495100000000
0!
0'
#495110000000
1!
1$
b1 %
1'
1*
b1 +
#495120000000
0!
0'
#495130000000
1!
b10 %
1'
b10 +
#495140000000
1"
1(
#495150000000
0!
0"
b100 &
0'
0(
b100 ,
#495160000000
1!
b11 %
1'
b11 +
#495170000000
0!
0'
#495180000000
1!
b100 %
1'
b100 +
#495190000000
0!
0'
#495200000000
1!
b101 %
1'
b101 +
#495210000000
0!
0'
#495220000000
1!
b110 %
1'
b110 +
#495230000000
0!
0'
#495240000000
1!
b111 %
1'
b111 +
#495250000000
0!
0'
#495260000000
1!
0$
b1000 %
1'
0*
b1000 +
#495270000000
0!
0'
#495280000000
1!
b1001 %
1'
b1001 +
#495290000000
0!
0'
#495300000000
1!
b0 %
1'
b0 +
#495310000000
0!
0'
#495320000000
1!
1$
b1 %
1'
1*
b1 +
#495330000000
0!
0'
#495340000000
1!
b10 %
1'
b10 +
#495350000000
0!
0'
#495360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#495370000000
0!
0'
#495380000000
1!
b100 %
1'
b100 +
#495390000000
0!
0'
#495400000000
1!
b101 %
1'
b101 +
#495410000000
0!
0'
#495420000000
1!
0$
b110 %
1'
0*
b110 +
#495430000000
0!
0'
#495440000000
1!
b111 %
1'
b111 +
#495450000000
0!
0'
#495460000000
1!
b1000 %
1'
b1000 +
#495470000000
0!
0'
#495480000000
1!
b1001 %
1'
b1001 +
#495490000000
0!
0'
#495500000000
1!
b0 %
1'
b0 +
#495510000000
0!
0'
#495520000000
1!
1$
b1 %
1'
1*
b1 +
#495530000000
0!
0'
#495540000000
1!
b10 %
1'
b10 +
#495550000000
0!
0'
#495560000000
1!
b11 %
1'
b11 +
#495570000000
1"
1(
#495580000000
0!
0"
b100 &
0'
0(
b100 ,
#495590000000
1!
b100 %
1'
b100 +
#495600000000
0!
0'
#495610000000
1!
b101 %
1'
b101 +
#495620000000
0!
0'
#495630000000
1!
b110 %
1'
b110 +
#495640000000
0!
0'
#495650000000
1!
b111 %
1'
b111 +
#495660000000
0!
0'
#495670000000
1!
0$
b1000 %
1'
0*
b1000 +
#495680000000
0!
0'
#495690000000
1!
b1001 %
1'
b1001 +
#495700000000
0!
0'
#495710000000
1!
b0 %
1'
b0 +
#495720000000
0!
0'
#495730000000
1!
1$
b1 %
1'
1*
b1 +
#495740000000
0!
0'
#495750000000
1!
b10 %
1'
b10 +
#495760000000
0!
0'
#495770000000
1!
b11 %
1'
b11 +
#495780000000
0!
0'
#495790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#495800000000
0!
0'
#495810000000
1!
b101 %
1'
b101 +
#495820000000
0!
0'
#495830000000
1!
0$
b110 %
1'
0*
b110 +
#495840000000
0!
0'
#495850000000
1!
b111 %
1'
b111 +
#495860000000
0!
0'
#495870000000
1!
b1000 %
1'
b1000 +
#495880000000
0!
0'
#495890000000
1!
b1001 %
1'
b1001 +
#495900000000
0!
0'
#495910000000
1!
b0 %
1'
b0 +
#495920000000
0!
0'
#495930000000
1!
1$
b1 %
1'
1*
b1 +
#495940000000
0!
0'
#495950000000
1!
b10 %
1'
b10 +
#495960000000
0!
0'
#495970000000
1!
b11 %
1'
b11 +
#495980000000
0!
0'
#495990000000
1!
b100 %
1'
b100 +
#496000000000
1"
1(
#496010000000
0!
0"
b100 &
0'
0(
b100 ,
#496020000000
1!
b101 %
1'
b101 +
#496030000000
0!
0'
#496040000000
1!
b110 %
1'
b110 +
#496050000000
0!
0'
#496060000000
1!
b111 %
1'
b111 +
#496070000000
0!
0'
#496080000000
1!
0$
b1000 %
1'
0*
b1000 +
#496090000000
0!
0'
#496100000000
1!
b1001 %
1'
b1001 +
#496110000000
0!
0'
#496120000000
1!
b0 %
1'
b0 +
#496130000000
0!
0'
#496140000000
1!
1$
b1 %
1'
1*
b1 +
#496150000000
0!
0'
#496160000000
1!
b10 %
1'
b10 +
#496170000000
0!
0'
#496180000000
1!
b11 %
1'
b11 +
#496190000000
0!
0'
#496200000000
1!
b100 %
1'
b100 +
#496210000000
0!
0'
#496220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#496230000000
0!
0'
#496240000000
1!
0$
b110 %
1'
0*
b110 +
#496250000000
0!
0'
#496260000000
1!
b111 %
1'
b111 +
#496270000000
0!
0'
#496280000000
1!
b1000 %
1'
b1000 +
#496290000000
0!
0'
#496300000000
1!
b1001 %
1'
b1001 +
#496310000000
0!
0'
#496320000000
1!
b0 %
1'
b0 +
#496330000000
0!
0'
#496340000000
1!
1$
b1 %
1'
1*
b1 +
#496350000000
0!
0'
#496360000000
1!
b10 %
1'
b10 +
#496370000000
0!
0'
#496380000000
1!
b11 %
1'
b11 +
#496390000000
0!
0'
#496400000000
1!
b100 %
1'
b100 +
#496410000000
0!
0'
#496420000000
1!
b101 %
1'
b101 +
#496430000000
1"
1(
#496440000000
0!
0"
b100 &
0'
0(
b100 ,
#496450000000
1!
b110 %
1'
b110 +
#496460000000
0!
0'
#496470000000
1!
b111 %
1'
b111 +
#496480000000
0!
0'
#496490000000
1!
0$
b1000 %
1'
0*
b1000 +
#496500000000
0!
0'
#496510000000
1!
b1001 %
1'
b1001 +
#496520000000
0!
0'
#496530000000
1!
b0 %
1'
b0 +
#496540000000
0!
0'
#496550000000
1!
1$
b1 %
1'
1*
b1 +
#496560000000
0!
0'
#496570000000
1!
b10 %
1'
b10 +
#496580000000
0!
0'
#496590000000
1!
b11 %
1'
b11 +
#496600000000
0!
0'
#496610000000
1!
b100 %
1'
b100 +
#496620000000
0!
0'
#496630000000
1!
b101 %
1'
b101 +
#496640000000
0!
0'
#496650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#496660000000
0!
0'
#496670000000
1!
b111 %
1'
b111 +
#496680000000
0!
0'
#496690000000
1!
b1000 %
1'
b1000 +
#496700000000
0!
0'
#496710000000
1!
b1001 %
1'
b1001 +
#496720000000
0!
0'
#496730000000
1!
b0 %
1'
b0 +
#496740000000
0!
0'
#496750000000
1!
1$
b1 %
1'
1*
b1 +
#496760000000
0!
0'
#496770000000
1!
b10 %
1'
b10 +
#496780000000
0!
0'
#496790000000
1!
b11 %
1'
b11 +
#496800000000
0!
0'
#496810000000
1!
b100 %
1'
b100 +
#496820000000
0!
0'
#496830000000
1!
b101 %
1'
b101 +
#496840000000
0!
0'
#496850000000
1!
0$
b110 %
1'
0*
b110 +
#496860000000
1"
1(
#496870000000
0!
0"
b100 &
0'
0(
b100 ,
#496880000000
1!
1$
b111 %
1'
1*
b111 +
#496890000000
0!
0'
#496900000000
1!
0$
b1000 %
1'
0*
b1000 +
#496910000000
0!
0'
#496920000000
1!
b1001 %
1'
b1001 +
#496930000000
0!
0'
#496940000000
1!
b0 %
1'
b0 +
#496950000000
0!
0'
#496960000000
1!
1$
b1 %
1'
1*
b1 +
#496970000000
0!
0'
#496980000000
1!
b10 %
1'
b10 +
#496990000000
0!
0'
#497000000000
1!
b11 %
1'
b11 +
#497010000000
0!
0'
#497020000000
1!
b100 %
1'
b100 +
#497030000000
0!
0'
#497040000000
1!
b101 %
1'
b101 +
#497050000000
0!
0'
#497060000000
1!
b110 %
1'
b110 +
#497070000000
0!
0'
#497080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#497090000000
0!
0'
#497100000000
1!
b1000 %
1'
b1000 +
#497110000000
0!
0'
#497120000000
1!
b1001 %
1'
b1001 +
#497130000000
0!
0'
#497140000000
1!
b0 %
1'
b0 +
#497150000000
0!
0'
#497160000000
1!
1$
b1 %
1'
1*
b1 +
#497170000000
0!
0'
#497180000000
1!
b10 %
1'
b10 +
#497190000000
0!
0'
#497200000000
1!
b11 %
1'
b11 +
#497210000000
0!
0'
#497220000000
1!
b100 %
1'
b100 +
#497230000000
0!
0'
#497240000000
1!
b101 %
1'
b101 +
#497250000000
0!
0'
#497260000000
1!
0$
b110 %
1'
0*
b110 +
#497270000000
0!
0'
#497280000000
1!
b111 %
1'
b111 +
#497290000000
1"
1(
#497300000000
0!
0"
b100 &
0'
0(
b100 ,
#497310000000
1!
b1000 %
1'
b1000 +
#497320000000
0!
0'
#497330000000
1!
b1001 %
1'
b1001 +
#497340000000
0!
0'
#497350000000
1!
b0 %
1'
b0 +
#497360000000
0!
0'
#497370000000
1!
1$
b1 %
1'
1*
b1 +
#497380000000
0!
0'
#497390000000
1!
b10 %
1'
b10 +
#497400000000
0!
0'
#497410000000
1!
b11 %
1'
b11 +
#497420000000
0!
0'
#497430000000
1!
b100 %
1'
b100 +
#497440000000
0!
0'
#497450000000
1!
b101 %
1'
b101 +
#497460000000
0!
0'
#497470000000
1!
b110 %
1'
b110 +
#497480000000
0!
0'
#497490000000
1!
b111 %
1'
b111 +
#497500000000
0!
0'
#497510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#497520000000
0!
0'
#497530000000
1!
b1001 %
1'
b1001 +
#497540000000
0!
0'
#497550000000
1!
b0 %
1'
b0 +
#497560000000
0!
0'
#497570000000
1!
1$
b1 %
1'
1*
b1 +
#497580000000
0!
0'
#497590000000
1!
b10 %
1'
b10 +
#497600000000
0!
0'
#497610000000
1!
b11 %
1'
b11 +
#497620000000
0!
0'
#497630000000
1!
b100 %
1'
b100 +
#497640000000
0!
0'
#497650000000
1!
b101 %
1'
b101 +
#497660000000
0!
0'
#497670000000
1!
0$
b110 %
1'
0*
b110 +
#497680000000
0!
0'
#497690000000
1!
b111 %
1'
b111 +
#497700000000
0!
0'
#497710000000
1!
b1000 %
1'
b1000 +
#497720000000
1"
1(
#497730000000
0!
0"
b100 &
0'
0(
b100 ,
#497740000000
1!
b1001 %
1'
b1001 +
#497750000000
0!
0'
#497760000000
1!
b0 %
1'
b0 +
#497770000000
0!
0'
#497780000000
1!
1$
b1 %
1'
1*
b1 +
#497790000000
0!
0'
#497800000000
1!
b10 %
1'
b10 +
#497810000000
0!
0'
#497820000000
1!
b11 %
1'
b11 +
#497830000000
0!
0'
#497840000000
1!
b100 %
1'
b100 +
#497850000000
0!
0'
#497860000000
1!
b101 %
1'
b101 +
#497870000000
0!
0'
#497880000000
1!
b110 %
1'
b110 +
#497890000000
0!
0'
#497900000000
1!
b111 %
1'
b111 +
#497910000000
0!
0'
#497920000000
1!
0$
b1000 %
1'
0*
b1000 +
#497930000000
0!
0'
#497940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#497950000000
0!
0'
#497960000000
1!
b0 %
1'
b0 +
#497970000000
0!
0'
#497980000000
1!
1$
b1 %
1'
1*
b1 +
#497990000000
0!
0'
#498000000000
1!
b10 %
1'
b10 +
#498010000000
0!
0'
#498020000000
1!
b11 %
1'
b11 +
#498030000000
0!
0'
#498040000000
1!
b100 %
1'
b100 +
#498050000000
0!
0'
#498060000000
1!
b101 %
1'
b101 +
#498070000000
0!
0'
#498080000000
1!
0$
b110 %
1'
0*
b110 +
#498090000000
0!
0'
#498100000000
1!
b111 %
1'
b111 +
#498110000000
0!
0'
#498120000000
1!
b1000 %
1'
b1000 +
#498130000000
0!
0'
#498140000000
1!
b1001 %
1'
b1001 +
#498150000000
1"
1(
#498160000000
0!
0"
b100 &
0'
0(
b100 ,
#498170000000
1!
b0 %
1'
b0 +
#498180000000
0!
0'
#498190000000
1!
1$
b1 %
1'
1*
b1 +
#498200000000
0!
0'
#498210000000
1!
b10 %
1'
b10 +
#498220000000
0!
0'
#498230000000
1!
b11 %
1'
b11 +
#498240000000
0!
0'
#498250000000
1!
b100 %
1'
b100 +
#498260000000
0!
0'
#498270000000
1!
b101 %
1'
b101 +
#498280000000
0!
0'
#498290000000
1!
b110 %
1'
b110 +
#498300000000
0!
0'
#498310000000
1!
b111 %
1'
b111 +
#498320000000
0!
0'
#498330000000
1!
0$
b1000 %
1'
0*
b1000 +
#498340000000
0!
0'
#498350000000
1!
b1001 %
1'
b1001 +
#498360000000
0!
0'
#498370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#498380000000
0!
0'
#498390000000
1!
1$
b1 %
1'
1*
b1 +
#498400000000
0!
0'
#498410000000
1!
b10 %
1'
b10 +
#498420000000
0!
0'
#498430000000
1!
b11 %
1'
b11 +
#498440000000
0!
0'
#498450000000
1!
b100 %
1'
b100 +
#498460000000
0!
0'
#498470000000
1!
b101 %
1'
b101 +
#498480000000
0!
0'
#498490000000
1!
0$
b110 %
1'
0*
b110 +
#498500000000
0!
0'
#498510000000
1!
b111 %
1'
b111 +
#498520000000
0!
0'
#498530000000
1!
b1000 %
1'
b1000 +
#498540000000
0!
0'
#498550000000
1!
b1001 %
1'
b1001 +
#498560000000
0!
0'
#498570000000
1!
b0 %
1'
b0 +
#498580000000
1"
1(
#498590000000
0!
0"
b100 &
0'
0(
b100 ,
#498600000000
1!
1$
b1 %
1'
1*
b1 +
#498610000000
0!
0'
#498620000000
1!
b10 %
1'
b10 +
#498630000000
0!
0'
#498640000000
1!
b11 %
1'
b11 +
#498650000000
0!
0'
#498660000000
1!
b100 %
1'
b100 +
#498670000000
0!
0'
#498680000000
1!
b101 %
1'
b101 +
#498690000000
0!
0'
#498700000000
1!
b110 %
1'
b110 +
#498710000000
0!
0'
#498720000000
1!
b111 %
1'
b111 +
#498730000000
0!
0'
#498740000000
1!
0$
b1000 %
1'
0*
b1000 +
#498750000000
0!
0'
#498760000000
1!
b1001 %
1'
b1001 +
#498770000000
0!
0'
#498780000000
1!
b0 %
1'
b0 +
#498790000000
0!
0'
#498800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#498810000000
0!
0'
#498820000000
1!
b10 %
1'
b10 +
#498830000000
0!
0'
#498840000000
1!
b11 %
1'
b11 +
#498850000000
0!
0'
#498860000000
1!
b100 %
1'
b100 +
#498870000000
0!
0'
#498880000000
1!
b101 %
1'
b101 +
#498890000000
0!
0'
#498900000000
1!
0$
b110 %
1'
0*
b110 +
#498910000000
0!
0'
#498920000000
1!
b111 %
1'
b111 +
#498930000000
0!
0'
#498940000000
1!
b1000 %
1'
b1000 +
#498950000000
0!
0'
#498960000000
1!
b1001 %
1'
b1001 +
#498970000000
0!
0'
#498980000000
1!
b0 %
1'
b0 +
#498990000000
0!
0'
#499000000000
1!
1$
b1 %
1'
1*
b1 +
#499010000000
1"
1(
#499020000000
0!
0"
b100 &
0'
0(
b100 ,
#499030000000
1!
b10 %
1'
b10 +
#499040000000
0!
0'
#499050000000
1!
b11 %
1'
b11 +
#499060000000
0!
0'
#499070000000
1!
b100 %
1'
b100 +
#499080000000
0!
0'
#499090000000
1!
b101 %
1'
b101 +
#499100000000
0!
0'
#499110000000
1!
b110 %
1'
b110 +
#499120000000
0!
0'
#499130000000
1!
b111 %
1'
b111 +
#499140000000
0!
0'
#499150000000
1!
0$
b1000 %
1'
0*
b1000 +
#499160000000
0!
0'
#499170000000
1!
b1001 %
1'
b1001 +
#499180000000
0!
0'
#499190000000
1!
b0 %
1'
b0 +
#499200000000
0!
0'
#499210000000
1!
1$
b1 %
1'
1*
b1 +
#499220000000
0!
0'
#499230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#499240000000
0!
0'
#499250000000
1!
b11 %
1'
b11 +
#499260000000
0!
0'
#499270000000
1!
b100 %
1'
b100 +
#499280000000
0!
0'
#499290000000
1!
b101 %
1'
b101 +
#499300000000
0!
0'
#499310000000
1!
0$
b110 %
1'
0*
b110 +
#499320000000
0!
0'
#499330000000
1!
b111 %
1'
b111 +
#499340000000
0!
0'
#499350000000
1!
b1000 %
1'
b1000 +
#499360000000
0!
0'
#499370000000
1!
b1001 %
1'
b1001 +
#499380000000
0!
0'
#499390000000
1!
b0 %
1'
b0 +
#499400000000
0!
0'
#499410000000
1!
1$
b1 %
1'
1*
b1 +
#499420000000
0!
0'
#499430000000
1!
b10 %
1'
b10 +
#499440000000
1"
1(
#499450000000
0!
0"
b100 &
0'
0(
b100 ,
#499460000000
1!
b11 %
1'
b11 +
#499470000000
0!
0'
#499480000000
1!
b100 %
1'
b100 +
#499490000000
0!
0'
#499500000000
1!
b101 %
1'
b101 +
#499510000000
0!
0'
#499520000000
1!
b110 %
1'
b110 +
#499530000000
0!
0'
#499540000000
1!
b111 %
1'
b111 +
#499550000000
0!
0'
#499560000000
1!
0$
b1000 %
1'
0*
b1000 +
#499570000000
0!
0'
#499580000000
1!
b1001 %
1'
b1001 +
#499590000000
0!
0'
#499600000000
1!
b0 %
1'
b0 +
#499610000000
0!
0'
#499620000000
1!
1$
b1 %
1'
1*
b1 +
#499630000000
0!
0'
#499640000000
1!
b10 %
1'
b10 +
#499650000000
0!
0'
#499660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#499670000000
0!
0'
#499680000000
1!
b100 %
1'
b100 +
#499690000000
0!
0'
#499700000000
1!
b101 %
1'
b101 +
#499710000000
0!
0'
#499720000000
1!
0$
b110 %
1'
0*
b110 +
#499730000000
0!
0'
#499740000000
1!
b111 %
1'
b111 +
#499750000000
0!
0'
#499760000000
1!
b1000 %
1'
b1000 +
#499770000000
0!
0'
#499780000000
1!
b1001 %
1'
b1001 +
#499790000000
0!
0'
#499800000000
1!
b0 %
1'
b0 +
#499810000000
0!
0'
#499820000000
1!
1$
b1 %
1'
1*
b1 +
#499830000000
0!
0'
#499840000000
1!
b10 %
1'
b10 +
#499850000000
0!
0'
#499860000000
1!
b11 %
1'
b11 +
#499870000000
1"
1(
#499880000000
0!
0"
b100 &
0'
0(
b100 ,
#499890000000
1!
b100 %
1'
b100 +
#499900000000
0!
0'
#499910000000
1!
b101 %
1'
b101 +
#499920000000
0!
0'
#499930000000
1!
b110 %
1'
b110 +
#499940000000
0!
0'
#499950000000
1!
b111 %
1'
b111 +
#499960000000
0!
0'
#499970000000
1!
0$
b1000 %
1'
0*
b1000 +
#499980000000
0!
0'
#499990000000
1!
b1001 %
1'
b1001 +
#500000000000
0!
0'
#500010000000
1!
b0 %
1'
b0 +
#500020000000
0!
0'
#500030000000
1!
1$
b1 %
1'
1*
b1 +
#500040000000
0!
0'
#500050000000
1!
b10 %
1'
b10 +
#500060000000
0!
0'
#500070000000
1!
b11 %
1'
b11 +
#500080000000
0!
0'
#500090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#500100000000
0!
0'
#500110000000
1!
b101 %
1'
b101 +
#500120000000
0!
0'
#500130000000
1!
0$
b110 %
1'
0*
b110 +
#500140000000
0!
0'
#500150000000
1!
b111 %
1'
b111 +
#500160000000
0!
0'
#500170000000
1!
b1000 %
1'
b1000 +
#500180000000
0!
0'
#500190000000
1!
b1001 %
1'
b1001 +
#500200000000
0!
0'
#500210000000
1!
b0 %
1'
b0 +
#500220000000
0!
0'
#500230000000
1!
1$
b1 %
1'
1*
b1 +
#500240000000
0!
0'
#500250000000
1!
b10 %
1'
b10 +
#500260000000
0!
0'
#500270000000
1!
b11 %
1'
b11 +
#500280000000
0!
0'
#500290000000
1!
b100 %
1'
b100 +
#500300000000
1"
1(
#500310000000
0!
0"
b100 &
0'
0(
b100 ,
#500320000000
1!
b101 %
1'
b101 +
#500330000000
0!
0'
#500340000000
1!
b110 %
1'
b110 +
#500350000000
0!
0'
#500360000000
1!
b111 %
1'
b111 +
#500370000000
0!
0'
#500380000000
1!
0$
b1000 %
1'
0*
b1000 +
#500390000000
0!
0'
#500400000000
1!
b1001 %
1'
b1001 +
#500410000000
0!
0'
#500420000000
1!
b0 %
1'
b0 +
#500430000000
0!
0'
#500440000000
1!
1$
b1 %
1'
1*
b1 +
#500450000000
0!
0'
#500460000000
1!
b10 %
1'
b10 +
#500470000000
0!
0'
#500480000000
1!
b11 %
1'
b11 +
#500490000000
0!
0'
#500500000000
1!
b100 %
1'
b100 +
#500510000000
0!
0'
#500520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#500530000000
0!
0'
#500540000000
1!
0$
b110 %
1'
0*
b110 +
#500550000000
0!
0'
#500560000000
1!
b111 %
1'
b111 +
#500570000000
0!
0'
#500580000000
1!
b1000 %
1'
b1000 +
#500590000000
0!
0'
#500600000000
1!
b1001 %
1'
b1001 +
#500610000000
0!
0'
#500620000000
1!
b0 %
1'
b0 +
#500630000000
0!
0'
#500640000000
1!
1$
b1 %
1'
1*
b1 +
#500650000000
0!
0'
#500660000000
1!
b10 %
1'
b10 +
#500670000000
0!
0'
#500680000000
1!
b11 %
1'
b11 +
#500690000000
0!
0'
#500700000000
1!
b100 %
1'
b100 +
#500710000000
0!
0'
#500720000000
1!
b101 %
1'
b101 +
#500730000000
1"
1(
#500740000000
0!
0"
b100 &
0'
0(
b100 ,
#500750000000
1!
b110 %
1'
b110 +
#500760000000
0!
0'
#500770000000
1!
b111 %
1'
b111 +
#500780000000
0!
0'
#500790000000
1!
0$
b1000 %
1'
0*
b1000 +
#500800000000
0!
0'
#500810000000
1!
b1001 %
1'
b1001 +
#500820000000
0!
0'
#500830000000
1!
b0 %
1'
b0 +
#500840000000
0!
0'
#500850000000
1!
1$
b1 %
1'
1*
b1 +
#500860000000
0!
0'
#500870000000
1!
b10 %
1'
b10 +
#500880000000
0!
0'
#500890000000
1!
b11 %
1'
b11 +
#500900000000
0!
0'
#500910000000
1!
b100 %
1'
b100 +
#500920000000
0!
0'
#500930000000
1!
b101 %
1'
b101 +
#500940000000
0!
0'
#500950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#500960000000
0!
0'
#500970000000
1!
b111 %
1'
b111 +
#500980000000
0!
0'
#500990000000
1!
b1000 %
1'
b1000 +
#501000000000
0!
0'
#501010000000
1!
b1001 %
1'
b1001 +
#501020000000
0!
0'
#501030000000
1!
b0 %
1'
b0 +
#501040000000
0!
0'
#501050000000
1!
1$
b1 %
1'
1*
b1 +
#501060000000
0!
0'
#501070000000
1!
b10 %
1'
b10 +
#501080000000
0!
0'
#501090000000
1!
b11 %
1'
b11 +
#501100000000
0!
0'
#501110000000
1!
b100 %
1'
b100 +
#501120000000
0!
0'
#501130000000
1!
b101 %
1'
b101 +
#501140000000
0!
0'
#501150000000
1!
0$
b110 %
1'
0*
b110 +
#501160000000
1"
1(
#501170000000
0!
0"
b100 &
0'
0(
b100 ,
#501180000000
1!
1$
b111 %
1'
1*
b111 +
#501190000000
0!
0'
#501200000000
1!
0$
b1000 %
1'
0*
b1000 +
#501210000000
0!
0'
#501220000000
1!
b1001 %
1'
b1001 +
#501230000000
0!
0'
#501240000000
1!
b0 %
1'
b0 +
#501250000000
0!
0'
#501260000000
1!
1$
b1 %
1'
1*
b1 +
#501270000000
0!
0'
#501280000000
1!
b10 %
1'
b10 +
#501290000000
0!
0'
#501300000000
1!
b11 %
1'
b11 +
#501310000000
0!
0'
#501320000000
1!
b100 %
1'
b100 +
#501330000000
0!
0'
#501340000000
1!
b101 %
1'
b101 +
#501350000000
0!
0'
#501360000000
1!
b110 %
1'
b110 +
#501370000000
0!
0'
#501380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#501390000000
0!
0'
#501400000000
1!
b1000 %
1'
b1000 +
#501410000000
0!
0'
#501420000000
1!
b1001 %
1'
b1001 +
#501430000000
0!
0'
#501440000000
1!
b0 %
1'
b0 +
#501450000000
0!
0'
#501460000000
1!
1$
b1 %
1'
1*
b1 +
#501470000000
0!
0'
#501480000000
1!
b10 %
1'
b10 +
#501490000000
0!
0'
#501500000000
1!
b11 %
1'
b11 +
#501510000000
0!
0'
#501520000000
1!
b100 %
1'
b100 +
#501530000000
0!
0'
#501540000000
1!
b101 %
1'
b101 +
#501550000000
0!
0'
#501560000000
1!
0$
b110 %
1'
0*
b110 +
#501570000000
0!
0'
#501580000000
1!
b111 %
1'
b111 +
#501590000000
1"
1(
#501600000000
0!
0"
b100 &
0'
0(
b100 ,
#501610000000
1!
b1000 %
1'
b1000 +
#501620000000
0!
0'
#501630000000
1!
b1001 %
1'
b1001 +
#501640000000
0!
0'
#501650000000
1!
b0 %
1'
b0 +
#501660000000
0!
0'
#501670000000
1!
1$
b1 %
1'
1*
b1 +
#501680000000
0!
0'
#501690000000
1!
b10 %
1'
b10 +
#501700000000
0!
0'
#501710000000
1!
b11 %
1'
b11 +
#501720000000
0!
0'
#501730000000
1!
b100 %
1'
b100 +
#501740000000
0!
0'
#501750000000
1!
b101 %
1'
b101 +
#501760000000
0!
0'
#501770000000
1!
b110 %
1'
b110 +
#501780000000
0!
0'
#501790000000
1!
b111 %
1'
b111 +
#501800000000
0!
0'
#501810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#501820000000
0!
0'
#501830000000
1!
b1001 %
1'
b1001 +
#501840000000
0!
0'
#501850000000
1!
b0 %
1'
b0 +
#501860000000
0!
0'
#501870000000
1!
1$
b1 %
1'
1*
b1 +
#501880000000
0!
0'
#501890000000
1!
b10 %
1'
b10 +
#501900000000
0!
0'
#501910000000
1!
b11 %
1'
b11 +
#501920000000
0!
0'
#501930000000
1!
b100 %
1'
b100 +
#501940000000
0!
0'
#501950000000
1!
b101 %
1'
b101 +
#501960000000
0!
0'
#501970000000
1!
0$
b110 %
1'
0*
b110 +
#501980000000
0!
0'
#501990000000
1!
b111 %
1'
b111 +
#502000000000
0!
0'
#502010000000
1!
b1000 %
1'
b1000 +
#502020000000
1"
1(
#502030000000
0!
0"
b100 &
0'
0(
b100 ,
#502040000000
1!
b1001 %
1'
b1001 +
#502050000000
0!
0'
#502060000000
1!
b0 %
1'
b0 +
#502070000000
0!
0'
#502080000000
1!
1$
b1 %
1'
1*
b1 +
#502090000000
0!
0'
#502100000000
1!
b10 %
1'
b10 +
#502110000000
0!
0'
#502120000000
1!
b11 %
1'
b11 +
#502130000000
0!
0'
#502140000000
1!
b100 %
1'
b100 +
#502150000000
0!
0'
#502160000000
1!
b101 %
1'
b101 +
#502170000000
0!
0'
#502180000000
1!
b110 %
1'
b110 +
#502190000000
0!
0'
#502200000000
1!
b111 %
1'
b111 +
#502210000000
0!
0'
#502220000000
1!
0$
b1000 %
1'
0*
b1000 +
#502230000000
0!
0'
#502240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#502250000000
0!
0'
#502260000000
1!
b0 %
1'
b0 +
#502270000000
0!
0'
#502280000000
1!
1$
b1 %
1'
1*
b1 +
#502290000000
0!
0'
#502300000000
1!
b10 %
1'
b10 +
#502310000000
0!
0'
#502320000000
1!
b11 %
1'
b11 +
#502330000000
0!
0'
#502340000000
1!
b100 %
1'
b100 +
#502350000000
0!
0'
#502360000000
1!
b101 %
1'
b101 +
#502370000000
0!
0'
#502380000000
1!
0$
b110 %
1'
0*
b110 +
#502390000000
0!
0'
#502400000000
1!
b111 %
1'
b111 +
#502410000000
0!
0'
#502420000000
1!
b1000 %
1'
b1000 +
#502430000000
0!
0'
#502440000000
1!
b1001 %
1'
b1001 +
#502450000000
1"
1(
#502460000000
0!
0"
b100 &
0'
0(
b100 ,
#502470000000
1!
b0 %
1'
b0 +
#502480000000
0!
0'
#502490000000
1!
1$
b1 %
1'
1*
b1 +
#502500000000
0!
0'
#502510000000
1!
b10 %
1'
b10 +
#502520000000
0!
0'
#502530000000
1!
b11 %
1'
b11 +
#502540000000
0!
0'
#502550000000
1!
b100 %
1'
b100 +
#502560000000
0!
0'
#502570000000
1!
b101 %
1'
b101 +
#502580000000
0!
0'
#502590000000
1!
b110 %
1'
b110 +
#502600000000
0!
0'
#502610000000
1!
b111 %
1'
b111 +
#502620000000
0!
0'
#502630000000
1!
0$
b1000 %
1'
0*
b1000 +
#502640000000
0!
0'
#502650000000
1!
b1001 %
1'
b1001 +
#502660000000
0!
0'
#502670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#502680000000
0!
0'
#502690000000
1!
1$
b1 %
1'
1*
b1 +
#502700000000
0!
0'
#502710000000
1!
b10 %
1'
b10 +
#502720000000
0!
0'
#502730000000
1!
b11 %
1'
b11 +
#502740000000
0!
0'
#502750000000
1!
b100 %
1'
b100 +
#502760000000
0!
0'
#502770000000
1!
b101 %
1'
b101 +
#502780000000
0!
0'
#502790000000
1!
0$
b110 %
1'
0*
b110 +
#502800000000
0!
0'
#502810000000
1!
b111 %
1'
b111 +
#502820000000
0!
0'
#502830000000
1!
b1000 %
1'
b1000 +
#502840000000
0!
0'
#502850000000
1!
b1001 %
1'
b1001 +
#502860000000
0!
0'
#502870000000
1!
b0 %
1'
b0 +
#502880000000
1"
1(
#502890000000
0!
0"
b100 &
0'
0(
b100 ,
#502900000000
1!
1$
b1 %
1'
1*
b1 +
#502910000000
0!
0'
#502920000000
1!
b10 %
1'
b10 +
#502930000000
0!
0'
#502940000000
1!
b11 %
1'
b11 +
#502950000000
0!
0'
#502960000000
1!
b100 %
1'
b100 +
#502970000000
0!
0'
#502980000000
1!
b101 %
1'
b101 +
#502990000000
0!
0'
#503000000000
1!
b110 %
1'
b110 +
#503010000000
0!
0'
#503020000000
1!
b111 %
1'
b111 +
#503030000000
0!
0'
#503040000000
1!
0$
b1000 %
1'
0*
b1000 +
#503050000000
0!
0'
#503060000000
1!
b1001 %
1'
b1001 +
#503070000000
0!
0'
#503080000000
1!
b0 %
1'
b0 +
#503090000000
0!
0'
#503100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#503110000000
0!
0'
#503120000000
1!
b10 %
1'
b10 +
#503130000000
0!
0'
#503140000000
1!
b11 %
1'
b11 +
#503150000000
0!
0'
#503160000000
1!
b100 %
1'
b100 +
#503170000000
0!
0'
#503180000000
1!
b101 %
1'
b101 +
#503190000000
0!
0'
#503200000000
1!
0$
b110 %
1'
0*
b110 +
#503210000000
0!
0'
#503220000000
1!
b111 %
1'
b111 +
#503230000000
0!
0'
#503240000000
1!
b1000 %
1'
b1000 +
#503250000000
0!
0'
#503260000000
1!
b1001 %
1'
b1001 +
#503270000000
0!
0'
#503280000000
1!
b0 %
1'
b0 +
#503290000000
0!
0'
#503300000000
1!
1$
b1 %
1'
1*
b1 +
#503310000000
1"
1(
#503320000000
0!
0"
b100 &
0'
0(
b100 ,
#503330000000
1!
b10 %
1'
b10 +
#503340000000
0!
0'
#503350000000
1!
b11 %
1'
b11 +
#503360000000
0!
0'
#503370000000
1!
b100 %
1'
b100 +
#503380000000
0!
0'
#503390000000
1!
b101 %
1'
b101 +
#503400000000
0!
0'
#503410000000
1!
b110 %
1'
b110 +
#503420000000
0!
0'
#503430000000
1!
b111 %
1'
b111 +
#503440000000
0!
0'
#503450000000
1!
0$
b1000 %
1'
0*
b1000 +
#503460000000
0!
0'
#503470000000
1!
b1001 %
1'
b1001 +
#503480000000
0!
0'
#503490000000
1!
b0 %
1'
b0 +
#503500000000
0!
0'
#503510000000
1!
1$
b1 %
1'
1*
b1 +
#503520000000
0!
0'
#503530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#503540000000
0!
0'
#503550000000
1!
b11 %
1'
b11 +
#503560000000
0!
0'
#503570000000
1!
b100 %
1'
b100 +
#503580000000
0!
0'
#503590000000
1!
b101 %
1'
b101 +
#503600000000
0!
0'
#503610000000
1!
0$
b110 %
1'
0*
b110 +
#503620000000
0!
0'
#503630000000
1!
b111 %
1'
b111 +
#503640000000
0!
0'
#503650000000
1!
b1000 %
1'
b1000 +
#503660000000
0!
0'
#503670000000
1!
b1001 %
1'
b1001 +
#503680000000
0!
0'
#503690000000
1!
b0 %
1'
b0 +
#503700000000
0!
0'
#503710000000
1!
1$
b1 %
1'
1*
b1 +
#503720000000
0!
0'
#503730000000
1!
b10 %
1'
b10 +
#503740000000
1"
1(
#503750000000
0!
0"
b100 &
0'
0(
b100 ,
#503760000000
1!
b11 %
1'
b11 +
#503770000000
0!
0'
#503780000000
1!
b100 %
1'
b100 +
#503790000000
0!
0'
#503800000000
1!
b101 %
1'
b101 +
#503810000000
0!
0'
#503820000000
1!
b110 %
1'
b110 +
#503830000000
0!
0'
#503840000000
1!
b111 %
1'
b111 +
#503850000000
0!
0'
#503860000000
1!
0$
b1000 %
1'
0*
b1000 +
#503870000000
0!
0'
#503880000000
1!
b1001 %
1'
b1001 +
#503890000000
0!
0'
#503900000000
1!
b0 %
1'
b0 +
#503910000000
0!
0'
#503920000000
1!
1$
b1 %
1'
1*
b1 +
#503930000000
0!
0'
#503940000000
1!
b10 %
1'
b10 +
#503950000000
0!
0'
#503960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#503970000000
0!
0'
#503980000000
1!
b100 %
1'
b100 +
#503990000000
0!
0'
#504000000000
1!
b101 %
1'
b101 +
#504010000000
0!
0'
#504020000000
1!
0$
b110 %
1'
0*
b110 +
#504030000000
0!
0'
#504040000000
1!
b111 %
1'
b111 +
#504050000000
0!
0'
#504060000000
1!
b1000 %
1'
b1000 +
#504070000000
0!
0'
#504080000000
1!
b1001 %
1'
b1001 +
#504090000000
0!
0'
#504100000000
1!
b0 %
1'
b0 +
#504110000000
0!
0'
#504120000000
1!
1$
b1 %
1'
1*
b1 +
#504130000000
0!
0'
#504140000000
1!
b10 %
1'
b10 +
#504150000000
0!
0'
#504160000000
1!
b11 %
1'
b11 +
#504170000000
1"
1(
#504180000000
0!
0"
b100 &
0'
0(
b100 ,
#504190000000
1!
b100 %
1'
b100 +
#504200000000
0!
0'
#504210000000
1!
b101 %
1'
b101 +
#504220000000
0!
0'
#504230000000
1!
b110 %
1'
b110 +
#504240000000
0!
0'
#504250000000
1!
b111 %
1'
b111 +
#504260000000
0!
0'
#504270000000
1!
0$
b1000 %
1'
0*
b1000 +
#504280000000
0!
0'
#504290000000
1!
b1001 %
1'
b1001 +
#504300000000
0!
0'
#504310000000
1!
b0 %
1'
b0 +
#504320000000
0!
0'
#504330000000
1!
1$
b1 %
1'
1*
b1 +
#504340000000
0!
0'
#504350000000
1!
b10 %
1'
b10 +
#504360000000
0!
0'
#504370000000
1!
b11 %
1'
b11 +
#504380000000
0!
0'
#504390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#504400000000
0!
0'
#504410000000
1!
b101 %
1'
b101 +
#504420000000
0!
0'
#504430000000
1!
0$
b110 %
1'
0*
b110 +
#504440000000
0!
0'
#504450000000
1!
b111 %
1'
b111 +
#504460000000
0!
0'
#504470000000
1!
b1000 %
1'
b1000 +
#504480000000
0!
0'
#504490000000
1!
b1001 %
1'
b1001 +
#504500000000
0!
0'
#504510000000
1!
b0 %
1'
b0 +
#504520000000
0!
0'
#504530000000
1!
1$
b1 %
1'
1*
b1 +
#504540000000
0!
0'
#504550000000
1!
b10 %
1'
b10 +
#504560000000
0!
0'
#504570000000
1!
b11 %
1'
b11 +
#504580000000
0!
0'
#504590000000
1!
b100 %
1'
b100 +
#504600000000
1"
1(
#504610000000
0!
0"
b100 &
0'
0(
b100 ,
#504620000000
1!
b101 %
1'
b101 +
#504630000000
0!
0'
#504640000000
1!
b110 %
1'
b110 +
#504650000000
0!
0'
#504660000000
1!
b111 %
1'
b111 +
#504670000000
0!
0'
#504680000000
1!
0$
b1000 %
1'
0*
b1000 +
#504690000000
0!
0'
#504700000000
1!
b1001 %
1'
b1001 +
#504710000000
0!
0'
#504720000000
1!
b0 %
1'
b0 +
#504730000000
0!
0'
#504740000000
1!
1$
b1 %
1'
1*
b1 +
#504750000000
0!
0'
#504760000000
1!
b10 %
1'
b10 +
#504770000000
0!
0'
#504780000000
1!
b11 %
1'
b11 +
#504790000000
0!
0'
#504800000000
1!
b100 %
1'
b100 +
#504810000000
0!
0'
#504820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#504830000000
0!
0'
#504840000000
1!
0$
b110 %
1'
0*
b110 +
#504850000000
0!
0'
#504860000000
1!
b111 %
1'
b111 +
#504870000000
0!
0'
#504880000000
1!
b1000 %
1'
b1000 +
#504890000000
0!
0'
#504900000000
1!
b1001 %
1'
b1001 +
#504910000000
0!
0'
#504920000000
1!
b0 %
1'
b0 +
#504930000000
0!
0'
#504940000000
1!
1$
b1 %
1'
1*
b1 +
#504950000000
0!
0'
#504960000000
1!
b10 %
1'
b10 +
#504970000000
0!
0'
#504980000000
1!
b11 %
1'
b11 +
#504990000000
0!
0'
#505000000000
1!
b100 %
1'
b100 +
#505010000000
0!
0'
#505020000000
1!
b101 %
1'
b101 +
#505030000000
1"
1(
#505040000000
0!
0"
b100 &
0'
0(
b100 ,
#505050000000
1!
b110 %
1'
b110 +
#505060000000
0!
0'
#505070000000
1!
b111 %
1'
b111 +
#505080000000
0!
0'
#505090000000
1!
0$
b1000 %
1'
0*
b1000 +
#505100000000
0!
0'
#505110000000
1!
b1001 %
1'
b1001 +
#505120000000
0!
0'
#505130000000
1!
b0 %
1'
b0 +
#505140000000
0!
0'
#505150000000
1!
1$
b1 %
1'
1*
b1 +
#505160000000
0!
0'
#505170000000
1!
b10 %
1'
b10 +
#505180000000
0!
0'
#505190000000
1!
b11 %
1'
b11 +
#505200000000
0!
0'
#505210000000
1!
b100 %
1'
b100 +
#505220000000
0!
0'
#505230000000
1!
b101 %
1'
b101 +
#505240000000
0!
0'
#505250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#505260000000
0!
0'
#505270000000
1!
b111 %
1'
b111 +
#505280000000
0!
0'
#505290000000
1!
b1000 %
1'
b1000 +
#505300000000
0!
0'
#505310000000
1!
b1001 %
1'
b1001 +
#505320000000
0!
0'
#505330000000
1!
b0 %
1'
b0 +
#505340000000
0!
0'
#505350000000
1!
1$
b1 %
1'
1*
b1 +
#505360000000
0!
0'
#505370000000
1!
b10 %
1'
b10 +
#505380000000
0!
0'
#505390000000
1!
b11 %
1'
b11 +
#505400000000
0!
0'
#505410000000
1!
b100 %
1'
b100 +
#505420000000
0!
0'
#505430000000
1!
b101 %
1'
b101 +
#505440000000
0!
0'
#505450000000
1!
0$
b110 %
1'
0*
b110 +
#505460000000
1"
1(
#505470000000
0!
0"
b100 &
0'
0(
b100 ,
#505480000000
1!
1$
b111 %
1'
1*
b111 +
#505490000000
0!
0'
#505500000000
1!
0$
b1000 %
1'
0*
b1000 +
#505510000000
0!
0'
#505520000000
1!
b1001 %
1'
b1001 +
#505530000000
0!
0'
#505540000000
1!
b0 %
1'
b0 +
#505550000000
0!
0'
#505560000000
1!
1$
b1 %
1'
1*
b1 +
#505570000000
0!
0'
#505580000000
1!
b10 %
1'
b10 +
#505590000000
0!
0'
#505600000000
1!
b11 %
1'
b11 +
#505610000000
0!
0'
#505620000000
1!
b100 %
1'
b100 +
#505630000000
0!
0'
#505640000000
1!
b101 %
1'
b101 +
#505650000000
0!
0'
#505660000000
1!
b110 %
1'
b110 +
#505670000000
0!
0'
#505680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#505690000000
0!
0'
#505700000000
1!
b1000 %
1'
b1000 +
#505710000000
0!
0'
#505720000000
1!
b1001 %
1'
b1001 +
#505730000000
0!
0'
#505740000000
1!
b0 %
1'
b0 +
#505750000000
0!
0'
#505760000000
1!
1$
b1 %
1'
1*
b1 +
#505770000000
0!
0'
#505780000000
1!
b10 %
1'
b10 +
#505790000000
0!
0'
#505800000000
1!
b11 %
1'
b11 +
#505810000000
0!
0'
#505820000000
1!
b100 %
1'
b100 +
#505830000000
0!
0'
#505840000000
1!
b101 %
1'
b101 +
#505850000000
0!
0'
#505860000000
1!
0$
b110 %
1'
0*
b110 +
#505870000000
0!
0'
#505880000000
1!
b111 %
1'
b111 +
#505890000000
1"
1(
#505900000000
0!
0"
b100 &
0'
0(
b100 ,
#505910000000
1!
b1000 %
1'
b1000 +
#505920000000
0!
0'
#505930000000
1!
b1001 %
1'
b1001 +
#505940000000
0!
0'
#505950000000
1!
b0 %
1'
b0 +
#505960000000
0!
0'
#505970000000
1!
1$
b1 %
1'
1*
b1 +
#505980000000
0!
0'
#505990000000
1!
b10 %
1'
b10 +
#506000000000
0!
0'
#506010000000
1!
b11 %
1'
b11 +
#506020000000
0!
0'
#506030000000
1!
b100 %
1'
b100 +
#506040000000
0!
0'
#506050000000
1!
b101 %
1'
b101 +
#506060000000
0!
0'
#506070000000
1!
b110 %
1'
b110 +
#506080000000
0!
0'
#506090000000
1!
b111 %
1'
b111 +
#506100000000
0!
0'
#506110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#506120000000
0!
0'
#506130000000
1!
b1001 %
1'
b1001 +
#506140000000
0!
0'
#506150000000
1!
b0 %
1'
b0 +
#506160000000
0!
0'
#506170000000
1!
1$
b1 %
1'
1*
b1 +
#506180000000
0!
0'
#506190000000
1!
b10 %
1'
b10 +
#506200000000
0!
0'
#506210000000
1!
b11 %
1'
b11 +
#506220000000
0!
0'
#506230000000
1!
b100 %
1'
b100 +
#506240000000
0!
0'
#506250000000
1!
b101 %
1'
b101 +
#506260000000
0!
0'
#506270000000
1!
0$
b110 %
1'
0*
b110 +
#506280000000
0!
0'
#506290000000
1!
b111 %
1'
b111 +
#506300000000
0!
0'
#506310000000
1!
b1000 %
1'
b1000 +
#506320000000
1"
1(
#506330000000
0!
0"
b100 &
0'
0(
b100 ,
#506340000000
1!
b1001 %
1'
b1001 +
#506350000000
0!
0'
#506360000000
1!
b0 %
1'
b0 +
#506370000000
0!
0'
#506380000000
1!
1$
b1 %
1'
1*
b1 +
#506390000000
0!
0'
#506400000000
1!
b10 %
1'
b10 +
#506410000000
0!
0'
#506420000000
1!
b11 %
1'
b11 +
#506430000000
0!
0'
#506440000000
1!
b100 %
1'
b100 +
#506450000000
0!
0'
#506460000000
1!
b101 %
1'
b101 +
#506470000000
0!
0'
#506480000000
1!
b110 %
1'
b110 +
#506490000000
0!
0'
#506500000000
1!
b111 %
1'
b111 +
#506510000000
0!
0'
#506520000000
1!
0$
b1000 %
1'
0*
b1000 +
#506530000000
0!
0'
#506540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#506550000000
0!
0'
#506560000000
1!
b0 %
1'
b0 +
#506570000000
0!
0'
#506580000000
1!
1$
b1 %
1'
1*
b1 +
#506590000000
0!
0'
#506600000000
1!
b10 %
1'
b10 +
#506610000000
0!
0'
#506620000000
1!
b11 %
1'
b11 +
#506630000000
0!
0'
#506640000000
1!
b100 %
1'
b100 +
#506650000000
0!
0'
#506660000000
1!
b101 %
1'
b101 +
#506670000000
0!
0'
#506680000000
1!
0$
b110 %
1'
0*
b110 +
#506690000000
0!
0'
#506700000000
1!
b111 %
1'
b111 +
#506710000000
0!
0'
#506720000000
1!
b1000 %
1'
b1000 +
#506730000000
0!
0'
#506740000000
1!
b1001 %
1'
b1001 +
#506750000000
1"
1(
#506760000000
0!
0"
b100 &
0'
0(
b100 ,
#506770000000
1!
b0 %
1'
b0 +
#506780000000
0!
0'
#506790000000
1!
1$
b1 %
1'
1*
b1 +
#506800000000
0!
0'
#506810000000
1!
b10 %
1'
b10 +
#506820000000
0!
0'
#506830000000
1!
b11 %
1'
b11 +
#506840000000
0!
0'
#506850000000
1!
b100 %
1'
b100 +
#506860000000
0!
0'
#506870000000
1!
b101 %
1'
b101 +
#506880000000
0!
0'
#506890000000
1!
b110 %
1'
b110 +
#506900000000
0!
0'
#506910000000
1!
b111 %
1'
b111 +
#506920000000
0!
0'
#506930000000
1!
0$
b1000 %
1'
0*
b1000 +
#506940000000
0!
0'
#506950000000
1!
b1001 %
1'
b1001 +
#506960000000
0!
0'
#506970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#506980000000
0!
0'
#506990000000
1!
1$
b1 %
1'
1*
b1 +
#507000000000
0!
0'
#507010000000
1!
b10 %
1'
b10 +
#507020000000
0!
0'
#507030000000
1!
b11 %
1'
b11 +
#507040000000
0!
0'
#507050000000
1!
b100 %
1'
b100 +
#507060000000
0!
0'
#507070000000
1!
b101 %
1'
b101 +
#507080000000
0!
0'
#507090000000
1!
0$
b110 %
1'
0*
b110 +
#507100000000
0!
0'
#507110000000
1!
b111 %
1'
b111 +
#507120000000
0!
0'
#507130000000
1!
b1000 %
1'
b1000 +
#507140000000
0!
0'
#507150000000
1!
b1001 %
1'
b1001 +
#507160000000
0!
0'
#507170000000
1!
b0 %
1'
b0 +
#507180000000
1"
1(
#507190000000
0!
0"
b100 &
0'
0(
b100 ,
#507200000000
1!
1$
b1 %
1'
1*
b1 +
#507210000000
0!
0'
#507220000000
1!
b10 %
1'
b10 +
#507230000000
0!
0'
#507240000000
1!
b11 %
1'
b11 +
#507250000000
0!
0'
#507260000000
1!
b100 %
1'
b100 +
#507270000000
0!
0'
#507280000000
1!
b101 %
1'
b101 +
#507290000000
0!
0'
#507300000000
1!
b110 %
1'
b110 +
#507310000000
0!
0'
#507320000000
1!
b111 %
1'
b111 +
#507330000000
0!
0'
#507340000000
1!
0$
b1000 %
1'
0*
b1000 +
#507350000000
0!
0'
#507360000000
1!
b1001 %
1'
b1001 +
#507370000000
0!
0'
#507380000000
1!
b0 %
1'
b0 +
#507390000000
0!
0'
#507400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#507410000000
0!
0'
#507420000000
1!
b10 %
1'
b10 +
#507430000000
0!
0'
#507440000000
1!
b11 %
1'
b11 +
#507450000000
0!
0'
#507460000000
1!
b100 %
1'
b100 +
#507470000000
0!
0'
#507480000000
1!
b101 %
1'
b101 +
#507490000000
0!
0'
#507500000000
1!
0$
b110 %
1'
0*
b110 +
#507510000000
0!
0'
#507520000000
1!
b111 %
1'
b111 +
#507530000000
0!
0'
#507540000000
1!
b1000 %
1'
b1000 +
#507550000000
0!
0'
#507560000000
1!
b1001 %
1'
b1001 +
#507570000000
0!
0'
#507580000000
1!
b0 %
1'
b0 +
#507590000000
0!
0'
#507600000000
1!
1$
b1 %
1'
1*
b1 +
#507610000000
1"
1(
#507620000000
0!
0"
b100 &
0'
0(
b100 ,
#507630000000
1!
b10 %
1'
b10 +
#507640000000
0!
0'
#507650000000
1!
b11 %
1'
b11 +
#507660000000
0!
0'
#507670000000
1!
b100 %
1'
b100 +
#507680000000
0!
0'
#507690000000
1!
b101 %
1'
b101 +
#507700000000
0!
0'
#507710000000
1!
b110 %
1'
b110 +
#507720000000
0!
0'
#507730000000
1!
b111 %
1'
b111 +
#507740000000
0!
0'
#507750000000
1!
0$
b1000 %
1'
0*
b1000 +
#507760000000
0!
0'
#507770000000
1!
b1001 %
1'
b1001 +
#507780000000
0!
0'
#507790000000
1!
b0 %
1'
b0 +
#507800000000
0!
0'
#507810000000
1!
1$
b1 %
1'
1*
b1 +
#507820000000
0!
0'
#507830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#507840000000
0!
0'
#507850000000
1!
b11 %
1'
b11 +
#507860000000
0!
0'
#507870000000
1!
b100 %
1'
b100 +
#507880000000
0!
0'
#507890000000
1!
b101 %
1'
b101 +
#507900000000
0!
0'
#507910000000
1!
0$
b110 %
1'
0*
b110 +
#507920000000
0!
0'
#507930000000
1!
b111 %
1'
b111 +
#507940000000
0!
0'
#507950000000
1!
b1000 %
1'
b1000 +
#507960000000
0!
0'
#507970000000
1!
b1001 %
1'
b1001 +
#507980000000
0!
0'
#507990000000
1!
b0 %
1'
b0 +
#508000000000
0!
0'
#508010000000
1!
1$
b1 %
1'
1*
b1 +
#508020000000
0!
0'
#508030000000
1!
b10 %
1'
b10 +
#508040000000
1"
1(
#508050000000
0!
0"
b100 &
0'
0(
b100 ,
#508060000000
1!
b11 %
1'
b11 +
#508070000000
0!
0'
#508080000000
1!
b100 %
1'
b100 +
#508090000000
0!
0'
#508100000000
1!
b101 %
1'
b101 +
#508110000000
0!
0'
#508120000000
1!
b110 %
1'
b110 +
#508130000000
0!
0'
#508140000000
1!
b111 %
1'
b111 +
#508150000000
0!
0'
#508160000000
1!
0$
b1000 %
1'
0*
b1000 +
#508170000000
0!
0'
#508180000000
1!
b1001 %
1'
b1001 +
#508190000000
0!
0'
#508200000000
1!
b0 %
1'
b0 +
#508210000000
0!
0'
#508220000000
1!
1$
b1 %
1'
1*
b1 +
#508230000000
0!
0'
#508240000000
1!
b10 %
1'
b10 +
#508250000000
0!
0'
#508260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#508270000000
0!
0'
#508280000000
1!
b100 %
1'
b100 +
#508290000000
0!
0'
#508300000000
1!
b101 %
1'
b101 +
#508310000000
0!
0'
#508320000000
1!
0$
b110 %
1'
0*
b110 +
#508330000000
0!
0'
#508340000000
1!
b111 %
1'
b111 +
#508350000000
0!
0'
#508360000000
1!
b1000 %
1'
b1000 +
#508370000000
0!
0'
#508380000000
1!
b1001 %
1'
b1001 +
#508390000000
0!
0'
#508400000000
1!
b0 %
1'
b0 +
#508410000000
0!
0'
#508420000000
1!
1$
b1 %
1'
1*
b1 +
#508430000000
0!
0'
#508440000000
1!
b10 %
1'
b10 +
#508450000000
0!
0'
#508460000000
1!
b11 %
1'
b11 +
#508470000000
1"
1(
#508480000000
0!
0"
b100 &
0'
0(
b100 ,
#508490000000
1!
b100 %
1'
b100 +
#508500000000
0!
0'
#508510000000
1!
b101 %
1'
b101 +
#508520000000
0!
0'
#508530000000
1!
b110 %
1'
b110 +
#508540000000
0!
0'
#508550000000
1!
b111 %
1'
b111 +
#508560000000
0!
0'
#508570000000
1!
0$
b1000 %
1'
0*
b1000 +
#508580000000
0!
0'
#508590000000
1!
b1001 %
1'
b1001 +
#508600000000
0!
0'
#508610000000
1!
b0 %
1'
b0 +
#508620000000
0!
0'
#508630000000
1!
1$
b1 %
1'
1*
b1 +
#508640000000
0!
0'
#508650000000
1!
b10 %
1'
b10 +
#508660000000
0!
0'
#508670000000
1!
b11 %
1'
b11 +
#508680000000
0!
0'
#508690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#508700000000
0!
0'
#508710000000
1!
b101 %
1'
b101 +
#508720000000
0!
0'
#508730000000
1!
0$
b110 %
1'
0*
b110 +
#508740000000
0!
0'
#508750000000
1!
b111 %
1'
b111 +
#508760000000
0!
0'
#508770000000
1!
b1000 %
1'
b1000 +
#508780000000
0!
0'
#508790000000
1!
b1001 %
1'
b1001 +
#508800000000
0!
0'
#508810000000
1!
b0 %
1'
b0 +
#508820000000
0!
0'
#508830000000
1!
1$
b1 %
1'
1*
b1 +
#508840000000
0!
0'
#508850000000
1!
b10 %
1'
b10 +
#508860000000
0!
0'
#508870000000
1!
b11 %
1'
b11 +
#508880000000
0!
0'
#508890000000
1!
b100 %
1'
b100 +
#508900000000
1"
1(
#508910000000
0!
0"
b100 &
0'
0(
b100 ,
#508920000000
1!
b101 %
1'
b101 +
#508930000000
0!
0'
#508940000000
1!
b110 %
1'
b110 +
#508950000000
0!
0'
#508960000000
1!
b111 %
1'
b111 +
#508970000000
0!
0'
#508980000000
1!
0$
b1000 %
1'
0*
b1000 +
#508990000000
0!
0'
#509000000000
1!
b1001 %
1'
b1001 +
#509010000000
0!
0'
#509020000000
1!
b0 %
1'
b0 +
#509030000000
0!
0'
#509040000000
1!
1$
b1 %
1'
1*
b1 +
#509050000000
0!
0'
#509060000000
1!
b10 %
1'
b10 +
#509070000000
0!
0'
#509080000000
1!
b11 %
1'
b11 +
#509090000000
0!
0'
#509100000000
1!
b100 %
1'
b100 +
#509110000000
0!
0'
#509120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#509130000000
0!
0'
#509140000000
1!
0$
b110 %
1'
0*
b110 +
#509150000000
0!
0'
#509160000000
1!
b111 %
1'
b111 +
#509170000000
0!
0'
#509180000000
1!
b1000 %
1'
b1000 +
#509190000000
0!
0'
#509200000000
1!
b1001 %
1'
b1001 +
#509210000000
0!
0'
#509220000000
1!
b0 %
1'
b0 +
#509230000000
0!
0'
#509240000000
1!
1$
b1 %
1'
1*
b1 +
#509250000000
0!
0'
#509260000000
1!
b10 %
1'
b10 +
#509270000000
0!
0'
#509280000000
1!
b11 %
1'
b11 +
#509290000000
0!
0'
#509300000000
1!
b100 %
1'
b100 +
#509310000000
0!
0'
#509320000000
1!
b101 %
1'
b101 +
#509330000000
1"
1(
#509340000000
0!
0"
b100 &
0'
0(
b100 ,
#509350000000
1!
b110 %
1'
b110 +
#509360000000
0!
0'
#509370000000
1!
b111 %
1'
b111 +
#509380000000
0!
0'
#509390000000
1!
0$
b1000 %
1'
0*
b1000 +
#509400000000
0!
0'
#509410000000
1!
b1001 %
1'
b1001 +
#509420000000
0!
0'
#509430000000
1!
b0 %
1'
b0 +
#509440000000
0!
0'
#509450000000
1!
1$
b1 %
1'
1*
b1 +
#509460000000
0!
0'
#509470000000
1!
b10 %
1'
b10 +
#509480000000
0!
0'
#509490000000
1!
b11 %
1'
b11 +
#509500000000
0!
0'
#509510000000
1!
b100 %
1'
b100 +
#509520000000
0!
0'
#509530000000
1!
b101 %
1'
b101 +
#509540000000
0!
0'
#509550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#509560000000
0!
0'
#509570000000
1!
b111 %
1'
b111 +
#509580000000
0!
0'
#509590000000
1!
b1000 %
1'
b1000 +
#509600000000
0!
0'
#509610000000
1!
b1001 %
1'
b1001 +
#509620000000
0!
0'
#509630000000
1!
b0 %
1'
b0 +
#509640000000
0!
0'
#509650000000
1!
1$
b1 %
1'
1*
b1 +
#509660000000
0!
0'
#509670000000
1!
b10 %
1'
b10 +
#509680000000
0!
0'
#509690000000
1!
b11 %
1'
b11 +
#509700000000
0!
0'
#509710000000
1!
b100 %
1'
b100 +
#509720000000
0!
0'
#509730000000
1!
b101 %
1'
b101 +
#509740000000
0!
0'
#509750000000
1!
0$
b110 %
1'
0*
b110 +
#509760000000
1"
1(
#509770000000
0!
0"
b100 &
0'
0(
b100 ,
#509780000000
1!
1$
b111 %
1'
1*
b111 +
#509790000000
0!
0'
#509800000000
1!
0$
b1000 %
1'
0*
b1000 +
#509810000000
0!
0'
#509820000000
1!
b1001 %
1'
b1001 +
#509830000000
0!
0'
#509840000000
1!
b0 %
1'
b0 +
#509850000000
0!
0'
#509860000000
1!
1$
b1 %
1'
1*
b1 +
#509870000000
0!
0'
#509880000000
1!
b10 %
1'
b10 +
#509890000000
0!
0'
#509900000000
1!
b11 %
1'
b11 +
#509910000000
0!
0'
#509920000000
1!
b100 %
1'
b100 +
#509930000000
0!
0'
#509940000000
1!
b101 %
1'
b101 +
#509950000000
0!
0'
#509960000000
1!
b110 %
1'
b110 +
#509970000000
0!
0'
#509980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#509990000000
0!
0'
#510000000000
1!
b1000 %
1'
b1000 +
#510010000000
0!
0'
#510020000000
1!
b1001 %
1'
b1001 +
#510030000000
0!
0'
#510040000000
1!
b0 %
1'
b0 +
#510050000000
0!
0'
#510060000000
1!
1$
b1 %
1'
1*
b1 +
#510070000000
0!
0'
#510080000000
1!
b10 %
1'
b10 +
#510090000000
0!
0'
#510100000000
1!
b11 %
1'
b11 +
#510110000000
0!
0'
#510120000000
1!
b100 %
1'
b100 +
#510130000000
0!
0'
#510140000000
1!
b101 %
1'
b101 +
#510150000000
0!
0'
#510160000000
1!
0$
b110 %
1'
0*
b110 +
#510170000000
0!
0'
#510180000000
1!
b111 %
1'
b111 +
#510190000000
1"
1(
#510200000000
0!
0"
b100 &
0'
0(
b100 ,
#510210000000
1!
b1000 %
1'
b1000 +
#510220000000
0!
0'
#510230000000
1!
b1001 %
1'
b1001 +
#510240000000
0!
0'
#510250000000
1!
b0 %
1'
b0 +
#510260000000
0!
0'
#510270000000
1!
1$
b1 %
1'
1*
b1 +
#510280000000
0!
0'
#510290000000
1!
b10 %
1'
b10 +
#510300000000
0!
0'
#510310000000
1!
b11 %
1'
b11 +
#510320000000
0!
0'
#510330000000
1!
b100 %
1'
b100 +
#510340000000
0!
0'
#510350000000
1!
b101 %
1'
b101 +
#510360000000
0!
0'
#510370000000
1!
b110 %
1'
b110 +
#510380000000
0!
0'
#510390000000
1!
b111 %
1'
b111 +
#510400000000
0!
0'
#510410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#510420000000
0!
0'
#510430000000
1!
b1001 %
1'
b1001 +
#510440000000
0!
0'
#510450000000
1!
b0 %
1'
b0 +
#510460000000
0!
0'
#510470000000
1!
1$
b1 %
1'
1*
b1 +
#510480000000
0!
0'
#510490000000
1!
b10 %
1'
b10 +
#510500000000
0!
0'
#510510000000
1!
b11 %
1'
b11 +
#510520000000
0!
0'
#510530000000
1!
b100 %
1'
b100 +
#510540000000
0!
0'
#510550000000
1!
b101 %
1'
b101 +
#510560000000
0!
0'
#510570000000
1!
0$
b110 %
1'
0*
b110 +
#510580000000
0!
0'
#510590000000
1!
b111 %
1'
b111 +
#510600000000
0!
0'
#510610000000
1!
b1000 %
1'
b1000 +
#510620000000
1"
1(
#510630000000
0!
0"
b100 &
0'
0(
b100 ,
#510640000000
1!
b1001 %
1'
b1001 +
#510650000000
0!
0'
#510660000000
1!
b0 %
1'
b0 +
#510670000000
0!
0'
#510680000000
1!
1$
b1 %
1'
1*
b1 +
#510690000000
0!
0'
#510700000000
1!
b10 %
1'
b10 +
#510710000000
0!
0'
#510720000000
1!
b11 %
1'
b11 +
#510730000000
0!
0'
#510740000000
1!
b100 %
1'
b100 +
#510750000000
0!
0'
#510760000000
1!
b101 %
1'
b101 +
#510770000000
0!
0'
#510780000000
1!
b110 %
1'
b110 +
#510790000000
0!
0'
#510800000000
1!
b111 %
1'
b111 +
#510810000000
0!
0'
#510820000000
1!
0$
b1000 %
1'
0*
b1000 +
#510830000000
0!
0'
#510840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#510850000000
0!
0'
#510860000000
1!
b0 %
1'
b0 +
#510870000000
0!
0'
#510880000000
1!
1$
b1 %
1'
1*
b1 +
#510890000000
0!
0'
#510900000000
1!
b10 %
1'
b10 +
#510910000000
0!
0'
#510920000000
1!
b11 %
1'
b11 +
#510930000000
0!
0'
#510940000000
1!
b100 %
1'
b100 +
#510950000000
0!
0'
#510960000000
1!
b101 %
1'
b101 +
#510970000000
0!
0'
#510980000000
1!
0$
b110 %
1'
0*
b110 +
#510990000000
0!
0'
#511000000000
1!
b111 %
1'
b111 +
#511010000000
0!
0'
#511020000000
1!
b1000 %
1'
b1000 +
#511030000000
0!
0'
#511040000000
1!
b1001 %
1'
b1001 +
#511050000000
1"
1(
#511060000000
0!
0"
b100 &
0'
0(
b100 ,
#511070000000
1!
b0 %
1'
b0 +
#511080000000
0!
0'
#511090000000
1!
1$
b1 %
1'
1*
b1 +
#511100000000
0!
0'
#511110000000
1!
b10 %
1'
b10 +
#511120000000
0!
0'
#511130000000
1!
b11 %
1'
b11 +
#511140000000
0!
0'
#511150000000
1!
b100 %
1'
b100 +
#511160000000
0!
0'
#511170000000
1!
b101 %
1'
b101 +
#511180000000
0!
0'
#511190000000
1!
b110 %
1'
b110 +
#511200000000
0!
0'
#511210000000
1!
b111 %
1'
b111 +
#511220000000
0!
0'
#511230000000
1!
0$
b1000 %
1'
0*
b1000 +
#511240000000
0!
0'
#511250000000
1!
b1001 %
1'
b1001 +
#511260000000
0!
0'
#511270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#511280000000
0!
0'
#511290000000
1!
1$
b1 %
1'
1*
b1 +
#511300000000
0!
0'
#511310000000
1!
b10 %
1'
b10 +
#511320000000
0!
0'
#511330000000
1!
b11 %
1'
b11 +
#511340000000
0!
0'
#511350000000
1!
b100 %
1'
b100 +
#511360000000
0!
0'
#511370000000
1!
b101 %
1'
b101 +
#511380000000
0!
0'
#511390000000
1!
0$
b110 %
1'
0*
b110 +
#511400000000
0!
0'
#511410000000
1!
b111 %
1'
b111 +
#511420000000
0!
0'
#511430000000
1!
b1000 %
1'
b1000 +
#511440000000
0!
0'
#511450000000
1!
b1001 %
1'
b1001 +
#511460000000
0!
0'
#511470000000
1!
b0 %
1'
b0 +
#511480000000
1"
1(
#511490000000
0!
0"
b100 &
0'
0(
b100 ,
#511500000000
1!
1$
b1 %
1'
1*
b1 +
#511510000000
0!
0'
#511520000000
1!
b10 %
1'
b10 +
#511530000000
0!
0'
#511540000000
1!
b11 %
1'
b11 +
#511550000000
0!
0'
#511560000000
1!
b100 %
1'
b100 +
#511570000000
0!
0'
#511580000000
1!
b101 %
1'
b101 +
#511590000000
0!
0'
#511600000000
1!
b110 %
1'
b110 +
#511610000000
0!
0'
#511620000000
1!
b111 %
1'
b111 +
#511630000000
0!
0'
#511640000000
1!
0$
b1000 %
1'
0*
b1000 +
#511650000000
0!
0'
#511660000000
1!
b1001 %
1'
b1001 +
#511670000000
0!
0'
#511680000000
1!
b0 %
1'
b0 +
#511690000000
0!
0'
#511700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#511710000000
0!
0'
#511720000000
1!
b10 %
1'
b10 +
#511730000000
0!
0'
#511740000000
1!
b11 %
1'
b11 +
#511750000000
0!
0'
#511760000000
1!
b100 %
1'
b100 +
#511770000000
0!
0'
#511780000000
1!
b101 %
1'
b101 +
#511790000000
0!
0'
#511800000000
1!
0$
b110 %
1'
0*
b110 +
#511810000000
0!
0'
#511820000000
1!
b111 %
1'
b111 +
#511830000000
0!
0'
#511840000000
1!
b1000 %
1'
b1000 +
#511850000000
0!
0'
#511860000000
1!
b1001 %
1'
b1001 +
#511870000000
0!
0'
#511880000000
1!
b0 %
1'
b0 +
#511890000000
0!
0'
#511900000000
1!
1$
b1 %
1'
1*
b1 +
#511910000000
1"
1(
#511920000000
0!
0"
b100 &
0'
0(
b100 ,
#511930000000
1!
b10 %
1'
b10 +
#511940000000
0!
0'
#511950000000
1!
b11 %
1'
b11 +
#511960000000
0!
0'
#511970000000
1!
b100 %
1'
b100 +
#511980000000
0!
0'
#511990000000
1!
b101 %
1'
b101 +
#512000000000
0!
0'
#512010000000
1!
b110 %
1'
b110 +
#512020000000
0!
0'
#512030000000
1!
b111 %
1'
b111 +
#512040000000
0!
0'
#512050000000
1!
0$
b1000 %
1'
0*
b1000 +
#512060000000
0!
0'
#512070000000
1!
b1001 %
1'
b1001 +
#512080000000
0!
0'
#512090000000
1!
b0 %
1'
b0 +
#512100000000
0!
0'
#512110000000
1!
1$
b1 %
1'
1*
b1 +
#512120000000
0!
0'
#512130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#512140000000
0!
0'
#512150000000
1!
b11 %
1'
b11 +
#512160000000
0!
0'
#512170000000
1!
b100 %
1'
b100 +
#512180000000
0!
0'
#512190000000
1!
b101 %
1'
b101 +
#512200000000
0!
0'
#512210000000
1!
0$
b110 %
1'
0*
b110 +
#512220000000
0!
0'
#512230000000
1!
b111 %
1'
b111 +
#512240000000
0!
0'
#512250000000
1!
b1000 %
1'
b1000 +
#512260000000
0!
0'
#512270000000
1!
b1001 %
1'
b1001 +
#512280000000
0!
0'
#512290000000
1!
b0 %
1'
b0 +
#512300000000
0!
0'
#512310000000
1!
1$
b1 %
1'
1*
b1 +
#512320000000
0!
0'
#512330000000
1!
b10 %
1'
b10 +
#512340000000
1"
1(
#512350000000
0!
0"
b100 &
0'
0(
b100 ,
#512360000000
1!
b11 %
1'
b11 +
#512370000000
0!
0'
#512380000000
1!
b100 %
1'
b100 +
#512390000000
0!
0'
#512400000000
1!
b101 %
1'
b101 +
#512410000000
0!
0'
#512420000000
1!
b110 %
1'
b110 +
#512430000000
0!
0'
#512440000000
1!
b111 %
1'
b111 +
#512450000000
0!
0'
#512460000000
1!
0$
b1000 %
1'
0*
b1000 +
#512470000000
0!
0'
#512480000000
1!
b1001 %
1'
b1001 +
#512490000000
0!
0'
#512500000000
1!
b0 %
1'
b0 +
#512510000000
0!
0'
#512520000000
1!
1$
b1 %
1'
1*
b1 +
#512530000000
0!
0'
#512540000000
1!
b10 %
1'
b10 +
#512550000000
0!
0'
#512560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#512570000000
0!
0'
#512580000000
1!
b100 %
1'
b100 +
#512590000000
0!
0'
#512600000000
1!
b101 %
1'
b101 +
#512610000000
0!
0'
#512620000000
1!
0$
b110 %
1'
0*
b110 +
#512630000000
0!
0'
#512640000000
1!
b111 %
1'
b111 +
#512650000000
0!
0'
#512660000000
1!
b1000 %
1'
b1000 +
#512670000000
0!
0'
#512680000000
1!
b1001 %
1'
b1001 +
#512690000000
0!
0'
#512700000000
1!
b0 %
1'
b0 +
#512710000000
0!
0'
#512720000000
1!
1$
b1 %
1'
1*
b1 +
#512730000000
0!
0'
#512740000000
1!
b10 %
1'
b10 +
#512750000000
0!
0'
#512760000000
1!
b11 %
1'
b11 +
#512770000000
1"
1(
#512780000000
0!
0"
b100 &
0'
0(
b100 ,
#512790000000
1!
b100 %
1'
b100 +
#512800000000
0!
0'
#512810000000
1!
b101 %
1'
b101 +
#512820000000
0!
0'
#512830000000
1!
b110 %
1'
b110 +
#512840000000
0!
0'
#512850000000
1!
b111 %
1'
b111 +
#512860000000
0!
0'
#512870000000
1!
0$
b1000 %
1'
0*
b1000 +
#512880000000
0!
0'
#512890000000
1!
b1001 %
1'
b1001 +
#512900000000
0!
0'
#512910000000
1!
b0 %
1'
b0 +
#512920000000
0!
0'
#512930000000
1!
1$
b1 %
1'
1*
b1 +
#512940000000
0!
0'
#512950000000
1!
b10 %
1'
b10 +
#512960000000
0!
0'
#512970000000
1!
b11 %
1'
b11 +
#512980000000
0!
0'
#512990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#513000000000
0!
0'
#513010000000
1!
b101 %
1'
b101 +
#513020000000
0!
0'
#513030000000
1!
0$
b110 %
1'
0*
b110 +
#513040000000
0!
0'
#513050000000
1!
b111 %
1'
b111 +
#513060000000
0!
0'
#513070000000
1!
b1000 %
1'
b1000 +
#513080000000
0!
0'
#513090000000
1!
b1001 %
1'
b1001 +
#513100000000
0!
0'
#513110000000
1!
b0 %
1'
b0 +
#513120000000
0!
0'
#513130000000
1!
1$
b1 %
1'
1*
b1 +
#513140000000
0!
0'
#513150000000
1!
b10 %
1'
b10 +
#513160000000
0!
0'
#513170000000
1!
b11 %
1'
b11 +
#513180000000
0!
0'
#513190000000
1!
b100 %
1'
b100 +
#513200000000
1"
1(
#513210000000
0!
0"
b100 &
0'
0(
b100 ,
#513220000000
1!
b101 %
1'
b101 +
#513230000000
0!
0'
#513240000000
1!
b110 %
1'
b110 +
#513250000000
0!
0'
#513260000000
1!
b111 %
1'
b111 +
#513270000000
0!
0'
#513280000000
1!
0$
b1000 %
1'
0*
b1000 +
#513290000000
0!
0'
#513300000000
1!
b1001 %
1'
b1001 +
#513310000000
0!
0'
#513320000000
1!
b0 %
1'
b0 +
#513330000000
0!
0'
#513340000000
1!
1$
b1 %
1'
1*
b1 +
#513350000000
0!
0'
#513360000000
1!
b10 %
1'
b10 +
#513370000000
0!
0'
#513380000000
1!
b11 %
1'
b11 +
#513390000000
0!
0'
#513400000000
1!
b100 %
1'
b100 +
#513410000000
0!
0'
#513420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#513430000000
0!
0'
#513440000000
1!
0$
b110 %
1'
0*
b110 +
#513450000000
0!
0'
#513460000000
1!
b111 %
1'
b111 +
#513470000000
0!
0'
#513480000000
1!
b1000 %
1'
b1000 +
#513490000000
0!
0'
#513500000000
1!
b1001 %
1'
b1001 +
#513510000000
0!
0'
#513520000000
1!
b0 %
1'
b0 +
#513530000000
0!
0'
#513540000000
1!
1$
b1 %
1'
1*
b1 +
#513550000000
0!
0'
#513560000000
1!
b10 %
1'
b10 +
#513570000000
0!
0'
#513580000000
1!
b11 %
1'
b11 +
#513590000000
0!
0'
#513600000000
1!
b100 %
1'
b100 +
#513610000000
0!
0'
#513620000000
1!
b101 %
1'
b101 +
#513630000000
1"
1(
#513640000000
0!
0"
b100 &
0'
0(
b100 ,
#513650000000
1!
b110 %
1'
b110 +
#513660000000
0!
0'
#513670000000
1!
b111 %
1'
b111 +
#513680000000
0!
0'
#513690000000
1!
0$
b1000 %
1'
0*
b1000 +
#513700000000
0!
0'
#513710000000
1!
b1001 %
1'
b1001 +
#513720000000
0!
0'
#513730000000
1!
b0 %
1'
b0 +
#513740000000
0!
0'
#513750000000
1!
1$
b1 %
1'
1*
b1 +
#513760000000
0!
0'
#513770000000
1!
b10 %
1'
b10 +
#513780000000
0!
0'
#513790000000
1!
b11 %
1'
b11 +
#513800000000
0!
0'
#513810000000
1!
b100 %
1'
b100 +
#513820000000
0!
0'
#513830000000
1!
b101 %
1'
b101 +
#513840000000
0!
0'
#513850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#513860000000
0!
0'
#513870000000
1!
b111 %
1'
b111 +
#513880000000
0!
0'
#513890000000
1!
b1000 %
1'
b1000 +
#513900000000
0!
0'
#513910000000
1!
b1001 %
1'
b1001 +
#513920000000
0!
0'
#513930000000
1!
b0 %
1'
b0 +
#513940000000
0!
0'
#513950000000
1!
1$
b1 %
1'
1*
b1 +
#513960000000
0!
0'
#513970000000
1!
b10 %
1'
b10 +
#513980000000
0!
0'
#513990000000
1!
b11 %
1'
b11 +
#514000000000
0!
0'
#514010000000
1!
b100 %
1'
b100 +
#514020000000
0!
0'
#514030000000
1!
b101 %
1'
b101 +
#514040000000
0!
0'
#514050000000
1!
0$
b110 %
1'
0*
b110 +
#514060000000
1"
1(
#514070000000
0!
0"
b100 &
0'
0(
b100 ,
#514080000000
1!
1$
b111 %
1'
1*
b111 +
#514090000000
0!
0'
#514100000000
1!
0$
b1000 %
1'
0*
b1000 +
#514110000000
0!
0'
#514120000000
1!
b1001 %
1'
b1001 +
#514130000000
0!
0'
#514140000000
1!
b0 %
1'
b0 +
#514150000000
0!
0'
#514160000000
1!
1$
b1 %
1'
1*
b1 +
#514170000000
0!
0'
#514180000000
1!
b10 %
1'
b10 +
#514190000000
0!
0'
#514200000000
1!
b11 %
1'
b11 +
#514210000000
0!
0'
#514220000000
1!
b100 %
1'
b100 +
#514230000000
0!
0'
#514240000000
1!
b101 %
1'
b101 +
#514250000000
0!
0'
#514260000000
1!
b110 %
1'
b110 +
#514270000000
0!
0'
#514280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#514290000000
0!
0'
#514300000000
1!
b1000 %
1'
b1000 +
#514310000000
0!
0'
#514320000000
1!
b1001 %
1'
b1001 +
#514330000000
0!
0'
#514340000000
1!
b0 %
1'
b0 +
#514350000000
0!
0'
#514360000000
1!
1$
b1 %
1'
1*
b1 +
#514370000000
0!
0'
#514380000000
1!
b10 %
1'
b10 +
#514390000000
0!
0'
#514400000000
1!
b11 %
1'
b11 +
#514410000000
0!
0'
#514420000000
1!
b100 %
1'
b100 +
#514430000000
0!
0'
#514440000000
1!
b101 %
1'
b101 +
#514450000000
0!
0'
#514460000000
1!
0$
b110 %
1'
0*
b110 +
#514470000000
0!
0'
#514480000000
1!
b111 %
1'
b111 +
#514490000000
1"
1(
#514500000000
0!
0"
b100 &
0'
0(
b100 ,
#514510000000
1!
b1000 %
1'
b1000 +
#514520000000
0!
0'
#514530000000
1!
b1001 %
1'
b1001 +
#514540000000
0!
0'
#514550000000
1!
b0 %
1'
b0 +
#514560000000
0!
0'
#514570000000
1!
1$
b1 %
1'
1*
b1 +
#514580000000
0!
0'
#514590000000
1!
b10 %
1'
b10 +
#514600000000
0!
0'
#514610000000
1!
b11 %
1'
b11 +
#514620000000
0!
0'
#514630000000
1!
b100 %
1'
b100 +
#514640000000
0!
0'
#514650000000
1!
b101 %
1'
b101 +
#514660000000
0!
0'
#514670000000
1!
b110 %
1'
b110 +
#514680000000
0!
0'
#514690000000
1!
b111 %
1'
b111 +
#514700000000
0!
0'
#514710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#514720000000
0!
0'
#514730000000
1!
b1001 %
1'
b1001 +
#514740000000
0!
0'
#514750000000
1!
b0 %
1'
b0 +
#514760000000
0!
0'
#514770000000
1!
1$
b1 %
1'
1*
b1 +
#514780000000
0!
0'
#514790000000
1!
b10 %
1'
b10 +
#514800000000
0!
0'
#514810000000
1!
b11 %
1'
b11 +
#514820000000
0!
0'
#514830000000
1!
b100 %
1'
b100 +
#514840000000
0!
0'
#514850000000
1!
b101 %
1'
b101 +
#514860000000
0!
0'
#514870000000
1!
0$
b110 %
1'
0*
b110 +
#514880000000
0!
0'
#514890000000
1!
b111 %
1'
b111 +
#514900000000
0!
0'
#514910000000
1!
b1000 %
1'
b1000 +
#514920000000
1"
1(
#514930000000
0!
0"
b100 &
0'
0(
b100 ,
#514940000000
1!
b1001 %
1'
b1001 +
#514950000000
0!
0'
#514960000000
1!
b0 %
1'
b0 +
#514970000000
0!
0'
#514980000000
1!
1$
b1 %
1'
1*
b1 +
#514990000000
0!
0'
#515000000000
1!
b10 %
1'
b10 +
#515010000000
0!
0'
#515020000000
1!
b11 %
1'
b11 +
#515030000000
0!
0'
#515040000000
1!
b100 %
1'
b100 +
#515050000000
0!
0'
#515060000000
1!
b101 %
1'
b101 +
#515070000000
0!
0'
#515080000000
1!
b110 %
1'
b110 +
#515090000000
0!
0'
#515100000000
1!
b111 %
1'
b111 +
#515110000000
0!
0'
#515120000000
1!
0$
b1000 %
1'
0*
b1000 +
#515130000000
0!
0'
#515140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#515150000000
0!
0'
#515160000000
1!
b0 %
1'
b0 +
#515170000000
0!
0'
#515180000000
1!
1$
b1 %
1'
1*
b1 +
#515190000000
0!
0'
#515200000000
1!
b10 %
1'
b10 +
#515210000000
0!
0'
#515220000000
1!
b11 %
1'
b11 +
#515230000000
0!
0'
#515240000000
1!
b100 %
1'
b100 +
#515250000000
0!
0'
#515260000000
1!
b101 %
1'
b101 +
#515270000000
0!
0'
#515280000000
1!
0$
b110 %
1'
0*
b110 +
#515290000000
0!
0'
#515300000000
1!
b111 %
1'
b111 +
#515310000000
0!
0'
#515320000000
1!
b1000 %
1'
b1000 +
#515330000000
0!
0'
#515340000000
1!
b1001 %
1'
b1001 +
#515350000000
1"
1(
#515360000000
0!
0"
b100 &
0'
0(
b100 ,
#515370000000
1!
b0 %
1'
b0 +
#515380000000
0!
0'
#515390000000
1!
1$
b1 %
1'
1*
b1 +
#515400000000
0!
0'
#515410000000
1!
b10 %
1'
b10 +
#515420000000
0!
0'
#515430000000
1!
b11 %
1'
b11 +
#515440000000
0!
0'
#515450000000
1!
b100 %
1'
b100 +
#515460000000
0!
0'
#515470000000
1!
b101 %
1'
b101 +
#515480000000
0!
0'
#515490000000
1!
b110 %
1'
b110 +
#515500000000
0!
0'
#515510000000
1!
b111 %
1'
b111 +
#515520000000
0!
0'
#515530000000
1!
0$
b1000 %
1'
0*
b1000 +
#515540000000
0!
0'
#515550000000
1!
b1001 %
1'
b1001 +
#515560000000
0!
0'
#515570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#515580000000
0!
0'
#515590000000
1!
1$
b1 %
1'
1*
b1 +
#515600000000
0!
0'
#515610000000
1!
b10 %
1'
b10 +
#515620000000
0!
0'
#515630000000
1!
b11 %
1'
b11 +
#515640000000
0!
0'
#515650000000
1!
b100 %
1'
b100 +
#515660000000
0!
0'
#515670000000
1!
b101 %
1'
b101 +
#515680000000
0!
0'
#515690000000
1!
0$
b110 %
1'
0*
b110 +
#515700000000
0!
0'
#515710000000
1!
b111 %
1'
b111 +
#515720000000
0!
0'
#515730000000
1!
b1000 %
1'
b1000 +
#515740000000
0!
0'
#515750000000
1!
b1001 %
1'
b1001 +
#515760000000
0!
0'
#515770000000
1!
b0 %
1'
b0 +
#515780000000
1"
1(
#515790000000
0!
0"
b100 &
0'
0(
b100 ,
#515800000000
1!
1$
b1 %
1'
1*
b1 +
#515810000000
0!
0'
#515820000000
1!
b10 %
1'
b10 +
#515830000000
0!
0'
#515840000000
1!
b11 %
1'
b11 +
#515850000000
0!
0'
#515860000000
1!
b100 %
1'
b100 +
#515870000000
0!
0'
#515880000000
1!
b101 %
1'
b101 +
#515890000000
0!
0'
#515900000000
1!
b110 %
1'
b110 +
#515910000000
0!
0'
#515920000000
1!
b111 %
1'
b111 +
#515930000000
0!
0'
#515940000000
1!
0$
b1000 %
1'
0*
b1000 +
#515950000000
0!
0'
#515960000000
1!
b1001 %
1'
b1001 +
#515970000000
0!
0'
#515980000000
1!
b0 %
1'
b0 +
#515990000000
0!
0'
#516000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#516010000000
0!
0'
#516020000000
1!
b10 %
1'
b10 +
#516030000000
0!
0'
#516040000000
1!
b11 %
1'
b11 +
#516050000000
0!
0'
#516060000000
1!
b100 %
1'
b100 +
#516070000000
0!
0'
#516080000000
1!
b101 %
1'
b101 +
#516090000000
0!
0'
#516100000000
1!
0$
b110 %
1'
0*
b110 +
#516110000000
0!
0'
#516120000000
1!
b111 %
1'
b111 +
#516130000000
0!
0'
#516140000000
1!
b1000 %
1'
b1000 +
#516150000000
0!
0'
#516160000000
1!
b1001 %
1'
b1001 +
#516170000000
0!
0'
#516180000000
1!
b0 %
1'
b0 +
#516190000000
0!
0'
#516200000000
1!
1$
b1 %
1'
1*
b1 +
#516210000000
1"
1(
#516220000000
0!
0"
b100 &
0'
0(
b100 ,
#516230000000
1!
b10 %
1'
b10 +
#516240000000
0!
0'
#516250000000
1!
b11 %
1'
b11 +
#516260000000
0!
0'
#516270000000
1!
b100 %
1'
b100 +
#516280000000
0!
0'
#516290000000
1!
b101 %
1'
b101 +
#516300000000
0!
0'
#516310000000
1!
b110 %
1'
b110 +
#516320000000
0!
0'
#516330000000
1!
b111 %
1'
b111 +
#516340000000
0!
0'
#516350000000
1!
0$
b1000 %
1'
0*
b1000 +
#516360000000
0!
0'
#516370000000
1!
b1001 %
1'
b1001 +
#516380000000
0!
0'
#516390000000
1!
b0 %
1'
b0 +
#516400000000
0!
0'
#516410000000
1!
1$
b1 %
1'
1*
b1 +
#516420000000
0!
0'
#516430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#516440000000
0!
0'
#516450000000
1!
b11 %
1'
b11 +
#516460000000
0!
0'
#516470000000
1!
b100 %
1'
b100 +
#516480000000
0!
0'
#516490000000
1!
b101 %
1'
b101 +
#516500000000
0!
0'
#516510000000
1!
0$
b110 %
1'
0*
b110 +
#516520000000
0!
0'
#516530000000
1!
b111 %
1'
b111 +
#516540000000
0!
0'
#516550000000
1!
b1000 %
1'
b1000 +
#516560000000
0!
0'
#516570000000
1!
b1001 %
1'
b1001 +
#516580000000
0!
0'
#516590000000
1!
b0 %
1'
b0 +
#516600000000
0!
0'
#516610000000
1!
1$
b1 %
1'
1*
b1 +
#516620000000
0!
0'
#516630000000
1!
b10 %
1'
b10 +
#516640000000
1"
1(
#516650000000
0!
0"
b100 &
0'
0(
b100 ,
#516660000000
1!
b11 %
1'
b11 +
#516670000000
0!
0'
#516680000000
1!
b100 %
1'
b100 +
#516690000000
0!
0'
#516700000000
1!
b101 %
1'
b101 +
#516710000000
0!
0'
#516720000000
1!
b110 %
1'
b110 +
#516730000000
0!
0'
#516740000000
1!
b111 %
1'
b111 +
#516750000000
0!
0'
#516760000000
1!
0$
b1000 %
1'
0*
b1000 +
#516770000000
0!
0'
#516780000000
1!
b1001 %
1'
b1001 +
#516790000000
0!
0'
#516800000000
1!
b0 %
1'
b0 +
#516810000000
0!
0'
#516820000000
1!
1$
b1 %
1'
1*
b1 +
#516830000000
0!
0'
#516840000000
1!
b10 %
1'
b10 +
#516850000000
0!
0'
#516860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#516870000000
0!
0'
#516880000000
1!
b100 %
1'
b100 +
#516890000000
0!
0'
#516900000000
1!
b101 %
1'
b101 +
#516910000000
0!
0'
#516920000000
1!
0$
b110 %
1'
0*
b110 +
#516930000000
0!
0'
#516940000000
1!
b111 %
1'
b111 +
#516950000000
0!
0'
#516960000000
1!
b1000 %
1'
b1000 +
#516970000000
0!
0'
#516980000000
1!
b1001 %
1'
b1001 +
#516990000000
0!
0'
#517000000000
1!
b0 %
1'
b0 +
#517010000000
0!
0'
#517020000000
1!
1$
b1 %
1'
1*
b1 +
#517030000000
0!
0'
#517040000000
1!
b10 %
1'
b10 +
#517050000000
0!
0'
#517060000000
1!
b11 %
1'
b11 +
#517070000000
1"
1(
#517080000000
0!
0"
b100 &
0'
0(
b100 ,
#517090000000
1!
b100 %
1'
b100 +
#517100000000
0!
0'
#517110000000
1!
b101 %
1'
b101 +
#517120000000
0!
0'
#517130000000
1!
b110 %
1'
b110 +
#517140000000
0!
0'
#517150000000
1!
b111 %
1'
b111 +
#517160000000
0!
0'
#517170000000
1!
0$
b1000 %
1'
0*
b1000 +
#517180000000
0!
0'
#517190000000
1!
b1001 %
1'
b1001 +
#517200000000
0!
0'
#517210000000
1!
b0 %
1'
b0 +
#517220000000
0!
0'
#517230000000
1!
1$
b1 %
1'
1*
b1 +
#517240000000
0!
0'
#517250000000
1!
b10 %
1'
b10 +
#517260000000
0!
0'
#517270000000
1!
b11 %
1'
b11 +
#517280000000
0!
0'
#517290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#517300000000
0!
0'
#517310000000
1!
b101 %
1'
b101 +
#517320000000
0!
0'
#517330000000
1!
0$
b110 %
1'
0*
b110 +
#517340000000
0!
0'
#517350000000
1!
b111 %
1'
b111 +
#517360000000
0!
0'
#517370000000
1!
b1000 %
1'
b1000 +
#517380000000
0!
0'
#517390000000
1!
b1001 %
1'
b1001 +
#517400000000
0!
0'
#517410000000
1!
b0 %
1'
b0 +
#517420000000
0!
0'
#517430000000
1!
1$
b1 %
1'
1*
b1 +
#517440000000
0!
0'
#517450000000
1!
b10 %
1'
b10 +
#517460000000
0!
0'
#517470000000
1!
b11 %
1'
b11 +
#517480000000
0!
0'
#517490000000
1!
b100 %
1'
b100 +
#517500000000
1"
1(
#517510000000
0!
0"
b100 &
0'
0(
b100 ,
#517520000000
1!
b101 %
1'
b101 +
#517530000000
0!
0'
#517540000000
1!
b110 %
1'
b110 +
#517550000000
0!
0'
#517560000000
1!
b111 %
1'
b111 +
#517570000000
0!
0'
#517580000000
1!
0$
b1000 %
1'
0*
b1000 +
#517590000000
0!
0'
#517600000000
1!
b1001 %
1'
b1001 +
#517610000000
0!
0'
#517620000000
1!
b0 %
1'
b0 +
#517630000000
0!
0'
#517640000000
1!
1$
b1 %
1'
1*
b1 +
#517650000000
0!
0'
#517660000000
1!
b10 %
1'
b10 +
#517670000000
0!
0'
#517680000000
1!
b11 %
1'
b11 +
#517690000000
0!
0'
#517700000000
1!
b100 %
1'
b100 +
#517710000000
0!
0'
#517720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#517730000000
0!
0'
#517740000000
1!
0$
b110 %
1'
0*
b110 +
#517750000000
0!
0'
#517760000000
1!
b111 %
1'
b111 +
#517770000000
0!
0'
#517780000000
1!
b1000 %
1'
b1000 +
#517790000000
0!
0'
#517800000000
1!
b1001 %
1'
b1001 +
#517810000000
0!
0'
#517820000000
1!
b0 %
1'
b0 +
#517830000000
0!
0'
#517840000000
1!
1$
b1 %
1'
1*
b1 +
#517850000000
0!
0'
#517860000000
1!
b10 %
1'
b10 +
#517870000000
0!
0'
#517880000000
1!
b11 %
1'
b11 +
#517890000000
0!
0'
#517900000000
1!
b100 %
1'
b100 +
#517910000000
0!
0'
#517920000000
1!
b101 %
1'
b101 +
#517930000000
1"
1(
#517940000000
0!
0"
b100 &
0'
0(
b100 ,
#517950000000
1!
b110 %
1'
b110 +
#517960000000
0!
0'
#517970000000
1!
b111 %
1'
b111 +
#517980000000
0!
0'
#517990000000
1!
0$
b1000 %
1'
0*
b1000 +
#518000000000
0!
0'
#518010000000
1!
b1001 %
1'
b1001 +
#518020000000
0!
0'
#518030000000
1!
b0 %
1'
b0 +
#518040000000
0!
0'
#518050000000
1!
1$
b1 %
1'
1*
b1 +
#518060000000
0!
0'
#518070000000
1!
b10 %
1'
b10 +
#518080000000
0!
0'
#518090000000
1!
b11 %
1'
b11 +
#518100000000
0!
0'
#518110000000
1!
b100 %
1'
b100 +
#518120000000
0!
0'
#518130000000
1!
b101 %
1'
b101 +
#518140000000
0!
0'
#518150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#518160000000
0!
0'
#518170000000
1!
b111 %
1'
b111 +
#518180000000
0!
0'
#518190000000
1!
b1000 %
1'
b1000 +
#518200000000
0!
0'
#518210000000
1!
b1001 %
1'
b1001 +
#518220000000
0!
0'
#518230000000
1!
b0 %
1'
b0 +
#518240000000
0!
0'
#518250000000
1!
1$
b1 %
1'
1*
b1 +
#518260000000
0!
0'
#518270000000
1!
b10 %
1'
b10 +
#518280000000
0!
0'
#518290000000
1!
b11 %
1'
b11 +
#518300000000
0!
0'
#518310000000
1!
b100 %
1'
b100 +
#518320000000
0!
0'
#518330000000
1!
b101 %
1'
b101 +
#518340000000
0!
0'
#518350000000
1!
0$
b110 %
1'
0*
b110 +
#518360000000
1"
1(
#518370000000
0!
0"
b100 &
0'
0(
b100 ,
#518380000000
1!
1$
b111 %
1'
1*
b111 +
#518390000000
0!
0'
#518400000000
1!
0$
b1000 %
1'
0*
b1000 +
#518410000000
0!
0'
#518420000000
1!
b1001 %
1'
b1001 +
#518430000000
0!
0'
#518440000000
1!
b0 %
1'
b0 +
#518450000000
0!
0'
#518460000000
1!
1$
b1 %
1'
1*
b1 +
#518470000000
0!
0'
#518480000000
1!
b10 %
1'
b10 +
#518490000000
0!
0'
#518500000000
1!
b11 %
1'
b11 +
#518510000000
0!
0'
#518520000000
1!
b100 %
1'
b100 +
#518530000000
0!
0'
#518540000000
1!
b101 %
1'
b101 +
#518550000000
0!
0'
#518560000000
1!
b110 %
1'
b110 +
#518570000000
0!
0'
#518580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#518590000000
0!
0'
#518600000000
1!
b1000 %
1'
b1000 +
#518610000000
0!
0'
#518620000000
1!
b1001 %
1'
b1001 +
#518630000000
0!
0'
#518640000000
1!
b0 %
1'
b0 +
#518650000000
0!
0'
#518660000000
1!
1$
b1 %
1'
1*
b1 +
#518670000000
0!
0'
#518680000000
1!
b10 %
1'
b10 +
#518690000000
0!
0'
#518700000000
1!
b11 %
1'
b11 +
#518710000000
0!
0'
#518720000000
1!
b100 %
1'
b100 +
#518730000000
0!
0'
#518740000000
1!
b101 %
1'
b101 +
#518750000000
0!
0'
#518760000000
1!
0$
b110 %
1'
0*
b110 +
#518770000000
0!
0'
#518780000000
1!
b111 %
1'
b111 +
#518790000000
1"
1(
#518800000000
0!
0"
b100 &
0'
0(
b100 ,
#518810000000
1!
b1000 %
1'
b1000 +
#518820000000
0!
0'
#518830000000
1!
b1001 %
1'
b1001 +
#518840000000
0!
0'
#518850000000
1!
b0 %
1'
b0 +
#518860000000
0!
0'
#518870000000
1!
1$
b1 %
1'
1*
b1 +
#518880000000
0!
0'
#518890000000
1!
b10 %
1'
b10 +
#518900000000
0!
0'
#518910000000
1!
b11 %
1'
b11 +
#518920000000
0!
0'
#518930000000
1!
b100 %
1'
b100 +
#518940000000
0!
0'
#518950000000
1!
b101 %
1'
b101 +
#518960000000
0!
0'
#518970000000
1!
b110 %
1'
b110 +
#518980000000
0!
0'
#518990000000
1!
b111 %
1'
b111 +
#519000000000
0!
0'
#519010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#519020000000
0!
0'
#519030000000
1!
b1001 %
1'
b1001 +
#519040000000
0!
0'
#519050000000
1!
b0 %
1'
b0 +
#519060000000
0!
0'
#519070000000
1!
1$
b1 %
1'
1*
b1 +
#519080000000
0!
0'
#519090000000
1!
b10 %
1'
b10 +
#519100000000
0!
0'
#519110000000
1!
b11 %
1'
b11 +
#519120000000
0!
0'
#519130000000
1!
b100 %
1'
b100 +
#519140000000
0!
0'
#519150000000
1!
b101 %
1'
b101 +
#519160000000
0!
0'
#519170000000
1!
0$
b110 %
1'
0*
b110 +
#519180000000
0!
0'
#519190000000
1!
b111 %
1'
b111 +
#519200000000
0!
0'
#519210000000
1!
b1000 %
1'
b1000 +
#519220000000
1"
1(
#519230000000
0!
0"
b100 &
0'
0(
b100 ,
#519240000000
1!
b1001 %
1'
b1001 +
#519250000000
0!
0'
#519260000000
1!
b0 %
1'
b0 +
#519270000000
0!
0'
#519280000000
1!
1$
b1 %
1'
1*
b1 +
#519290000000
0!
0'
#519300000000
1!
b10 %
1'
b10 +
#519310000000
0!
0'
#519320000000
1!
b11 %
1'
b11 +
#519330000000
0!
0'
#519340000000
1!
b100 %
1'
b100 +
#519350000000
0!
0'
#519360000000
1!
b101 %
1'
b101 +
#519370000000
0!
0'
#519380000000
1!
b110 %
1'
b110 +
#519390000000
0!
0'
#519400000000
1!
b111 %
1'
b111 +
#519410000000
0!
0'
#519420000000
1!
0$
b1000 %
1'
0*
b1000 +
#519430000000
0!
0'
#519440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#519450000000
0!
0'
#519460000000
1!
b0 %
1'
b0 +
#519470000000
0!
0'
#519480000000
1!
1$
b1 %
1'
1*
b1 +
#519490000000
0!
0'
#519500000000
1!
b10 %
1'
b10 +
#519510000000
0!
0'
#519520000000
1!
b11 %
1'
b11 +
#519530000000
0!
0'
#519540000000
1!
b100 %
1'
b100 +
#519550000000
0!
0'
#519560000000
1!
b101 %
1'
b101 +
#519570000000
0!
0'
#519580000000
1!
0$
b110 %
1'
0*
b110 +
#519590000000
0!
0'
#519600000000
1!
b111 %
1'
b111 +
#519610000000
0!
0'
#519620000000
1!
b1000 %
1'
b1000 +
#519630000000
0!
0'
#519640000000
1!
b1001 %
1'
b1001 +
#519650000000
1"
1(
#519660000000
0!
0"
b100 &
0'
0(
b100 ,
#519670000000
1!
b0 %
1'
b0 +
#519680000000
0!
0'
#519690000000
1!
1$
b1 %
1'
1*
b1 +
#519700000000
0!
0'
#519710000000
1!
b10 %
1'
b10 +
#519720000000
0!
0'
#519730000000
1!
b11 %
1'
b11 +
#519740000000
0!
0'
#519750000000
1!
b100 %
1'
b100 +
#519760000000
0!
0'
#519770000000
1!
b101 %
1'
b101 +
#519780000000
0!
0'
#519790000000
1!
b110 %
1'
b110 +
#519800000000
0!
0'
#519810000000
1!
b111 %
1'
b111 +
#519820000000
0!
0'
#519830000000
1!
0$
b1000 %
1'
0*
b1000 +
#519840000000
0!
0'
#519850000000
1!
b1001 %
1'
b1001 +
#519860000000
0!
0'
#519870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#519880000000
0!
0'
#519890000000
1!
1$
b1 %
1'
1*
b1 +
#519900000000
0!
0'
#519910000000
1!
b10 %
1'
b10 +
#519920000000
0!
0'
#519930000000
1!
b11 %
1'
b11 +
#519940000000
0!
0'
#519950000000
1!
b100 %
1'
b100 +
#519960000000
0!
0'
#519970000000
1!
b101 %
1'
b101 +
#519980000000
0!
0'
#519990000000
1!
0$
b110 %
1'
0*
b110 +
#520000000000
0!
0'
#520010000000
1!
b111 %
1'
b111 +
#520020000000
0!
0'
#520030000000
1!
b1000 %
1'
b1000 +
#520040000000
0!
0'
#520050000000
1!
b1001 %
1'
b1001 +
#520060000000
0!
0'
#520070000000
1!
b0 %
1'
b0 +
#520080000000
1"
1(
#520090000000
0!
0"
b100 &
0'
0(
b100 ,
#520100000000
1!
1$
b1 %
1'
1*
b1 +
#520110000000
0!
0'
#520120000000
1!
b10 %
1'
b10 +
#520130000000
0!
0'
#520140000000
1!
b11 %
1'
b11 +
#520150000000
0!
0'
#520160000000
1!
b100 %
1'
b100 +
#520170000000
0!
0'
#520180000000
1!
b101 %
1'
b101 +
#520190000000
0!
0'
#520200000000
1!
b110 %
1'
b110 +
#520210000000
0!
0'
#520220000000
1!
b111 %
1'
b111 +
#520230000000
0!
0'
#520240000000
1!
0$
b1000 %
1'
0*
b1000 +
#520250000000
0!
0'
#520260000000
1!
b1001 %
1'
b1001 +
#520270000000
0!
0'
#520280000000
1!
b0 %
1'
b0 +
#520290000000
0!
0'
#520300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#520310000000
0!
0'
#520320000000
1!
b10 %
1'
b10 +
#520330000000
0!
0'
#520340000000
1!
b11 %
1'
b11 +
#520350000000
0!
0'
#520360000000
1!
b100 %
1'
b100 +
#520370000000
0!
0'
#520380000000
1!
b101 %
1'
b101 +
#520390000000
0!
0'
#520400000000
1!
0$
b110 %
1'
0*
b110 +
#520410000000
0!
0'
#520420000000
1!
b111 %
1'
b111 +
#520430000000
0!
0'
#520440000000
1!
b1000 %
1'
b1000 +
#520450000000
0!
0'
#520460000000
1!
b1001 %
1'
b1001 +
#520470000000
0!
0'
#520480000000
1!
b0 %
1'
b0 +
#520490000000
0!
0'
#520500000000
1!
1$
b1 %
1'
1*
b1 +
#520510000000
1"
1(
#520520000000
0!
0"
b100 &
0'
0(
b100 ,
#520530000000
1!
b10 %
1'
b10 +
#520540000000
0!
0'
#520550000000
1!
b11 %
1'
b11 +
#520560000000
0!
0'
#520570000000
1!
b100 %
1'
b100 +
#520580000000
0!
0'
#520590000000
1!
b101 %
1'
b101 +
#520600000000
0!
0'
#520610000000
1!
b110 %
1'
b110 +
#520620000000
0!
0'
#520630000000
1!
b111 %
1'
b111 +
#520640000000
0!
0'
#520650000000
1!
0$
b1000 %
1'
0*
b1000 +
#520660000000
0!
0'
#520670000000
1!
b1001 %
1'
b1001 +
#520680000000
0!
0'
#520690000000
1!
b0 %
1'
b0 +
#520700000000
0!
0'
#520710000000
1!
1$
b1 %
1'
1*
b1 +
#520720000000
0!
0'
#520730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#520740000000
0!
0'
#520750000000
1!
b11 %
1'
b11 +
#520760000000
0!
0'
#520770000000
1!
b100 %
1'
b100 +
#520780000000
0!
0'
#520790000000
1!
b101 %
1'
b101 +
#520800000000
0!
0'
#520810000000
1!
0$
b110 %
1'
0*
b110 +
#520820000000
0!
0'
#520830000000
1!
b111 %
1'
b111 +
#520840000000
0!
0'
#520850000000
1!
b1000 %
1'
b1000 +
#520860000000
0!
0'
#520870000000
1!
b1001 %
1'
b1001 +
#520880000000
0!
0'
#520890000000
1!
b0 %
1'
b0 +
#520900000000
0!
0'
#520910000000
1!
1$
b1 %
1'
1*
b1 +
#520920000000
0!
0'
#520930000000
1!
b10 %
1'
b10 +
#520940000000
1"
1(
#520950000000
0!
0"
b100 &
0'
0(
b100 ,
#520960000000
1!
b11 %
1'
b11 +
#520970000000
0!
0'
#520980000000
1!
b100 %
1'
b100 +
#520990000000
0!
0'
#521000000000
1!
b101 %
1'
b101 +
#521010000000
0!
0'
#521020000000
1!
b110 %
1'
b110 +
#521030000000
0!
0'
#521040000000
1!
b111 %
1'
b111 +
#521050000000
0!
0'
#521060000000
1!
0$
b1000 %
1'
0*
b1000 +
#521070000000
0!
0'
#521080000000
1!
b1001 %
1'
b1001 +
#521090000000
0!
0'
#521100000000
1!
b0 %
1'
b0 +
#521110000000
0!
0'
#521120000000
1!
1$
b1 %
1'
1*
b1 +
#521130000000
0!
0'
#521140000000
1!
b10 %
1'
b10 +
#521150000000
0!
0'
#521160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#521170000000
0!
0'
#521180000000
1!
b100 %
1'
b100 +
#521190000000
0!
0'
#521200000000
1!
b101 %
1'
b101 +
#521210000000
0!
0'
#521220000000
1!
0$
b110 %
1'
0*
b110 +
#521230000000
0!
0'
#521240000000
1!
b111 %
1'
b111 +
#521250000000
0!
0'
#521260000000
1!
b1000 %
1'
b1000 +
#521270000000
0!
0'
#521280000000
1!
b1001 %
1'
b1001 +
#521290000000
0!
0'
#521300000000
1!
b0 %
1'
b0 +
#521310000000
0!
0'
#521320000000
1!
1$
b1 %
1'
1*
b1 +
#521330000000
0!
0'
#521340000000
1!
b10 %
1'
b10 +
#521350000000
0!
0'
#521360000000
1!
b11 %
1'
b11 +
#521370000000
1"
1(
#521380000000
0!
0"
b100 &
0'
0(
b100 ,
#521390000000
1!
b100 %
1'
b100 +
#521400000000
0!
0'
#521410000000
1!
b101 %
1'
b101 +
#521420000000
0!
0'
#521430000000
1!
b110 %
1'
b110 +
#521440000000
0!
0'
#521450000000
1!
b111 %
1'
b111 +
#521460000000
0!
0'
#521470000000
1!
0$
b1000 %
1'
0*
b1000 +
#521480000000
0!
0'
#521490000000
1!
b1001 %
1'
b1001 +
#521500000000
0!
0'
#521510000000
1!
b0 %
1'
b0 +
#521520000000
0!
0'
#521530000000
1!
1$
b1 %
1'
1*
b1 +
#521540000000
0!
0'
#521550000000
1!
b10 %
1'
b10 +
#521560000000
0!
0'
#521570000000
1!
b11 %
1'
b11 +
#521580000000
0!
0'
#521590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#521600000000
0!
0'
#521610000000
1!
b101 %
1'
b101 +
#521620000000
0!
0'
#521630000000
1!
0$
b110 %
1'
0*
b110 +
#521640000000
0!
0'
#521650000000
1!
b111 %
1'
b111 +
#521660000000
0!
0'
#521670000000
1!
b1000 %
1'
b1000 +
#521680000000
0!
0'
#521690000000
1!
b1001 %
1'
b1001 +
#521700000000
0!
0'
#521710000000
1!
b0 %
1'
b0 +
#521720000000
0!
0'
#521730000000
1!
1$
b1 %
1'
1*
b1 +
#521740000000
0!
0'
#521750000000
1!
b10 %
1'
b10 +
#521760000000
0!
0'
#521770000000
1!
b11 %
1'
b11 +
#521780000000
0!
0'
#521790000000
1!
b100 %
1'
b100 +
#521800000000
1"
1(
#521810000000
0!
0"
b100 &
0'
0(
b100 ,
#521820000000
1!
b101 %
1'
b101 +
#521830000000
0!
0'
#521840000000
1!
b110 %
1'
b110 +
#521850000000
0!
0'
#521860000000
1!
b111 %
1'
b111 +
#521870000000
0!
0'
#521880000000
1!
0$
b1000 %
1'
0*
b1000 +
#521890000000
0!
0'
#521900000000
1!
b1001 %
1'
b1001 +
#521910000000
0!
0'
#521920000000
1!
b0 %
1'
b0 +
#521930000000
0!
0'
#521940000000
1!
1$
b1 %
1'
1*
b1 +
#521950000000
0!
0'
#521960000000
1!
b10 %
1'
b10 +
#521970000000
0!
0'
#521980000000
1!
b11 %
1'
b11 +
#521990000000
0!
0'
#522000000000
1!
b100 %
1'
b100 +
#522010000000
0!
0'
#522020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#522030000000
0!
0'
#522040000000
1!
0$
b110 %
1'
0*
b110 +
#522050000000
0!
0'
#522060000000
1!
b111 %
1'
b111 +
#522070000000
0!
0'
#522080000000
1!
b1000 %
1'
b1000 +
#522090000000
0!
0'
#522100000000
1!
b1001 %
1'
b1001 +
#522110000000
0!
0'
#522120000000
1!
b0 %
1'
b0 +
#522130000000
0!
0'
#522140000000
1!
1$
b1 %
1'
1*
b1 +
#522150000000
0!
0'
#522160000000
1!
b10 %
1'
b10 +
#522170000000
0!
0'
#522180000000
1!
b11 %
1'
b11 +
#522190000000
0!
0'
#522200000000
1!
b100 %
1'
b100 +
#522210000000
0!
0'
#522220000000
1!
b101 %
1'
b101 +
#522230000000
1"
1(
#522240000000
0!
0"
b100 &
0'
0(
b100 ,
#522250000000
1!
b110 %
1'
b110 +
#522260000000
0!
0'
#522270000000
1!
b111 %
1'
b111 +
#522280000000
0!
0'
#522290000000
1!
0$
b1000 %
1'
0*
b1000 +
#522300000000
0!
0'
#522310000000
1!
b1001 %
1'
b1001 +
#522320000000
0!
0'
#522330000000
1!
b0 %
1'
b0 +
#522340000000
0!
0'
#522350000000
1!
1$
b1 %
1'
1*
b1 +
#522360000000
0!
0'
#522370000000
1!
b10 %
1'
b10 +
#522380000000
0!
0'
#522390000000
1!
b11 %
1'
b11 +
#522400000000
0!
0'
#522410000000
1!
b100 %
1'
b100 +
#522420000000
0!
0'
#522430000000
1!
b101 %
1'
b101 +
#522440000000
0!
0'
#522450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#522460000000
0!
0'
#522470000000
1!
b111 %
1'
b111 +
#522480000000
0!
0'
#522490000000
1!
b1000 %
1'
b1000 +
#522500000000
0!
0'
#522510000000
1!
b1001 %
1'
b1001 +
#522520000000
0!
0'
#522530000000
1!
b0 %
1'
b0 +
#522540000000
0!
0'
#522550000000
1!
1$
b1 %
1'
1*
b1 +
#522560000000
0!
0'
#522570000000
1!
b10 %
1'
b10 +
#522580000000
0!
0'
#522590000000
1!
b11 %
1'
b11 +
#522600000000
0!
0'
#522610000000
1!
b100 %
1'
b100 +
#522620000000
0!
0'
#522630000000
1!
b101 %
1'
b101 +
#522640000000
0!
0'
#522650000000
1!
0$
b110 %
1'
0*
b110 +
#522660000000
1"
1(
#522670000000
0!
0"
b100 &
0'
0(
b100 ,
#522680000000
1!
1$
b111 %
1'
1*
b111 +
#522690000000
0!
0'
#522700000000
1!
0$
b1000 %
1'
0*
b1000 +
#522710000000
0!
0'
#522720000000
1!
b1001 %
1'
b1001 +
#522730000000
0!
0'
#522740000000
1!
b0 %
1'
b0 +
#522750000000
0!
0'
#522760000000
1!
1$
b1 %
1'
1*
b1 +
#522770000000
0!
0'
#522780000000
1!
b10 %
1'
b10 +
#522790000000
0!
0'
#522800000000
1!
b11 %
1'
b11 +
#522810000000
0!
0'
#522820000000
1!
b100 %
1'
b100 +
#522830000000
0!
0'
#522840000000
1!
b101 %
1'
b101 +
#522850000000
0!
0'
#522860000000
1!
b110 %
1'
b110 +
#522870000000
0!
0'
#522880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#522890000000
0!
0'
#522900000000
1!
b1000 %
1'
b1000 +
#522910000000
0!
0'
#522920000000
1!
b1001 %
1'
b1001 +
#522930000000
0!
0'
#522940000000
1!
b0 %
1'
b0 +
#522950000000
0!
0'
#522960000000
1!
1$
b1 %
1'
1*
b1 +
#522970000000
0!
0'
#522980000000
1!
b10 %
1'
b10 +
#522990000000
0!
0'
#523000000000
1!
b11 %
1'
b11 +
#523010000000
0!
0'
#523020000000
1!
b100 %
1'
b100 +
#523030000000
0!
0'
#523040000000
1!
b101 %
1'
b101 +
#523050000000
0!
0'
#523060000000
1!
0$
b110 %
1'
0*
b110 +
#523070000000
0!
0'
#523080000000
1!
b111 %
1'
b111 +
#523090000000
1"
1(
#523100000000
0!
0"
b100 &
0'
0(
b100 ,
#523110000000
1!
b1000 %
1'
b1000 +
#523120000000
0!
0'
#523130000000
1!
b1001 %
1'
b1001 +
#523140000000
0!
0'
#523150000000
1!
b0 %
1'
b0 +
#523160000000
0!
0'
#523170000000
1!
1$
b1 %
1'
1*
b1 +
#523180000000
0!
0'
#523190000000
1!
b10 %
1'
b10 +
#523200000000
0!
0'
#523210000000
1!
b11 %
1'
b11 +
#523220000000
0!
0'
#523230000000
1!
b100 %
1'
b100 +
#523240000000
0!
0'
#523250000000
1!
b101 %
1'
b101 +
#523260000000
0!
0'
#523270000000
1!
b110 %
1'
b110 +
#523280000000
0!
0'
#523290000000
1!
b111 %
1'
b111 +
#523300000000
0!
0'
#523310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#523320000000
0!
0'
#523330000000
1!
b1001 %
1'
b1001 +
#523340000000
0!
0'
#523350000000
1!
b0 %
1'
b0 +
#523360000000
0!
0'
#523370000000
1!
1$
b1 %
1'
1*
b1 +
#523380000000
0!
0'
#523390000000
1!
b10 %
1'
b10 +
#523400000000
0!
0'
#523410000000
1!
b11 %
1'
b11 +
#523420000000
0!
0'
#523430000000
1!
b100 %
1'
b100 +
#523440000000
0!
0'
#523450000000
1!
b101 %
1'
b101 +
#523460000000
0!
0'
#523470000000
1!
0$
b110 %
1'
0*
b110 +
#523480000000
0!
0'
#523490000000
1!
b111 %
1'
b111 +
#523500000000
0!
0'
#523510000000
1!
b1000 %
1'
b1000 +
#523520000000
1"
1(
#523530000000
0!
0"
b100 &
0'
0(
b100 ,
#523540000000
1!
b1001 %
1'
b1001 +
#523550000000
0!
0'
#523560000000
1!
b0 %
1'
b0 +
#523570000000
0!
0'
#523580000000
1!
1$
b1 %
1'
1*
b1 +
#523590000000
0!
0'
#523600000000
1!
b10 %
1'
b10 +
#523610000000
0!
0'
#523620000000
1!
b11 %
1'
b11 +
#523630000000
0!
0'
#523640000000
1!
b100 %
1'
b100 +
#523650000000
0!
0'
#523660000000
1!
b101 %
1'
b101 +
#523670000000
0!
0'
#523680000000
1!
b110 %
1'
b110 +
#523690000000
0!
0'
#523700000000
1!
b111 %
1'
b111 +
#523710000000
0!
0'
#523720000000
1!
0$
b1000 %
1'
0*
b1000 +
#523730000000
0!
0'
#523740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#523750000000
0!
0'
#523760000000
1!
b0 %
1'
b0 +
#523770000000
0!
0'
#523780000000
1!
1$
b1 %
1'
1*
b1 +
#523790000000
0!
0'
#523800000000
1!
b10 %
1'
b10 +
#523810000000
0!
0'
#523820000000
1!
b11 %
1'
b11 +
#523830000000
0!
0'
#523840000000
1!
b100 %
1'
b100 +
#523850000000
0!
0'
#523860000000
1!
b101 %
1'
b101 +
#523870000000
0!
0'
#523880000000
1!
0$
b110 %
1'
0*
b110 +
#523890000000
0!
0'
#523900000000
1!
b111 %
1'
b111 +
#523910000000
0!
0'
#523920000000
1!
b1000 %
1'
b1000 +
#523930000000
0!
0'
#523940000000
1!
b1001 %
1'
b1001 +
#523950000000
1"
1(
#523960000000
0!
0"
b100 &
0'
0(
b100 ,
#523970000000
1!
b0 %
1'
b0 +
#523980000000
0!
0'
#523990000000
1!
1$
b1 %
1'
1*
b1 +
#524000000000
0!
0'
#524010000000
1!
b10 %
1'
b10 +
#524020000000
0!
0'
#524030000000
1!
b11 %
1'
b11 +
#524040000000
0!
0'
#524050000000
1!
b100 %
1'
b100 +
#524060000000
0!
0'
#524070000000
1!
b101 %
1'
b101 +
#524080000000
0!
0'
#524090000000
1!
b110 %
1'
b110 +
#524100000000
0!
0'
#524110000000
1!
b111 %
1'
b111 +
#524120000000
0!
0'
#524130000000
1!
0$
b1000 %
1'
0*
b1000 +
#524140000000
0!
0'
#524150000000
1!
b1001 %
1'
b1001 +
#524160000000
0!
0'
#524170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#524180000000
0!
0'
#524190000000
1!
1$
b1 %
1'
1*
b1 +
#524200000000
0!
0'
#524210000000
1!
b10 %
1'
b10 +
#524220000000
0!
0'
#524230000000
1!
b11 %
1'
b11 +
#524240000000
0!
0'
#524250000000
1!
b100 %
1'
b100 +
#524260000000
0!
0'
#524270000000
1!
b101 %
1'
b101 +
#524280000000
0!
0'
#524290000000
1!
0$
b110 %
1'
0*
b110 +
#524300000000
0!
0'
#524310000000
1!
b111 %
1'
b111 +
#524320000000
0!
0'
#524330000000
1!
b1000 %
1'
b1000 +
#524340000000
0!
0'
#524350000000
1!
b1001 %
1'
b1001 +
#524360000000
0!
0'
#524370000000
1!
b0 %
1'
b0 +
#524380000000
1"
1(
#524390000000
0!
0"
b100 &
0'
0(
b100 ,
#524400000000
1!
1$
b1 %
1'
1*
b1 +
#524410000000
0!
0'
#524420000000
1!
b10 %
1'
b10 +
#524430000000
0!
0'
#524440000000
1!
b11 %
1'
b11 +
#524450000000
0!
0'
#524460000000
1!
b100 %
1'
b100 +
#524470000000
0!
0'
#524480000000
1!
b101 %
1'
b101 +
#524490000000
0!
0'
#524500000000
1!
b110 %
1'
b110 +
#524510000000
0!
0'
#524520000000
1!
b111 %
1'
b111 +
#524530000000
0!
0'
#524540000000
1!
0$
b1000 %
1'
0*
b1000 +
#524550000000
0!
0'
#524560000000
1!
b1001 %
1'
b1001 +
#524570000000
0!
0'
#524580000000
1!
b0 %
1'
b0 +
#524590000000
0!
0'
#524600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#524610000000
0!
0'
#524620000000
1!
b10 %
1'
b10 +
#524630000000
0!
0'
#524640000000
1!
b11 %
1'
b11 +
#524650000000
0!
0'
#524660000000
1!
b100 %
1'
b100 +
#524670000000
0!
0'
#524680000000
1!
b101 %
1'
b101 +
#524690000000
0!
0'
#524700000000
1!
0$
b110 %
1'
0*
b110 +
#524710000000
0!
0'
#524720000000
1!
b111 %
1'
b111 +
#524730000000
0!
0'
#524740000000
1!
b1000 %
1'
b1000 +
#524750000000
0!
0'
#524760000000
1!
b1001 %
1'
b1001 +
#524770000000
0!
0'
#524780000000
1!
b0 %
1'
b0 +
#524790000000
0!
0'
#524800000000
1!
1$
b1 %
1'
1*
b1 +
#524810000000
1"
1(
#524820000000
0!
0"
b100 &
0'
0(
b100 ,
#524830000000
1!
b10 %
1'
b10 +
#524840000000
0!
0'
#524850000000
1!
b11 %
1'
b11 +
#524860000000
0!
0'
#524870000000
1!
b100 %
1'
b100 +
#524880000000
0!
0'
#524890000000
1!
b101 %
1'
b101 +
#524900000000
0!
0'
#524910000000
1!
b110 %
1'
b110 +
#524920000000
0!
0'
#524930000000
1!
b111 %
1'
b111 +
#524940000000
0!
0'
#524950000000
1!
0$
b1000 %
1'
0*
b1000 +
#524960000000
0!
0'
#524970000000
1!
b1001 %
1'
b1001 +
#524980000000
0!
0'
#524990000000
1!
b0 %
1'
b0 +
#525000000000
0!
0'
#525010000000
1!
1$
b1 %
1'
1*
b1 +
#525020000000
0!
0'
#525030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#525040000000
0!
0'
#525050000000
1!
b11 %
1'
b11 +
#525060000000
0!
0'
#525070000000
1!
b100 %
1'
b100 +
#525080000000
0!
0'
#525090000000
1!
b101 %
1'
b101 +
#525100000000
0!
0'
#525110000000
1!
0$
b110 %
1'
0*
b110 +
#525120000000
0!
0'
#525130000000
1!
b111 %
1'
b111 +
#525140000000
0!
0'
#525150000000
1!
b1000 %
1'
b1000 +
#525160000000
0!
0'
#525170000000
1!
b1001 %
1'
b1001 +
#525180000000
0!
0'
#525190000000
1!
b0 %
1'
b0 +
#525200000000
0!
0'
#525210000000
1!
1$
b1 %
1'
1*
b1 +
#525220000000
0!
0'
#525230000000
1!
b10 %
1'
b10 +
#525240000000
1"
1(
#525250000000
0!
0"
b100 &
0'
0(
b100 ,
#525260000000
1!
b11 %
1'
b11 +
#525270000000
0!
0'
#525280000000
1!
b100 %
1'
b100 +
#525290000000
0!
0'
#525300000000
1!
b101 %
1'
b101 +
#525310000000
0!
0'
#525320000000
1!
b110 %
1'
b110 +
#525330000000
0!
0'
#525340000000
1!
b111 %
1'
b111 +
#525350000000
0!
0'
#525360000000
1!
0$
b1000 %
1'
0*
b1000 +
#525370000000
0!
0'
#525380000000
1!
b1001 %
1'
b1001 +
#525390000000
0!
0'
#525400000000
1!
b0 %
1'
b0 +
#525410000000
0!
0'
#525420000000
1!
1$
b1 %
1'
1*
b1 +
#525430000000
0!
0'
#525440000000
1!
b10 %
1'
b10 +
#525450000000
0!
0'
#525460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#525470000000
0!
0'
#525480000000
1!
b100 %
1'
b100 +
#525490000000
0!
0'
#525500000000
1!
b101 %
1'
b101 +
#525510000000
0!
0'
#525520000000
1!
0$
b110 %
1'
0*
b110 +
#525530000000
0!
0'
#525540000000
1!
b111 %
1'
b111 +
#525550000000
0!
0'
#525560000000
1!
b1000 %
1'
b1000 +
#525570000000
0!
0'
#525580000000
1!
b1001 %
1'
b1001 +
#525590000000
0!
0'
#525600000000
1!
b0 %
1'
b0 +
#525610000000
0!
0'
#525620000000
1!
1$
b1 %
1'
1*
b1 +
#525630000000
0!
0'
#525640000000
1!
b10 %
1'
b10 +
#525650000000
0!
0'
#525660000000
1!
b11 %
1'
b11 +
#525670000000
1"
1(
#525680000000
0!
0"
b100 &
0'
0(
b100 ,
#525690000000
1!
b100 %
1'
b100 +
#525700000000
0!
0'
#525710000000
1!
b101 %
1'
b101 +
#525720000000
0!
0'
#525730000000
1!
b110 %
1'
b110 +
#525740000000
0!
0'
#525750000000
1!
b111 %
1'
b111 +
#525760000000
0!
0'
#525770000000
1!
0$
b1000 %
1'
0*
b1000 +
#525780000000
0!
0'
#525790000000
1!
b1001 %
1'
b1001 +
#525800000000
0!
0'
#525810000000
1!
b0 %
1'
b0 +
#525820000000
0!
0'
#525830000000
1!
1$
b1 %
1'
1*
b1 +
#525840000000
0!
0'
#525850000000
1!
b10 %
1'
b10 +
#525860000000
0!
0'
#525870000000
1!
b11 %
1'
b11 +
#525880000000
0!
0'
#525890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#525900000000
0!
0'
#525910000000
1!
b101 %
1'
b101 +
#525920000000
0!
0'
#525930000000
1!
0$
b110 %
1'
0*
b110 +
#525940000000
0!
0'
#525950000000
1!
b111 %
1'
b111 +
#525960000000
0!
0'
#525970000000
1!
b1000 %
1'
b1000 +
#525980000000
0!
0'
#525990000000
1!
b1001 %
1'
b1001 +
#526000000000
0!
0'
#526010000000
1!
b0 %
1'
b0 +
#526020000000
0!
0'
#526030000000
1!
1$
b1 %
1'
1*
b1 +
#526040000000
0!
0'
#526050000000
1!
b10 %
1'
b10 +
#526060000000
0!
0'
#526070000000
1!
b11 %
1'
b11 +
#526080000000
0!
0'
#526090000000
1!
b100 %
1'
b100 +
#526100000000
1"
1(
#526110000000
0!
0"
b100 &
0'
0(
b100 ,
#526120000000
1!
b101 %
1'
b101 +
#526130000000
0!
0'
#526140000000
1!
b110 %
1'
b110 +
#526150000000
0!
0'
#526160000000
1!
b111 %
1'
b111 +
#526170000000
0!
0'
#526180000000
1!
0$
b1000 %
1'
0*
b1000 +
#526190000000
0!
0'
#526200000000
1!
b1001 %
1'
b1001 +
#526210000000
0!
0'
#526220000000
1!
b0 %
1'
b0 +
#526230000000
0!
0'
#526240000000
1!
1$
b1 %
1'
1*
b1 +
#526250000000
0!
0'
#526260000000
1!
b10 %
1'
b10 +
#526270000000
0!
0'
#526280000000
1!
b11 %
1'
b11 +
#526290000000
0!
0'
#526300000000
1!
b100 %
1'
b100 +
#526310000000
0!
0'
#526320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#526330000000
0!
0'
#526340000000
1!
0$
b110 %
1'
0*
b110 +
#526350000000
0!
0'
#526360000000
1!
b111 %
1'
b111 +
#526370000000
0!
0'
#526380000000
1!
b1000 %
1'
b1000 +
#526390000000
0!
0'
#526400000000
1!
b1001 %
1'
b1001 +
#526410000000
0!
0'
#526420000000
1!
b0 %
1'
b0 +
#526430000000
0!
0'
#526440000000
1!
1$
b1 %
1'
1*
b1 +
#526450000000
0!
0'
#526460000000
1!
b10 %
1'
b10 +
#526470000000
0!
0'
#526480000000
1!
b11 %
1'
b11 +
#526490000000
0!
0'
#526500000000
1!
b100 %
1'
b100 +
#526510000000
0!
0'
#526520000000
1!
b101 %
1'
b101 +
#526530000000
1"
1(
#526540000000
0!
0"
b100 &
0'
0(
b100 ,
#526550000000
1!
b110 %
1'
b110 +
#526560000000
0!
0'
#526570000000
1!
b111 %
1'
b111 +
#526580000000
0!
0'
#526590000000
1!
0$
b1000 %
1'
0*
b1000 +
#526600000000
0!
0'
#526610000000
1!
b1001 %
1'
b1001 +
#526620000000
0!
0'
#526630000000
1!
b0 %
1'
b0 +
#526640000000
0!
0'
#526650000000
1!
1$
b1 %
1'
1*
b1 +
#526660000000
0!
0'
#526670000000
1!
b10 %
1'
b10 +
#526680000000
0!
0'
#526690000000
1!
b11 %
1'
b11 +
#526700000000
0!
0'
#526710000000
1!
b100 %
1'
b100 +
#526720000000
0!
0'
#526730000000
1!
b101 %
1'
b101 +
#526740000000
0!
0'
#526750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#526760000000
0!
0'
#526770000000
1!
b111 %
1'
b111 +
#526780000000
0!
0'
#526790000000
1!
b1000 %
1'
b1000 +
#526800000000
0!
0'
#526810000000
1!
b1001 %
1'
b1001 +
#526820000000
0!
0'
#526830000000
1!
b0 %
1'
b0 +
#526840000000
0!
0'
#526850000000
1!
1$
b1 %
1'
1*
b1 +
#526860000000
0!
0'
#526870000000
1!
b10 %
1'
b10 +
#526880000000
0!
0'
#526890000000
1!
b11 %
1'
b11 +
#526900000000
0!
0'
#526910000000
1!
b100 %
1'
b100 +
#526920000000
0!
0'
#526930000000
1!
b101 %
1'
b101 +
#526940000000
0!
0'
#526950000000
1!
0$
b110 %
1'
0*
b110 +
#526960000000
1"
1(
#526970000000
0!
0"
b100 &
0'
0(
b100 ,
#526980000000
1!
1$
b111 %
1'
1*
b111 +
#526990000000
0!
0'
#527000000000
1!
0$
b1000 %
1'
0*
b1000 +
#527010000000
0!
0'
#527020000000
1!
b1001 %
1'
b1001 +
#527030000000
0!
0'
#527040000000
1!
b0 %
1'
b0 +
#527050000000
0!
0'
#527060000000
1!
1$
b1 %
1'
1*
b1 +
#527070000000
0!
0'
#527080000000
1!
b10 %
1'
b10 +
#527090000000
0!
0'
#527100000000
1!
b11 %
1'
b11 +
#527110000000
0!
0'
#527120000000
1!
b100 %
1'
b100 +
#527130000000
0!
0'
#527140000000
1!
b101 %
1'
b101 +
#527150000000
0!
0'
#527160000000
1!
b110 %
1'
b110 +
#527170000000
0!
0'
#527180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#527190000000
0!
0'
#527200000000
1!
b1000 %
1'
b1000 +
#527210000000
0!
0'
#527220000000
1!
b1001 %
1'
b1001 +
#527230000000
0!
0'
#527240000000
1!
b0 %
1'
b0 +
#527250000000
0!
0'
#527260000000
1!
1$
b1 %
1'
1*
b1 +
#527270000000
0!
0'
#527280000000
1!
b10 %
1'
b10 +
#527290000000
0!
0'
#527300000000
1!
b11 %
1'
b11 +
#527310000000
0!
0'
#527320000000
1!
b100 %
1'
b100 +
#527330000000
0!
0'
#527340000000
1!
b101 %
1'
b101 +
#527350000000
0!
0'
#527360000000
1!
0$
b110 %
1'
0*
b110 +
#527370000000
0!
0'
#527380000000
1!
b111 %
1'
b111 +
#527390000000
1"
1(
#527400000000
0!
0"
b100 &
0'
0(
b100 ,
#527410000000
1!
b1000 %
1'
b1000 +
#527420000000
0!
0'
#527430000000
1!
b1001 %
1'
b1001 +
#527440000000
0!
0'
#527450000000
1!
b0 %
1'
b0 +
#527460000000
0!
0'
#527470000000
1!
1$
b1 %
1'
1*
b1 +
#527480000000
0!
0'
#527490000000
1!
b10 %
1'
b10 +
#527500000000
0!
0'
#527510000000
1!
b11 %
1'
b11 +
#527520000000
0!
0'
#527530000000
1!
b100 %
1'
b100 +
#527540000000
0!
0'
#527550000000
1!
b101 %
1'
b101 +
#527560000000
0!
0'
#527570000000
1!
b110 %
1'
b110 +
#527580000000
0!
0'
#527590000000
1!
b111 %
1'
b111 +
#527600000000
0!
0'
#527610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#527620000000
0!
0'
#527630000000
1!
b1001 %
1'
b1001 +
#527640000000
0!
0'
#527650000000
1!
b0 %
1'
b0 +
#527660000000
0!
0'
#527670000000
1!
1$
b1 %
1'
1*
b1 +
#527680000000
0!
0'
#527690000000
1!
b10 %
1'
b10 +
#527700000000
0!
0'
#527710000000
1!
b11 %
1'
b11 +
#527720000000
0!
0'
#527730000000
1!
b100 %
1'
b100 +
#527740000000
0!
0'
#527750000000
1!
b101 %
1'
b101 +
#527760000000
0!
0'
#527770000000
1!
0$
b110 %
1'
0*
b110 +
#527780000000
0!
0'
#527790000000
1!
b111 %
1'
b111 +
#527800000000
0!
0'
#527810000000
1!
b1000 %
1'
b1000 +
#527820000000
1"
1(
#527830000000
0!
0"
b100 &
0'
0(
b100 ,
#527840000000
1!
b1001 %
1'
b1001 +
#527850000000
0!
0'
#527860000000
1!
b0 %
1'
b0 +
#527870000000
0!
0'
#527880000000
1!
1$
b1 %
1'
1*
b1 +
#527890000000
0!
0'
#527900000000
1!
b10 %
1'
b10 +
#527910000000
0!
0'
#527920000000
1!
b11 %
1'
b11 +
#527930000000
0!
0'
#527940000000
1!
b100 %
1'
b100 +
#527950000000
0!
0'
#527960000000
1!
b101 %
1'
b101 +
#527970000000
0!
0'
#527980000000
1!
b110 %
1'
b110 +
#527990000000
0!
0'
#528000000000
1!
b111 %
1'
b111 +
#528010000000
0!
0'
#528020000000
1!
0$
b1000 %
1'
0*
b1000 +
#528030000000
0!
0'
#528040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#528050000000
0!
0'
#528060000000
1!
b0 %
1'
b0 +
#528070000000
0!
0'
#528080000000
1!
1$
b1 %
1'
1*
b1 +
#528090000000
0!
0'
#528100000000
1!
b10 %
1'
b10 +
#528110000000
0!
0'
#528120000000
1!
b11 %
1'
b11 +
#528130000000
0!
0'
#528140000000
1!
b100 %
1'
b100 +
#528150000000
0!
0'
#528160000000
1!
b101 %
1'
b101 +
#528170000000
0!
0'
#528180000000
1!
0$
b110 %
1'
0*
b110 +
#528190000000
0!
0'
#528200000000
1!
b111 %
1'
b111 +
#528210000000
0!
0'
#528220000000
1!
b1000 %
1'
b1000 +
#528230000000
0!
0'
#528240000000
1!
b1001 %
1'
b1001 +
#528250000000
1"
1(
#528260000000
0!
0"
b100 &
0'
0(
b100 ,
#528270000000
1!
b0 %
1'
b0 +
#528280000000
0!
0'
#528290000000
1!
1$
b1 %
1'
1*
b1 +
#528300000000
0!
0'
#528310000000
1!
b10 %
1'
b10 +
#528320000000
0!
0'
#528330000000
1!
b11 %
1'
b11 +
#528340000000
0!
0'
#528350000000
1!
b100 %
1'
b100 +
#528360000000
0!
0'
#528370000000
1!
b101 %
1'
b101 +
#528380000000
0!
0'
#528390000000
1!
b110 %
1'
b110 +
#528400000000
0!
0'
#528410000000
1!
b111 %
1'
b111 +
#528420000000
0!
0'
#528430000000
1!
0$
b1000 %
1'
0*
b1000 +
#528440000000
0!
0'
#528450000000
1!
b1001 %
1'
b1001 +
#528460000000
0!
0'
#528470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#528480000000
0!
0'
#528490000000
1!
1$
b1 %
1'
1*
b1 +
#528500000000
0!
0'
#528510000000
1!
b10 %
1'
b10 +
#528520000000
0!
0'
#528530000000
1!
b11 %
1'
b11 +
#528540000000
0!
0'
#528550000000
1!
b100 %
1'
b100 +
#528560000000
0!
0'
#528570000000
1!
b101 %
1'
b101 +
#528580000000
0!
0'
#528590000000
1!
0$
b110 %
1'
0*
b110 +
#528600000000
0!
0'
#528610000000
1!
b111 %
1'
b111 +
#528620000000
0!
0'
#528630000000
1!
b1000 %
1'
b1000 +
#528640000000
0!
0'
#528650000000
1!
b1001 %
1'
b1001 +
#528660000000
0!
0'
#528670000000
1!
b0 %
1'
b0 +
#528680000000
1"
1(
#528690000000
0!
0"
b100 &
0'
0(
b100 ,
#528700000000
1!
1$
b1 %
1'
1*
b1 +
#528710000000
0!
0'
#528720000000
1!
b10 %
1'
b10 +
#528730000000
0!
0'
#528740000000
1!
b11 %
1'
b11 +
#528750000000
0!
0'
#528760000000
1!
b100 %
1'
b100 +
#528770000000
0!
0'
#528780000000
1!
b101 %
1'
b101 +
#528790000000
0!
0'
#528800000000
1!
b110 %
1'
b110 +
#528810000000
0!
0'
#528820000000
1!
b111 %
1'
b111 +
#528830000000
0!
0'
#528840000000
1!
0$
b1000 %
1'
0*
b1000 +
#528850000000
0!
0'
#528860000000
1!
b1001 %
1'
b1001 +
#528870000000
0!
0'
#528880000000
1!
b0 %
1'
b0 +
#528890000000
0!
0'
#528900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#528910000000
0!
0'
#528920000000
1!
b10 %
1'
b10 +
#528930000000
0!
0'
#528940000000
1!
b11 %
1'
b11 +
#528950000000
0!
0'
#528960000000
1!
b100 %
1'
b100 +
#528970000000
0!
0'
#528980000000
1!
b101 %
1'
b101 +
#528990000000
0!
0'
#529000000000
1!
0$
b110 %
1'
0*
b110 +
#529010000000
0!
0'
#529020000000
1!
b111 %
1'
b111 +
#529030000000
0!
0'
#529040000000
1!
b1000 %
1'
b1000 +
#529050000000
0!
0'
#529060000000
1!
b1001 %
1'
b1001 +
#529070000000
0!
0'
#529080000000
1!
b0 %
1'
b0 +
#529090000000
0!
0'
#529100000000
1!
1$
b1 %
1'
1*
b1 +
#529110000000
1"
1(
#529120000000
0!
0"
b100 &
0'
0(
b100 ,
#529130000000
1!
b10 %
1'
b10 +
#529140000000
0!
0'
#529150000000
1!
b11 %
1'
b11 +
#529160000000
0!
0'
#529170000000
1!
b100 %
1'
b100 +
#529180000000
0!
0'
#529190000000
1!
b101 %
1'
b101 +
#529200000000
0!
0'
#529210000000
1!
b110 %
1'
b110 +
#529220000000
0!
0'
#529230000000
1!
b111 %
1'
b111 +
#529240000000
0!
0'
#529250000000
1!
0$
b1000 %
1'
0*
b1000 +
#529260000000
0!
0'
#529270000000
1!
b1001 %
1'
b1001 +
#529280000000
0!
0'
#529290000000
1!
b0 %
1'
b0 +
#529300000000
0!
0'
#529310000000
1!
1$
b1 %
1'
1*
b1 +
#529320000000
0!
0'
#529330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#529340000000
0!
0'
#529350000000
1!
b11 %
1'
b11 +
#529360000000
0!
0'
#529370000000
1!
b100 %
1'
b100 +
#529380000000
0!
0'
#529390000000
1!
b101 %
1'
b101 +
#529400000000
0!
0'
#529410000000
1!
0$
b110 %
1'
0*
b110 +
#529420000000
0!
0'
#529430000000
1!
b111 %
1'
b111 +
#529440000000
0!
0'
#529450000000
1!
b1000 %
1'
b1000 +
#529460000000
0!
0'
#529470000000
1!
b1001 %
1'
b1001 +
#529480000000
0!
0'
#529490000000
1!
b0 %
1'
b0 +
#529500000000
0!
0'
#529510000000
1!
1$
b1 %
1'
1*
b1 +
#529520000000
0!
0'
#529530000000
1!
b10 %
1'
b10 +
#529540000000
1"
1(
#529550000000
0!
0"
b100 &
0'
0(
b100 ,
#529560000000
1!
b11 %
1'
b11 +
#529570000000
0!
0'
#529580000000
1!
b100 %
1'
b100 +
#529590000000
0!
0'
#529600000000
1!
b101 %
1'
b101 +
#529610000000
0!
0'
#529620000000
1!
b110 %
1'
b110 +
#529630000000
0!
0'
#529640000000
1!
b111 %
1'
b111 +
#529650000000
0!
0'
#529660000000
1!
0$
b1000 %
1'
0*
b1000 +
#529670000000
0!
0'
#529680000000
1!
b1001 %
1'
b1001 +
#529690000000
0!
0'
#529700000000
1!
b0 %
1'
b0 +
#529710000000
0!
0'
#529720000000
1!
1$
b1 %
1'
1*
b1 +
#529730000000
0!
0'
#529740000000
1!
b10 %
1'
b10 +
#529750000000
0!
0'
#529760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#529770000000
0!
0'
#529780000000
1!
b100 %
1'
b100 +
#529790000000
0!
0'
#529800000000
1!
b101 %
1'
b101 +
#529810000000
0!
0'
#529820000000
1!
0$
b110 %
1'
0*
b110 +
#529830000000
0!
0'
#529840000000
1!
b111 %
1'
b111 +
#529850000000
0!
0'
#529860000000
1!
b1000 %
1'
b1000 +
#529870000000
0!
0'
#529880000000
1!
b1001 %
1'
b1001 +
#529890000000
0!
0'
#529900000000
1!
b0 %
1'
b0 +
#529910000000
0!
0'
#529920000000
1!
1$
b1 %
1'
1*
b1 +
#529930000000
0!
0'
#529940000000
1!
b10 %
1'
b10 +
#529950000000
0!
0'
#529960000000
1!
b11 %
1'
b11 +
#529970000000
1"
1(
#529980000000
0!
0"
b100 &
0'
0(
b100 ,
#529990000000
1!
b100 %
1'
b100 +
#530000000000
0!
0'
#530010000000
1!
b101 %
1'
b101 +
#530020000000
0!
0'
#530030000000
1!
b110 %
1'
b110 +
#530040000000
0!
0'
#530050000000
1!
b111 %
1'
b111 +
#530060000000
0!
0'
#530070000000
1!
0$
b1000 %
1'
0*
b1000 +
#530080000000
0!
0'
#530090000000
1!
b1001 %
1'
b1001 +
#530100000000
0!
0'
#530110000000
1!
b0 %
1'
b0 +
#530120000000
0!
0'
#530130000000
1!
1$
b1 %
1'
1*
b1 +
#530140000000
0!
0'
#530150000000
1!
b10 %
1'
b10 +
#530160000000
0!
0'
#530170000000
1!
b11 %
1'
b11 +
#530180000000
0!
0'
#530190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#530200000000
0!
0'
#530210000000
1!
b101 %
1'
b101 +
#530220000000
0!
0'
#530230000000
1!
0$
b110 %
1'
0*
b110 +
#530240000000
0!
0'
#530250000000
1!
b111 %
1'
b111 +
#530260000000
0!
0'
#530270000000
1!
b1000 %
1'
b1000 +
#530280000000
0!
0'
#530290000000
1!
b1001 %
1'
b1001 +
#530300000000
0!
0'
#530310000000
1!
b0 %
1'
b0 +
#530320000000
0!
0'
#530330000000
1!
1$
b1 %
1'
1*
b1 +
#530340000000
0!
0'
#530350000000
1!
b10 %
1'
b10 +
#530360000000
0!
0'
#530370000000
1!
b11 %
1'
b11 +
#530380000000
0!
0'
#530390000000
1!
b100 %
1'
b100 +
#530400000000
1"
1(
#530410000000
0!
0"
b100 &
0'
0(
b100 ,
#530420000000
1!
b101 %
1'
b101 +
#530430000000
0!
0'
#530440000000
1!
b110 %
1'
b110 +
#530450000000
0!
0'
#530460000000
1!
b111 %
1'
b111 +
#530470000000
0!
0'
#530480000000
1!
0$
b1000 %
1'
0*
b1000 +
#530490000000
0!
0'
#530500000000
1!
b1001 %
1'
b1001 +
#530510000000
0!
0'
#530520000000
1!
b0 %
1'
b0 +
#530530000000
0!
0'
#530540000000
1!
1$
b1 %
1'
1*
b1 +
#530550000000
0!
0'
#530560000000
1!
b10 %
1'
b10 +
#530570000000
0!
0'
#530580000000
1!
b11 %
1'
b11 +
#530590000000
0!
0'
#530600000000
1!
b100 %
1'
b100 +
#530610000000
0!
0'
#530620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#530630000000
0!
0'
#530640000000
1!
0$
b110 %
1'
0*
b110 +
#530650000000
0!
0'
#530660000000
1!
b111 %
1'
b111 +
#530670000000
0!
0'
#530680000000
1!
b1000 %
1'
b1000 +
#530690000000
0!
0'
#530700000000
1!
b1001 %
1'
b1001 +
#530710000000
0!
0'
#530720000000
1!
b0 %
1'
b0 +
#530730000000
0!
0'
#530740000000
1!
1$
b1 %
1'
1*
b1 +
#530750000000
0!
0'
#530760000000
1!
b10 %
1'
b10 +
#530770000000
0!
0'
#530780000000
1!
b11 %
1'
b11 +
#530790000000
0!
0'
#530800000000
1!
b100 %
1'
b100 +
#530810000000
0!
0'
#530820000000
1!
b101 %
1'
b101 +
#530830000000
1"
1(
#530840000000
0!
0"
b100 &
0'
0(
b100 ,
#530850000000
1!
b110 %
1'
b110 +
#530860000000
0!
0'
#530870000000
1!
b111 %
1'
b111 +
#530880000000
0!
0'
#530890000000
1!
0$
b1000 %
1'
0*
b1000 +
#530900000000
0!
0'
#530910000000
1!
b1001 %
1'
b1001 +
#530920000000
0!
0'
#530930000000
1!
b0 %
1'
b0 +
#530940000000
0!
0'
#530950000000
1!
1$
b1 %
1'
1*
b1 +
#530960000000
0!
0'
#530970000000
1!
b10 %
1'
b10 +
#530980000000
0!
0'
#530990000000
1!
b11 %
1'
b11 +
#531000000000
0!
0'
#531010000000
1!
b100 %
1'
b100 +
#531020000000
0!
0'
#531030000000
1!
b101 %
1'
b101 +
#531040000000
0!
0'
#531050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#531060000000
0!
0'
#531070000000
1!
b111 %
1'
b111 +
#531080000000
0!
0'
#531090000000
1!
b1000 %
1'
b1000 +
#531100000000
0!
0'
#531110000000
1!
b1001 %
1'
b1001 +
#531120000000
0!
0'
#531130000000
1!
b0 %
1'
b0 +
#531140000000
0!
0'
#531150000000
1!
1$
b1 %
1'
1*
b1 +
#531160000000
0!
0'
#531170000000
1!
b10 %
1'
b10 +
#531180000000
0!
0'
#531190000000
1!
b11 %
1'
b11 +
#531200000000
0!
0'
#531210000000
1!
b100 %
1'
b100 +
#531220000000
0!
0'
#531230000000
1!
b101 %
1'
b101 +
#531240000000
0!
0'
#531250000000
1!
0$
b110 %
1'
0*
b110 +
#531260000000
1"
1(
#531270000000
0!
0"
b100 &
0'
0(
b100 ,
#531280000000
1!
1$
b111 %
1'
1*
b111 +
#531290000000
0!
0'
#531300000000
1!
0$
b1000 %
1'
0*
b1000 +
#531310000000
0!
0'
#531320000000
1!
b1001 %
1'
b1001 +
#531330000000
0!
0'
#531340000000
1!
b0 %
1'
b0 +
#531350000000
0!
0'
#531360000000
1!
1$
b1 %
1'
1*
b1 +
#531370000000
0!
0'
#531380000000
1!
b10 %
1'
b10 +
#531390000000
0!
0'
#531400000000
1!
b11 %
1'
b11 +
#531410000000
0!
0'
#531420000000
1!
b100 %
1'
b100 +
#531430000000
0!
0'
#531440000000
1!
b101 %
1'
b101 +
#531450000000
0!
0'
#531460000000
1!
b110 %
1'
b110 +
#531470000000
0!
0'
#531480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#531490000000
0!
0'
#531500000000
1!
b1000 %
1'
b1000 +
#531510000000
0!
0'
#531520000000
1!
b1001 %
1'
b1001 +
#531530000000
0!
0'
#531540000000
1!
b0 %
1'
b0 +
#531550000000
0!
0'
#531560000000
1!
1$
b1 %
1'
1*
b1 +
#531570000000
0!
0'
#531580000000
1!
b10 %
1'
b10 +
#531590000000
0!
0'
#531600000000
1!
b11 %
1'
b11 +
#531610000000
0!
0'
#531620000000
1!
b100 %
1'
b100 +
#531630000000
0!
0'
#531640000000
1!
b101 %
1'
b101 +
#531650000000
0!
0'
#531660000000
1!
0$
b110 %
1'
0*
b110 +
#531670000000
0!
0'
#531680000000
1!
b111 %
1'
b111 +
#531690000000
1"
1(
#531700000000
0!
0"
b100 &
0'
0(
b100 ,
#531710000000
1!
b1000 %
1'
b1000 +
#531720000000
0!
0'
#531730000000
1!
b1001 %
1'
b1001 +
#531740000000
0!
0'
#531750000000
1!
b0 %
1'
b0 +
#531760000000
0!
0'
#531770000000
1!
1$
b1 %
1'
1*
b1 +
#531780000000
0!
0'
#531790000000
1!
b10 %
1'
b10 +
#531800000000
0!
0'
#531810000000
1!
b11 %
1'
b11 +
#531820000000
0!
0'
#531830000000
1!
b100 %
1'
b100 +
#531840000000
0!
0'
#531850000000
1!
b101 %
1'
b101 +
#531860000000
0!
0'
#531870000000
1!
b110 %
1'
b110 +
#531880000000
0!
0'
#531890000000
1!
b111 %
1'
b111 +
#531900000000
0!
0'
#531910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#531920000000
0!
0'
#531930000000
1!
b1001 %
1'
b1001 +
#531940000000
0!
0'
#531950000000
1!
b0 %
1'
b0 +
#531960000000
0!
0'
#531970000000
1!
1$
b1 %
1'
1*
b1 +
#531980000000
0!
0'
#531990000000
1!
b10 %
1'
b10 +
#532000000000
0!
0'
#532010000000
1!
b11 %
1'
b11 +
#532020000000
0!
0'
#532030000000
1!
b100 %
1'
b100 +
#532040000000
0!
0'
#532050000000
1!
b101 %
1'
b101 +
#532060000000
0!
0'
#532070000000
1!
0$
b110 %
1'
0*
b110 +
#532080000000
0!
0'
#532090000000
1!
b111 %
1'
b111 +
#532100000000
0!
0'
#532110000000
1!
b1000 %
1'
b1000 +
#532120000000
1"
1(
#532130000000
0!
0"
b100 &
0'
0(
b100 ,
#532140000000
1!
b1001 %
1'
b1001 +
#532150000000
0!
0'
#532160000000
1!
b0 %
1'
b0 +
#532170000000
0!
0'
#532180000000
1!
1$
b1 %
1'
1*
b1 +
#532190000000
0!
0'
#532200000000
1!
b10 %
1'
b10 +
#532210000000
0!
0'
#532220000000
1!
b11 %
1'
b11 +
#532230000000
0!
0'
#532240000000
1!
b100 %
1'
b100 +
#532250000000
0!
0'
#532260000000
1!
b101 %
1'
b101 +
#532270000000
0!
0'
#532280000000
1!
b110 %
1'
b110 +
#532290000000
0!
0'
#532300000000
1!
b111 %
1'
b111 +
#532310000000
0!
0'
#532320000000
1!
0$
b1000 %
1'
0*
b1000 +
#532330000000
0!
0'
#532340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#532350000000
0!
0'
#532360000000
1!
b0 %
1'
b0 +
#532370000000
0!
0'
#532380000000
1!
1$
b1 %
1'
1*
b1 +
#532390000000
0!
0'
#532400000000
1!
b10 %
1'
b10 +
#532410000000
0!
0'
#532420000000
1!
b11 %
1'
b11 +
#532430000000
0!
0'
#532440000000
1!
b100 %
1'
b100 +
#532450000000
0!
0'
#532460000000
1!
b101 %
1'
b101 +
#532470000000
0!
0'
#532480000000
1!
0$
b110 %
1'
0*
b110 +
#532490000000
0!
0'
#532500000000
1!
b111 %
1'
b111 +
#532510000000
0!
0'
#532520000000
1!
b1000 %
1'
b1000 +
#532530000000
0!
0'
#532540000000
1!
b1001 %
1'
b1001 +
#532550000000
1"
1(
#532560000000
0!
0"
b100 &
0'
0(
b100 ,
#532570000000
1!
b0 %
1'
b0 +
#532580000000
0!
0'
#532590000000
1!
1$
b1 %
1'
1*
b1 +
#532600000000
0!
0'
#532610000000
1!
b10 %
1'
b10 +
#532620000000
0!
0'
#532630000000
1!
b11 %
1'
b11 +
#532640000000
0!
0'
#532650000000
1!
b100 %
1'
b100 +
#532660000000
0!
0'
#532670000000
1!
b101 %
1'
b101 +
#532680000000
0!
0'
#532690000000
1!
b110 %
1'
b110 +
#532700000000
0!
0'
#532710000000
1!
b111 %
1'
b111 +
#532720000000
0!
0'
#532730000000
1!
0$
b1000 %
1'
0*
b1000 +
#532740000000
0!
0'
#532750000000
1!
b1001 %
1'
b1001 +
#532760000000
0!
0'
#532770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#532780000000
0!
0'
#532790000000
1!
1$
b1 %
1'
1*
b1 +
#532800000000
0!
0'
#532810000000
1!
b10 %
1'
b10 +
#532820000000
0!
0'
#532830000000
1!
b11 %
1'
b11 +
#532840000000
0!
0'
#532850000000
1!
b100 %
1'
b100 +
#532860000000
0!
0'
#532870000000
1!
b101 %
1'
b101 +
#532880000000
0!
0'
#532890000000
1!
0$
b110 %
1'
0*
b110 +
#532900000000
0!
0'
#532910000000
1!
b111 %
1'
b111 +
#532920000000
0!
0'
#532930000000
1!
b1000 %
1'
b1000 +
#532940000000
0!
0'
#532950000000
1!
b1001 %
1'
b1001 +
#532960000000
0!
0'
#532970000000
1!
b0 %
1'
b0 +
#532980000000
1"
1(
#532990000000
0!
0"
b100 &
0'
0(
b100 ,
#533000000000
1!
1$
b1 %
1'
1*
b1 +
#533010000000
0!
0'
#533020000000
1!
b10 %
1'
b10 +
#533030000000
0!
0'
#533040000000
1!
b11 %
1'
b11 +
#533050000000
0!
0'
#533060000000
1!
b100 %
1'
b100 +
#533070000000
0!
0'
#533080000000
1!
b101 %
1'
b101 +
#533090000000
0!
0'
#533100000000
1!
b110 %
1'
b110 +
#533110000000
0!
0'
#533120000000
1!
b111 %
1'
b111 +
#533130000000
0!
0'
#533140000000
1!
0$
b1000 %
1'
0*
b1000 +
#533150000000
0!
0'
#533160000000
1!
b1001 %
1'
b1001 +
#533170000000
0!
0'
#533180000000
1!
b0 %
1'
b0 +
#533190000000
0!
0'
#533200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#533210000000
0!
0'
#533220000000
1!
b10 %
1'
b10 +
#533230000000
0!
0'
#533240000000
1!
b11 %
1'
b11 +
#533250000000
0!
0'
#533260000000
1!
b100 %
1'
b100 +
#533270000000
0!
0'
#533280000000
1!
b101 %
1'
b101 +
#533290000000
0!
0'
#533300000000
1!
0$
b110 %
1'
0*
b110 +
#533310000000
0!
0'
#533320000000
1!
b111 %
1'
b111 +
#533330000000
0!
0'
#533340000000
1!
b1000 %
1'
b1000 +
#533350000000
0!
0'
#533360000000
1!
b1001 %
1'
b1001 +
#533370000000
0!
0'
#533380000000
1!
b0 %
1'
b0 +
#533390000000
0!
0'
#533400000000
1!
1$
b1 %
1'
1*
b1 +
#533410000000
1"
1(
#533420000000
0!
0"
b100 &
0'
0(
b100 ,
#533430000000
1!
b10 %
1'
b10 +
#533440000000
0!
0'
#533450000000
1!
b11 %
1'
b11 +
#533460000000
0!
0'
#533470000000
1!
b100 %
1'
b100 +
#533480000000
0!
0'
#533490000000
1!
b101 %
1'
b101 +
#533500000000
0!
0'
#533510000000
1!
b110 %
1'
b110 +
#533520000000
0!
0'
#533530000000
1!
b111 %
1'
b111 +
#533540000000
0!
0'
#533550000000
1!
0$
b1000 %
1'
0*
b1000 +
#533560000000
0!
0'
#533570000000
1!
b1001 %
1'
b1001 +
#533580000000
0!
0'
#533590000000
1!
b0 %
1'
b0 +
#533600000000
0!
0'
#533610000000
1!
1$
b1 %
1'
1*
b1 +
#533620000000
0!
0'
#533630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#533640000000
0!
0'
#533650000000
1!
b11 %
1'
b11 +
#533660000000
0!
0'
#533670000000
1!
b100 %
1'
b100 +
#533680000000
0!
0'
#533690000000
1!
b101 %
1'
b101 +
#533700000000
0!
0'
#533710000000
1!
0$
b110 %
1'
0*
b110 +
#533720000000
0!
0'
#533730000000
1!
b111 %
1'
b111 +
#533740000000
0!
0'
#533750000000
1!
b1000 %
1'
b1000 +
#533760000000
0!
0'
#533770000000
1!
b1001 %
1'
b1001 +
#533780000000
0!
0'
#533790000000
1!
b0 %
1'
b0 +
#533800000000
0!
0'
#533810000000
1!
1$
b1 %
1'
1*
b1 +
#533820000000
0!
0'
#533830000000
1!
b10 %
1'
b10 +
#533840000000
1"
1(
#533850000000
0!
0"
b100 &
0'
0(
b100 ,
#533860000000
1!
b11 %
1'
b11 +
#533870000000
0!
0'
#533880000000
1!
b100 %
1'
b100 +
#533890000000
0!
0'
#533900000000
1!
b101 %
1'
b101 +
#533910000000
0!
0'
#533920000000
1!
b110 %
1'
b110 +
#533930000000
0!
0'
#533940000000
1!
b111 %
1'
b111 +
#533950000000
0!
0'
#533960000000
1!
0$
b1000 %
1'
0*
b1000 +
#533970000000
0!
0'
#533980000000
1!
b1001 %
1'
b1001 +
#533990000000
0!
0'
#534000000000
1!
b0 %
1'
b0 +
#534010000000
0!
0'
#534020000000
1!
1$
b1 %
1'
1*
b1 +
#534030000000
0!
0'
#534040000000
1!
b10 %
1'
b10 +
#534050000000
0!
0'
#534060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#534070000000
0!
0'
#534080000000
1!
b100 %
1'
b100 +
#534090000000
0!
0'
#534100000000
1!
b101 %
1'
b101 +
#534110000000
0!
0'
#534120000000
1!
0$
b110 %
1'
0*
b110 +
#534130000000
0!
0'
#534140000000
1!
b111 %
1'
b111 +
#534150000000
0!
0'
#534160000000
1!
b1000 %
1'
b1000 +
#534170000000
0!
0'
#534180000000
1!
b1001 %
1'
b1001 +
#534190000000
0!
0'
#534200000000
1!
b0 %
1'
b0 +
#534210000000
0!
0'
#534220000000
1!
1$
b1 %
1'
1*
b1 +
#534230000000
0!
0'
#534240000000
1!
b10 %
1'
b10 +
#534250000000
0!
0'
#534260000000
1!
b11 %
1'
b11 +
#534270000000
1"
1(
#534280000000
0!
0"
b100 &
0'
0(
b100 ,
#534290000000
1!
b100 %
1'
b100 +
#534300000000
0!
0'
#534310000000
1!
b101 %
1'
b101 +
#534320000000
0!
0'
#534330000000
1!
b110 %
1'
b110 +
#534340000000
0!
0'
#534350000000
1!
b111 %
1'
b111 +
#534360000000
0!
0'
#534370000000
1!
0$
b1000 %
1'
0*
b1000 +
#534380000000
0!
0'
#534390000000
1!
b1001 %
1'
b1001 +
#534400000000
0!
0'
#534410000000
1!
b0 %
1'
b0 +
#534420000000
0!
0'
#534430000000
1!
1$
b1 %
1'
1*
b1 +
#534440000000
0!
0'
#534450000000
1!
b10 %
1'
b10 +
#534460000000
0!
0'
#534470000000
1!
b11 %
1'
b11 +
#534480000000
0!
0'
#534490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#534500000000
0!
0'
#534510000000
1!
b101 %
1'
b101 +
#534520000000
0!
0'
#534530000000
1!
0$
b110 %
1'
0*
b110 +
#534540000000
0!
0'
#534550000000
1!
b111 %
1'
b111 +
#534560000000
0!
0'
#534570000000
1!
b1000 %
1'
b1000 +
#534580000000
0!
0'
#534590000000
1!
b1001 %
1'
b1001 +
#534600000000
0!
0'
#534610000000
1!
b0 %
1'
b0 +
#534620000000
0!
0'
#534630000000
1!
1$
b1 %
1'
1*
b1 +
#534640000000
0!
0'
#534650000000
1!
b10 %
1'
b10 +
#534660000000
0!
0'
#534670000000
1!
b11 %
1'
b11 +
#534680000000
0!
0'
#534690000000
1!
b100 %
1'
b100 +
#534700000000
1"
1(
#534710000000
0!
0"
b100 &
0'
0(
b100 ,
#534720000000
1!
b101 %
1'
b101 +
#534730000000
0!
0'
#534740000000
1!
b110 %
1'
b110 +
#534750000000
0!
0'
#534760000000
1!
b111 %
1'
b111 +
#534770000000
0!
0'
#534780000000
1!
0$
b1000 %
1'
0*
b1000 +
#534790000000
0!
0'
#534800000000
1!
b1001 %
1'
b1001 +
#534810000000
0!
0'
#534820000000
1!
b0 %
1'
b0 +
#534830000000
0!
0'
#534840000000
1!
1$
b1 %
1'
1*
b1 +
#534850000000
0!
0'
#534860000000
1!
b10 %
1'
b10 +
#534870000000
0!
0'
#534880000000
1!
b11 %
1'
b11 +
#534890000000
0!
0'
#534900000000
1!
b100 %
1'
b100 +
#534910000000
0!
0'
#534920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#534930000000
0!
0'
#534940000000
1!
0$
b110 %
1'
0*
b110 +
#534950000000
0!
0'
#534960000000
1!
b111 %
1'
b111 +
#534970000000
0!
0'
#534980000000
1!
b1000 %
1'
b1000 +
#534990000000
0!
0'
#535000000000
1!
b1001 %
1'
b1001 +
#535010000000
0!
0'
#535020000000
1!
b0 %
1'
b0 +
#535030000000
0!
0'
#535040000000
1!
1$
b1 %
1'
1*
b1 +
#535050000000
0!
0'
#535060000000
1!
b10 %
1'
b10 +
#535070000000
0!
0'
#535080000000
1!
b11 %
1'
b11 +
#535090000000
0!
0'
#535100000000
1!
b100 %
1'
b100 +
#535110000000
0!
0'
#535120000000
1!
b101 %
1'
b101 +
#535130000000
1"
1(
#535140000000
0!
0"
b100 &
0'
0(
b100 ,
#535150000000
1!
b110 %
1'
b110 +
#535160000000
0!
0'
#535170000000
1!
b111 %
1'
b111 +
#535180000000
0!
0'
#535190000000
1!
0$
b1000 %
1'
0*
b1000 +
#535200000000
0!
0'
#535210000000
1!
b1001 %
1'
b1001 +
#535220000000
0!
0'
#535230000000
1!
b0 %
1'
b0 +
#535240000000
0!
0'
#535250000000
1!
1$
b1 %
1'
1*
b1 +
#535260000000
0!
0'
#535270000000
1!
b10 %
1'
b10 +
#535280000000
0!
0'
#535290000000
1!
b11 %
1'
b11 +
#535300000000
0!
0'
#535310000000
1!
b100 %
1'
b100 +
#535320000000
0!
0'
#535330000000
1!
b101 %
1'
b101 +
#535340000000
0!
0'
#535350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#535360000000
0!
0'
#535370000000
1!
b111 %
1'
b111 +
#535380000000
0!
0'
#535390000000
1!
b1000 %
1'
b1000 +
#535400000000
0!
0'
#535410000000
1!
b1001 %
1'
b1001 +
#535420000000
0!
0'
#535430000000
1!
b0 %
1'
b0 +
#535440000000
0!
0'
#535450000000
1!
1$
b1 %
1'
1*
b1 +
#535460000000
0!
0'
#535470000000
1!
b10 %
1'
b10 +
#535480000000
0!
0'
#535490000000
1!
b11 %
1'
b11 +
#535500000000
0!
0'
#535510000000
1!
b100 %
1'
b100 +
#535520000000
0!
0'
#535530000000
1!
b101 %
1'
b101 +
#535540000000
0!
0'
#535550000000
1!
0$
b110 %
1'
0*
b110 +
#535560000000
1"
1(
#535570000000
0!
0"
b100 &
0'
0(
b100 ,
#535580000000
1!
1$
b111 %
1'
1*
b111 +
#535590000000
0!
0'
#535600000000
1!
0$
b1000 %
1'
0*
b1000 +
#535610000000
0!
0'
#535620000000
1!
b1001 %
1'
b1001 +
#535630000000
0!
0'
#535640000000
1!
b0 %
1'
b0 +
#535650000000
0!
0'
#535660000000
1!
1$
b1 %
1'
1*
b1 +
#535670000000
0!
0'
#535680000000
1!
b10 %
1'
b10 +
#535690000000
0!
0'
#535700000000
1!
b11 %
1'
b11 +
#535710000000
0!
0'
#535720000000
1!
b100 %
1'
b100 +
#535730000000
0!
0'
#535740000000
1!
b101 %
1'
b101 +
#535750000000
0!
0'
#535760000000
1!
b110 %
1'
b110 +
#535770000000
0!
0'
#535780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#535790000000
0!
0'
#535800000000
1!
b1000 %
1'
b1000 +
#535810000000
0!
0'
#535820000000
1!
b1001 %
1'
b1001 +
#535830000000
0!
0'
#535840000000
1!
b0 %
1'
b0 +
#535850000000
0!
0'
#535860000000
1!
1$
b1 %
1'
1*
b1 +
#535870000000
0!
0'
#535880000000
1!
b10 %
1'
b10 +
#535890000000
0!
0'
#535900000000
1!
b11 %
1'
b11 +
#535910000000
0!
0'
#535920000000
1!
b100 %
1'
b100 +
#535930000000
0!
0'
#535940000000
1!
b101 %
1'
b101 +
#535950000000
0!
0'
#535960000000
1!
0$
b110 %
1'
0*
b110 +
#535970000000
0!
0'
#535980000000
1!
b111 %
1'
b111 +
#535990000000
1"
1(
#536000000000
0!
0"
b100 &
0'
0(
b100 ,
#536010000000
1!
b1000 %
1'
b1000 +
#536020000000
0!
0'
#536030000000
1!
b1001 %
1'
b1001 +
#536040000000
0!
0'
#536050000000
1!
b0 %
1'
b0 +
#536060000000
0!
0'
#536070000000
1!
1$
b1 %
1'
1*
b1 +
#536080000000
0!
0'
#536090000000
1!
b10 %
1'
b10 +
#536100000000
0!
0'
#536110000000
1!
b11 %
1'
b11 +
#536120000000
0!
0'
#536130000000
1!
b100 %
1'
b100 +
#536140000000
0!
0'
#536150000000
1!
b101 %
1'
b101 +
#536160000000
0!
0'
#536170000000
1!
b110 %
1'
b110 +
#536180000000
0!
0'
#536190000000
1!
b111 %
1'
b111 +
#536200000000
0!
0'
#536210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#536220000000
0!
0'
#536230000000
1!
b1001 %
1'
b1001 +
#536240000000
0!
0'
#536250000000
1!
b0 %
1'
b0 +
#536260000000
0!
0'
#536270000000
1!
1$
b1 %
1'
1*
b1 +
#536280000000
0!
0'
#536290000000
1!
b10 %
1'
b10 +
#536300000000
0!
0'
#536310000000
1!
b11 %
1'
b11 +
#536320000000
0!
0'
#536330000000
1!
b100 %
1'
b100 +
#536340000000
0!
0'
#536350000000
1!
b101 %
1'
b101 +
#536360000000
0!
0'
#536370000000
1!
0$
b110 %
1'
0*
b110 +
#536380000000
0!
0'
#536390000000
1!
b111 %
1'
b111 +
#536400000000
0!
0'
#536410000000
1!
b1000 %
1'
b1000 +
#536420000000
1"
1(
#536430000000
0!
0"
b100 &
0'
0(
b100 ,
#536440000000
1!
b1001 %
1'
b1001 +
#536450000000
0!
0'
#536460000000
1!
b0 %
1'
b0 +
#536470000000
0!
0'
#536480000000
1!
1$
b1 %
1'
1*
b1 +
#536490000000
0!
0'
#536500000000
1!
b10 %
1'
b10 +
#536510000000
0!
0'
#536520000000
1!
b11 %
1'
b11 +
#536530000000
0!
0'
#536540000000
1!
b100 %
1'
b100 +
#536550000000
0!
0'
#536560000000
1!
b101 %
1'
b101 +
#536570000000
0!
0'
#536580000000
1!
b110 %
1'
b110 +
#536590000000
0!
0'
#536600000000
1!
b111 %
1'
b111 +
#536610000000
0!
0'
#536620000000
1!
0$
b1000 %
1'
0*
b1000 +
#536630000000
0!
0'
#536640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#536650000000
0!
0'
#536660000000
1!
b0 %
1'
b0 +
#536670000000
0!
0'
#536680000000
1!
1$
b1 %
1'
1*
b1 +
#536690000000
0!
0'
#536700000000
1!
b10 %
1'
b10 +
#536710000000
0!
0'
#536720000000
1!
b11 %
1'
b11 +
#536730000000
0!
0'
#536740000000
1!
b100 %
1'
b100 +
#536750000000
0!
0'
#536760000000
1!
b101 %
1'
b101 +
#536770000000
0!
0'
#536780000000
1!
0$
b110 %
1'
0*
b110 +
#536790000000
0!
0'
#536800000000
1!
b111 %
1'
b111 +
#536810000000
0!
0'
#536820000000
1!
b1000 %
1'
b1000 +
#536830000000
0!
0'
#536840000000
1!
b1001 %
1'
b1001 +
#536850000000
1"
1(
#536860000000
0!
0"
b100 &
0'
0(
b100 ,
#536870000000
1!
b0 %
1'
b0 +
#536880000000
0!
0'
#536890000000
1!
1$
b1 %
1'
1*
b1 +
#536900000000
0!
0'
#536910000000
1!
b10 %
1'
b10 +
#536920000000
0!
0'
#536930000000
1!
b11 %
1'
b11 +
#536940000000
0!
0'
#536950000000
1!
b100 %
1'
b100 +
#536960000000
0!
0'
#536970000000
1!
b101 %
1'
b101 +
#536980000000
0!
0'
#536990000000
1!
b110 %
1'
b110 +
#537000000000
0!
0'
#537010000000
1!
b111 %
1'
b111 +
#537020000000
0!
0'
#537030000000
1!
0$
b1000 %
1'
0*
b1000 +
#537040000000
0!
0'
#537050000000
1!
b1001 %
1'
b1001 +
#537060000000
0!
0'
#537070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#537080000000
0!
0'
#537090000000
1!
1$
b1 %
1'
1*
b1 +
#537100000000
0!
0'
#537110000000
1!
b10 %
1'
b10 +
#537120000000
0!
0'
#537130000000
1!
b11 %
1'
b11 +
#537140000000
0!
0'
#537150000000
1!
b100 %
1'
b100 +
#537160000000
0!
0'
#537170000000
1!
b101 %
1'
b101 +
#537180000000
0!
0'
#537190000000
1!
0$
b110 %
1'
0*
b110 +
#537200000000
0!
0'
#537210000000
1!
b111 %
1'
b111 +
#537220000000
0!
0'
#537230000000
1!
b1000 %
1'
b1000 +
#537240000000
0!
0'
#537250000000
1!
b1001 %
1'
b1001 +
#537260000000
0!
0'
#537270000000
1!
b0 %
1'
b0 +
#537280000000
1"
1(
#537290000000
0!
0"
b100 &
0'
0(
b100 ,
#537300000000
1!
1$
b1 %
1'
1*
b1 +
#537310000000
0!
0'
#537320000000
1!
b10 %
1'
b10 +
#537330000000
0!
0'
#537340000000
1!
b11 %
1'
b11 +
#537350000000
0!
0'
#537360000000
1!
b100 %
1'
b100 +
#537370000000
0!
0'
#537380000000
1!
b101 %
1'
b101 +
#537390000000
0!
0'
#537400000000
1!
b110 %
1'
b110 +
#537410000000
0!
0'
#537420000000
1!
b111 %
1'
b111 +
#537430000000
0!
0'
#537440000000
1!
0$
b1000 %
1'
0*
b1000 +
#537450000000
0!
0'
#537460000000
1!
b1001 %
1'
b1001 +
#537470000000
0!
0'
#537480000000
1!
b0 %
1'
b0 +
#537490000000
0!
0'
#537500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#537510000000
0!
0'
#537520000000
1!
b10 %
1'
b10 +
#537530000000
0!
0'
#537540000000
1!
b11 %
1'
b11 +
#537550000000
0!
0'
#537560000000
1!
b100 %
1'
b100 +
#537570000000
0!
0'
#537580000000
1!
b101 %
1'
b101 +
#537590000000
0!
0'
#537600000000
1!
0$
b110 %
1'
0*
b110 +
#537610000000
0!
0'
#537620000000
1!
b111 %
1'
b111 +
#537630000000
0!
0'
#537640000000
1!
b1000 %
1'
b1000 +
#537650000000
0!
0'
#537660000000
1!
b1001 %
1'
b1001 +
#537670000000
0!
0'
#537680000000
1!
b0 %
1'
b0 +
#537690000000
0!
0'
#537700000000
1!
1$
b1 %
1'
1*
b1 +
#537710000000
1"
1(
#537720000000
0!
0"
b100 &
0'
0(
b100 ,
#537730000000
1!
b10 %
1'
b10 +
#537740000000
0!
0'
#537750000000
1!
b11 %
1'
b11 +
#537760000000
0!
0'
#537770000000
1!
b100 %
1'
b100 +
#537780000000
0!
0'
#537790000000
1!
b101 %
1'
b101 +
#537800000000
0!
0'
#537810000000
1!
b110 %
1'
b110 +
#537820000000
0!
0'
#537830000000
1!
b111 %
1'
b111 +
#537840000000
0!
0'
#537850000000
1!
0$
b1000 %
1'
0*
b1000 +
#537860000000
0!
0'
#537870000000
1!
b1001 %
1'
b1001 +
#537880000000
0!
0'
#537890000000
1!
b0 %
1'
b0 +
#537900000000
0!
0'
#537910000000
1!
1$
b1 %
1'
1*
b1 +
#537920000000
0!
0'
#537930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#537940000000
0!
0'
#537950000000
1!
b11 %
1'
b11 +
#537960000000
0!
0'
#537970000000
1!
b100 %
1'
b100 +
#537980000000
0!
0'
#537990000000
1!
b101 %
1'
b101 +
#538000000000
0!
0'
#538010000000
1!
0$
b110 %
1'
0*
b110 +
#538020000000
0!
0'
#538030000000
1!
b111 %
1'
b111 +
#538040000000
0!
0'
#538050000000
1!
b1000 %
1'
b1000 +
#538060000000
0!
0'
#538070000000
1!
b1001 %
1'
b1001 +
#538080000000
0!
0'
#538090000000
1!
b0 %
1'
b0 +
#538100000000
0!
0'
#538110000000
1!
1$
b1 %
1'
1*
b1 +
#538120000000
0!
0'
#538130000000
1!
b10 %
1'
b10 +
#538140000000
1"
1(
#538150000000
0!
0"
b100 &
0'
0(
b100 ,
#538160000000
1!
b11 %
1'
b11 +
#538170000000
0!
0'
#538180000000
1!
b100 %
1'
b100 +
#538190000000
0!
0'
#538200000000
1!
b101 %
1'
b101 +
#538210000000
0!
0'
#538220000000
1!
b110 %
1'
b110 +
#538230000000
0!
0'
#538240000000
1!
b111 %
1'
b111 +
#538250000000
0!
0'
#538260000000
1!
0$
b1000 %
1'
0*
b1000 +
#538270000000
0!
0'
#538280000000
1!
b1001 %
1'
b1001 +
#538290000000
0!
0'
#538300000000
1!
b0 %
1'
b0 +
#538310000000
0!
0'
#538320000000
1!
1$
b1 %
1'
1*
b1 +
#538330000000
0!
0'
#538340000000
1!
b10 %
1'
b10 +
#538350000000
0!
0'
#538360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#538370000000
0!
0'
#538380000000
1!
b100 %
1'
b100 +
#538390000000
0!
0'
#538400000000
1!
b101 %
1'
b101 +
#538410000000
0!
0'
#538420000000
1!
0$
b110 %
1'
0*
b110 +
#538430000000
0!
0'
#538440000000
1!
b111 %
1'
b111 +
#538450000000
0!
0'
#538460000000
1!
b1000 %
1'
b1000 +
#538470000000
0!
0'
#538480000000
1!
b1001 %
1'
b1001 +
#538490000000
0!
0'
#538500000000
1!
b0 %
1'
b0 +
#538510000000
0!
0'
#538520000000
1!
1$
b1 %
1'
1*
b1 +
#538530000000
0!
0'
#538540000000
1!
b10 %
1'
b10 +
#538550000000
0!
0'
#538560000000
1!
b11 %
1'
b11 +
#538570000000
1"
1(
#538580000000
0!
0"
b100 &
0'
0(
b100 ,
#538590000000
1!
b100 %
1'
b100 +
#538600000000
0!
0'
#538610000000
1!
b101 %
1'
b101 +
#538620000000
0!
0'
#538630000000
1!
b110 %
1'
b110 +
#538640000000
0!
0'
#538650000000
1!
b111 %
1'
b111 +
#538660000000
0!
0'
#538670000000
1!
0$
b1000 %
1'
0*
b1000 +
#538680000000
0!
0'
#538690000000
1!
b1001 %
1'
b1001 +
#538700000000
0!
0'
#538710000000
1!
b0 %
1'
b0 +
#538720000000
0!
0'
#538730000000
1!
1$
b1 %
1'
1*
b1 +
#538740000000
0!
0'
#538750000000
1!
b10 %
1'
b10 +
#538760000000
0!
0'
#538770000000
1!
b11 %
1'
b11 +
#538780000000
0!
0'
#538790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#538800000000
0!
0'
#538810000000
1!
b101 %
1'
b101 +
#538820000000
0!
0'
#538830000000
1!
0$
b110 %
1'
0*
b110 +
#538840000000
0!
0'
#538850000000
1!
b111 %
1'
b111 +
#538860000000
0!
0'
#538870000000
1!
b1000 %
1'
b1000 +
#538880000000
0!
0'
#538890000000
1!
b1001 %
1'
b1001 +
#538900000000
0!
0'
#538910000000
1!
b0 %
1'
b0 +
#538920000000
0!
0'
#538930000000
1!
1$
b1 %
1'
1*
b1 +
#538940000000
0!
0'
#538950000000
1!
b10 %
1'
b10 +
#538960000000
0!
0'
#538970000000
1!
b11 %
1'
b11 +
#538980000000
0!
0'
#538990000000
1!
b100 %
1'
b100 +
#539000000000
1"
1(
#539010000000
0!
0"
b100 &
0'
0(
b100 ,
#539020000000
1!
b101 %
1'
b101 +
#539030000000
0!
0'
#539040000000
1!
b110 %
1'
b110 +
#539050000000
0!
0'
#539060000000
1!
b111 %
1'
b111 +
#539070000000
0!
0'
#539080000000
1!
0$
b1000 %
1'
0*
b1000 +
#539090000000
0!
0'
#539100000000
1!
b1001 %
1'
b1001 +
#539110000000
0!
0'
#539120000000
1!
b0 %
1'
b0 +
#539130000000
0!
0'
#539140000000
1!
1$
b1 %
1'
1*
b1 +
#539150000000
0!
0'
#539160000000
1!
b10 %
1'
b10 +
#539170000000
0!
0'
#539180000000
1!
b11 %
1'
b11 +
#539190000000
0!
0'
#539200000000
1!
b100 %
1'
b100 +
#539210000000
0!
0'
#539220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#539230000000
0!
0'
#539240000000
1!
0$
b110 %
1'
0*
b110 +
#539250000000
0!
0'
#539260000000
1!
b111 %
1'
b111 +
#539270000000
0!
0'
#539280000000
1!
b1000 %
1'
b1000 +
#539290000000
0!
0'
#539300000000
1!
b1001 %
1'
b1001 +
#539310000000
0!
0'
#539320000000
1!
b0 %
1'
b0 +
#539330000000
0!
0'
#539340000000
1!
1$
b1 %
1'
1*
b1 +
#539350000000
0!
0'
#539360000000
1!
b10 %
1'
b10 +
#539370000000
0!
0'
#539380000000
1!
b11 %
1'
b11 +
#539390000000
0!
0'
#539400000000
1!
b100 %
1'
b100 +
#539410000000
0!
0'
#539420000000
1!
b101 %
1'
b101 +
#539430000000
1"
1(
#539440000000
0!
0"
b100 &
0'
0(
b100 ,
#539450000000
1!
b110 %
1'
b110 +
#539460000000
0!
0'
#539470000000
1!
b111 %
1'
b111 +
#539480000000
0!
0'
#539490000000
1!
0$
b1000 %
1'
0*
b1000 +
#539500000000
0!
0'
#539510000000
1!
b1001 %
1'
b1001 +
#539520000000
0!
0'
#539530000000
1!
b0 %
1'
b0 +
#539540000000
0!
0'
#539550000000
1!
1$
b1 %
1'
1*
b1 +
#539560000000
0!
0'
#539570000000
1!
b10 %
1'
b10 +
#539580000000
0!
0'
#539590000000
1!
b11 %
1'
b11 +
#539600000000
0!
0'
#539610000000
1!
b100 %
1'
b100 +
#539620000000
0!
0'
#539630000000
1!
b101 %
1'
b101 +
#539640000000
0!
0'
#539650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#539660000000
0!
0'
#539670000000
1!
b111 %
1'
b111 +
#539680000000
0!
0'
#539690000000
1!
b1000 %
1'
b1000 +
#539700000000
0!
0'
#539710000000
1!
b1001 %
1'
b1001 +
#539720000000
0!
0'
#539730000000
1!
b0 %
1'
b0 +
#539740000000
0!
0'
#539750000000
1!
1$
b1 %
1'
1*
b1 +
#539760000000
0!
0'
#539770000000
1!
b10 %
1'
b10 +
#539780000000
0!
0'
#539790000000
1!
b11 %
1'
b11 +
#539800000000
0!
0'
#539810000000
1!
b100 %
1'
b100 +
#539820000000
0!
0'
#539830000000
1!
b101 %
1'
b101 +
#539840000000
0!
0'
#539850000000
1!
0$
b110 %
1'
0*
b110 +
#539860000000
1"
1(
#539870000000
0!
0"
b100 &
0'
0(
b100 ,
#539880000000
1!
1$
b111 %
1'
1*
b111 +
#539890000000
0!
0'
#539900000000
1!
0$
b1000 %
1'
0*
b1000 +
#539910000000
0!
0'
#539920000000
1!
b1001 %
1'
b1001 +
#539930000000
0!
0'
#539940000000
1!
b0 %
1'
b0 +
#539950000000
0!
0'
#539960000000
1!
1$
b1 %
1'
1*
b1 +
#539970000000
0!
0'
#539980000000
1!
b10 %
1'
b10 +
#539990000000
0!
0'
#540000000000
1!
b11 %
1'
b11 +
#540010000000
0!
0'
#540020000000
1!
b100 %
1'
b100 +
#540030000000
0!
0'
#540040000000
1!
b101 %
1'
b101 +
#540050000000
0!
0'
#540060000000
1!
b110 %
1'
b110 +
#540070000000
0!
0'
#540080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#540090000000
0!
0'
#540100000000
1!
b1000 %
1'
b1000 +
#540110000000
0!
0'
#540120000000
1!
b1001 %
1'
b1001 +
#540130000000
0!
0'
#540140000000
1!
b0 %
1'
b0 +
#540150000000
0!
0'
#540160000000
1!
1$
b1 %
1'
1*
b1 +
#540170000000
0!
0'
#540180000000
1!
b10 %
1'
b10 +
#540190000000
0!
0'
#540200000000
1!
b11 %
1'
b11 +
#540210000000
0!
0'
#540220000000
1!
b100 %
1'
b100 +
#540230000000
0!
0'
#540240000000
1!
b101 %
1'
b101 +
#540250000000
0!
0'
#540260000000
1!
0$
b110 %
1'
0*
b110 +
#540270000000
0!
0'
#540280000000
1!
b111 %
1'
b111 +
#540290000000
1"
1(
#540300000000
0!
0"
b100 &
0'
0(
b100 ,
#540310000000
1!
b1000 %
1'
b1000 +
#540320000000
0!
0'
#540330000000
1!
b1001 %
1'
b1001 +
#540340000000
0!
0'
#540350000000
1!
b0 %
1'
b0 +
#540360000000
0!
0'
#540370000000
1!
1$
b1 %
1'
1*
b1 +
#540380000000
0!
0'
#540390000000
1!
b10 %
1'
b10 +
#540400000000
0!
0'
#540410000000
1!
b11 %
1'
b11 +
#540420000000
0!
0'
#540430000000
1!
b100 %
1'
b100 +
#540440000000
0!
0'
#540450000000
1!
b101 %
1'
b101 +
#540460000000
0!
0'
#540470000000
1!
b110 %
1'
b110 +
#540480000000
0!
0'
#540490000000
1!
b111 %
1'
b111 +
#540500000000
0!
0'
#540510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#540520000000
0!
0'
#540530000000
1!
b1001 %
1'
b1001 +
#540540000000
0!
0'
#540550000000
1!
b0 %
1'
b0 +
#540560000000
0!
0'
#540570000000
1!
1$
b1 %
1'
1*
b1 +
#540580000000
0!
0'
#540590000000
1!
b10 %
1'
b10 +
#540600000000
0!
0'
#540610000000
1!
b11 %
1'
b11 +
#540620000000
0!
0'
#540630000000
1!
b100 %
1'
b100 +
#540640000000
0!
0'
#540650000000
1!
b101 %
1'
b101 +
#540660000000
0!
0'
#540670000000
1!
0$
b110 %
1'
0*
b110 +
#540680000000
0!
0'
#540690000000
1!
b111 %
1'
b111 +
#540700000000
0!
0'
#540710000000
1!
b1000 %
1'
b1000 +
#540720000000
1"
1(
#540730000000
0!
0"
b100 &
0'
0(
b100 ,
#540740000000
1!
b1001 %
1'
b1001 +
#540750000000
0!
0'
#540760000000
1!
b0 %
1'
b0 +
#540770000000
0!
0'
#540780000000
1!
1$
b1 %
1'
1*
b1 +
#540790000000
0!
0'
#540800000000
1!
b10 %
1'
b10 +
#540810000000
0!
0'
#540820000000
1!
b11 %
1'
b11 +
#540830000000
0!
0'
#540840000000
1!
b100 %
1'
b100 +
#540850000000
0!
0'
#540860000000
1!
b101 %
1'
b101 +
#540870000000
0!
0'
#540880000000
1!
b110 %
1'
b110 +
#540890000000
0!
0'
#540900000000
1!
b111 %
1'
b111 +
#540910000000
0!
0'
#540920000000
1!
0$
b1000 %
1'
0*
b1000 +
#540930000000
0!
0'
#540940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#540950000000
0!
0'
#540960000000
1!
b0 %
1'
b0 +
#540970000000
0!
0'
#540980000000
1!
1$
b1 %
1'
1*
b1 +
#540990000000
0!
0'
#541000000000
1!
b10 %
1'
b10 +
#541010000000
0!
0'
#541020000000
1!
b11 %
1'
b11 +
#541030000000
0!
0'
#541040000000
1!
b100 %
1'
b100 +
#541050000000
0!
0'
#541060000000
1!
b101 %
1'
b101 +
#541070000000
0!
0'
#541080000000
1!
0$
b110 %
1'
0*
b110 +
#541090000000
0!
0'
#541100000000
1!
b111 %
1'
b111 +
#541110000000
0!
0'
#541120000000
1!
b1000 %
1'
b1000 +
#541130000000
0!
0'
#541140000000
1!
b1001 %
1'
b1001 +
#541150000000
1"
1(
#541160000000
0!
0"
b100 &
0'
0(
b100 ,
#541170000000
1!
b0 %
1'
b0 +
#541180000000
0!
0'
#541190000000
1!
1$
b1 %
1'
1*
b1 +
#541200000000
0!
0'
#541210000000
1!
b10 %
1'
b10 +
#541220000000
0!
0'
#541230000000
1!
b11 %
1'
b11 +
#541240000000
0!
0'
#541250000000
1!
b100 %
1'
b100 +
#541260000000
0!
0'
#541270000000
1!
b101 %
1'
b101 +
#541280000000
0!
0'
#541290000000
1!
b110 %
1'
b110 +
#541300000000
0!
0'
#541310000000
1!
b111 %
1'
b111 +
#541320000000
0!
0'
#541330000000
1!
0$
b1000 %
1'
0*
b1000 +
#541340000000
0!
0'
#541350000000
1!
b1001 %
1'
b1001 +
#541360000000
0!
0'
#541370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#541380000000
0!
0'
#541390000000
1!
1$
b1 %
1'
1*
b1 +
#541400000000
0!
0'
#541410000000
1!
b10 %
1'
b10 +
#541420000000
0!
0'
#541430000000
1!
b11 %
1'
b11 +
#541440000000
0!
0'
#541450000000
1!
b100 %
1'
b100 +
#541460000000
0!
0'
#541470000000
1!
b101 %
1'
b101 +
#541480000000
0!
0'
#541490000000
1!
0$
b110 %
1'
0*
b110 +
#541500000000
0!
0'
#541510000000
1!
b111 %
1'
b111 +
#541520000000
0!
0'
#541530000000
1!
b1000 %
1'
b1000 +
#541540000000
0!
0'
#541550000000
1!
b1001 %
1'
b1001 +
#541560000000
0!
0'
#541570000000
1!
b0 %
1'
b0 +
#541580000000
1"
1(
#541590000000
0!
0"
b100 &
0'
0(
b100 ,
#541600000000
1!
1$
b1 %
1'
1*
b1 +
#541610000000
0!
0'
#541620000000
1!
b10 %
1'
b10 +
#541630000000
0!
0'
#541640000000
1!
b11 %
1'
b11 +
#541650000000
0!
0'
#541660000000
1!
b100 %
1'
b100 +
#541670000000
0!
0'
#541680000000
1!
b101 %
1'
b101 +
#541690000000
0!
0'
#541700000000
1!
b110 %
1'
b110 +
#541710000000
0!
0'
#541720000000
1!
b111 %
1'
b111 +
#541730000000
0!
0'
#541740000000
1!
0$
b1000 %
1'
0*
b1000 +
#541750000000
0!
0'
#541760000000
1!
b1001 %
1'
b1001 +
#541770000000
0!
0'
#541780000000
1!
b0 %
1'
b0 +
#541790000000
0!
0'
#541800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#541810000000
0!
0'
#541820000000
1!
b10 %
1'
b10 +
#541830000000
0!
0'
#541840000000
1!
b11 %
1'
b11 +
#541850000000
0!
0'
#541860000000
1!
b100 %
1'
b100 +
#541870000000
0!
0'
#541880000000
1!
b101 %
1'
b101 +
#541890000000
0!
0'
#541900000000
1!
0$
b110 %
1'
0*
b110 +
#541910000000
0!
0'
#541920000000
1!
b111 %
1'
b111 +
#541930000000
0!
0'
#541940000000
1!
b1000 %
1'
b1000 +
#541950000000
0!
0'
#541960000000
1!
b1001 %
1'
b1001 +
#541970000000
0!
0'
#541980000000
1!
b0 %
1'
b0 +
#541990000000
0!
0'
#542000000000
1!
1$
b1 %
1'
1*
b1 +
#542010000000
1"
1(
#542020000000
0!
0"
b100 &
0'
0(
b100 ,
#542030000000
1!
b10 %
1'
b10 +
#542040000000
0!
0'
#542050000000
1!
b11 %
1'
b11 +
#542060000000
0!
0'
#542070000000
1!
b100 %
1'
b100 +
#542080000000
0!
0'
#542090000000
1!
b101 %
1'
b101 +
#542100000000
0!
0'
#542110000000
1!
b110 %
1'
b110 +
#542120000000
0!
0'
#542130000000
1!
b111 %
1'
b111 +
#542140000000
0!
0'
#542150000000
1!
0$
b1000 %
1'
0*
b1000 +
#542160000000
0!
0'
#542170000000
1!
b1001 %
1'
b1001 +
#542180000000
0!
0'
#542190000000
1!
b0 %
1'
b0 +
#542200000000
0!
0'
#542210000000
1!
1$
b1 %
1'
1*
b1 +
#542220000000
0!
0'
#542230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#542240000000
0!
0'
#542250000000
1!
b11 %
1'
b11 +
#542260000000
0!
0'
#542270000000
1!
b100 %
1'
b100 +
#542280000000
0!
0'
#542290000000
1!
b101 %
1'
b101 +
#542300000000
0!
0'
#542310000000
1!
0$
b110 %
1'
0*
b110 +
#542320000000
0!
0'
#542330000000
1!
b111 %
1'
b111 +
#542340000000
0!
0'
#542350000000
1!
b1000 %
1'
b1000 +
#542360000000
0!
0'
#542370000000
1!
b1001 %
1'
b1001 +
#542380000000
0!
0'
#542390000000
1!
b0 %
1'
b0 +
#542400000000
0!
0'
#542410000000
1!
1$
b1 %
1'
1*
b1 +
#542420000000
0!
0'
#542430000000
1!
b10 %
1'
b10 +
#542440000000
1"
1(
#542450000000
0!
0"
b100 &
0'
0(
b100 ,
#542460000000
1!
b11 %
1'
b11 +
#542470000000
0!
0'
#542480000000
1!
b100 %
1'
b100 +
#542490000000
0!
0'
#542500000000
1!
b101 %
1'
b101 +
#542510000000
0!
0'
#542520000000
1!
b110 %
1'
b110 +
#542530000000
0!
0'
#542540000000
1!
b111 %
1'
b111 +
#542550000000
0!
0'
#542560000000
1!
0$
b1000 %
1'
0*
b1000 +
#542570000000
0!
0'
#542580000000
1!
b1001 %
1'
b1001 +
#542590000000
0!
0'
#542600000000
1!
b0 %
1'
b0 +
#542610000000
0!
0'
#542620000000
1!
1$
b1 %
1'
1*
b1 +
#542630000000
0!
0'
#542640000000
1!
b10 %
1'
b10 +
#542650000000
0!
0'
#542660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#542670000000
0!
0'
#542680000000
1!
b100 %
1'
b100 +
#542690000000
0!
0'
#542700000000
1!
b101 %
1'
b101 +
#542710000000
0!
0'
#542720000000
1!
0$
b110 %
1'
0*
b110 +
#542730000000
0!
0'
#542740000000
1!
b111 %
1'
b111 +
#542750000000
0!
0'
#542760000000
1!
b1000 %
1'
b1000 +
#542770000000
0!
0'
#542780000000
1!
b1001 %
1'
b1001 +
#542790000000
0!
0'
#542800000000
1!
b0 %
1'
b0 +
#542810000000
0!
0'
#542820000000
1!
1$
b1 %
1'
1*
b1 +
#542830000000
0!
0'
#542840000000
1!
b10 %
1'
b10 +
#542850000000
0!
0'
#542860000000
1!
b11 %
1'
b11 +
#542870000000
1"
1(
#542880000000
0!
0"
b100 &
0'
0(
b100 ,
#542890000000
1!
b100 %
1'
b100 +
#542900000000
0!
0'
#542910000000
1!
b101 %
1'
b101 +
#542920000000
0!
0'
#542930000000
1!
b110 %
1'
b110 +
#542940000000
0!
0'
#542950000000
1!
b111 %
1'
b111 +
#542960000000
0!
0'
#542970000000
1!
0$
b1000 %
1'
0*
b1000 +
#542980000000
0!
0'
#542990000000
1!
b1001 %
1'
b1001 +
#543000000000
0!
0'
#543010000000
1!
b0 %
1'
b0 +
#543020000000
0!
0'
#543030000000
1!
1$
b1 %
1'
1*
b1 +
#543040000000
0!
0'
#543050000000
1!
b10 %
1'
b10 +
#543060000000
0!
0'
#543070000000
1!
b11 %
1'
b11 +
#543080000000
0!
0'
#543090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#543100000000
0!
0'
#543110000000
1!
b101 %
1'
b101 +
#543120000000
0!
0'
#543130000000
1!
0$
b110 %
1'
0*
b110 +
#543140000000
0!
0'
#543150000000
1!
b111 %
1'
b111 +
#543160000000
0!
0'
#543170000000
1!
b1000 %
1'
b1000 +
#543180000000
0!
0'
#543190000000
1!
b1001 %
1'
b1001 +
#543200000000
0!
0'
#543210000000
1!
b0 %
1'
b0 +
#543220000000
0!
0'
#543230000000
1!
1$
b1 %
1'
1*
b1 +
#543240000000
0!
0'
#543250000000
1!
b10 %
1'
b10 +
#543260000000
0!
0'
#543270000000
1!
b11 %
1'
b11 +
#543280000000
0!
0'
#543290000000
1!
b100 %
1'
b100 +
#543300000000
1"
1(
#543310000000
0!
0"
b100 &
0'
0(
b100 ,
#543320000000
1!
b101 %
1'
b101 +
#543330000000
0!
0'
#543340000000
1!
b110 %
1'
b110 +
#543350000000
0!
0'
#543360000000
1!
b111 %
1'
b111 +
#543370000000
0!
0'
#543380000000
1!
0$
b1000 %
1'
0*
b1000 +
#543390000000
0!
0'
#543400000000
1!
b1001 %
1'
b1001 +
#543410000000
0!
0'
#543420000000
1!
b0 %
1'
b0 +
#543430000000
0!
0'
#543440000000
1!
1$
b1 %
1'
1*
b1 +
#543450000000
0!
0'
#543460000000
1!
b10 %
1'
b10 +
#543470000000
0!
0'
#543480000000
1!
b11 %
1'
b11 +
#543490000000
0!
0'
#543500000000
1!
b100 %
1'
b100 +
#543510000000
0!
0'
#543520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#543530000000
0!
0'
#543540000000
1!
0$
b110 %
1'
0*
b110 +
#543550000000
0!
0'
#543560000000
1!
b111 %
1'
b111 +
#543570000000
0!
0'
#543580000000
1!
b1000 %
1'
b1000 +
#543590000000
0!
0'
#543600000000
1!
b1001 %
1'
b1001 +
#543610000000
0!
0'
#543620000000
1!
b0 %
1'
b0 +
#543630000000
0!
0'
#543640000000
1!
1$
b1 %
1'
1*
b1 +
#543650000000
0!
0'
#543660000000
1!
b10 %
1'
b10 +
#543670000000
0!
0'
#543680000000
1!
b11 %
1'
b11 +
#543690000000
0!
0'
#543700000000
1!
b100 %
1'
b100 +
#543710000000
0!
0'
#543720000000
1!
b101 %
1'
b101 +
#543730000000
1"
1(
#543740000000
0!
0"
b100 &
0'
0(
b100 ,
#543750000000
1!
b110 %
1'
b110 +
#543760000000
0!
0'
#543770000000
1!
b111 %
1'
b111 +
#543780000000
0!
0'
#543790000000
1!
0$
b1000 %
1'
0*
b1000 +
#543800000000
0!
0'
#543810000000
1!
b1001 %
1'
b1001 +
#543820000000
0!
0'
#543830000000
1!
b0 %
1'
b0 +
#543840000000
0!
0'
#543850000000
1!
1$
b1 %
1'
1*
b1 +
#543860000000
0!
0'
#543870000000
1!
b10 %
1'
b10 +
#543880000000
0!
0'
#543890000000
1!
b11 %
1'
b11 +
#543900000000
0!
0'
#543910000000
1!
b100 %
1'
b100 +
#543920000000
0!
0'
#543930000000
1!
b101 %
1'
b101 +
#543940000000
0!
0'
#543950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#543960000000
0!
0'
#543970000000
1!
b111 %
1'
b111 +
#543980000000
0!
0'
#543990000000
1!
b1000 %
1'
b1000 +
#544000000000
0!
0'
#544010000000
1!
b1001 %
1'
b1001 +
#544020000000
0!
0'
#544030000000
1!
b0 %
1'
b0 +
#544040000000
0!
0'
#544050000000
1!
1$
b1 %
1'
1*
b1 +
#544060000000
0!
0'
#544070000000
1!
b10 %
1'
b10 +
#544080000000
0!
0'
#544090000000
1!
b11 %
1'
b11 +
#544100000000
0!
0'
#544110000000
1!
b100 %
1'
b100 +
#544120000000
0!
0'
#544130000000
1!
b101 %
1'
b101 +
#544140000000
0!
0'
#544150000000
1!
0$
b110 %
1'
0*
b110 +
#544160000000
1"
1(
#544170000000
0!
0"
b100 &
0'
0(
b100 ,
#544180000000
1!
1$
b111 %
1'
1*
b111 +
#544190000000
0!
0'
#544200000000
1!
0$
b1000 %
1'
0*
b1000 +
#544210000000
0!
0'
#544220000000
1!
b1001 %
1'
b1001 +
#544230000000
0!
0'
#544240000000
1!
b0 %
1'
b0 +
#544250000000
0!
0'
#544260000000
1!
1$
b1 %
1'
1*
b1 +
#544270000000
0!
0'
#544280000000
1!
b10 %
1'
b10 +
#544290000000
0!
0'
#544300000000
1!
b11 %
1'
b11 +
#544310000000
0!
0'
#544320000000
1!
b100 %
1'
b100 +
#544330000000
0!
0'
#544340000000
1!
b101 %
1'
b101 +
#544350000000
0!
0'
#544360000000
1!
b110 %
1'
b110 +
#544370000000
0!
0'
#544380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#544390000000
0!
0'
#544400000000
1!
b1000 %
1'
b1000 +
#544410000000
0!
0'
#544420000000
1!
b1001 %
1'
b1001 +
#544430000000
0!
0'
#544440000000
1!
b0 %
1'
b0 +
#544450000000
0!
0'
#544460000000
1!
1$
b1 %
1'
1*
b1 +
#544470000000
0!
0'
#544480000000
1!
b10 %
1'
b10 +
#544490000000
0!
0'
#544500000000
1!
b11 %
1'
b11 +
#544510000000
0!
0'
#544520000000
1!
b100 %
1'
b100 +
#544530000000
0!
0'
#544540000000
1!
b101 %
1'
b101 +
#544550000000
0!
0'
#544560000000
1!
0$
b110 %
1'
0*
b110 +
#544570000000
0!
0'
#544580000000
1!
b111 %
1'
b111 +
#544590000000
1"
1(
#544600000000
0!
0"
b100 &
0'
0(
b100 ,
#544610000000
1!
b1000 %
1'
b1000 +
#544620000000
0!
0'
#544630000000
1!
b1001 %
1'
b1001 +
#544640000000
0!
0'
#544650000000
1!
b0 %
1'
b0 +
#544660000000
0!
0'
#544670000000
1!
1$
b1 %
1'
1*
b1 +
#544680000000
0!
0'
#544690000000
1!
b10 %
1'
b10 +
#544700000000
0!
0'
#544710000000
1!
b11 %
1'
b11 +
#544720000000
0!
0'
#544730000000
1!
b100 %
1'
b100 +
#544740000000
0!
0'
#544750000000
1!
b101 %
1'
b101 +
#544760000000
0!
0'
#544770000000
1!
b110 %
1'
b110 +
#544780000000
0!
0'
#544790000000
1!
b111 %
1'
b111 +
#544800000000
0!
0'
#544810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#544820000000
0!
0'
#544830000000
1!
b1001 %
1'
b1001 +
#544840000000
0!
0'
#544850000000
1!
b0 %
1'
b0 +
#544860000000
0!
0'
#544870000000
1!
1$
b1 %
1'
1*
b1 +
#544880000000
0!
0'
#544890000000
1!
b10 %
1'
b10 +
#544900000000
0!
0'
#544910000000
1!
b11 %
1'
b11 +
#544920000000
0!
0'
#544930000000
1!
b100 %
1'
b100 +
#544940000000
0!
0'
#544950000000
1!
b101 %
1'
b101 +
#544960000000
0!
0'
#544970000000
1!
0$
b110 %
1'
0*
b110 +
#544980000000
0!
0'
#544990000000
1!
b111 %
1'
b111 +
#545000000000
0!
0'
#545010000000
1!
b1000 %
1'
b1000 +
#545020000000
1"
1(
#545030000000
0!
0"
b100 &
0'
0(
b100 ,
#545040000000
1!
b1001 %
1'
b1001 +
#545050000000
0!
0'
#545060000000
1!
b0 %
1'
b0 +
#545070000000
0!
0'
#545080000000
1!
1$
b1 %
1'
1*
b1 +
#545090000000
0!
0'
#545100000000
1!
b10 %
1'
b10 +
#545110000000
0!
0'
#545120000000
1!
b11 %
1'
b11 +
#545130000000
0!
0'
#545140000000
1!
b100 %
1'
b100 +
#545150000000
0!
0'
#545160000000
1!
b101 %
1'
b101 +
#545170000000
0!
0'
#545180000000
1!
b110 %
1'
b110 +
#545190000000
0!
0'
#545200000000
1!
b111 %
1'
b111 +
#545210000000
0!
0'
#545220000000
1!
0$
b1000 %
1'
0*
b1000 +
#545230000000
0!
0'
#545240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#545250000000
0!
0'
#545260000000
1!
b0 %
1'
b0 +
#545270000000
0!
0'
#545280000000
1!
1$
b1 %
1'
1*
b1 +
#545290000000
0!
0'
#545300000000
1!
b10 %
1'
b10 +
#545310000000
0!
0'
#545320000000
1!
b11 %
1'
b11 +
#545330000000
0!
0'
#545340000000
1!
b100 %
1'
b100 +
#545350000000
0!
0'
#545360000000
1!
b101 %
1'
b101 +
#545370000000
0!
0'
#545380000000
1!
0$
b110 %
1'
0*
b110 +
#545390000000
0!
0'
#545400000000
1!
b111 %
1'
b111 +
#545410000000
0!
0'
#545420000000
1!
b1000 %
1'
b1000 +
#545430000000
0!
0'
#545440000000
1!
b1001 %
1'
b1001 +
#545450000000
1"
1(
#545460000000
0!
0"
b100 &
0'
0(
b100 ,
#545470000000
1!
b0 %
1'
b0 +
#545480000000
0!
0'
#545490000000
1!
1$
b1 %
1'
1*
b1 +
#545500000000
0!
0'
#545510000000
1!
b10 %
1'
b10 +
#545520000000
0!
0'
#545530000000
1!
b11 %
1'
b11 +
#545540000000
0!
0'
#545550000000
1!
b100 %
1'
b100 +
#545560000000
0!
0'
#545570000000
1!
b101 %
1'
b101 +
#545580000000
0!
0'
#545590000000
1!
b110 %
1'
b110 +
#545600000000
0!
0'
#545610000000
1!
b111 %
1'
b111 +
#545620000000
0!
0'
#545630000000
1!
0$
b1000 %
1'
0*
b1000 +
#545640000000
0!
0'
#545650000000
1!
b1001 %
1'
b1001 +
#545660000000
0!
0'
#545670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#545680000000
0!
0'
#545690000000
1!
1$
b1 %
1'
1*
b1 +
#545700000000
0!
0'
#545710000000
1!
b10 %
1'
b10 +
#545720000000
0!
0'
#545730000000
1!
b11 %
1'
b11 +
#545740000000
0!
0'
#545750000000
1!
b100 %
1'
b100 +
#545760000000
0!
0'
#545770000000
1!
b101 %
1'
b101 +
#545780000000
0!
0'
#545790000000
1!
0$
b110 %
1'
0*
b110 +
#545800000000
0!
0'
#545810000000
1!
b111 %
1'
b111 +
#545820000000
0!
0'
#545830000000
1!
b1000 %
1'
b1000 +
#545840000000
0!
0'
#545850000000
1!
b1001 %
1'
b1001 +
#545860000000
0!
0'
#545870000000
1!
b0 %
1'
b0 +
#545880000000
1"
1(
#545890000000
0!
0"
b100 &
0'
0(
b100 ,
#545900000000
1!
1$
b1 %
1'
1*
b1 +
#545910000000
0!
0'
#545920000000
1!
b10 %
1'
b10 +
#545930000000
0!
0'
#545940000000
1!
b11 %
1'
b11 +
#545950000000
0!
0'
#545960000000
1!
b100 %
1'
b100 +
#545970000000
0!
0'
#545980000000
1!
b101 %
1'
b101 +
#545990000000
0!
0'
#546000000000
1!
b110 %
1'
b110 +
#546010000000
0!
0'
#546020000000
1!
b111 %
1'
b111 +
#546030000000
0!
0'
#546040000000
1!
0$
b1000 %
1'
0*
b1000 +
#546050000000
0!
0'
#546060000000
1!
b1001 %
1'
b1001 +
#546070000000
0!
0'
#546080000000
1!
b0 %
1'
b0 +
#546090000000
0!
0'
#546100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#546110000000
0!
0'
#546120000000
1!
b10 %
1'
b10 +
#546130000000
0!
0'
#546140000000
1!
b11 %
1'
b11 +
#546150000000
0!
0'
#546160000000
1!
b100 %
1'
b100 +
#546170000000
0!
0'
#546180000000
1!
b101 %
1'
b101 +
#546190000000
0!
0'
#546200000000
1!
0$
b110 %
1'
0*
b110 +
#546210000000
0!
0'
#546220000000
1!
b111 %
1'
b111 +
#546230000000
0!
0'
#546240000000
1!
b1000 %
1'
b1000 +
#546250000000
0!
0'
#546260000000
1!
b1001 %
1'
b1001 +
#546270000000
0!
0'
#546280000000
1!
b0 %
1'
b0 +
#546290000000
0!
0'
#546300000000
1!
1$
b1 %
1'
1*
b1 +
#546310000000
1"
1(
#546320000000
0!
0"
b100 &
0'
0(
b100 ,
#546330000000
1!
b10 %
1'
b10 +
#546340000000
0!
0'
#546350000000
1!
b11 %
1'
b11 +
#546360000000
0!
0'
#546370000000
1!
b100 %
1'
b100 +
#546380000000
0!
0'
#546390000000
1!
b101 %
1'
b101 +
#546400000000
0!
0'
#546410000000
1!
b110 %
1'
b110 +
#546420000000
0!
0'
#546430000000
1!
b111 %
1'
b111 +
#546440000000
0!
0'
#546450000000
1!
0$
b1000 %
1'
0*
b1000 +
#546460000000
0!
0'
#546470000000
1!
b1001 %
1'
b1001 +
#546480000000
0!
0'
#546490000000
1!
b0 %
1'
b0 +
#546500000000
0!
0'
#546510000000
1!
1$
b1 %
1'
1*
b1 +
#546520000000
0!
0'
#546530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#546540000000
0!
0'
#546550000000
1!
b11 %
1'
b11 +
#546560000000
0!
0'
#546570000000
1!
b100 %
1'
b100 +
#546580000000
0!
0'
#546590000000
1!
b101 %
1'
b101 +
#546600000000
0!
0'
#546610000000
1!
0$
b110 %
1'
0*
b110 +
#546620000000
0!
0'
#546630000000
1!
b111 %
1'
b111 +
#546640000000
0!
0'
#546650000000
1!
b1000 %
1'
b1000 +
#546660000000
0!
0'
#546670000000
1!
b1001 %
1'
b1001 +
#546680000000
0!
0'
#546690000000
1!
b0 %
1'
b0 +
#546700000000
0!
0'
#546710000000
1!
1$
b1 %
1'
1*
b1 +
#546720000000
0!
0'
#546730000000
1!
b10 %
1'
b10 +
#546740000000
1"
1(
#546750000000
0!
0"
b100 &
0'
0(
b100 ,
#546760000000
1!
b11 %
1'
b11 +
#546770000000
0!
0'
#546780000000
1!
b100 %
1'
b100 +
#546790000000
0!
0'
#546800000000
1!
b101 %
1'
b101 +
#546810000000
0!
0'
#546820000000
1!
b110 %
1'
b110 +
#546830000000
0!
0'
#546840000000
1!
b111 %
1'
b111 +
#546850000000
0!
0'
#546860000000
1!
0$
b1000 %
1'
0*
b1000 +
#546870000000
0!
0'
#546880000000
1!
b1001 %
1'
b1001 +
#546890000000
0!
0'
#546900000000
1!
b0 %
1'
b0 +
#546910000000
0!
0'
#546920000000
1!
1$
b1 %
1'
1*
b1 +
#546930000000
0!
0'
#546940000000
1!
b10 %
1'
b10 +
#546950000000
0!
0'
#546960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#546970000000
0!
0'
#546980000000
1!
b100 %
1'
b100 +
#546990000000
0!
0'
#547000000000
1!
b101 %
1'
b101 +
#547010000000
0!
0'
#547020000000
1!
0$
b110 %
1'
0*
b110 +
#547030000000
0!
0'
#547040000000
1!
b111 %
1'
b111 +
#547050000000
0!
0'
#547060000000
1!
b1000 %
1'
b1000 +
#547070000000
0!
0'
#547080000000
1!
b1001 %
1'
b1001 +
#547090000000
0!
0'
#547100000000
1!
b0 %
1'
b0 +
#547110000000
0!
0'
#547120000000
1!
1$
b1 %
1'
1*
b1 +
#547130000000
0!
0'
#547140000000
1!
b10 %
1'
b10 +
#547150000000
0!
0'
#547160000000
1!
b11 %
1'
b11 +
#547170000000
1"
1(
#547180000000
0!
0"
b100 &
0'
0(
b100 ,
#547190000000
1!
b100 %
1'
b100 +
#547200000000
0!
0'
#547210000000
1!
b101 %
1'
b101 +
#547220000000
0!
0'
#547230000000
1!
b110 %
1'
b110 +
#547240000000
0!
0'
#547250000000
1!
b111 %
1'
b111 +
#547260000000
0!
0'
#547270000000
1!
0$
b1000 %
1'
0*
b1000 +
#547280000000
0!
0'
#547290000000
1!
b1001 %
1'
b1001 +
#547300000000
0!
0'
#547310000000
1!
b0 %
1'
b0 +
#547320000000
0!
0'
#547330000000
1!
1$
b1 %
1'
1*
b1 +
#547340000000
0!
0'
#547350000000
1!
b10 %
1'
b10 +
#547360000000
0!
0'
#547370000000
1!
b11 %
1'
b11 +
#547380000000
0!
0'
#547390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#547400000000
0!
0'
#547410000000
1!
b101 %
1'
b101 +
#547420000000
0!
0'
#547430000000
1!
0$
b110 %
1'
0*
b110 +
#547440000000
0!
0'
#547450000000
1!
b111 %
1'
b111 +
#547460000000
0!
0'
#547470000000
1!
b1000 %
1'
b1000 +
#547480000000
0!
0'
#547490000000
1!
b1001 %
1'
b1001 +
#547500000000
0!
0'
#547510000000
1!
b0 %
1'
b0 +
#547520000000
0!
0'
#547530000000
1!
1$
b1 %
1'
1*
b1 +
#547540000000
0!
0'
#547550000000
1!
b10 %
1'
b10 +
#547560000000
0!
0'
#547570000000
1!
b11 %
1'
b11 +
#547580000000
0!
0'
#547590000000
1!
b100 %
1'
b100 +
#547600000000
1"
1(
#547610000000
0!
0"
b100 &
0'
0(
b100 ,
#547620000000
1!
b101 %
1'
b101 +
#547630000000
0!
0'
#547640000000
1!
b110 %
1'
b110 +
#547650000000
0!
0'
#547660000000
1!
b111 %
1'
b111 +
#547670000000
0!
0'
#547680000000
1!
0$
b1000 %
1'
0*
b1000 +
#547690000000
0!
0'
#547700000000
1!
b1001 %
1'
b1001 +
#547710000000
0!
0'
#547720000000
1!
b0 %
1'
b0 +
#547730000000
0!
0'
#547740000000
1!
1$
b1 %
1'
1*
b1 +
#547750000000
0!
0'
#547760000000
1!
b10 %
1'
b10 +
#547770000000
0!
0'
#547780000000
1!
b11 %
1'
b11 +
#547790000000
0!
0'
#547800000000
1!
b100 %
1'
b100 +
#547810000000
0!
0'
#547820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#547830000000
0!
0'
#547840000000
1!
0$
b110 %
1'
0*
b110 +
#547850000000
0!
0'
#547860000000
1!
b111 %
1'
b111 +
#547870000000
0!
0'
#547880000000
1!
b1000 %
1'
b1000 +
#547890000000
0!
0'
#547900000000
1!
b1001 %
1'
b1001 +
#547910000000
0!
0'
#547920000000
1!
b0 %
1'
b0 +
#547930000000
0!
0'
#547940000000
1!
1$
b1 %
1'
1*
b1 +
#547950000000
0!
0'
#547960000000
1!
b10 %
1'
b10 +
#547970000000
0!
0'
#547980000000
1!
b11 %
1'
b11 +
#547990000000
0!
0'
#548000000000
1!
b100 %
1'
b100 +
#548010000000
0!
0'
#548020000000
1!
b101 %
1'
b101 +
#548030000000
1"
1(
#548040000000
0!
0"
b100 &
0'
0(
b100 ,
#548050000000
1!
b110 %
1'
b110 +
#548060000000
0!
0'
#548070000000
1!
b111 %
1'
b111 +
#548080000000
0!
0'
#548090000000
1!
0$
b1000 %
1'
0*
b1000 +
#548100000000
0!
0'
#548110000000
1!
b1001 %
1'
b1001 +
#548120000000
0!
0'
#548130000000
1!
b0 %
1'
b0 +
#548140000000
0!
0'
#548150000000
1!
1$
b1 %
1'
1*
b1 +
#548160000000
0!
0'
#548170000000
1!
b10 %
1'
b10 +
#548180000000
0!
0'
#548190000000
1!
b11 %
1'
b11 +
#548200000000
0!
0'
#548210000000
1!
b100 %
1'
b100 +
#548220000000
0!
0'
#548230000000
1!
b101 %
1'
b101 +
#548240000000
0!
0'
#548250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#548260000000
0!
0'
#548270000000
1!
b111 %
1'
b111 +
#548280000000
0!
0'
#548290000000
1!
b1000 %
1'
b1000 +
#548300000000
0!
0'
#548310000000
1!
b1001 %
1'
b1001 +
#548320000000
0!
0'
#548330000000
1!
b0 %
1'
b0 +
#548340000000
0!
0'
#548350000000
1!
1$
b1 %
1'
1*
b1 +
#548360000000
0!
0'
#548370000000
1!
b10 %
1'
b10 +
#548380000000
0!
0'
#548390000000
1!
b11 %
1'
b11 +
#548400000000
0!
0'
#548410000000
1!
b100 %
1'
b100 +
#548420000000
0!
0'
#548430000000
1!
b101 %
1'
b101 +
#548440000000
0!
0'
#548450000000
1!
0$
b110 %
1'
0*
b110 +
#548460000000
1"
1(
#548470000000
0!
0"
b100 &
0'
0(
b100 ,
#548480000000
1!
1$
b111 %
1'
1*
b111 +
#548490000000
0!
0'
#548500000000
1!
0$
b1000 %
1'
0*
b1000 +
#548510000000
0!
0'
#548520000000
1!
b1001 %
1'
b1001 +
#548530000000
0!
0'
#548540000000
1!
b0 %
1'
b0 +
#548550000000
0!
0'
#548560000000
1!
1$
b1 %
1'
1*
b1 +
#548570000000
0!
0'
#548580000000
1!
b10 %
1'
b10 +
#548590000000
0!
0'
#548600000000
1!
b11 %
1'
b11 +
#548610000000
0!
0'
#548620000000
1!
b100 %
1'
b100 +
#548630000000
0!
0'
#548640000000
1!
b101 %
1'
b101 +
#548650000000
0!
0'
#548660000000
1!
b110 %
1'
b110 +
#548670000000
0!
0'
#548680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#548690000000
0!
0'
#548700000000
1!
b1000 %
1'
b1000 +
#548710000000
0!
0'
#548720000000
1!
b1001 %
1'
b1001 +
#548730000000
0!
0'
#548740000000
1!
b0 %
1'
b0 +
#548750000000
0!
0'
#548760000000
1!
1$
b1 %
1'
1*
b1 +
#548770000000
0!
0'
#548780000000
1!
b10 %
1'
b10 +
#548790000000
0!
0'
#548800000000
1!
b11 %
1'
b11 +
#548810000000
0!
0'
#548820000000
1!
b100 %
1'
b100 +
#548830000000
0!
0'
#548840000000
1!
b101 %
1'
b101 +
#548850000000
0!
0'
#548860000000
1!
0$
b110 %
1'
0*
b110 +
#548870000000
0!
0'
#548880000000
1!
b111 %
1'
b111 +
#548890000000
1"
1(
#548900000000
0!
0"
b100 &
0'
0(
b100 ,
#548910000000
1!
b1000 %
1'
b1000 +
#548920000000
0!
0'
#548930000000
1!
b1001 %
1'
b1001 +
#548940000000
0!
0'
#548950000000
1!
b0 %
1'
b0 +
#548960000000
0!
0'
#548970000000
1!
1$
b1 %
1'
1*
b1 +
#548980000000
0!
0'
#548990000000
1!
b10 %
1'
b10 +
#549000000000
0!
0'
#549010000000
1!
b11 %
1'
b11 +
#549020000000
0!
0'
#549030000000
1!
b100 %
1'
b100 +
#549040000000
0!
0'
#549050000000
1!
b101 %
1'
b101 +
#549060000000
0!
0'
#549070000000
1!
b110 %
1'
b110 +
#549080000000
0!
0'
#549090000000
1!
b111 %
1'
b111 +
#549100000000
0!
0'
#549110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#549120000000
0!
0'
#549130000000
1!
b1001 %
1'
b1001 +
#549140000000
0!
0'
#549150000000
1!
b0 %
1'
b0 +
#549160000000
0!
0'
#549170000000
1!
1$
b1 %
1'
1*
b1 +
#549180000000
0!
0'
#549190000000
1!
b10 %
1'
b10 +
#549200000000
0!
0'
#549210000000
1!
b11 %
1'
b11 +
#549220000000
0!
0'
#549230000000
1!
b100 %
1'
b100 +
#549240000000
0!
0'
#549250000000
1!
b101 %
1'
b101 +
#549260000000
0!
0'
#549270000000
1!
0$
b110 %
1'
0*
b110 +
#549280000000
0!
0'
#549290000000
1!
b111 %
1'
b111 +
#549300000000
0!
0'
#549310000000
1!
b1000 %
1'
b1000 +
#549320000000
1"
1(
#549330000000
0!
0"
b100 &
0'
0(
b100 ,
#549340000000
1!
b1001 %
1'
b1001 +
#549350000000
0!
0'
#549360000000
1!
b0 %
1'
b0 +
#549370000000
0!
0'
#549380000000
1!
1$
b1 %
1'
1*
b1 +
#549390000000
0!
0'
#549400000000
1!
b10 %
1'
b10 +
#549410000000
0!
0'
#549420000000
1!
b11 %
1'
b11 +
#549430000000
0!
0'
#549440000000
1!
b100 %
1'
b100 +
#549450000000
0!
0'
#549460000000
1!
b101 %
1'
b101 +
#549470000000
0!
0'
#549480000000
1!
b110 %
1'
b110 +
#549490000000
0!
0'
#549500000000
1!
b111 %
1'
b111 +
#549510000000
0!
0'
#549520000000
1!
0$
b1000 %
1'
0*
b1000 +
#549530000000
0!
0'
#549540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#549550000000
0!
0'
#549560000000
1!
b0 %
1'
b0 +
#549570000000
0!
0'
#549580000000
1!
1$
b1 %
1'
1*
b1 +
#549590000000
0!
0'
#549600000000
1!
b10 %
1'
b10 +
#549610000000
0!
0'
#549620000000
1!
b11 %
1'
b11 +
#549630000000
0!
0'
#549640000000
1!
b100 %
1'
b100 +
#549650000000
0!
0'
#549660000000
1!
b101 %
1'
b101 +
#549670000000
0!
0'
#549680000000
1!
0$
b110 %
1'
0*
b110 +
#549690000000
0!
0'
#549700000000
1!
b111 %
1'
b111 +
#549710000000
0!
0'
#549720000000
1!
b1000 %
1'
b1000 +
#549730000000
0!
0'
#549740000000
1!
b1001 %
1'
b1001 +
#549750000000
1"
1(
#549760000000
0!
0"
b100 &
0'
0(
b100 ,
#549770000000
1!
b0 %
1'
b0 +
#549780000000
0!
0'
#549790000000
1!
1$
b1 %
1'
1*
b1 +
#549800000000
0!
0'
#549810000000
1!
b10 %
1'
b10 +
#549820000000
0!
0'
#549830000000
1!
b11 %
1'
b11 +
#549840000000
0!
0'
#549850000000
1!
b100 %
1'
b100 +
#549860000000
0!
0'
#549870000000
1!
b101 %
1'
b101 +
#549880000000
0!
0'
#549890000000
1!
b110 %
1'
b110 +
#549900000000
0!
0'
#549910000000
1!
b111 %
1'
b111 +
#549920000000
0!
0'
#549930000000
1!
0$
b1000 %
1'
0*
b1000 +
#549940000000
0!
0'
#549950000000
1!
b1001 %
1'
b1001 +
#549960000000
0!
0'
#549970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#549980000000
0!
0'
#549990000000
1!
1$
b1 %
1'
1*
b1 +
#550000000000
0!
0'
#550010000000
1!
b10 %
1'
b10 +
#550020000000
0!
0'
#550030000000
1!
b11 %
1'
b11 +
#550040000000
0!
0'
#550050000000
1!
b100 %
1'
b100 +
#550060000000
0!
0'
#550070000000
1!
b101 %
1'
b101 +
#550080000000
0!
0'
#550090000000
1!
0$
b110 %
1'
0*
b110 +
#550100000000
0!
0'
#550110000000
1!
b111 %
1'
b111 +
#550120000000
0!
0'
#550130000000
1!
b1000 %
1'
b1000 +
#550140000000
0!
0'
#550150000000
1!
b1001 %
1'
b1001 +
#550160000000
0!
0'
#550170000000
1!
b0 %
1'
b0 +
#550180000000
1"
1(
#550190000000
0!
0"
b100 &
0'
0(
b100 ,
#550200000000
1!
1$
b1 %
1'
1*
b1 +
#550210000000
0!
0'
#550220000000
1!
b10 %
1'
b10 +
#550230000000
0!
0'
#550240000000
1!
b11 %
1'
b11 +
#550250000000
0!
0'
#550260000000
1!
b100 %
1'
b100 +
#550270000000
0!
0'
#550280000000
1!
b101 %
1'
b101 +
#550290000000
0!
0'
#550300000000
1!
b110 %
1'
b110 +
#550310000000
0!
0'
#550320000000
1!
b111 %
1'
b111 +
#550330000000
0!
0'
#550340000000
1!
0$
b1000 %
1'
0*
b1000 +
#550350000000
0!
0'
#550360000000
1!
b1001 %
1'
b1001 +
#550370000000
0!
0'
#550380000000
1!
b0 %
1'
b0 +
#550390000000
0!
0'
#550400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#550410000000
0!
0'
#550420000000
1!
b10 %
1'
b10 +
#550430000000
0!
0'
#550440000000
1!
b11 %
1'
b11 +
#550450000000
0!
0'
#550460000000
1!
b100 %
1'
b100 +
#550470000000
0!
0'
#550480000000
1!
b101 %
1'
b101 +
#550490000000
0!
0'
#550500000000
1!
0$
b110 %
1'
0*
b110 +
#550510000000
0!
0'
#550520000000
1!
b111 %
1'
b111 +
#550530000000
0!
0'
#550540000000
1!
b1000 %
1'
b1000 +
#550550000000
0!
0'
#550560000000
1!
b1001 %
1'
b1001 +
#550570000000
0!
0'
#550580000000
1!
b0 %
1'
b0 +
#550590000000
0!
0'
#550600000000
1!
1$
b1 %
1'
1*
b1 +
#550610000000
1"
1(
#550620000000
0!
0"
b100 &
0'
0(
b100 ,
#550630000000
1!
b10 %
1'
b10 +
#550640000000
0!
0'
#550650000000
1!
b11 %
1'
b11 +
#550660000000
0!
0'
#550670000000
1!
b100 %
1'
b100 +
#550680000000
0!
0'
#550690000000
1!
b101 %
1'
b101 +
#550700000000
0!
0'
#550710000000
1!
b110 %
1'
b110 +
#550720000000
0!
0'
#550730000000
1!
b111 %
1'
b111 +
#550740000000
0!
0'
#550750000000
1!
0$
b1000 %
1'
0*
b1000 +
#550760000000
0!
0'
#550770000000
1!
b1001 %
1'
b1001 +
#550780000000
0!
0'
#550790000000
1!
b0 %
1'
b0 +
#550800000000
0!
0'
#550810000000
1!
1$
b1 %
1'
1*
b1 +
#550820000000
0!
0'
#550830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#550840000000
0!
0'
#550850000000
1!
b11 %
1'
b11 +
#550860000000
0!
0'
#550870000000
1!
b100 %
1'
b100 +
#550880000000
0!
0'
#550890000000
1!
b101 %
1'
b101 +
#550900000000
0!
0'
#550910000000
1!
0$
b110 %
1'
0*
b110 +
#550920000000
0!
0'
#550930000000
1!
b111 %
1'
b111 +
#550940000000
0!
0'
#550950000000
1!
b1000 %
1'
b1000 +
#550960000000
0!
0'
#550970000000
1!
b1001 %
1'
b1001 +
#550980000000
0!
0'
#550990000000
1!
b0 %
1'
b0 +
#551000000000
0!
0'
#551010000000
1!
1$
b1 %
1'
1*
b1 +
#551020000000
0!
0'
#551030000000
1!
b10 %
1'
b10 +
#551040000000
1"
1(
#551050000000
0!
0"
b100 &
0'
0(
b100 ,
#551060000000
1!
b11 %
1'
b11 +
#551070000000
0!
0'
#551080000000
1!
b100 %
1'
b100 +
#551090000000
0!
0'
#551100000000
1!
b101 %
1'
b101 +
#551110000000
0!
0'
#551120000000
1!
b110 %
1'
b110 +
#551130000000
0!
0'
#551140000000
1!
b111 %
1'
b111 +
#551150000000
0!
0'
#551160000000
1!
0$
b1000 %
1'
0*
b1000 +
#551170000000
0!
0'
#551180000000
1!
b1001 %
1'
b1001 +
#551190000000
0!
0'
#551200000000
1!
b0 %
1'
b0 +
#551210000000
0!
0'
#551220000000
1!
1$
b1 %
1'
1*
b1 +
#551230000000
0!
0'
#551240000000
1!
b10 %
1'
b10 +
#551250000000
0!
0'
#551260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#551270000000
0!
0'
#551280000000
1!
b100 %
1'
b100 +
#551290000000
0!
0'
#551300000000
1!
b101 %
1'
b101 +
#551310000000
0!
0'
#551320000000
1!
0$
b110 %
1'
0*
b110 +
#551330000000
0!
0'
#551340000000
1!
b111 %
1'
b111 +
#551350000000
0!
0'
#551360000000
1!
b1000 %
1'
b1000 +
#551370000000
0!
0'
#551380000000
1!
b1001 %
1'
b1001 +
#551390000000
0!
0'
#551400000000
1!
b0 %
1'
b0 +
#551410000000
0!
0'
#551420000000
1!
1$
b1 %
1'
1*
b1 +
#551430000000
0!
0'
#551440000000
1!
b10 %
1'
b10 +
#551450000000
0!
0'
#551460000000
1!
b11 %
1'
b11 +
#551470000000
1"
1(
#551480000000
0!
0"
b100 &
0'
0(
b100 ,
#551490000000
1!
b100 %
1'
b100 +
#551500000000
0!
0'
#551510000000
1!
b101 %
1'
b101 +
#551520000000
0!
0'
#551530000000
1!
b110 %
1'
b110 +
#551540000000
0!
0'
#551550000000
1!
b111 %
1'
b111 +
#551560000000
0!
0'
#551570000000
1!
0$
b1000 %
1'
0*
b1000 +
#551580000000
0!
0'
#551590000000
1!
b1001 %
1'
b1001 +
#551600000000
0!
0'
#551610000000
1!
b0 %
1'
b0 +
#551620000000
0!
0'
#551630000000
1!
1$
b1 %
1'
1*
b1 +
#551640000000
0!
0'
#551650000000
1!
b10 %
1'
b10 +
#551660000000
0!
0'
#551670000000
1!
b11 %
1'
b11 +
#551680000000
0!
0'
#551690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#551700000000
0!
0'
#551710000000
1!
b101 %
1'
b101 +
#551720000000
0!
0'
#551730000000
1!
0$
b110 %
1'
0*
b110 +
#551740000000
0!
0'
#551750000000
1!
b111 %
1'
b111 +
#551760000000
0!
0'
#551770000000
1!
b1000 %
1'
b1000 +
#551780000000
0!
0'
#551790000000
1!
b1001 %
1'
b1001 +
#551800000000
0!
0'
#551810000000
1!
b0 %
1'
b0 +
#551820000000
0!
0'
#551830000000
1!
1$
b1 %
1'
1*
b1 +
#551840000000
0!
0'
#551850000000
1!
b10 %
1'
b10 +
#551860000000
0!
0'
#551870000000
1!
b11 %
1'
b11 +
#551880000000
0!
0'
#551890000000
1!
b100 %
1'
b100 +
#551900000000
1"
1(
#551910000000
0!
0"
b100 &
0'
0(
b100 ,
#551920000000
1!
b101 %
1'
b101 +
#551930000000
0!
0'
#551940000000
1!
b110 %
1'
b110 +
#551950000000
0!
0'
#551960000000
1!
b111 %
1'
b111 +
#551970000000
0!
0'
#551980000000
1!
0$
b1000 %
1'
0*
b1000 +
#551990000000
0!
0'
#552000000000
1!
b1001 %
1'
b1001 +
#552010000000
0!
0'
#552020000000
1!
b0 %
1'
b0 +
#552030000000
0!
0'
#552040000000
1!
1$
b1 %
1'
1*
b1 +
#552050000000
0!
0'
#552060000000
1!
b10 %
1'
b10 +
#552070000000
0!
0'
#552080000000
1!
b11 %
1'
b11 +
#552090000000
0!
0'
#552100000000
1!
b100 %
1'
b100 +
#552110000000
0!
0'
#552120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#552130000000
0!
0'
#552140000000
1!
0$
b110 %
1'
0*
b110 +
#552150000000
0!
0'
#552160000000
1!
b111 %
1'
b111 +
#552170000000
0!
0'
#552180000000
1!
b1000 %
1'
b1000 +
#552190000000
0!
0'
#552200000000
1!
b1001 %
1'
b1001 +
#552210000000
0!
0'
#552220000000
1!
b0 %
1'
b0 +
#552230000000
0!
0'
#552240000000
1!
1$
b1 %
1'
1*
b1 +
#552250000000
0!
0'
#552260000000
1!
b10 %
1'
b10 +
#552270000000
0!
0'
#552280000000
1!
b11 %
1'
b11 +
#552290000000
0!
0'
#552300000000
1!
b100 %
1'
b100 +
#552310000000
0!
0'
#552320000000
1!
b101 %
1'
b101 +
#552330000000
1"
1(
#552340000000
0!
0"
b100 &
0'
0(
b100 ,
#552350000000
1!
b110 %
1'
b110 +
#552360000000
0!
0'
#552370000000
1!
b111 %
1'
b111 +
#552380000000
0!
0'
#552390000000
1!
0$
b1000 %
1'
0*
b1000 +
#552400000000
0!
0'
#552410000000
1!
b1001 %
1'
b1001 +
#552420000000
0!
0'
#552430000000
1!
b0 %
1'
b0 +
#552440000000
0!
0'
#552450000000
1!
1$
b1 %
1'
1*
b1 +
#552460000000
0!
0'
#552470000000
1!
b10 %
1'
b10 +
#552480000000
0!
0'
#552490000000
1!
b11 %
1'
b11 +
#552500000000
0!
0'
#552510000000
1!
b100 %
1'
b100 +
#552520000000
0!
0'
#552530000000
1!
b101 %
1'
b101 +
#552540000000
0!
0'
#552550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#552560000000
0!
0'
#552570000000
1!
b111 %
1'
b111 +
#552580000000
0!
0'
#552590000000
1!
b1000 %
1'
b1000 +
#552600000000
0!
0'
#552610000000
1!
b1001 %
1'
b1001 +
#552620000000
0!
0'
#552630000000
1!
b0 %
1'
b0 +
#552640000000
0!
0'
#552650000000
1!
1$
b1 %
1'
1*
b1 +
#552660000000
0!
0'
#552670000000
1!
b10 %
1'
b10 +
#552680000000
0!
0'
#552690000000
1!
b11 %
1'
b11 +
#552700000000
0!
0'
#552710000000
1!
b100 %
1'
b100 +
#552720000000
0!
0'
#552730000000
1!
b101 %
1'
b101 +
#552740000000
0!
0'
#552750000000
1!
0$
b110 %
1'
0*
b110 +
#552760000000
1"
1(
#552770000000
0!
0"
b100 &
0'
0(
b100 ,
#552780000000
1!
1$
b111 %
1'
1*
b111 +
#552790000000
0!
0'
#552800000000
1!
0$
b1000 %
1'
0*
b1000 +
#552810000000
0!
0'
#552820000000
1!
b1001 %
1'
b1001 +
#552830000000
0!
0'
#552840000000
1!
b0 %
1'
b0 +
#552850000000
0!
0'
#552860000000
1!
1$
b1 %
1'
1*
b1 +
#552870000000
0!
0'
#552880000000
1!
b10 %
1'
b10 +
#552890000000
0!
0'
#552900000000
1!
b11 %
1'
b11 +
#552910000000
0!
0'
#552920000000
1!
b100 %
1'
b100 +
#552930000000
0!
0'
#552940000000
1!
b101 %
1'
b101 +
#552950000000
0!
0'
#552960000000
1!
b110 %
1'
b110 +
#552970000000
0!
0'
#552980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#552990000000
0!
0'
#553000000000
1!
b1000 %
1'
b1000 +
#553010000000
0!
0'
#553020000000
1!
b1001 %
1'
b1001 +
#553030000000
0!
0'
#553040000000
1!
b0 %
1'
b0 +
#553050000000
0!
0'
#553060000000
1!
1$
b1 %
1'
1*
b1 +
#553070000000
0!
0'
#553080000000
1!
b10 %
1'
b10 +
#553090000000
0!
0'
#553100000000
1!
b11 %
1'
b11 +
#553110000000
0!
0'
#553120000000
1!
b100 %
1'
b100 +
#553130000000
0!
0'
#553140000000
1!
b101 %
1'
b101 +
#553150000000
0!
0'
#553160000000
1!
0$
b110 %
1'
0*
b110 +
#553170000000
0!
0'
#553180000000
1!
b111 %
1'
b111 +
#553190000000
1"
1(
#553200000000
0!
0"
b100 &
0'
0(
b100 ,
#553210000000
1!
b1000 %
1'
b1000 +
#553220000000
0!
0'
#553230000000
1!
b1001 %
1'
b1001 +
#553240000000
0!
0'
#553250000000
1!
b0 %
1'
b0 +
#553260000000
0!
0'
#553270000000
1!
1$
b1 %
1'
1*
b1 +
#553280000000
0!
0'
#553290000000
1!
b10 %
1'
b10 +
#553300000000
0!
0'
#553310000000
1!
b11 %
1'
b11 +
#553320000000
0!
0'
#553330000000
1!
b100 %
1'
b100 +
#553340000000
0!
0'
#553350000000
1!
b101 %
1'
b101 +
#553360000000
0!
0'
#553370000000
1!
b110 %
1'
b110 +
#553380000000
0!
0'
#553390000000
1!
b111 %
1'
b111 +
#553400000000
0!
0'
#553410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#553420000000
0!
0'
#553430000000
1!
b1001 %
1'
b1001 +
#553440000000
0!
0'
#553450000000
1!
b0 %
1'
b0 +
#553460000000
0!
0'
#553470000000
1!
1$
b1 %
1'
1*
b1 +
#553480000000
0!
0'
#553490000000
1!
b10 %
1'
b10 +
#553500000000
0!
0'
#553510000000
1!
b11 %
1'
b11 +
#553520000000
0!
0'
#553530000000
1!
b100 %
1'
b100 +
#553540000000
0!
0'
#553550000000
1!
b101 %
1'
b101 +
#553560000000
0!
0'
#553570000000
1!
0$
b110 %
1'
0*
b110 +
#553580000000
0!
0'
#553590000000
1!
b111 %
1'
b111 +
#553600000000
0!
0'
#553610000000
1!
b1000 %
1'
b1000 +
#553620000000
1"
1(
#553630000000
0!
0"
b100 &
0'
0(
b100 ,
#553640000000
1!
b1001 %
1'
b1001 +
#553650000000
0!
0'
#553660000000
1!
b0 %
1'
b0 +
#553670000000
0!
0'
#553680000000
1!
1$
b1 %
1'
1*
b1 +
#553690000000
0!
0'
#553700000000
1!
b10 %
1'
b10 +
#553710000000
0!
0'
#553720000000
1!
b11 %
1'
b11 +
#553730000000
0!
0'
#553740000000
1!
b100 %
1'
b100 +
#553750000000
0!
0'
#553760000000
1!
b101 %
1'
b101 +
#553770000000
0!
0'
#553780000000
1!
b110 %
1'
b110 +
#553790000000
0!
0'
#553800000000
1!
b111 %
1'
b111 +
#553810000000
0!
0'
#553820000000
1!
0$
b1000 %
1'
0*
b1000 +
#553830000000
0!
0'
#553840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#553850000000
0!
0'
#553860000000
1!
b0 %
1'
b0 +
#553870000000
0!
0'
#553880000000
1!
1$
b1 %
1'
1*
b1 +
#553890000000
0!
0'
#553900000000
1!
b10 %
1'
b10 +
#553910000000
0!
0'
#553920000000
1!
b11 %
1'
b11 +
#553930000000
0!
0'
#553940000000
1!
b100 %
1'
b100 +
#553950000000
0!
0'
#553960000000
1!
b101 %
1'
b101 +
#553970000000
0!
0'
#553980000000
1!
0$
b110 %
1'
0*
b110 +
#553990000000
0!
0'
#554000000000
1!
b111 %
1'
b111 +
#554010000000
0!
0'
#554020000000
1!
b1000 %
1'
b1000 +
#554030000000
0!
0'
#554040000000
1!
b1001 %
1'
b1001 +
#554050000000
1"
1(
#554060000000
0!
0"
b100 &
0'
0(
b100 ,
#554070000000
1!
b0 %
1'
b0 +
#554080000000
0!
0'
#554090000000
1!
1$
b1 %
1'
1*
b1 +
#554100000000
0!
0'
#554110000000
1!
b10 %
1'
b10 +
#554120000000
0!
0'
#554130000000
1!
b11 %
1'
b11 +
#554140000000
0!
0'
#554150000000
1!
b100 %
1'
b100 +
#554160000000
0!
0'
#554170000000
1!
b101 %
1'
b101 +
#554180000000
0!
0'
#554190000000
1!
b110 %
1'
b110 +
#554200000000
0!
0'
#554210000000
1!
b111 %
1'
b111 +
#554220000000
0!
0'
#554230000000
1!
0$
b1000 %
1'
0*
b1000 +
#554240000000
0!
0'
#554250000000
1!
b1001 %
1'
b1001 +
#554260000000
0!
0'
#554270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#554280000000
0!
0'
#554290000000
1!
1$
b1 %
1'
1*
b1 +
#554300000000
0!
0'
#554310000000
1!
b10 %
1'
b10 +
#554320000000
0!
0'
#554330000000
1!
b11 %
1'
b11 +
#554340000000
0!
0'
#554350000000
1!
b100 %
1'
b100 +
#554360000000
0!
0'
#554370000000
1!
b101 %
1'
b101 +
#554380000000
0!
0'
#554390000000
1!
0$
b110 %
1'
0*
b110 +
#554400000000
0!
0'
#554410000000
1!
b111 %
1'
b111 +
#554420000000
0!
0'
#554430000000
1!
b1000 %
1'
b1000 +
#554440000000
0!
0'
#554450000000
1!
b1001 %
1'
b1001 +
#554460000000
0!
0'
#554470000000
1!
b0 %
1'
b0 +
#554480000000
1"
1(
#554490000000
0!
0"
b100 &
0'
0(
b100 ,
#554500000000
1!
1$
b1 %
1'
1*
b1 +
#554510000000
0!
0'
#554520000000
1!
b10 %
1'
b10 +
#554530000000
0!
0'
#554540000000
1!
b11 %
1'
b11 +
#554550000000
0!
0'
#554560000000
1!
b100 %
1'
b100 +
#554570000000
0!
0'
#554580000000
1!
b101 %
1'
b101 +
#554590000000
0!
0'
#554600000000
1!
b110 %
1'
b110 +
#554610000000
0!
0'
#554620000000
1!
b111 %
1'
b111 +
#554630000000
0!
0'
#554640000000
1!
0$
b1000 %
1'
0*
b1000 +
#554650000000
0!
0'
#554660000000
1!
b1001 %
1'
b1001 +
#554670000000
0!
0'
#554680000000
1!
b0 %
1'
b0 +
#554690000000
0!
0'
#554700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#554710000000
0!
0'
#554720000000
1!
b10 %
1'
b10 +
#554730000000
0!
0'
#554740000000
1!
b11 %
1'
b11 +
#554750000000
0!
0'
#554760000000
1!
b100 %
1'
b100 +
#554770000000
0!
0'
#554780000000
1!
b101 %
1'
b101 +
#554790000000
0!
0'
#554800000000
1!
0$
b110 %
1'
0*
b110 +
#554810000000
0!
0'
#554820000000
1!
b111 %
1'
b111 +
#554830000000
0!
0'
#554840000000
1!
b1000 %
1'
b1000 +
#554850000000
0!
0'
#554860000000
1!
b1001 %
1'
b1001 +
#554870000000
0!
0'
#554880000000
1!
b0 %
1'
b0 +
#554890000000
0!
0'
#554900000000
1!
1$
b1 %
1'
1*
b1 +
#554910000000
1"
1(
#554920000000
0!
0"
b100 &
0'
0(
b100 ,
#554930000000
1!
b10 %
1'
b10 +
#554940000000
0!
0'
#554950000000
1!
b11 %
1'
b11 +
#554960000000
0!
0'
#554970000000
1!
b100 %
1'
b100 +
#554980000000
0!
0'
#554990000000
1!
b101 %
1'
b101 +
#555000000000
0!
0'
#555010000000
1!
b110 %
1'
b110 +
#555020000000
0!
0'
#555030000000
1!
b111 %
1'
b111 +
#555040000000
0!
0'
#555050000000
1!
0$
b1000 %
1'
0*
b1000 +
#555060000000
0!
0'
#555070000000
1!
b1001 %
1'
b1001 +
#555080000000
0!
0'
#555090000000
1!
b0 %
1'
b0 +
#555100000000
0!
0'
#555110000000
1!
1$
b1 %
1'
1*
b1 +
#555120000000
0!
0'
#555130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#555140000000
0!
0'
#555150000000
1!
b11 %
1'
b11 +
#555160000000
0!
0'
#555170000000
1!
b100 %
1'
b100 +
#555180000000
0!
0'
#555190000000
1!
b101 %
1'
b101 +
#555200000000
0!
0'
#555210000000
1!
0$
b110 %
1'
0*
b110 +
#555220000000
0!
0'
#555230000000
1!
b111 %
1'
b111 +
#555240000000
0!
0'
#555250000000
1!
b1000 %
1'
b1000 +
#555260000000
0!
0'
#555270000000
1!
b1001 %
1'
b1001 +
#555280000000
0!
0'
#555290000000
1!
b0 %
1'
b0 +
#555300000000
0!
0'
#555310000000
1!
1$
b1 %
1'
1*
b1 +
#555320000000
0!
0'
#555330000000
1!
b10 %
1'
b10 +
#555340000000
1"
1(
#555350000000
0!
0"
b100 &
0'
0(
b100 ,
#555360000000
1!
b11 %
1'
b11 +
#555370000000
0!
0'
#555380000000
1!
b100 %
1'
b100 +
#555390000000
0!
0'
#555400000000
1!
b101 %
1'
b101 +
#555410000000
0!
0'
#555420000000
1!
b110 %
1'
b110 +
#555430000000
0!
0'
#555440000000
1!
b111 %
1'
b111 +
#555450000000
0!
0'
#555460000000
1!
0$
b1000 %
1'
0*
b1000 +
#555470000000
0!
0'
#555480000000
1!
b1001 %
1'
b1001 +
#555490000000
0!
0'
#555500000000
1!
b0 %
1'
b0 +
#555510000000
0!
0'
#555520000000
1!
1$
b1 %
1'
1*
b1 +
#555530000000
0!
0'
#555540000000
1!
b10 %
1'
b10 +
#555550000000
0!
0'
#555560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#555570000000
0!
0'
#555580000000
1!
b100 %
1'
b100 +
#555590000000
0!
0'
#555600000000
1!
b101 %
1'
b101 +
#555610000000
0!
0'
#555620000000
1!
0$
b110 %
1'
0*
b110 +
#555630000000
0!
0'
#555640000000
1!
b111 %
1'
b111 +
#555650000000
0!
0'
#555660000000
1!
b1000 %
1'
b1000 +
#555670000000
0!
0'
#555680000000
1!
b1001 %
1'
b1001 +
#555690000000
0!
0'
#555700000000
1!
b0 %
1'
b0 +
#555710000000
0!
0'
#555720000000
1!
1$
b1 %
1'
1*
b1 +
#555730000000
0!
0'
#555740000000
1!
b10 %
1'
b10 +
#555750000000
0!
0'
#555760000000
1!
b11 %
1'
b11 +
#555770000000
1"
1(
#555780000000
0!
0"
b100 &
0'
0(
b100 ,
#555790000000
1!
b100 %
1'
b100 +
#555800000000
0!
0'
#555810000000
1!
b101 %
1'
b101 +
#555820000000
0!
0'
#555830000000
1!
b110 %
1'
b110 +
#555840000000
0!
0'
#555850000000
1!
b111 %
1'
b111 +
#555860000000
0!
0'
#555870000000
1!
0$
b1000 %
1'
0*
b1000 +
#555880000000
0!
0'
#555890000000
1!
b1001 %
1'
b1001 +
#555900000000
0!
0'
#555910000000
1!
b0 %
1'
b0 +
#555920000000
0!
0'
#555930000000
1!
1$
b1 %
1'
1*
b1 +
#555940000000
0!
0'
#555950000000
1!
b10 %
1'
b10 +
#555960000000
0!
0'
#555970000000
1!
b11 %
1'
b11 +
#555980000000
0!
0'
#555990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#556000000000
0!
0'
#556010000000
1!
b101 %
1'
b101 +
#556020000000
0!
0'
#556030000000
1!
0$
b110 %
1'
0*
b110 +
#556040000000
0!
0'
#556050000000
1!
b111 %
1'
b111 +
#556060000000
0!
0'
#556070000000
1!
b1000 %
1'
b1000 +
#556080000000
0!
0'
#556090000000
1!
b1001 %
1'
b1001 +
#556100000000
0!
0'
#556110000000
1!
b0 %
1'
b0 +
#556120000000
0!
0'
#556130000000
1!
1$
b1 %
1'
1*
b1 +
#556140000000
0!
0'
#556150000000
1!
b10 %
1'
b10 +
#556160000000
0!
0'
#556170000000
1!
b11 %
1'
b11 +
#556180000000
0!
0'
#556190000000
1!
b100 %
1'
b100 +
#556200000000
1"
1(
#556210000000
0!
0"
b100 &
0'
0(
b100 ,
#556220000000
1!
b101 %
1'
b101 +
#556230000000
0!
0'
#556240000000
1!
b110 %
1'
b110 +
#556250000000
0!
0'
#556260000000
1!
b111 %
1'
b111 +
#556270000000
0!
0'
#556280000000
1!
0$
b1000 %
1'
0*
b1000 +
#556290000000
0!
0'
#556300000000
1!
b1001 %
1'
b1001 +
#556310000000
0!
0'
#556320000000
1!
b0 %
1'
b0 +
#556330000000
0!
0'
#556340000000
1!
1$
b1 %
1'
1*
b1 +
#556350000000
0!
0'
#556360000000
1!
b10 %
1'
b10 +
#556370000000
0!
0'
#556380000000
1!
b11 %
1'
b11 +
#556390000000
0!
0'
#556400000000
1!
b100 %
1'
b100 +
#556410000000
0!
0'
#556420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#556430000000
0!
0'
#556440000000
1!
0$
b110 %
1'
0*
b110 +
#556450000000
0!
0'
#556460000000
1!
b111 %
1'
b111 +
#556470000000
0!
0'
#556480000000
1!
b1000 %
1'
b1000 +
#556490000000
0!
0'
#556500000000
1!
b1001 %
1'
b1001 +
#556510000000
0!
0'
#556520000000
1!
b0 %
1'
b0 +
#556530000000
0!
0'
#556540000000
1!
1$
b1 %
1'
1*
b1 +
#556550000000
0!
0'
#556560000000
1!
b10 %
1'
b10 +
#556570000000
0!
0'
#556580000000
1!
b11 %
1'
b11 +
#556590000000
0!
0'
#556600000000
1!
b100 %
1'
b100 +
#556610000000
0!
0'
#556620000000
1!
b101 %
1'
b101 +
#556630000000
1"
1(
#556640000000
0!
0"
b100 &
0'
0(
b100 ,
#556650000000
1!
b110 %
1'
b110 +
#556660000000
0!
0'
#556670000000
1!
b111 %
1'
b111 +
#556680000000
0!
0'
#556690000000
1!
0$
b1000 %
1'
0*
b1000 +
#556700000000
0!
0'
#556710000000
1!
b1001 %
1'
b1001 +
#556720000000
0!
0'
#556730000000
1!
b0 %
1'
b0 +
#556740000000
0!
0'
#556750000000
1!
1$
b1 %
1'
1*
b1 +
#556760000000
0!
0'
#556770000000
1!
b10 %
1'
b10 +
#556780000000
0!
0'
#556790000000
1!
b11 %
1'
b11 +
#556800000000
0!
0'
#556810000000
1!
b100 %
1'
b100 +
#556820000000
0!
0'
#556830000000
1!
b101 %
1'
b101 +
#556840000000
0!
0'
#556850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#556860000000
0!
0'
#556870000000
1!
b111 %
1'
b111 +
#556880000000
0!
0'
#556890000000
1!
b1000 %
1'
b1000 +
#556900000000
0!
0'
#556910000000
1!
b1001 %
1'
b1001 +
#556920000000
0!
0'
#556930000000
1!
b0 %
1'
b0 +
#556940000000
0!
0'
#556950000000
1!
1$
b1 %
1'
1*
b1 +
#556960000000
0!
0'
#556970000000
1!
b10 %
1'
b10 +
#556980000000
0!
0'
#556990000000
1!
b11 %
1'
b11 +
#557000000000
0!
0'
#557010000000
1!
b100 %
1'
b100 +
#557020000000
0!
0'
#557030000000
1!
b101 %
1'
b101 +
#557040000000
0!
0'
#557050000000
1!
0$
b110 %
1'
0*
b110 +
#557060000000
1"
1(
#557070000000
0!
0"
b100 &
0'
0(
b100 ,
#557080000000
1!
1$
b111 %
1'
1*
b111 +
#557090000000
0!
0'
#557100000000
1!
0$
b1000 %
1'
0*
b1000 +
#557110000000
0!
0'
#557120000000
1!
b1001 %
1'
b1001 +
#557130000000
0!
0'
#557140000000
1!
b0 %
1'
b0 +
#557150000000
0!
0'
#557160000000
1!
1$
b1 %
1'
1*
b1 +
#557170000000
0!
0'
#557180000000
1!
b10 %
1'
b10 +
#557190000000
0!
0'
#557200000000
1!
b11 %
1'
b11 +
#557210000000
0!
0'
#557220000000
1!
b100 %
1'
b100 +
#557230000000
0!
0'
#557240000000
1!
b101 %
1'
b101 +
#557250000000
0!
0'
#557260000000
1!
b110 %
1'
b110 +
#557270000000
0!
0'
#557280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#557290000000
0!
0'
#557300000000
1!
b1000 %
1'
b1000 +
#557310000000
0!
0'
#557320000000
1!
b1001 %
1'
b1001 +
#557330000000
0!
0'
#557340000000
1!
b0 %
1'
b0 +
#557350000000
0!
0'
#557360000000
1!
1$
b1 %
1'
1*
b1 +
#557370000000
0!
0'
#557380000000
1!
b10 %
1'
b10 +
#557390000000
0!
0'
#557400000000
1!
b11 %
1'
b11 +
#557410000000
0!
0'
#557420000000
1!
b100 %
1'
b100 +
#557430000000
0!
0'
#557440000000
1!
b101 %
1'
b101 +
#557450000000
0!
0'
#557460000000
1!
0$
b110 %
1'
0*
b110 +
#557470000000
0!
0'
#557480000000
1!
b111 %
1'
b111 +
#557490000000
1"
1(
#557500000000
0!
0"
b100 &
0'
0(
b100 ,
#557510000000
1!
b1000 %
1'
b1000 +
#557520000000
0!
0'
#557530000000
1!
b1001 %
1'
b1001 +
#557540000000
0!
0'
#557550000000
1!
b0 %
1'
b0 +
#557560000000
0!
0'
#557570000000
1!
1$
b1 %
1'
1*
b1 +
#557580000000
0!
0'
#557590000000
1!
b10 %
1'
b10 +
#557600000000
0!
0'
#557610000000
1!
b11 %
1'
b11 +
#557620000000
0!
0'
#557630000000
1!
b100 %
1'
b100 +
#557640000000
0!
0'
#557650000000
1!
b101 %
1'
b101 +
#557660000000
0!
0'
#557670000000
1!
b110 %
1'
b110 +
#557680000000
0!
0'
#557690000000
1!
b111 %
1'
b111 +
#557700000000
0!
0'
#557710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#557720000000
0!
0'
#557730000000
1!
b1001 %
1'
b1001 +
#557740000000
0!
0'
#557750000000
1!
b0 %
1'
b0 +
#557760000000
0!
0'
#557770000000
1!
1$
b1 %
1'
1*
b1 +
#557780000000
0!
0'
#557790000000
1!
b10 %
1'
b10 +
#557800000000
0!
0'
#557810000000
1!
b11 %
1'
b11 +
#557820000000
0!
0'
#557830000000
1!
b100 %
1'
b100 +
#557840000000
0!
0'
#557850000000
1!
b101 %
1'
b101 +
#557860000000
0!
0'
#557870000000
1!
0$
b110 %
1'
0*
b110 +
#557880000000
0!
0'
#557890000000
1!
b111 %
1'
b111 +
#557900000000
0!
0'
#557910000000
1!
b1000 %
1'
b1000 +
#557920000000
1"
1(
#557930000000
0!
0"
b100 &
0'
0(
b100 ,
#557940000000
1!
b1001 %
1'
b1001 +
#557950000000
0!
0'
#557960000000
1!
b0 %
1'
b0 +
#557970000000
0!
0'
#557980000000
1!
1$
b1 %
1'
1*
b1 +
#557990000000
0!
0'
#558000000000
1!
b10 %
1'
b10 +
#558010000000
0!
0'
#558020000000
1!
b11 %
1'
b11 +
#558030000000
0!
0'
#558040000000
1!
b100 %
1'
b100 +
#558050000000
0!
0'
#558060000000
1!
b101 %
1'
b101 +
#558070000000
0!
0'
#558080000000
1!
b110 %
1'
b110 +
#558090000000
0!
0'
#558100000000
1!
b111 %
1'
b111 +
#558110000000
0!
0'
#558120000000
1!
0$
b1000 %
1'
0*
b1000 +
#558130000000
0!
0'
#558140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#558150000000
0!
0'
#558160000000
1!
b0 %
1'
b0 +
#558170000000
0!
0'
#558180000000
1!
1$
b1 %
1'
1*
b1 +
#558190000000
0!
0'
#558200000000
1!
b10 %
1'
b10 +
#558210000000
0!
0'
#558220000000
1!
b11 %
1'
b11 +
#558230000000
0!
0'
#558240000000
1!
b100 %
1'
b100 +
#558250000000
0!
0'
#558260000000
1!
b101 %
1'
b101 +
#558270000000
0!
0'
#558280000000
1!
0$
b110 %
1'
0*
b110 +
#558290000000
0!
0'
#558300000000
1!
b111 %
1'
b111 +
#558310000000
0!
0'
#558320000000
1!
b1000 %
1'
b1000 +
#558330000000
0!
0'
#558340000000
1!
b1001 %
1'
b1001 +
#558350000000
1"
1(
#558360000000
0!
0"
b100 &
0'
0(
b100 ,
#558370000000
1!
b0 %
1'
b0 +
#558380000000
0!
0'
#558390000000
1!
1$
b1 %
1'
1*
b1 +
#558400000000
0!
0'
#558410000000
1!
b10 %
1'
b10 +
#558420000000
0!
0'
#558430000000
1!
b11 %
1'
b11 +
#558440000000
0!
0'
#558450000000
1!
b100 %
1'
b100 +
#558460000000
0!
0'
#558470000000
1!
b101 %
1'
b101 +
#558480000000
0!
0'
#558490000000
1!
b110 %
1'
b110 +
#558500000000
0!
0'
#558510000000
1!
b111 %
1'
b111 +
#558520000000
0!
0'
#558530000000
1!
0$
b1000 %
1'
0*
b1000 +
#558540000000
0!
0'
#558550000000
1!
b1001 %
1'
b1001 +
#558560000000
0!
0'
#558570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#558580000000
0!
0'
#558590000000
1!
1$
b1 %
1'
1*
b1 +
#558600000000
0!
0'
#558610000000
1!
b10 %
1'
b10 +
#558620000000
0!
0'
#558630000000
1!
b11 %
1'
b11 +
#558640000000
0!
0'
#558650000000
1!
b100 %
1'
b100 +
#558660000000
0!
0'
#558670000000
1!
b101 %
1'
b101 +
#558680000000
0!
0'
#558690000000
1!
0$
b110 %
1'
0*
b110 +
#558700000000
0!
0'
#558710000000
1!
b111 %
1'
b111 +
#558720000000
0!
0'
#558730000000
1!
b1000 %
1'
b1000 +
#558740000000
0!
0'
#558750000000
1!
b1001 %
1'
b1001 +
#558760000000
0!
0'
#558770000000
1!
b0 %
1'
b0 +
#558780000000
1"
1(
#558790000000
0!
0"
b100 &
0'
0(
b100 ,
#558800000000
1!
1$
b1 %
1'
1*
b1 +
#558810000000
0!
0'
#558820000000
1!
b10 %
1'
b10 +
#558830000000
0!
0'
#558840000000
1!
b11 %
1'
b11 +
#558850000000
0!
0'
#558860000000
1!
b100 %
1'
b100 +
#558870000000
0!
0'
#558880000000
1!
b101 %
1'
b101 +
#558890000000
0!
0'
#558900000000
1!
b110 %
1'
b110 +
#558910000000
0!
0'
#558920000000
1!
b111 %
1'
b111 +
#558930000000
0!
0'
#558940000000
1!
0$
b1000 %
1'
0*
b1000 +
#558950000000
0!
0'
#558960000000
1!
b1001 %
1'
b1001 +
#558970000000
0!
0'
#558980000000
1!
b0 %
1'
b0 +
#558990000000
0!
0'
#559000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#559010000000
0!
0'
#559020000000
1!
b10 %
1'
b10 +
#559030000000
0!
0'
#559040000000
1!
b11 %
1'
b11 +
#559050000000
0!
0'
#559060000000
1!
b100 %
1'
b100 +
#559070000000
0!
0'
#559080000000
1!
b101 %
1'
b101 +
#559090000000
0!
0'
#559100000000
1!
0$
b110 %
1'
0*
b110 +
#559110000000
0!
0'
#559120000000
1!
b111 %
1'
b111 +
#559130000000
0!
0'
#559140000000
1!
b1000 %
1'
b1000 +
#559150000000
0!
0'
#559160000000
1!
b1001 %
1'
b1001 +
#559170000000
0!
0'
#559180000000
1!
b0 %
1'
b0 +
#559190000000
0!
0'
#559200000000
1!
1$
b1 %
1'
1*
b1 +
#559210000000
1"
1(
#559220000000
0!
0"
b100 &
0'
0(
b100 ,
#559230000000
1!
b10 %
1'
b10 +
#559240000000
0!
0'
#559250000000
1!
b11 %
1'
b11 +
#559260000000
0!
0'
#559270000000
1!
b100 %
1'
b100 +
#559280000000
0!
0'
#559290000000
1!
b101 %
1'
b101 +
#559300000000
0!
0'
#559310000000
1!
b110 %
1'
b110 +
#559320000000
0!
0'
#559330000000
1!
b111 %
1'
b111 +
#559340000000
0!
0'
#559350000000
1!
0$
b1000 %
1'
0*
b1000 +
#559360000000
0!
0'
#559370000000
1!
b1001 %
1'
b1001 +
#559380000000
0!
0'
#559390000000
1!
b0 %
1'
b0 +
#559400000000
0!
0'
#559410000000
1!
1$
b1 %
1'
1*
b1 +
#559420000000
0!
0'
#559430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#559440000000
0!
0'
#559450000000
1!
b11 %
1'
b11 +
#559460000000
0!
0'
#559470000000
1!
b100 %
1'
b100 +
#559480000000
0!
0'
#559490000000
1!
b101 %
1'
b101 +
#559500000000
0!
0'
#559510000000
1!
0$
b110 %
1'
0*
b110 +
#559520000000
0!
0'
#559530000000
1!
b111 %
1'
b111 +
#559540000000
0!
0'
#559550000000
1!
b1000 %
1'
b1000 +
#559560000000
0!
0'
#559570000000
1!
b1001 %
1'
b1001 +
#559580000000
0!
0'
#559590000000
1!
b0 %
1'
b0 +
#559600000000
0!
0'
#559610000000
1!
1$
b1 %
1'
1*
b1 +
#559620000000
0!
0'
#559630000000
1!
b10 %
1'
b10 +
#559640000000
1"
1(
#559650000000
0!
0"
b100 &
0'
0(
b100 ,
#559660000000
1!
b11 %
1'
b11 +
#559670000000
0!
0'
#559680000000
1!
b100 %
1'
b100 +
#559690000000
0!
0'
#559700000000
1!
b101 %
1'
b101 +
#559710000000
0!
0'
#559720000000
1!
b110 %
1'
b110 +
#559730000000
0!
0'
#559740000000
1!
b111 %
1'
b111 +
#559750000000
0!
0'
#559760000000
1!
0$
b1000 %
1'
0*
b1000 +
#559770000000
0!
0'
#559780000000
1!
b1001 %
1'
b1001 +
#559790000000
0!
0'
#559800000000
1!
b0 %
1'
b0 +
#559810000000
0!
0'
#559820000000
1!
1$
b1 %
1'
1*
b1 +
#559830000000
0!
0'
#559840000000
1!
b10 %
1'
b10 +
#559850000000
0!
0'
#559860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#559870000000
0!
0'
#559880000000
1!
b100 %
1'
b100 +
#559890000000
0!
0'
#559900000000
1!
b101 %
1'
b101 +
#559910000000
0!
0'
#559920000000
1!
0$
b110 %
1'
0*
b110 +
#559930000000
0!
0'
#559940000000
1!
b111 %
1'
b111 +
#559950000000
0!
0'
#559960000000
1!
b1000 %
1'
b1000 +
#559970000000
0!
0'
#559980000000
1!
b1001 %
1'
b1001 +
#559990000000
0!
0'
#560000000000
1!
b0 %
1'
b0 +
#560010000000
0!
0'
#560020000000
1!
1$
b1 %
1'
1*
b1 +
#560030000000
0!
0'
#560040000000
1!
b10 %
1'
b10 +
#560050000000
0!
0'
#560060000000
1!
b11 %
1'
b11 +
#560070000000
1"
1(
#560080000000
0!
0"
b100 &
0'
0(
b100 ,
#560090000000
1!
b100 %
1'
b100 +
#560100000000
0!
0'
#560110000000
1!
b101 %
1'
b101 +
#560120000000
0!
0'
#560130000000
1!
b110 %
1'
b110 +
#560140000000
0!
0'
#560150000000
1!
b111 %
1'
b111 +
#560160000000
0!
0'
#560170000000
1!
0$
b1000 %
1'
0*
b1000 +
#560180000000
0!
0'
#560190000000
1!
b1001 %
1'
b1001 +
#560200000000
0!
0'
#560210000000
1!
b0 %
1'
b0 +
#560220000000
0!
0'
#560230000000
1!
1$
b1 %
1'
1*
b1 +
#560240000000
0!
0'
#560250000000
1!
b10 %
1'
b10 +
#560260000000
0!
0'
#560270000000
1!
b11 %
1'
b11 +
#560280000000
0!
0'
#560290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#560300000000
0!
0'
#560310000000
1!
b101 %
1'
b101 +
#560320000000
0!
0'
#560330000000
1!
0$
b110 %
1'
0*
b110 +
#560340000000
0!
0'
#560350000000
1!
b111 %
1'
b111 +
#560360000000
0!
0'
#560370000000
1!
b1000 %
1'
b1000 +
#560380000000
0!
0'
#560390000000
1!
b1001 %
1'
b1001 +
#560400000000
0!
0'
#560410000000
1!
b0 %
1'
b0 +
#560420000000
0!
0'
#560430000000
1!
1$
b1 %
1'
1*
b1 +
#560440000000
0!
0'
#560450000000
1!
b10 %
1'
b10 +
#560460000000
0!
0'
#560470000000
1!
b11 %
1'
b11 +
#560480000000
0!
0'
#560490000000
1!
b100 %
1'
b100 +
#560500000000
1"
1(
#560510000000
0!
0"
b100 &
0'
0(
b100 ,
#560520000000
1!
b101 %
1'
b101 +
#560530000000
0!
0'
#560540000000
1!
b110 %
1'
b110 +
#560550000000
0!
0'
#560560000000
1!
b111 %
1'
b111 +
#560570000000
0!
0'
#560580000000
1!
0$
b1000 %
1'
0*
b1000 +
#560590000000
0!
0'
#560600000000
1!
b1001 %
1'
b1001 +
#560610000000
0!
0'
#560620000000
1!
b0 %
1'
b0 +
#560630000000
0!
0'
#560640000000
1!
1$
b1 %
1'
1*
b1 +
#560650000000
0!
0'
#560660000000
1!
b10 %
1'
b10 +
#560670000000
0!
0'
#560680000000
1!
b11 %
1'
b11 +
#560690000000
0!
0'
#560700000000
1!
b100 %
1'
b100 +
#560710000000
0!
0'
#560720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#560730000000
0!
0'
#560740000000
1!
0$
b110 %
1'
0*
b110 +
#560750000000
0!
0'
#560760000000
1!
b111 %
1'
b111 +
#560770000000
0!
0'
#560780000000
1!
b1000 %
1'
b1000 +
#560790000000
0!
0'
#560800000000
1!
b1001 %
1'
b1001 +
#560810000000
0!
0'
#560820000000
1!
b0 %
1'
b0 +
#560830000000
0!
0'
#560840000000
1!
1$
b1 %
1'
1*
b1 +
#560850000000
0!
0'
#560860000000
1!
b10 %
1'
b10 +
#560870000000
0!
0'
#560880000000
1!
b11 %
1'
b11 +
#560890000000
0!
0'
#560900000000
1!
b100 %
1'
b100 +
#560910000000
0!
0'
#560920000000
1!
b101 %
1'
b101 +
#560930000000
1"
1(
#560940000000
0!
0"
b100 &
0'
0(
b100 ,
#560950000000
1!
b110 %
1'
b110 +
#560960000000
0!
0'
#560970000000
1!
b111 %
1'
b111 +
#560980000000
0!
0'
#560990000000
1!
0$
b1000 %
1'
0*
b1000 +
#561000000000
0!
0'
#561010000000
1!
b1001 %
1'
b1001 +
#561020000000
0!
0'
#561030000000
1!
b0 %
1'
b0 +
#561040000000
0!
0'
#561050000000
1!
1$
b1 %
1'
1*
b1 +
#561060000000
0!
0'
#561070000000
1!
b10 %
1'
b10 +
#561080000000
0!
0'
#561090000000
1!
b11 %
1'
b11 +
#561100000000
0!
0'
#561110000000
1!
b100 %
1'
b100 +
#561120000000
0!
0'
#561130000000
1!
b101 %
1'
b101 +
#561140000000
0!
0'
#561150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#561160000000
0!
0'
#561170000000
1!
b111 %
1'
b111 +
#561180000000
0!
0'
#561190000000
1!
b1000 %
1'
b1000 +
#561200000000
0!
0'
#561210000000
1!
b1001 %
1'
b1001 +
#561220000000
0!
0'
#561230000000
1!
b0 %
1'
b0 +
#561240000000
0!
0'
#561250000000
1!
1$
b1 %
1'
1*
b1 +
#561260000000
0!
0'
#561270000000
1!
b10 %
1'
b10 +
#561280000000
0!
0'
#561290000000
1!
b11 %
1'
b11 +
#561300000000
0!
0'
#561310000000
1!
b100 %
1'
b100 +
#561320000000
0!
0'
#561330000000
1!
b101 %
1'
b101 +
#561340000000
0!
0'
#561350000000
1!
0$
b110 %
1'
0*
b110 +
#561360000000
1"
1(
#561370000000
0!
0"
b100 &
0'
0(
b100 ,
#561380000000
1!
1$
b111 %
1'
1*
b111 +
#561390000000
0!
0'
#561400000000
1!
0$
b1000 %
1'
0*
b1000 +
#561410000000
0!
0'
#561420000000
1!
b1001 %
1'
b1001 +
#561430000000
0!
0'
#561440000000
1!
b0 %
1'
b0 +
#561450000000
0!
0'
#561460000000
1!
1$
b1 %
1'
1*
b1 +
#561470000000
0!
0'
#561480000000
1!
b10 %
1'
b10 +
#561490000000
0!
0'
#561500000000
1!
b11 %
1'
b11 +
#561510000000
0!
0'
#561520000000
1!
b100 %
1'
b100 +
#561530000000
0!
0'
#561540000000
1!
b101 %
1'
b101 +
#561550000000
0!
0'
#561560000000
1!
b110 %
1'
b110 +
#561570000000
0!
0'
#561580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#561590000000
0!
0'
#561600000000
1!
b1000 %
1'
b1000 +
#561610000000
0!
0'
#561620000000
1!
b1001 %
1'
b1001 +
#561630000000
0!
0'
#561640000000
1!
b0 %
1'
b0 +
#561650000000
0!
0'
#561660000000
1!
1$
b1 %
1'
1*
b1 +
#561670000000
0!
0'
#561680000000
1!
b10 %
1'
b10 +
#561690000000
0!
0'
#561700000000
1!
b11 %
1'
b11 +
#561710000000
0!
0'
#561720000000
1!
b100 %
1'
b100 +
#561730000000
0!
0'
#561740000000
1!
b101 %
1'
b101 +
#561750000000
0!
0'
#561760000000
1!
0$
b110 %
1'
0*
b110 +
#561770000000
0!
0'
#561780000000
1!
b111 %
1'
b111 +
#561790000000
1"
1(
#561800000000
0!
0"
b100 &
0'
0(
b100 ,
#561810000000
1!
b1000 %
1'
b1000 +
#561820000000
0!
0'
#561830000000
1!
b1001 %
1'
b1001 +
#561840000000
0!
0'
#561850000000
1!
b0 %
1'
b0 +
#561860000000
0!
0'
#561870000000
1!
1$
b1 %
1'
1*
b1 +
#561880000000
0!
0'
#561890000000
1!
b10 %
1'
b10 +
#561900000000
0!
0'
#561910000000
1!
b11 %
1'
b11 +
#561920000000
0!
0'
#561930000000
1!
b100 %
1'
b100 +
#561940000000
0!
0'
#561950000000
1!
b101 %
1'
b101 +
#561960000000
0!
0'
#561970000000
1!
b110 %
1'
b110 +
#561980000000
0!
0'
#561990000000
1!
b111 %
1'
b111 +
#562000000000
0!
0'
#562010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#562020000000
0!
0'
#562030000000
1!
b1001 %
1'
b1001 +
#562040000000
0!
0'
#562050000000
1!
b0 %
1'
b0 +
#562060000000
0!
0'
#562070000000
1!
1$
b1 %
1'
1*
b1 +
#562080000000
0!
0'
#562090000000
1!
b10 %
1'
b10 +
#562100000000
0!
0'
#562110000000
1!
b11 %
1'
b11 +
#562120000000
0!
0'
#562130000000
1!
b100 %
1'
b100 +
#562140000000
0!
0'
#562150000000
1!
b101 %
1'
b101 +
#562160000000
0!
0'
#562170000000
1!
0$
b110 %
1'
0*
b110 +
#562180000000
0!
0'
#562190000000
1!
b111 %
1'
b111 +
#562200000000
0!
0'
#562210000000
1!
b1000 %
1'
b1000 +
#562220000000
1"
1(
#562230000000
0!
0"
b100 &
0'
0(
b100 ,
#562240000000
1!
b1001 %
1'
b1001 +
#562250000000
0!
0'
#562260000000
1!
b0 %
1'
b0 +
#562270000000
0!
0'
#562280000000
1!
1$
b1 %
1'
1*
b1 +
#562290000000
0!
0'
#562300000000
1!
b10 %
1'
b10 +
#562310000000
0!
0'
#562320000000
1!
b11 %
1'
b11 +
#562330000000
0!
0'
#562340000000
1!
b100 %
1'
b100 +
#562350000000
0!
0'
#562360000000
1!
b101 %
1'
b101 +
#562370000000
0!
0'
#562380000000
1!
b110 %
1'
b110 +
#562390000000
0!
0'
#562400000000
1!
b111 %
1'
b111 +
#562410000000
0!
0'
#562420000000
1!
0$
b1000 %
1'
0*
b1000 +
#562430000000
0!
0'
#562440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#562450000000
0!
0'
#562460000000
1!
b0 %
1'
b0 +
#562470000000
0!
0'
#562480000000
1!
1$
b1 %
1'
1*
b1 +
#562490000000
0!
0'
#562500000000
1!
b10 %
1'
b10 +
#562510000000
0!
0'
#562520000000
1!
b11 %
1'
b11 +
#562530000000
0!
0'
#562540000000
1!
b100 %
1'
b100 +
#562550000000
0!
0'
#562560000000
1!
b101 %
1'
b101 +
#562570000000
0!
0'
#562580000000
1!
0$
b110 %
1'
0*
b110 +
#562590000000
0!
0'
#562600000000
1!
b111 %
1'
b111 +
#562610000000
0!
0'
#562620000000
1!
b1000 %
1'
b1000 +
#562630000000
0!
0'
#562640000000
1!
b1001 %
1'
b1001 +
#562650000000
1"
1(
#562660000000
0!
0"
b100 &
0'
0(
b100 ,
#562670000000
1!
b0 %
1'
b0 +
#562680000000
0!
0'
#562690000000
1!
1$
b1 %
1'
1*
b1 +
#562700000000
0!
0'
#562710000000
1!
b10 %
1'
b10 +
#562720000000
0!
0'
#562730000000
1!
b11 %
1'
b11 +
#562740000000
0!
0'
#562750000000
1!
b100 %
1'
b100 +
#562760000000
0!
0'
#562770000000
1!
b101 %
1'
b101 +
#562780000000
0!
0'
#562790000000
1!
b110 %
1'
b110 +
#562800000000
0!
0'
#562810000000
1!
b111 %
1'
b111 +
#562820000000
0!
0'
#562830000000
1!
0$
b1000 %
1'
0*
b1000 +
#562840000000
0!
0'
#562850000000
1!
b1001 %
1'
b1001 +
#562860000000
0!
0'
#562870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#562880000000
0!
0'
#562890000000
1!
1$
b1 %
1'
1*
b1 +
#562900000000
0!
0'
#562910000000
1!
b10 %
1'
b10 +
#562920000000
0!
0'
#562930000000
1!
b11 %
1'
b11 +
#562940000000
0!
0'
#562950000000
1!
b100 %
1'
b100 +
#562960000000
0!
0'
#562970000000
1!
b101 %
1'
b101 +
#562980000000
0!
0'
#562990000000
1!
0$
b110 %
1'
0*
b110 +
#563000000000
0!
0'
#563010000000
1!
b111 %
1'
b111 +
#563020000000
0!
0'
#563030000000
1!
b1000 %
1'
b1000 +
#563040000000
0!
0'
#563050000000
1!
b1001 %
1'
b1001 +
#563060000000
0!
0'
#563070000000
1!
b0 %
1'
b0 +
#563080000000
1"
1(
#563090000000
0!
0"
b100 &
0'
0(
b100 ,
#563100000000
1!
1$
b1 %
1'
1*
b1 +
#563110000000
0!
0'
#563120000000
1!
b10 %
1'
b10 +
#563130000000
0!
0'
#563140000000
1!
b11 %
1'
b11 +
#563150000000
0!
0'
#563160000000
1!
b100 %
1'
b100 +
#563170000000
0!
0'
#563180000000
1!
b101 %
1'
b101 +
#563190000000
0!
0'
#563200000000
1!
b110 %
1'
b110 +
#563210000000
0!
0'
#563220000000
1!
b111 %
1'
b111 +
#563230000000
0!
0'
#563240000000
1!
0$
b1000 %
1'
0*
b1000 +
#563250000000
0!
0'
#563260000000
1!
b1001 %
1'
b1001 +
#563270000000
0!
0'
#563280000000
1!
b0 %
1'
b0 +
#563290000000
0!
0'
#563300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#563310000000
0!
0'
#563320000000
1!
b10 %
1'
b10 +
#563330000000
0!
0'
#563340000000
1!
b11 %
1'
b11 +
#563350000000
0!
0'
#563360000000
1!
b100 %
1'
b100 +
#563370000000
0!
0'
#563380000000
1!
b101 %
1'
b101 +
#563390000000
0!
0'
#563400000000
1!
0$
b110 %
1'
0*
b110 +
#563410000000
0!
0'
#563420000000
1!
b111 %
1'
b111 +
#563430000000
0!
0'
#563440000000
1!
b1000 %
1'
b1000 +
#563450000000
0!
0'
#563460000000
1!
b1001 %
1'
b1001 +
#563470000000
0!
0'
#563480000000
1!
b0 %
1'
b0 +
#563490000000
0!
0'
#563500000000
1!
1$
b1 %
1'
1*
b1 +
#563510000000
1"
1(
#563520000000
0!
0"
b100 &
0'
0(
b100 ,
#563530000000
1!
b10 %
1'
b10 +
#563540000000
0!
0'
#563550000000
1!
b11 %
1'
b11 +
#563560000000
0!
0'
#563570000000
1!
b100 %
1'
b100 +
#563580000000
0!
0'
#563590000000
1!
b101 %
1'
b101 +
#563600000000
0!
0'
#563610000000
1!
b110 %
1'
b110 +
#563620000000
0!
0'
#563630000000
1!
b111 %
1'
b111 +
#563640000000
0!
0'
#563650000000
1!
0$
b1000 %
1'
0*
b1000 +
#563660000000
0!
0'
#563670000000
1!
b1001 %
1'
b1001 +
#563680000000
0!
0'
#563690000000
1!
b0 %
1'
b0 +
#563700000000
0!
0'
#563710000000
1!
1$
b1 %
1'
1*
b1 +
#563720000000
0!
0'
#563730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#563740000000
0!
0'
#563750000000
1!
b11 %
1'
b11 +
#563760000000
0!
0'
#563770000000
1!
b100 %
1'
b100 +
#563780000000
0!
0'
#563790000000
1!
b101 %
1'
b101 +
#563800000000
0!
0'
#563810000000
1!
0$
b110 %
1'
0*
b110 +
#563820000000
0!
0'
#563830000000
1!
b111 %
1'
b111 +
#563840000000
0!
0'
#563850000000
1!
b1000 %
1'
b1000 +
#563860000000
0!
0'
#563870000000
1!
b1001 %
1'
b1001 +
#563880000000
0!
0'
#563890000000
1!
b0 %
1'
b0 +
#563900000000
0!
0'
#563910000000
1!
1$
b1 %
1'
1*
b1 +
#563920000000
0!
0'
#563930000000
1!
b10 %
1'
b10 +
#563940000000
1"
1(
#563950000000
0!
0"
b100 &
0'
0(
b100 ,
#563960000000
1!
b11 %
1'
b11 +
#563970000000
0!
0'
#563980000000
1!
b100 %
1'
b100 +
#563990000000
0!
0'
#564000000000
1!
b101 %
1'
b101 +
#564010000000
0!
0'
#564020000000
1!
b110 %
1'
b110 +
#564030000000
0!
0'
#564040000000
1!
b111 %
1'
b111 +
#564050000000
0!
0'
#564060000000
1!
0$
b1000 %
1'
0*
b1000 +
#564070000000
0!
0'
#564080000000
1!
b1001 %
1'
b1001 +
#564090000000
0!
0'
#564100000000
1!
b0 %
1'
b0 +
#564110000000
0!
0'
#564120000000
1!
1$
b1 %
1'
1*
b1 +
#564130000000
0!
0'
#564140000000
1!
b10 %
1'
b10 +
#564150000000
0!
0'
#564160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#564170000000
0!
0'
#564180000000
1!
b100 %
1'
b100 +
#564190000000
0!
0'
#564200000000
1!
b101 %
1'
b101 +
#564210000000
0!
0'
#564220000000
1!
0$
b110 %
1'
0*
b110 +
#564230000000
0!
0'
#564240000000
1!
b111 %
1'
b111 +
#564250000000
0!
0'
#564260000000
1!
b1000 %
1'
b1000 +
#564270000000
0!
0'
#564280000000
1!
b1001 %
1'
b1001 +
#564290000000
0!
0'
#564300000000
1!
b0 %
1'
b0 +
#564310000000
0!
0'
#564320000000
1!
1$
b1 %
1'
1*
b1 +
#564330000000
0!
0'
#564340000000
1!
b10 %
1'
b10 +
#564350000000
0!
0'
#564360000000
1!
b11 %
1'
b11 +
#564370000000
1"
1(
#564380000000
0!
0"
b100 &
0'
0(
b100 ,
#564390000000
1!
b100 %
1'
b100 +
#564400000000
0!
0'
#564410000000
1!
b101 %
1'
b101 +
#564420000000
0!
0'
#564430000000
1!
b110 %
1'
b110 +
#564440000000
0!
0'
#564450000000
1!
b111 %
1'
b111 +
#564460000000
0!
0'
#564470000000
1!
0$
b1000 %
1'
0*
b1000 +
#564480000000
0!
0'
#564490000000
1!
b1001 %
1'
b1001 +
#564500000000
0!
0'
#564510000000
1!
b0 %
1'
b0 +
#564520000000
0!
0'
#564530000000
1!
1$
b1 %
1'
1*
b1 +
#564540000000
0!
0'
#564550000000
1!
b10 %
1'
b10 +
#564560000000
0!
0'
#564570000000
1!
b11 %
1'
b11 +
#564580000000
0!
0'
#564590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#564600000000
0!
0'
#564610000000
1!
b101 %
1'
b101 +
#564620000000
0!
0'
#564630000000
1!
0$
b110 %
1'
0*
b110 +
#564640000000
0!
0'
#564650000000
1!
b111 %
1'
b111 +
#564660000000
0!
0'
#564670000000
1!
b1000 %
1'
b1000 +
#564680000000
0!
0'
#564690000000
1!
b1001 %
1'
b1001 +
#564700000000
0!
0'
#564710000000
1!
b0 %
1'
b0 +
#564720000000
0!
0'
#564730000000
1!
1$
b1 %
1'
1*
b1 +
#564740000000
0!
0'
#564750000000
1!
b10 %
1'
b10 +
#564760000000
0!
0'
#564770000000
1!
b11 %
1'
b11 +
#564780000000
0!
0'
#564790000000
1!
b100 %
1'
b100 +
#564800000000
1"
1(
#564810000000
0!
0"
b100 &
0'
0(
b100 ,
#564820000000
1!
b101 %
1'
b101 +
#564830000000
0!
0'
#564840000000
1!
b110 %
1'
b110 +
#564850000000
0!
0'
#564860000000
1!
b111 %
1'
b111 +
#564870000000
0!
0'
#564880000000
1!
0$
b1000 %
1'
0*
b1000 +
#564890000000
0!
0'
#564900000000
1!
b1001 %
1'
b1001 +
#564910000000
0!
0'
#564920000000
1!
b0 %
1'
b0 +
#564930000000
0!
0'
#564940000000
1!
1$
b1 %
1'
1*
b1 +
#564950000000
0!
0'
#564960000000
1!
b10 %
1'
b10 +
#564970000000
0!
0'
#564980000000
1!
b11 %
1'
b11 +
#564990000000
0!
0'
#565000000000
1!
b100 %
1'
b100 +
#565010000000
0!
0'
#565020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#565030000000
0!
0'
#565040000000
1!
0$
b110 %
1'
0*
b110 +
#565050000000
0!
0'
#565060000000
1!
b111 %
1'
b111 +
#565070000000
0!
0'
#565080000000
1!
b1000 %
1'
b1000 +
#565090000000
0!
0'
#565100000000
1!
b1001 %
1'
b1001 +
#565110000000
0!
0'
#565120000000
1!
b0 %
1'
b0 +
#565130000000
0!
0'
#565140000000
1!
1$
b1 %
1'
1*
b1 +
#565150000000
0!
0'
#565160000000
1!
b10 %
1'
b10 +
#565170000000
0!
0'
#565180000000
1!
b11 %
1'
b11 +
#565190000000
0!
0'
#565200000000
1!
b100 %
1'
b100 +
#565210000000
0!
0'
#565220000000
1!
b101 %
1'
b101 +
#565230000000
1"
1(
#565240000000
0!
0"
b100 &
0'
0(
b100 ,
#565250000000
1!
b110 %
1'
b110 +
#565260000000
0!
0'
#565270000000
1!
b111 %
1'
b111 +
#565280000000
0!
0'
#565290000000
1!
0$
b1000 %
1'
0*
b1000 +
#565300000000
0!
0'
#565310000000
1!
b1001 %
1'
b1001 +
#565320000000
0!
0'
#565330000000
1!
b0 %
1'
b0 +
#565340000000
0!
0'
#565350000000
1!
1$
b1 %
1'
1*
b1 +
#565360000000
0!
0'
#565370000000
1!
b10 %
1'
b10 +
#565380000000
0!
0'
#565390000000
1!
b11 %
1'
b11 +
#565400000000
0!
0'
#565410000000
1!
b100 %
1'
b100 +
#565420000000
0!
0'
#565430000000
1!
b101 %
1'
b101 +
#565440000000
0!
0'
#565450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#565460000000
0!
0'
#565470000000
1!
b111 %
1'
b111 +
#565480000000
0!
0'
#565490000000
1!
b1000 %
1'
b1000 +
#565500000000
0!
0'
#565510000000
1!
b1001 %
1'
b1001 +
#565520000000
0!
0'
#565530000000
1!
b0 %
1'
b0 +
#565540000000
0!
0'
#565550000000
1!
1$
b1 %
1'
1*
b1 +
#565560000000
0!
0'
#565570000000
1!
b10 %
1'
b10 +
#565580000000
0!
0'
#565590000000
1!
b11 %
1'
b11 +
#565600000000
0!
0'
#565610000000
1!
b100 %
1'
b100 +
#565620000000
0!
0'
#565630000000
1!
b101 %
1'
b101 +
#565640000000
0!
0'
#565650000000
1!
0$
b110 %
1'
0*
b110 +
#565660000000
1"
1(
#565670000000
0!
0"
b100 &
0'
0(
b100 ,
#565680000000
1!
1$
b111 %
1'
1*
b111 +
#565690000000
0!
0'
#565700000000
1!
0$
b1000 %
1'
0*
b1000 +
#565710000000
0!
0'
#565720000000
1!
b1001 %
1'
b1001 +
#565730000000
0!
0'
#565740000000
1!
b0 %
1'
b0 +
#565750000000
0!
0'
#565760000000
1!
1$
b1 %
1'
1*
b1 +
#565770000000
0!
0'
#565780000000
1!
b10 %
1'
b10 +
#565790000000
0!
0'
#565800000000
1!
b11 %
1'
b11 +
#565810000000
0!
0'
#565820000000
1!
b100 %
1'
b100 +
#565830000000
0!
0'
#565840000000
1!
b101 %
1'
b101 +
#565850000000
0!
0'
#565860000000
1!
b110 %
1'
b110 +
#565870000000
0!
0'
#565880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#565890000000
0!
0'
#565900000000
1!
b1000 %
1'
b1000 +
#565910000000
0!
0'
#565920000000
1!
b1001 %
1'
b1001 +
#565930000000
0!
0'
#565940000000
1!
b0 %
1'
b0 +
#565950000000
0!
0'
#565960000000
1!
1$
b1 %
1'
1*
b1 +
#565970000000
0!
0'
#565980000000
1!
b10 %
1'
b10 +
#565990000000
0!
0'
#566000000000
1!
b11 %
1'
b11 +
#566010000000
0!
0'
#566020000000
1!
b100 %
1'
b100 +
#566030000000
0!
0'
#566040000000
1!
b101 %
1'
b101 +
#566050000000
0!
0'
#566060000000
1!
0$
b110 %
1'
0*
b110 +
#566070000000
0!
0'
#566080000000
1!
b111 %
1'
b111 +
#566090000000
1"
1(
#566100000000
0!
0"
b100 &
0'
0(
b100 ,
#566110000000
1!
b1000 %
1'
b1000 +
#566120000000
0!
0'
#566130000000
1!
b1001 %
1'
b1001 +
#566140000000
0!
0'
#566150000000
1!
b0 %
1'
b0 +
#566160000000
0!
0'
#566170000000
1!
1$
b1 %
1'
1*
b1 +
#566180000000
0!
0'
#566190000000
1!
b10 %
1'
b10 +
#566200000000
0!
0'
#566210000000
1!
b11 %
1'
b11 +
#566220000000
0!
0'
#566230000000
1!
b100 %
1'
b100 +
#566240000000
0!
0'
#566250000000
1!
b101 %
1'
b101 +
#566260000000
0!
0'
#566270000000
1!
b110 %
1'
b110 +
#566280000000
0!
0'
#566290000000
1!
b111 %
1'
b111 +
#566300000000
0!
0'
#566310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#566320000000
0!
0'
#566330000000
1!
b1001 %
1'
b1001 +
#566340000000
0!
0'
#566350000000
1!
b0 %
1'
b0 +
#566360000000
0!
0'
#566370000000
1!
1$
b1 %
1'
1*
b1 +
#566380000000
0!
0'
#566390000000
1!
b10 %
1'
b10 +
#566400000000
0!
0'
#566410000000
1!
b11 %
1'
b11 +
#566420000000
0!
0'
#566430000000
1!
b100 %
1'
b100 +
#566440000000
0!
0'
#566450000000
1!
b101 %
1'
b101 +
#566460000000
0!
0'
#566470000000
1!
0$
b110 %
1'
0*
b110 +
#566480000000
0!
0'
#566490000000
1!
b111 %
1'
b111 +
#566500000000
0!
0'
#566510000000
1!
b1000 %
1'
b1000 +
#566520000000
1"
1(
#566530000000
0!
0"
b100 &
0'
0(
b100 ,
#566540000000
1!
b1001 %
1'
b1001 +
#566550000000
0!
0'
#566560000000
1!
b0 %
1'
b0 +
#566570000000
0!
0'
#566580000000
1!
1$
b1 %
1'
1*
b1 +
#566590000000
0!
0'
#566600000000
1!
b10 %
1'
b10 +
#566610000000
0!
0'
#566620000000
1!
b11 %
1'
b11 +
#566630000000
0!
0'
#566640000000
1!
b100 %
1'
b100 +
#566650000000
0!
0'
#566660000000
1!
b101 %
1'
b101 +
#566670000000
0!
0'
#566680000000
1!
b110 %
1'
b110 +
#566690000000
0!
0'
#566700000000
1!
b111 %
1'
b111 +
#566710000000
0!
0'
#566720000000
1!
0$
b1000 %
1'
0*
b1000 +
#566730000000
0!
0'
#566740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#566750000000
0!
0'
#566760000000
1!
b0 %
1'
b0 +
#566770000000
0!
0'
#566780000000
1!
1$
b1 %
1'
1*
b1 +
#566790000000
0!
0'
#566800000000
1!
b10 %
1'
b10 +
#566810000000
0!
0'
#566820000000
1!
b11 %
1'
b11 +
#566830000000
0!
0'
#566840000000
1!
b100 %
1'
b100 +
#566850000000
0!
0'
#566860000000
1!
b101 %
1'
b101 +
#566870000000
0!
0'
#566880000000
1!
0$
b110 %
1'
0*
b110 +
#566890000000
0!
0'
#566900000000
1!
b111 %
1'
b111 +
#566910000000
0!
0'
#566920000000
1!
b1000 %
1'
b1000 +
#566930000000
0!
0'
#566940000000
1!
b1001 %
1'
b1001 +
#566950000000
1"
1(
#566960000000
0!
0"
b100 &
0'
0(
b100 ,
#566970000000
1!
b0 %
1'
b0 +
#566980000000
0!
0'
#566990000000
1!
1$
b1 %
1'
1*
b1 +
#567000000000
0!
0'
#567010000000
1!
b10 %
1'
b10 +
#567020000000
0!
0'
#567030000000
1!
b11 %
1'
b11 +
#567040000000
0!
0'
#567050000000
1!
b100 %
1'
b100 +
#567060000000
0!
0'
#567070000000
1!
b101 %
1'
b101 +
#567080000000
0!
0'
#567090000000
1!
b110 %
1'
b110 +
#567100000000
0!
0'
#567110000000
1!
b111 %
1'
b111 +
#567120000000
0!
0'
#567130000000
1!
0$
b1000 %
1'
0*
b1000 +
#567140000000
0!
0'
#567150000000
1!
b1001 %
1'
b1001 +
#567160000000
0!
0'
#567170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#567180000000
0!
0'
#567190000000
1!
1$
b1 %
1'
1*
b1 +
#567200000000
0!
0'
#567210000000
1!
b10 %
1'
b10 +
#567220000000
0!
0'
#567230000000
1!
b11 %
1'
b11 +
#567240000000
0!
0'
#567250000000
1!
b100 %
1'
b100 +
#567260000000
0!
0'
#567270000000
1!
b101 %
1'
b101 +
#567280000000
0!
0'
#567290000000
1!
0$
b110 %
1'
0*
b110 +
#567300000000
0!
0'
#567310000000
1!
b111 %
1'
b111 +
#567320000000
0!
0'
#567330000000
1!
b1000 %
1'
b1000 +
#567340000000
0!
0'
#567350000000
1!
b1001 %
1'
b1001 +
#567360000000
0!
0'
#567370000000
1!
b0 %
1'
b0 +
#567380000000
1"
1(
#567390000000
0!
0"
b100 &
0'
0(
b100 ,
#567400000000
1!
1$
b1 %
1'
1*
b1 +
#567410000000
0!
0'
#567420000000
1!
b10 %
1'
b10 +
#567430000000
0!
0'
#567440000000
1!
b11 %
1'
b11 +
#567450000000
0!
0'
#567460000000
1!
b100 %
1'
b100 +
#567470000000
0!
0'
#567480000000
1!
b101 %
1'
b101 +
#567490000000
0!
0'
#567500000000
1!
b110 %
1'
b110 +
#567510000000
0!
0'
#567520000000
1!
b111 %
1'
b111 +
#567530000000
0!
0'
#567540000000
1!
0$
b1000 %
1'
0*
b1000 +
#567550000000
0!
0'
#567560000000
1!
b1001 %
1'
b1001 +
#567570000000
0!
0'
#567580000000
1!
b0 %
1'
b0 +
#567590000000
0!
0'
#567600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#567610000000
0!
0'
#567620000000
1!
b10 %
1'
b10 +
#567630000000
0!
0'
#567640000000
1!
b11 %
1'
b11 +
#567650000000
0!
0'
#567660000000
1!
b100 %
1'
b100 +
#567670000000
0!
0'
#567680000000
1!
b101 %
1'
b101 +
#567690000000
0!
0'
#567700000000
1!
0$
b110 %
1'
0*
b110 +
#567710000000
0!
0'
#567720000000
1!
b111 %
1'
b111 +
#567730000000
0!
0'
#567740000000
1!
b1000 %
1'
b1000 +
#567750000000
0!
0'
#567760000000
1!
b1001 %
1'
b1001 +
#567770000000
0!
0'
#567780000000
1!
b0 %
1'
b0 +
#567790000000
0!
0'
#567800000000
1!
1$
b1 %
1'
1*
b1 +
#567810000000
1"
1(
#567820000000
0!
0"
b100 &
0'
0(
b100 ,
#567830000000
1!
b10 %
1'
b10 +
#567840000000
0!
0'
#567850000000
1!
b11 %
1'
b11 +
#567860000000
0!
0'
#567870000000
1!
b100 %
1'
b100 +
#567880000000
0!
0'
#567890000000
1!
b101 %
1'
b101 +
#567900000000
0!
0'
#567910000000
1!
b110 %
1'
b110 +
#567920000000
0!
0'
#567930000000
1!
b111 %
1'
b111 +
#567940000000
0!
0'
#567950000000
1!
0$
b1000 %
1'
0*
b1000 +
#567960000000
0!
0'
#567970000000
1!
b1001 %
1'
b1001 +
#567980000000
0!
0'
#567990000000
1!
b0 %
1'
b0 +
#568000000000
0!
0'
#568010000000
1!
1$
b1 %
1'
1*
b1 +
#568020000000
0!
0'
#568030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#568040000000
0!
0'
#568050000000
1!
b11 %
1'
b11 +
#568060000000
0!
0'
#568070000000
1!
b100 %
1'
b100 +
#568080000000
0!
0'
#568090000000
1!
b101 %
1'
b101 +
#568100000000
0!
0'
#568110000000
1!
0$
b110 %
1'
0*
b110 +
#568120000000
0!
0'
#568130000000
1!
b111 %
1'
b111 +
#568140000000
0!
0'
#568150000000
1!
b1000 %
1'
b1000 +
#568160000000
0!
0'
#568170000000
1!
b1001 %
1'
b1001 +
#568180000000
0!
0'
#568190000000
1!
b0 %
1'
b0 +
#568200000000
0!
0'
#568210000000
1!
1$
b1 %
1'
1*
b1 +
#568220000000
0!
0'
#568230000000
1!
b10 %
1'
b10 +
#568240000000
1"
1(
#568250000000
0!
0"
b100 &
0'
0(
b100 ,
#568260000000
1!
b11 %
1'
b11 +
#568270000000
0!
0'
#568280000000
1!
b100 %
1'
b100 +
#568290000000
0!
0'
#568300000000
1!
b101 %
1'
b101 +
#568310000000
0!
0'
#568320000000
1!
b110 %
1'
b110 +
#568330000000
0!
0'
#568340000000
1!
b111 %
1'
b111 +
#568350000000
0!
0'
#568360000000
1!
0$
b1000 %
1'
0*
b1000 +
#568370000000
0!
0'
#568380000000
1!
b1001 %
1'
b1001 +
#568390000000
0!
0'
#568400000000
1!
b0 %
1'
b0 +
#568410000000
0!
0'
#568420000000
1!
1$
b1 %
1'
1*
b1 +
#568430000000
0!
0'
#568440000000
1!
b10 %
1'
b10 +
#568450000000
0!
0'
#568460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#568470000000
0!
0'
#568480000000
1!
b100 %
1'
b100 +
#568490000000
0!
0'
#568500000000
1!
b101 %
1'
b101 +
#568510000000
0!
0'
#568520000000
1!
0$
b110 %
1'
0*
b110 +
#568530000000
0!
0'
#568540000000
1!
b111 %
1'
b111 +
#568550000000
0!
0'
#568560000000
1!
b1000 %
1'
b1000 +
#568570000000
0!
0'
#568580000000
1!
b1001 %
1'
b1001 +
#568590000000
0!
0'
#568600000000
1!
b0 %
1'
b0 +
#568610000000
0!
0'
#568620000000
1!
1$
b1 %
1'
1*
b1 +
#568630000000
0!
0'
#568640000000
1!
b10 %
1'
b10 +
#568650000000
0!
0'
#568660000000
1!
b11 %
1'
b11 +
#568670000000
1"
1(
#568680000000
0!
0"
b100 &
0'
0(
b100 ,
#568690000000
1!
b100 %
1'
b100 +
#568700000000
0!
0'
#568710000000
1!
b101 %
1'
b101 +
#568720000000
0!
0'
#568730000000
1!
b110 %
1'
b110 +
#568740000000
0!
0'
#568750000000
1!
b111 %
1'
b111 +
#568760000000
0!
0'
#568770000000
1!
0$
b1000 %
1'
0*
b1000 +
#568780000000
0!
0'
#568790000000
1!
b1001 %
1'
b1001 +
#568800000000
0!
0'
#568810000000
1!
b0 %
1'
b0 +
#568820000000
0!
0'
#568830000000
1!
1$
b1 %
1'
1*
b1 +
#568840000000
0!
0'
#568850000000
1!
b10 %
1'
b10 +
#568860000000
0!
0'
#568870000000
1!
b11 %
1'
b11 +
#568880000000
0!
0'
#568890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#568900000000
0!
0'
#568910000000
1!
b101 %
1'
b101 +
#568920000000
0!
0'
#568930000000
1!
0$
b110 %
1'
0*
b110 +
#568940000000
0!
0'
#568950000000
1!
b111 %
1'
b111 +
#568960000000
0!
0'
#568970000000
1!
b1000 %
1'
b1000 +
#568980000000
0!
0'
#568990000000
1!
b1001 %
1'
b1001 +
#569000000000
0!
0'
#569010000000
1!
b0 %
1'
b0 +
#569020000000
0!
0'
#569030000000
1!
1$
b1 %
1'
1*
b1 +
#569040000000
0!
0'
#569050000000
1!
b10 %
1'
b10 +
#569060000000
0!
0'
#569070000000
1!
b11 %
1'
b11 +
#569080000000
0!
0'
#569090000000
1!
b100 %
1'
b100 +
#569100000000
1"
1(
#569110000000
0!
0"
b100 &
0'
0(
b100 ,
#569120000000
1!
b101 %
1'
b101 +
#569130000000
0!
0'
#569140000000
1!
b110 %
1'
b110 +
#569150000000
0!
0'
#569160000000
1!
b111 %
1'
b111 +
#569170000000
0!
0'
#569180000000
1!
0$
b1000 %
1'
0*
b1000 +
#569190000000
0!
0'
#569200000000
1!
b1001 %
1'
b1001 +
#569210000000
0!
0'
#569220000000
1!
b0 %
1'
b0 +
#569230000000
0!
0'
#569240000000
1!
1$
b1 %
1'
1*
b1 +
#569250000000
0!
0'
#569260000000
1!
b10 %
1'
b10 +
#569270000000
0!
0'
#569280000000
1!
b11 %
1'
b11 +
#569290000000
0!
0'
#569300000000
1!
b100 %
1'
b100 +
#569310000000
0!
0'
#569320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#569330000000
0!
0'
#569340000000
1!
0$
b110 %
1'
0*
b110 +
#569350000000
0!
0'
#569360000000
1!
b111 %
1'
b111 +
#569370000000
0!
0'
#569380000000
1!
b1000 %
1'
b1000 +
#569390000000
0!
0'
#569400000000
1!
b1001 %
1'
b1001 +
#569410000000
0!
0'
#569420000000
1!
b0 %
1'
b0 +
#569430000000
0!
0'
#569440000000
1!
1$
b1 %
1'
1*
b1 +
#569450000000
0!
0'
#569460000000
1!
b10 %
1'
b10 +
#569470000000
0!
0'
#569480000000
1!
b11 %
1'
b11 +
#569490000000
0!
0'
#569500000000
1!
b100 %
1'
b100 +
#569510000000
0!
0'
#569520000000
1!
b101 %
1'
b101 +
#569530000000
1"
1(
#569540000000
0!
0"
b100 &
0'
0(
b100 ,
#569550000000
1!
b110 %
1'
b110 +
#569560000000
0!
0'
#569570000000
1!
b111 %
1'
b111 +
#569580000000
0!
0'
#569590000000
1!
0$
b1000 %
1'
0*
b1000 +
#569600000000
0!
0'
#569610000000
1!
b1001 %
1'
b1001 +
#569620000000
0!
0'
#569630000000
1!
b0 %
1'
b0 +
#569640000000
0!
0'
#569650000000
1!
1$
b1 %
1'
1*
b1 +
#569660000000
0!
0'
#569670000000
1!
b10 %
1'
b10 +
#569680000000
0!
0'
#569690000000
1!
b11 %
1'
b11 +
#569700000000
0!
0'
#569710000000
1!
b100 %
1'
b100 +
#569720000000
0!
0'
#569730000000
1!
b101 %
1'
b101 +
#569740000000
0!
0'
#569750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#569760000000
0!
0'
#569770000000
1!
b111 %
1'
b111 +
#569780000000
0!
0'
#569790000000
1!
b1000 %
1'
b1000 +
#569800000000
0!
0'
#569810000000
1!
b1001 %
1'
b1001 +
#569820000000
0!
0'
#569830000000
1!
b0 %
1'
b0 +
#569840000000
0!
0'
#569850000000
1!
1$
b1 %
1'
1*
b1 +
#569860000000
0!
0'
#569870000000
1!
b10 %
1'
b10 +
#569880000000
0!
0'
#569890000000
1!
b11 %
1'
b11 +
#569900000000
0!
0'
#569910000000
1!
b100 %
1'
b100 +
#569920000000
0!
0'
#569930000000
1!
b101 %
1'
b101 +
#569940000000
0!
0'
#569950000000
1!
0$
b110 %
1'
0*
b110 +
#569960000000
1"
1(
#569970000000
0!
0"
b100 &
0'
0(
b100 ,
#569980000000
1!
1$
b111 %
1'
1*
b111 +
#569990000000
0!
0'
#570000000000
1!
0$
b1000 %
1'
0*
b1000 +
#570010000000
0!
0'
#570020000000
1!
b1001 %
1'
b1001 +
#570030000000
0!
0'
#570040000000
1!
b0 %
1'
b0 +
#570050000000
0!
0'
#570060000000
1!
1$
b1 %
1'
1*
b1 +
#570070000000
0!
0'
#570080000000
1!
b10 %
1'
b10 +
#570090000000
0!
0'
#570100000000
1!
b11 %
1'
b11 +
#570110000000
0!
0'
#570120000000
1!
b100 %
1'
b100 +
#570130000000
0!
0'
#570140000000
1!
b101 %
1'
b101 +
#570150000000
0!
0'
#570160000000
1!
b110 %
1'
b110 +
#570170000000
0!
0'
#570180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#570190000000
0!
0'
#570200000000
1!
b1000 %
1'
b1000 +
#570210000000
0!
0'
#570220000000
1!
b1001 %
1'
b1001 +
#570230000000
0!
0'
#570240000000
1!
b0 %
1'
b0 +
#570250000000
0!
0'
#570260000000
1!
1$
b1 %
1'
1*
b1 +
#570270000000
0!
0'
#570280000000
1!
b10 %
1'
b10 +
#570290000000
0!
0'
#570300000000
1!
b11 %
1'
b11 +
#570310000000
0!
0'
#570320000000
1!
b100 %
1'
b100 +
#570330000000
0!
0'
#570340000000
1!
b101 %
1'
b101 +
#570350000000
0!
0'
#570360000000
1!
0$
b110 %
1'
0*
b110 +
#570370000000
0!
0'
#570380000000
1!
b111 %
1'
b111 +
#570390000000
1"
1(
#570400000000
0!
0"
b100 &
0'
0(
b100 ,
#570410000000
1!
b1000 %
1'
b1000 +
#570420000000
0!
0'
#570430000000
1!
b1001 %
1'
b1001 +
#570440000000
0!
0'
#570450000000
1!
b0 %
1'
b0 +
#570460000000
0!
0'
#570470000000
1!
1$
b1 %
1'
1*
b1 +
#570480000000
0!
0'
#570490000000
1!
b10 %
1'
b10 +
#570500000000
0!
0'
#570510000000
1!
b11 %
1'
b11 +
#570520000000
0!
0'
#570530000000
1!
b100 %
1'
b100 +
#570540000000
0!
0'
#570550000000
1!
b101 %
1'
b101 +
#570560000000
0!
0'
#570570000000
1!
b110 %
1'
b110 +
#570580000000
0!
0'
#570590000000
1!
b111 %
1'
b111 +
#570600000000
0!
0'
#570610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#570620000000
0!
0'
#570630000000
1!
b1001 %
1'
b1001 +
#570640000000
0!
0'
#570650000000
1!
b0 %
1'
b0 +
#570660000000
0!
0'
#570670000000
1!
1$
b1 %
1'
1*
b1 +
#570680000000
0!
0'
#570690000000
1!
b10 %
1'
b10 +
#570700000000
0!
0'
#570710000000
1!
b11 %
1'
b11 +
#570720000000
0!
0'
#570730000000
1!
b100 %
1'
b100 +
#570740000000
0!
0'
#570750000000
1!
b101 %
1'
b101 +
#570760000000
0!
0'
#570770000000
1!
0$
b110 %
1'
0*
b110 +
#570780000000
0!
0'
#570790000000
1!
b111 %
1'
b111 +
#570800000000
0!
0'
#570810000000
1!
b1000 %
1'
b1000 +
#570820000000
1"
1(
#570830000000
0!
0"
b100 &
0'
0(
b100 ,
#570840000000
1!
b1001 %
1'
b1001 +
#570850000000
0!
0'
#570860000000
1!
b0 %
1'
b0 +
#570870000000
0!
0'
#570880000000
1!
1$
b1 %
1'
1*
b1 +
#570890000000
0!
0'
#570900000000
1!
b10 %
1'
b10 +
#570910000000
0!
0'
#570920000000
1!
b11 %
1'
b11 +
#570930000000
0!
0'
#570940000000
1!
b100 %
1'
b100 +
#570950000000
0!
0'
#570960000000
1!
b101 %
1'
b101 +
#570970000000
0!
0'
#570980000000
1!
b110 %
1'
b110 +
#570990000000
0!
0'
#571000000000
1!
b111 %
1'
b111 +
#571010000000
0!
0'
#571020000000
1!
0$
b1000 %
1'
0*
b1000 +
#571030000000
0!
0'
#571040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#571050000000
0!
0'
#571060000000
1!
b0 %
1'
b0 +
#571070000000
0!
0'
#571080000000
1!
1$
b1 %
1'
1*
b1 +
#571090000000
0!
0'
#571100000000
1!
b10 %
1'
b10 +
#571110000000
0!
0'
#571120000000
1!
b11 %
1'
b11 +
#571130000000
0!
0'
#571140000000
1!
b100 %
1'
b100 +
#571150000000
0!
0'
#571160000000
1!
b101 %
1'
b101 +
#571170000000
0!
0'
#571180000000
1!
0$
b110 %
1'
0*
b110 +
#571190000000
0!
0'
#571200000000
1!
b111 %
1'
b111 +
#571210000000
0!
0'
#571220000000
1!
b1000 %
1'
b1000 +
#571230000000
0!
0'
#571240000000
1!
b1001 %
1'
b1001 +
#571250000000
1"
1(
#571260000000
0!
0"
b100 &
0'
0(
b100 ,
#571270000000
1!
b0 %
1'
b0 +
#571280000000
0!
0'
#571290000000
1!
1$
b1 %
1'
1*
b1 +
#571300000000
0!
0'
#571310000000
1!
b10 %
1'
b10 +
#571320000000
0!
0'
#571330000000
1!
b11 %
1'
b11 +
#571340000000
0!
0'
#571350000000
1!
b100 %
1'
b100 +
#571360000000
0!
0'
#571370000000
1!
b101 %
1'
b101 +
#571380000000
0!
0'
#571390000000
1!
b110 %
1'
b110 +
#571400000000
0!
0'
#571410000000
1!
b111 %
1'
b111 +
#571420000000
0!
0'
#571430000000
1!
0$
b1000 %
1'
0*
b1000 +
#571440000000
0!
0'
#571450000000
1!
b1001 %
1'
b1001 +
#571460000000
0!
0'
#571470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#571480000000
0!
0'
#571490000000
1!
1$
b1 %
1'
1*
b1 +
#571500000000
0!
0'
#571510000000
1!
b10 %
1'
b10 +
#571520000000
0!
0'
#571530000000
1!
b11 %
1'
b11 +
#571540000000
0!
0'
#571550000000
1!
b100 %
1'
b100 +
#571560000000
0!
0'
#571570000000
1!
b101 %
1'
b101 +
#571580000000
0!
0'
#571590000000
1!
0$
b110 %
1'
0*
b110 +
#571600000000
0!
0'
#571610000000
1!
b111 %
1'
b111 +
#571620000000
0!
0'
#571630000000
1!
b1000 %
1'
b1000 +
#571640000000
0!
0'
#571650000000
1!
b1001 %
1'
b1001 +
#571660000000
0!
0'
#571670000000
1!
b0 %
1'
b0 +
#571680000000
1"
1(
#571690000000
0!
0"
b100 &
0'
0(
b100 ,
#571700000000
1!
1$
b1 %
1'
1*
b1 +
#571710000000
0!
0'
#571720000000
1!
b10 %
1'
b10 +
#571730000000
0!
0'
#571740000000
1!
b11 %
1'
b11 +
#571750000000
0!
0'
#571760000000
1!
b100 %
1'
b100 +
#571770000000
0!
0'
#571780000000
1!
b101 %
1'
b101 +
#571790000000
0!
0'
#571800000000
1!
b110 %
1'
b110 +
#571810000000
0!
0'
#571820000000
1!
b111 %
1'
b111 +
#571830000000
0!
0'
#571840000000
1!
0$
b1000 %
1'
0*
b1000 +
#571850000000
0!
0'
#571860000000
1!
b1001 %
1'
b1001 +
#571870000000
0!
0'
#571880000000
1!
b0 %
1'
b0 +
#571890000000
0!
0'
#571900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#571910000000
0!
0'
#571920000000
1!
b10 %
1'
b10 +
#571930000000
0!
0'
#571940000000
1!
b11 %
1'
b11 +
#571950000000
0!
0'
#571960000000
1!
b100 %
1'
b100 +
#571970000000
0!
0'
#571980000000
1!
b101 %
1'
b101 +
#571990000000
0!
0'
#572000000000
1!
0$
b110 %
1'
0*
b110 +
#572010000000
0!
0'
#572020000000
1!
b111 %
1'
b111 +
#572030000000
0!
0'
#572040000000
1!
b1000 %
1'
b1000 +
#572050000000
0!
0'
#572060000000
1!
b1001 %
1'
b1001 +
#572070000000
0!
0'
#572080000000
1!
b0 %
1'
b0 +
#572090000000
0!
0'
#572100000000
1!
1$
b1 %
1'
1*
b1 +
#572110000000
1"
1(
#572120000000
0!
0"
b100 &
0'
0(
b100 ,
#572130000000
1!
b10 %
1'
b10 +
#572140000000
0!
0'
#572150000000
1!
b11 %
1'
b11 +
#572160000000
0!
0'
#572170000000
1!
b100 %
1'
b100 +
#572180000000
0!
0'
#572190000000
1!
b101 %
1'
b101 +
#572200000000
0!
0'
#572210000000
1!
b110 %
1'
b110 +
#572220000000
0!
0'
#572230000000
1!
b111 %
1'
b111 +
#572240000000
0!
0'
#572250000000
1!
0$
b1000 %
1'
0*
b1000 +
#572260000000
0!
0'
#572270000000
1!
b1001 %
1'
b1001 +
#572280000000
0!
0'
#572290000000
1!
b0 %
1'
b0 +
#572300000000
0!
0'
#572310000000
1!
1$
b1 %
1'
1*
b1 +
#572320000000
0!
0'
#572330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#572340000000
0!
0'
#572350000000
1!
b11 %
1'
b11 +
#572360000000
0!
0'
#572370000000
1!
b100 %
1'
b100 +
#572380000000
0!
0'
#572390000000
1!
b101 %
1'
b101 +
#572400000000
0!
0'
#572410000000
1!
0$
b110 %
1'
0*
b110 +
#572420000000
0!
0'
#572430000000
1!
b111 %
1'
b111 +
#572440000000
0!
0'
#572450000000
1!
b1000 %
1'
b1000 +
#572460000000
0!
0'
#572470000000
1!
b1001 %
1'
b1001 +
#572480000000
0!
0'
#572490000000
1!
b0 %
1'
b0 +
#572500000000
0!
0'
#572510000000
1!
1$
b1 %
1'
1*
b1 +
#572520000000
0!
0'
#572530000000
1!
b10 %
1'
b10 +
#572540000000
1"
1(
#572550000000
0!
0"
b100 &
0'
0(
b100 ,
#572560000000
1!
b11 %
1'
b11 +
#572570000000
0!
0'
#572580000000
1!
b100 %
1'
b100 +
#572590000000
0!
0'
#572600000000
1!
b101 %
1'
b101 +
#572610000000
0!
0'
#572620000000
1!
b110 %
1'
b110 +
#572630000000
0!
0'
#572640000000
1!
b111 %
1'
b111 +
#572650000000
0!
0'
#572660000000
1!
0$
b1000 %
1'
0*
b1000 +
#572670000000
0!
0'
#572680000000
1!
b1001 %
1'
b1001 +
#572690000000
0!
0'
#572700000000
1!
b0 %
1'
b0 +
#572710000000
0!
0'
#572720000000
1!
1$
b1 %
1'
1*
b1 +
#572730000000
0!
0'
#572740000000
1!
b10 %
1'
b10 +
#572750000000
0!
0'
#572760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#572770000000
0!
0'
#572780000000
1!
b100 %
1'
b100 +
#572790000000
0!
0'
#572800000000
1!
b101 %
1'
b101 +
#572810000000
0!
0'
#572820000000
1!
0$
b110 %
1'
0*
b110 +
#572830000000
0!
0'
#572840000000
1!
b111 %
1'
b111 +
#572850000000
0!
0'
#572860000000
1!
b1000 %
1'
b1000 +
#572870000000
0!
0'
#572880000000
1!
b1001 %
1'
b1001 +
#572890000000
0!
0'
#572900000000
1!
b0 %
1'
b0 +
#572910000000
0!
0'
#572920000000
1!
1$
b1 %
1'
1*
b1 +
#572930000000
0!
0'
#572940000000
1!
b10 %
1'
b10 +
#572950000000
0!
0'
#572960000000
1!
b11 %
1'
b11 +
#572970000000
1"
1(
#572980000000
0!
0"
b100 &
0'
0(
b100 ,
#572990000000
1!
b100 %
1'
b100 +
#573000000000
0!
0'
#573010000000
1!
b101 %
1'
b101 +
#573020000000
0!
0'
#573030000000
1!
b110 %
1'
b110 +
#573040000000
0!
0'
#573050000000
1!
b111 %
1'
b111 +
#573060000000
0!
0'
#573070000000
1!
0$
b1000 %
1'
0*
b1000 +
#573080000000
0!
0'
#573090000000
1!
b1001 %
1'
b1001 +
#573100000000
0!
0'
#573110000000
1!
b0 %
1'
b0 +
#573120000000
0!
0'
#573130000000
1!
1$
b1 %
1'
1*
b1 +
#573140000000
0!
0'
#573150000000
1!
b10 %
1'
b10 +
#573160000000
0!
0'
#573170000000
1!
b11 %
1'
b11 +
#573180000000
0!
0'
#573190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#573200000000
0!
0'
#573210000000
1!
b101 %
1'
b101 +
#573220000000
0!
0'
#573230000000
1!
0$
b110 %
1'
0*
b110 +
#573240000000
0!
0'
#573250000000
1!
b111 %
1'
b111 +
#573260000000
0!
0'
#573270000000
1!
b1000 %
1'
b1000 +
#573280000000
0!
0'
#573290000000
1!
b1001 %
1'
b1001 +
#573300000000
0!
0'
#573310000000
1!
b0 %
1'
b0 +
#573320000000
0!
0'
#573330000000
1!
1$
b1 %
1'
1*
b1 +
#573340000000
0!
0'
#573350000000
1!
b10 %
1'
b10 +
#573360000000
0!
0'
#573370000000
1!
b11 %
1'
b11 +
#573380000000
0!
0'
#573390000000
1!
b100 %
1'
b100 +
#573400000000
1"
1(
#573410000000
0!
0"
b100 &
0'
0(
b100 ,
#573420000000
1!
b101 %
1'
b101 +
#573430000000
0!
0'
#573440000000
1!
b110 %
1'
b110 +
#573450000000
0!
0'
#573460000000
1!
b111 %
1'
b111 +
#573470000000
0!
0'
#573480000000
1!
0$
b1000 %
1'
0*
b1000 +
#573490000000
0!
0'
#573500000000
1!
b1001 %
1'
b1001 +
#573510000000
0!
0'
#573520000000
1!
b0 %
1'
b0 +
#573530000000
0!
0'
#573540000000
1!
1$
b1 %
1'
1*
b1 +
#573550000000
0!
0'
#573560000000
1!
b10 %
1'
b10 +
#573570000000
0!
0'
#573580000000
1!
b11 %
1'
b11 +
#573590000000
0!
0'
#573600000000
1!
b100 %
1'
b100 +
#573610000000
0!
0'
#573620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#573630000000
0!
0'
#573640000000
1!
0$
b110 %
1'
0*
b110 +
#573650000000
0!
0'
#573660000000
1!
b111 %
1'
b111 +
#573670000000
0!
0'
#573680000000
1!
b1000 %
1'
b1000 +
#573690000000
0!
0'
#573700000000
1!
b1001 %
1'
b1001 +
#573710000000
0!
0'
#573720000000
1!
b0 %
1'
b0 +
#573730000000
0!
0'
#573740000000
1!
1$
b1 %
1'
1*
b1 +
#573750000000
0!
0'
#573760000000
1!
b10 %
1'
b10 +
#573770000000
0!
0'
#573780000000
1!
b11 %
1'
b11 +
#573790000000
0!
0'
#573800000000
1!
b100 %
1'
b100 +
#573810000000
0!
0'
#573820000000
1!
b101 %
1'
b101 +
#573830000000
1"
1(
#573840000000
0!
0"
b100 &
0'
0(
b100 ,
#573850000000
1!
b110 %
1'
b110 +
#573860000000
0!
0'
#573870000000
1!
b111 %
1'
b111 +
#573880000000
0!
0'
#573890000000
1!
0$
b1000 %
1'
0*
b1000 +
#573900000000
0!
0'
#573910000000
1!
b1001 %
1'
b1001 +
#573920000000
0!
0'
#573930000000
1!
b0 %
1'
b0 +
#573940000000
0!
0'
#573950000000
1!
1$
b1 %
1'
1*
b1 +
#573960000000
0!
0'
#573970000000
1!
b10 %
1'
b10 +
#573980000000
0!
0'
#573990000000
1!
b11 %
1'
b11 +
#574000000000
0!
0'
#574010000000
1!
b100 %
1'
b100 +
#574020000000
0!
0'
#574030000000
1!
b101 %
1'
b101 +
#574040000000
0!
0'
#574050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#574060000000
0!
0'
#574070000000
1!
b111 %
1'
b111 +
#574080000000
0!
0'
#574090000000
1!
b1000 %
1'
b1000 +
#574100000000
0!
0'
#574110000000
1!
b1001 %
1'
b1001 +
#574120000000
0!
0'
#574130000000
1!
b0 %
1'
b0 +
#574140000000
0!
0'
#574150000000
1!
1$
b1 %
1'
1*
b1 +
#574160000000
0!
0'
#574170000000
1!
b10 %
1'
b10 +
#574180000000
0!
0'
#574190000000
1!
b11 %
1'
b11 +
#574200000000
0!
0'
#574210000000
1!
b100 %
1'
b100 +
#574220000000
0!
0'
#574230000000
1!
b101 %
1'
b101 +
#574240000000
0!
0'
#574250000000
1!
0$
b110 %
1'
0*
b110 +
#574260000000
1"
1(
#574270000000
0!
0"
b100 &
0'
0(
b100 ,
#574280000000
1!
1$
b111 %
1'
1*
b111 +
#574290000000
0!
0'
#574300000000
1!
0$
b1000 %
1'
0*
b1000 +
#574310000000
0!
0'
#574320000000
1!
b1001 %
1'
b1001 +
#574330000000
0!
0'
#574340000000
1!
b0 %
1'
b0 +
#574350000000
0!
0'
#574360000000
1!
1$
b1 %
1'
1*
b1 +
#574370000000
0!
0'
#574380000000
1!
b10 %
1'
b10 +
#574390000000
0!
0'
#574400000000
1!
b11 %
1'
b11 +
#574410000000
0!
0'
#574420000000
1!
b100 %
1'
b100 +
#574430000000
0!
0'
#574440000000
1!
b101 %
1'
b101 +
#574450000000
0!
0'
#574460000000
1!
b110 %
1'
b110 +
#574470000000
0!
0'
#574480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#574490000000
0!
0'
#574500000000
1!
b1000 %
1'
b1000 +
#574510000000
0!
0'
#574520000000
1!
b1001 %
1'
b1001 +
#574530000000
0!
0'
#574540000000
1!
b0 %
1'
b0 +
#574550000000
0!
0'
#574560000000
1!
1$
b1 %
1'
1*
b1 +
#574570000000
0!
0'
#574580000000
1!
b10 %
1'
b10 +
#574590000000
0!
0'
#574600000000
1!
b11 %
1'
b11 +
#574610000000
0!
0'
#574620000000
1!
b100 %
1'
b100 +
#574630000000
0!
0'
#574640000000
1!
b101 %
1'
b101 +
#574650000000
0!
0'
#574660000000
1!
0$
b110 %
1'
0*
b110 +
#574670000000
0!
0'
#574680000000
1!
b111 %
1'
b111 +
#574690000000
1"
1(
#574700000000
0!
0"
b100 &
0'
0(
b100 ,
#574710000000
1!
b1000 %
1'
b1000 +
#574720000000
0!
0'
#574730000000
1!
b1001 %
1'
b1001 +
#574740000000
0!
0'
#574750000000
1!
b0 %
1'
b0 +
#574760000000
0!
0'
#574770000000
1!
1$
b1 %
1'
1*
b1 +
#574780000000
0!
0'
#574790000000
1!
b10 %
1'
b10 +
#574800000000
0!
0'
#574810000000
1!
b11 %
1'
b11 +
#574820000000
0!
0'
#574830000000
1!
b100 %
1'
b100 +
#574840000000
0!
0'
#574850000000
1!
b101 %
1'
b101 +
#574860000000
0!
0'
#574870000000
1!
b110 %
1'
b110 +
#574880000000
0!
0'
#574890000000
1!
b111 %
1'
b111 +
#574900000000
0!
0'
#574910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#574920000000
0!
0'
#574930000000
1!
b1001 %
1'
b1001 +
#574940000000
0!
0'
#574950000000
1!
b0 %
1'
b0 +
#574960000000
0!
0'
#574970000000
1!
1$
b1 %
1'
1*
b1 +
#574980000000
0!
0'
#574990000000
1!
b10 %
1'
b10 +
#575000000000
0!
0'
#575010000000
1!
b11 %
1'
b11 +
#575020000000
0!
0'
#575030000000
1!
b100 %
1'
b100 +
#575040000000
0!
0'
#575050000000
1!
b101 %
1'
b101 +
#575060000000
0!
0'
#575070000000
1!
0$
b110 %
1'
0*
b110 +
#575080000000
0!
0'
#575090000000
1!
b111 %
1'
b111 +
#575100000000
0!
0'
#575110000000
1!
b1000 %
1'
b1000 +
#575120000000
1"
1(
#575130000000
0!
0"
b100 &
0'
0(
b100 ,
#575140000000
1!
b1001 %
1'
b1001 +
#575150000000
0!
0'
#575160000000
1!
b0 %
1'
b0 +
#575170000000
0!
0'
#575180000000
1!
1$
b1 %
1'
1*
b1 +
#575190000000
0!
0'
#575200000000
1!
b10 %
1'
b10 +
#575210000000
0!
0'
#575220000000
1!
b11 %
1'
b11 +
#575230000000
0!
0'
#575240000000
1!
b100 %
1'
b100 +
#575250000000
0!
0'
#575260000000
1!
b101 %
1'
b101 +
#575270000000
0!
0'
#575280000000
1!
b110 %
1'
b110 +
#575290000000
0!
0'
#575300000000
1!
b111 %
1'
b111 +
#575310000000
0!
0'
#575320000000
1!
0$
b1000 %
1'
0*
b1000 +
#575330000000
0!
0'
#575340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#575350000000
0!
0'
#575360000000
1!
b0 %
1'
b0 +
#575370000000
0!
0'
#575380000000
1!
1$
b1 %
1'
1*
b1 +
#575390000000
0!
0'
#575400000000
1!
b10 %
1'
b10 +
#575410000000
0!
0'
#575420000000
1!
b11 %
1'
b11 +
#575430000000
0!
0'
#575440000000
1!
b100 %
1'
b100 +
#575450000000
0!
0'
#575460000000
1!
b101 %
1'
b101 +
#575470000000
0!
0'
#575480000000
1!
0$
b110 %
1'
0*
b110 +
#575490000000
0!
0'
#575500000000
1!
b111 %
1'
b111 +
#575510000000
0!
0'
#575520000000
1!
b1000 %
1'
b1000 +
#575530000000
0!
0'
#575540000000
1!
b1001 %
1'
b1001 +
#575550000000
1"
1(
#575560000000
0!
0"
b100 &
0'
0(
b100 ,
#575570000000
1!
b0 %
1'
b0 +
#575580000000
0!
0'
#575590000000
1!
1$
b1 %
1'
1*
b1 +
#575600000000
0!
0'
#575610000000
1!
b10 %
1'
b10 +
#575620000000
0!
0'
#575630000000
1!
b11 %
1'
b11 +
#575640000000
0!
0'
#575650000000
1!
b100 %
1'
b100 +
#575660000000
0!
0'
#575670000000
1!
b101 %
1'
b101 +
#575680000000
0!
0'
#575690000000
1!
b110 %
1'
b110 +
#575700000000
0!
0'
#575710000000
1!
b111 %
1'
b111 +
#575720000000
0!
0'
#575730000000
1!
0$
b1000 %
1'
0*
b1000 +
#575740000000
0!
0'
#575750000000
1!
b1001 %
1'
b1001 +
#575760000000
0!
0'
#575770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#575780000000
0!
0'
#575790000000
1!
1$
b1 %
1'
1*
b1 +
#575800000000
0!
0'
#575810000000
1!
b10 %
1'
b10 +
#575820000000
0!
0'
#575830000000
1!
b11 %
1'
b11 +
#575840000000
0!
0'
#575850000000
1!
b100 %
1'
b100 +
#575860000000
0!
0'
#575870000000
1!
b101 %
1'
b101 +
#575880000000
0!
0'
#575890000000
1!
0$
b110 %
1'
0*
b110 +
#575900000000
0!
0'
#575910000000
1!
b111 %
1'
b111 +
#575920000000
0!
0'
#575930000000
1!
b1000 %
1'
b1000 +
#575940000000
0!
0'
#575950000000
1!
b1001 %
1'
b1001 +
#575960000000
0!
0'
#575970000000
1!
b0 %
1'
b0 +
#575980000000
1"
1(
#575990000000
0!
0"
b100 &
0'
0(
b100 ,
#576000000000
1!
1$
b1 %
1'
1*
b1 +
#576010000000
0!
0'
#576020000000
1!
b10 %
1'
b10 +
#576030000000
0!
0'
#576040000000
1!
b11 %
1'
b11 +
#576050000000
0!
0'
#576060000000
1!
b100 %
1'
b100 +
#576070000000
0!
0'
#576080000000
1!
b101 %
1'
b101 +
#576090000000
0!
0'
#576100000000
1!
b110 %
1'
b110 +
#576110000000
0!
0'
#576120000000
1!
b111 %
1'
b111 +
#576130000000
0!
0'
#576140000000
1!
0$
b1000 %
1'
0*
b1000 +
#576150000000
0!
0'
#576160000000
1!
b1001 %
1'
b1001 +
#576170000000
0!
0'
#576180000000
1!
b0 %
1'
b0 +
#576190000000
0!
0'
#576200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#576210000000
0!
0'
#576220000000
1!
b10 %
1'
b10 +
#576230000000
0!
0'
#576240000000
1!
b11 %
1'
b11 +
#576250000000
0!
0'
#576260000000
1!
b100 %
1'
b100 +
#576270000000
0!
0'
#576280000000
1!
b101 %
1'
b101 +
#576290000000
0!
0'
#576300000000
1!
0$
b110 %
1'
0*
b110 +
#576310000000
0!
0'
#576320000000
1!
b111 %
1'
b111 +
#576330000000
0!
0'
#576340000000
1!
b1000 %
1'
b1000 +
#576350000000
0!
0'
#576360000000
1!
b1001 %
1'
b1001 +
#576370000000
0!
0'
#576380000000
1!
b0 %
1'
b0 +
#576390000000
0!
0'
#576400000000
1!
1$
b1 %
1'
1*
b1 +
#576410000000
1"
1(
#576420000000
0!
0"
b100 &
0'
0(
b100 ,
#576430000000
1!
b10 %
1'
b10 +
#576440000000
0!
0'
#576450000000
1!
b11 %
1'
b11 +
#576460000000
0!
0'
#576470000000
1!
b100 %
1'
b100 +
#576480000000
0!
0'
#576490000000
1!
b101 %
1'
b101 +
#576500000000
0!
0'
#576510000000
1!
b110 %
1'
b110 +
#576520000000
0!
0'
#576530000000
1!
b111 %
1'
b111 +
#576540000000
0!
0'
#576550000000
1!
0$
b1000 %
1'
0*
b1000 +
#576560000000
0!
0'
#576570000000
1!
b1001 %
1'
b1001 +
#576580000000
0!
0'
#576590000000
1!
b0 %
1'
b0 +
#576600000000
0!
0'
#576610000000
1!
1$
b1 %
1'
1*
b1 +
#576620000000
0!
0'
#576630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#576640000000
0!
0'
#576650000000
1!
b11 %
1'
b11 +
#576660000000
0!
0'
#576670000000
1!
b100 %
1'
b100 +
#576680000000
0!
0'
#576690000000
1!
b101 %
1'
b101 +
#576700000000
0!
0'
#576710000000
1!
0$
b110 %
1'
0*
b110 +
#576720000000
0!
0'
#576730000000
1!
b111 %
1'
b111 +
#576740000000
0!
0'
#576750000000
1!
b1000 %
1'
b1000 +
#576760000000
0!
0'
#576770000000
1!
b1001 %
1'
b1001 +
#576780000000
0!
0'
#576790000000
1!
b0 %
1'
b0 +
#576800000000
0!
0'
#576810000000
1!
1$
b1 %
1'
1*
b1 +
#576820000000
0!
0'
#576830000000
1!
b10 %
1'
b10 +
#576840000000
1"
1(
#576850000000
0!
0"
b100 &
0'
0(
b100 ,
#576860000000
1!
b11 %
1'
b11 +
#576870000000
0!
0'
#576880000000
1!
b100 %
1'
b100 +
#576890000000
0!
0'
#576900000000
1!
b101 %
1'
b101 +
#576910000000
0!
0'
#576920000000
1!
b110 %
1'
b110 +
#576930000000
0!
0'
#576940000000
1!
b111 %
1'
b111 +
#576950000000
0!
0'
#576960000000
1!
0$
b1000 %
1'
0*
b1000 +
#576970000000
0!
0'
#576980000000
1!
b1001 %
1'
b1001 +
#576990000000
0!
0'
#577000000000
1!
b0 %
1'
b0 +
#577010000000
0!
0'
#577020000000
1!
1$
b1 %
1'
1*
b1 +
#577030000000
0!
0'
#577040000000
1!
b10 %
1'
b10 +
#577050000000
0!
0'
#577060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#577070000000
0!
0'
#577080000000
1!
b100 %
1'
b100 +
#577090000000
0!
0'
#577100000000
1!
b101 %
1'
b101 +
#577110000000
0!
0'
#577120000000
1!
0$
b110 %
1'
0*
b110 +
#577130000000
0!
0'
#577140000000
1!
b111 %
1'
b111 +
#577150000000
0!
0'
#577160000000
1!
b1000 %
1'
b1000 +
#577170000000
0!
0'
#577180000000
1!
b1001 %
1'
b1001 +
#577190000000
0!
0'
#577200000000
1!
b0 %
1'
b0 +
#577210000000
0!
0'
#577220000000
1!
1$
b1 %
1'
1*
b1 +
#577230000000
0!
0'
#577240000000
1!
b10 %
1'
b10 +
#577250000000
0!
0'
#577260000000
1!
b11 %
1'
b11 +
#577270000000
1"
1(
#577280000000
0!
0"
b100 &
0'
0(
b100 ,
#577290000000
1!
b100 %
1'
b100 +
#577300000000
0!
0'
#577310000000
1!
b101 %
1'
b101 +
#577320000000
0!
0'
#577330000000
1!
b110 %
1'
b110 +
#577340000000
0!
0'
#577350000000
1!
b111 %
1'
b111 +
#577360000000
0!
0'
#577370000000
1!
0$
b1000 %
1'
0*
b1000 +
#577380000000
0!
0'
#577390000000
1!
b1001 %
1'
b1001 +
#577400000000
0!
0'
#577410000000
1!
b0 %
1'
b0 +
#577420000000
0!
0'
#577430000000
1!
1$
b1 %
1'
1*
b1 +
#577440000000
0!
0'
#577450000000
1!
b10 %
1'
b10 +
#577460000000
0!
0'
#577470000000
1!
b11 %
1'
b11 +
#577480000000
0!
0'
#577490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#577500000000
0!
0'
#577510000000
1!
b101 %
1'
b101 +
#577520000000
0!
0'
#577530000000
1!
0$
b110 %
1'
0*
b110 +
#577540000000
0!
0'
#577550000000
1!
b111 %
1'
b111 +
#577560000000
0!
0'
#577570000000
1!
b1000 %
1'
b1000 +
#577580000000
0!
0'
#577590000000
1!
b1001 %
1'
b1001 +
#577600000000
0!
0'
#577610000000
1!
b0 %
1'
b0 +
#577620000000
0!
0'
#577630000000
1!
1$
b1 %
1'
1*
b1 +
#577640000000
0!
0'
#577650000000
1!
b10 %
1'
b10 +
#577660000000
0!
0'
#577670000000
1!
b11 %
1'
b11 +
#577680000000
0!
0'
#577690000000
1!
b100 %
1'
b100 +
#577700000000
1"
1(
#577710000000
0!
0"
b100 &
0'
0(
b100 ,
#577720000000
1!
b101 %
1'
b101 +
#577730000000
0!
0'
#577740000000
1!
b110 %
1'
b110 +
#577750000000
0!
0'
#577760000000
1!
b111 %
1'
b111 +
#577770000000
0!
0'
#577780000000
1!
0$
b1000 %
1'
0*
b1000 +
#577790000000
0!
0'
#577800000000
1!
b1001 %
1'
b1001 +
#577810000000
0!
0'
#577820000000
1!
b0 %
1'
b0 +
#577830000000
0!
0'
#577840000000
1!
1$
b1 %
1'
1*
b1 +
#577850000000
0!
0'
#577860000000
1!
b10 %
1'
b10 +
#577870000000
0!
0'
#577880000000
1!
b11 %
1'
b11 +
#577890000000
0!
0'
#577900000000
1!
b100 %
1'
b100 +
#577910000000
0!
0'
#577920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#577930000000
0!
0'
#577940000000
1!
0$
b110 %
1'
0*
b110 +
#577950000000
0!
0'
#577960000000
1!
b111 %
1'
b111 +
#577970000000
0!
0'
#577980000000
1!
b1000 %
1'
b1000 +
#577990000000
0!
0'
#578000000000
1!
b1001 %
1'
b1001 +
#578010000000
0!
0'
#578020000000
1!
b0 %
1'
b0 +
#578030000000
0!
0'
#578040000000
1!
1$
b1 %
1'
1*
b1 +
#578050000000
0!
0'
#578060000000
1!
b10 %
1'
b10 +
#578070000000
0!
0'
#578080000000
1!
b11 %
1'
b11 +
#578090000000
0!
0'
#578100000000
1!
b100 %
1'
b100 +
#578110000000
0!
0'
#578120000000
1!
b101 %
1'
b101 +
#578130000000
1"
1(
#578140000000
0!
0"
b100 &
0'
0(
b100 ,
#578150000000
1!
b110 %
1'
b110 +
#578160000000
0!
0'
#578170000000
1!
b111 %
1'
b111 +
#578180000000
0!
0'
#578190000000
1!
0$
b1000 %
1'
0*
b1000 +
#578200000000
0!
0'
#578210000000
1!
b1001 %
1'
b1001 +
#578220000000
0!
0'
#578230000000
1!
b0 %
1'
b0 +
#578240000000
0!
0'
#578250000000
1!
1$
b1 %
1'
1*
b1 +
#578260000000
0!
0'
#578270000000
1!
b10 %
1'
b10 +
#578280000000
0!
0'
#578290000000
1!
b11 %
1'
b11 +
#578300000000
0!
0'
#578310000000
1!
b100 %
1'
b100 +
#578320000000
0!
0'
#578330000000
1!
b101 %
1'
b101 +
#578340000000
0!
0'
#578350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#578360000000
0!
0'
#578370000000
1!
b111 %
1'
b111 +
#578380000000
0!
0'
#578390000000
1!
b1000 %
1'
b1000 +
#578400000000
0!
0'
#578410000000
1!
b1001 %
1'
b1001 +
#578420000000
0!
0'
#578430000000
1!
b0 %
1'
b0 +
#578440000000
0!
0'
#578450000000
1!
1$
b1 %
1'
1*
b1 +
#578460000000
0!
0'
#578470000000
1!
b10 %
1'
b10 +
#578480000000
0!
0'
#578490000000
1!
b11 %
1'
b11 +
#578500000000
0!
0'
#578510000000
1!
b100 %
1'
b100 +
#578520000000
0!
0'
#578530000000
1!
b101 %
1'
b101 +
#578540000000
0!
0'
#578550000000
1!
0$
b110 %
1'
0*
b110 +
#578560000000
1"
1(
#578570000000
0!
0"
b100 &
0'
0(
b100 ,
#578580000000
1!
1$
b111 %
1'
1*
b111 +
#578590000000
0!
0'
#578600000000
1!
0$
b1000 %
1'
0*
b1000 +
#578610000000
0!
0'
#578620000000
1!
b1001 %
1'
b1001 +
#578630000000
0!
0'
#578640000000
1!
b0 %
1'
b0 +
#578650000000
0!
0'
#578660000000
1!
1$
b1 %
1'
1*
b1 +
#578670000000
0!
0'
#578680000000
1!
b10 %
1'
b10 +
#578690000000
0!
0'
#578700000000
1!
b11 %
1'
b11 +
#578710000000
0!
0'
#578720000000
1!
b100 %
1'
b100 +
#578730000000
0!
0'
#578740000000
1!
b101 %
1'
b101 +
#578750000000
0!
0'
#578760000000
1!
b110 %
1'
b110 +
#578770000000
0!
0'
#578780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#578790000000
0!
0'
#578800000000
1!
b1000 %
1'
b1000 +
#578810000000
0!
0'
#578820000000
1!
b1001 %
1'
b1001 +
#578830000000
0!
0'
#578840000000
1!
b0 %
1'
b0 +
#578850000000
0!
0'
#578860000000
1!
1$
b1 %
1'
1*
b1 +
#578870000000
0!
0'
#578880000000
1!
b10 %
1'
b10 +
#578890000000
0!
0'
#578900000000
1!
b11 %
1'
b11 +
#578910000000
0!
0'
#578920000000
1!
b100 %
1'
b100 +
#578930000000
0!
0'
#578940000000
1!
b101 %
1'
b101 +
#578950000000
0!
0'
#578960000000
1!
0$
b110 %
1'
0*
b110 +
#578970000000
0!
0'
#578980000000
1!
b111 %
1'
b111 +
#578990000000
1"
1(
#579000000000
0!
0"
b100 &
0'
0(
b100 ,
#579010000000
1!
b1000 %
1'
b1000 +
#579020000000
0!
0'
#579030000000
1!
b1001 %
1'
b1001 +
#579040000000
0!
0'
#579050000000
1!
b0 %
1'
b0 +
#579060000000
0!
0'
#579070000000
1!
1$
b1 %
1'
1*
b1 +
#579080000000
0!
0'
#579090000000
1!
b10 %
1'
b10 +
#579100000000
0!
0'
#579110000000
1!
b11 %
1'
b11 +
#579120000000
0!
0'
#579130000000
1!
b100 %
1'
b100 +
#579140000000
0!
0'
#579150000000
1!
b101 %
1'
b101 +
#579160000000
0!
0'
#579170000000
1!
b110 %
1'
b110 +
#579180000000
0!
0'
#579190000000
1!
b111 %
1'
b111 +
#579200000000
0!
0'
#579210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#579220000000
0!
0'
#579230000000
1!
b1001 %
1'
b1001 +
#579240000000
0!
0'
#579250000000
1!
b0 %
1'
b0 +
#579260000000
0!
0'
#579270000000
1!
1$
b1 %
1'
1*
b1 +
#579280000000
0!
0'
#579290000000
1!
b10 %
1'
b10 +
#579300000000
0!
0'
#579310000000
1!
b11 %
1'
b11 +
#579320000000
0!
0'
#579330000000
1!
b100 %
1'
b100 +
#579340000000
0!
0'
#579350000000
1!
b101 %
1'
b101 +
#579360000000
0!
0'
#579370000000
1!
0$
b110 %
1'
0*
b110 +
#579380000000
0!
0'
#579390000000
1!
b111 %
1'
b111 +
#579400000000
0!
0'
#579410000000
1!
b1000 %
1'
b1000 +
#579420000000
1"
1(
#579430000000
0!
0"
b100 &
0'
0(
b100 ,
#579440000000
1!
b1001 %
1'
b1001 +
#579450000000
0!
0'
#579460000000
1!
b0 %
1'
b0 +
#579470000000
0!
0'
#579480000000
1!
1$
b1 %
1'
1*
b1 +
#579490000000
0!
0'
#579500000000
1!
b10 %
1'
b10 +
#579510000000
0!
0'
#579520000000
1!
b11 %
1'
b11 +
#579530000000
0!
0'
#579540000000
1!
b100 %
1'
b100 +
#579550000000
0!
0'
#579560000000
1!
b101 %
1'
b101 +
#579570000000
0!
0'
#579580000000
1!
b110 %
1'
b110 +
#579590000000
0!
0'
#579600000000
1!
b111 %
1'
b111 +
#579610000000
0!
0'
#579620000000
1!
0$
b1000 %
1'
0*
b1000 +
#579630000000
0!
0'
#579640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#579650000000
0!
0'
#579660000000
1!
b0 %
1'
b0 +
#579670000000
0!
0'
#579680000000
1!
1$
b1 %
1'
1*
b1 +
#579690000000
0!
0'
#579700000000
1!
b10 %
1'
b10 +
#579710000000
0!
0'
#579720000000
1!
b11 %
1'
b11 +
#579730000000
0!
0'
#579740000000
1!
b100 %
1'
b100 +
#579750000000
0!
0'
#579760000000
1!
b101 %
1'
b101 +
#579770000000
0!
0'
#579780000000
1!
0$
b110 %
1'
0*
b110 +
#579790000000
0!
0'
#579800000000
1!
b111 %
1'
b111 +
#579810000000
0!
0'
#579820000000
1!
b1000 %
1'
b1000 +
#579830000000
0!
0'
#579840000000
1!
b1001 %
1'
b1001 +
#579850000000
1"
1(
#579860000000
0!
0"
b100 &
0'
0(
b100 ,
#579870000000
1!
b0 %
1'
b0 +
#579880000000
0!
0'
#579890000000
1!
1$
b1 %
1'
1*
b1 +
#579900000000
0!
0'
#579910000000
1!
b10 %
1'
b10 +
#579920000000
0!
0'
#579930000000
1!
b11 %
1'
b11 +
#579940000000
0!
0'
#579950000000
1!
b100 %
1'
b100 +
#579960000000
0!
0'
#579970000000
1!
b101 %
1'
b101 +
#579980000000
0!
0'
#579990000000
1!
b110 %
1'
b110 +
#580000000000
0!
0'
#580010000000
1!
b111 %
1'
b111 +
#580020000000
0!
0'
#580030000000
1!
0$
b1000 %
1'
0*
b1000 +
#580040000000
0!
0'
#580050000000
1!
b1001 %
1'
b1001 +
#580060000000
0!
0'
#580070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#580080000000
0!
0'
#580090000000
1!
1$
b1 %
1'
1*
b1 +
#580100000000
0!
0'
#580110000000
1!
b10 %
1'
b10 +
#580120000000
0!
0'
#580130000000
1!
b11 %
1'
b11 +
#580140000000
0!
0'
#580150000000
1!
b100 %
1'
b100 +
#580160000000
0!
0'
#580170000000
1!
b101 %
1'
b101 +
#580180000000
0!
0'
#580190000000
1!
0$
b110 %
1'
0*
b110 +
#580200000000
0!
0'
#580210000000
1!
b111 %
1'
b111 +
#580220000000
0!
0'
#580230000000
1!
b1000 %
1'
b1000 +
#580240000000
0!
0'
#580250000000
1!
b1001 %
1'
b1001 +
#580260000000
0!
0'
#580270000000
1!
b0 %
1'
b0 +
#580280000000
1"
1(
#580290000000
0!
0"
b100 &
0'
0(
b100 ,
#580300000000
1!
1$
b1 %
1'
1*
b1 +
#580310000000
0!
0'
#580320000000
1!
b10 %
1'
b10 +
#580330000000
0!
0'
#580340000000
1!
b11 %
1'
b11 +
#580350000000
0!
0'
#580360000000
1!
b100 %
1'
b100 +
#580370000000
0!
0'
#580380000000
1!
b101 %
1'
b101 +
#580390000000
0!
0'
#580400000000
1!
b110 %
1'
b110 +
#580410000000
0!
0'
#580420000000
1!
b111 %
1'
b111 +
#580430000000
0!
0'
#580440000000
1!
0$
b1000 %
1'
0*
b1000 +
#580450000000
0!
0'
#580460000000
1!
b1001 %
1'
b1001 +
#580470000000
0!
0'
#580480000000
1!
b0 %
1'
b0 +
#580490000000
0!
0'
#580500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#580510000000
0!
0'
#580520000000
1!
b10 %
1'
b10 +
#580530000000
0!
0'
#580540000000
1!
b11 %
1'
b11 +
#580550000000
0!
0'
#580560000000
1!
b100 %
1'
b100 +
#580570000000
0!
0'
#580580000000
1!
b101 %
1'
b101 +
#580590000000
0!
0'
#580600000000
1!
0$
b110 %
1'
0*
b110 +
#580610000000
0!
0'
#580620000000
1!
b111 %
1'
b111 +
#580630000000
0!
0'
#580640000000
1!
b1000 %
1'
b1000 +
#580650000000
0!
0'
#580660000000
1!
b1001 %
1'
b1001 +
#580670000000
0!
0'
#580680000000
1!
b0 %
1'
b0 +
#580690000000
0!
0'
#580700000000
1!
1$
b1 %
1'
1*
b1 +
#580710000000
1"
1(
#580720000000
0!
0"
b100 &
0'
0(
b100 ,
#580730000000
1!
b10 %
1'
b10 +
#580740000000
0!
0'
#580750000000
1!
b11 %
1'
b11 +
#580760000000
0!
0'
#580770000000
1!
b100 %
1'
b100 +
#580780000000
0!
0'
#580790000000
1!
b101 %
1'
b101 +
#580800000000
0!
0'
#580810000000
1!
b110 %
1'
b110 +
#580820000000
0!
0'
#580830000000
1!
b111 %
1'
b111 +
#580840000000
0!
0'
#580850000000
1!
0$
b1000 %
1'
0*
b1000 +
#580860000000
0!
0'
#580870000000
1!
b1001 %
1'
b1001 +
#580880000000
0!
0'
#580890000000
1!
b0 %
1'
b0 +
#580900000000
0!
0'
#580910000000
1!
1$
b1 %
1'
1*
b1 +
#580920000000
0!
0'
#580930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#580940000000
0!
0'
#580950000000
1!
b11 %
1'
b11 +
#580960000000
0!
0'
#580970000000
1!
b100 %
1'
b100 +
#580980000000
0!
0'
#580990000000
1!
b101 %
1'
b101 +
#581000000000
0!
0'
#581010000000
1!
0$
b110 %
1'
0*
b110 +
#581020000000
0!
0'
#581030000000
1!
b111 %
1'
b111 +
#581040000000
0!
0'
#581050000000
1!
b1000 %
1'
b1000 +
#581060000000
0!
0'
#581070000000
1!
b1001 %
1'
b1001 +
#581080000000
0!
0'
#581090000000
1!
b0 %
1'
b0 +
#581100000000
0!
0'
#581110000000
1!
1$
b1 %
1'
1*
b1 +
#581120000000
0!
0'
#581130000000
1!
b10 %
1'
b10 +
#581140000000
1"
1(
#581150000000
0!
0"
b100 &
0'
0(
b100 ,
#581160000000
1!
b11 %
1'
b11 +
#581170000000
0!
0'
#581180000000
1!
b100 %
1'
b100 +
#581190000000
0!
0'
#581200000000
1!
b101 %
1'
b101 +
#581210000000
0!
0'
#581220000000
1!
b110 %
1'
b110 +
#581230000000
0!
0'
#581240000000
1!
b111 %
1'
b111 +
#581250000000
0!
0'
#581260000000
1!
0$
b1000 %
1'
0*
b1000 +
#581270000000
0!
0'
#581280000000
1!
b1001 %
1'
b1001 +
#581290000000
0!
0'
#581300000000
1!
b0 %
1'
b0 +
#581310000000
0!
0'
#581320000000
1!
1$
b1 %
1'
1*
b1 +
#581330000000
0!
0'
#581340000000
1!
b10 %
1'
b10 +
#581350000000
0!
0'
#581360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#581370000000
0!
0'
#581380000000
1!
b100 %
1'
b100 +
#581390000000
0!
0'
#581400000000
1!
b101 %
1'
b101 +
#581410000000
0!
0'
#581420000000
1!
0$
b110 %
1'
0*
b110 +
#581430000000
0!
0'
#581440000000
1!
b111 %
1'
b111 +
#581450000000
0!
0'
#581460000000
1!
b1000 %
1'
b1000 +
#581470000000
0!
0'
#581480000000
1!
b1001 %
1'
b1001 +
#581490000000
0!
0'
#581500000000
1!
b0 %
1'
b0 +
#581510000000
0!
0'
#581520000000
1!
1$
b1 %
1'
1*
b1 +
#581530000000
0!
0'
#581540000000
1!
b10 %
1'
b10 +
#581550000000
0!
0'
#581560000000
1!
b11 %
1'
b11 +
#581570000000
1"
1(
#581580000000
0!
0"
b100 &
0'
0(
b100 ,
#581590000000
1!
b100 %
1'
b100 +
#581600000000
0!
0'
#581610000000
1!
b101 %
1'
b101 +
#581620000000
0!
0'
#581630000000
1!
b110 %
1'
b110 +
#581640000000
0!
0'
#581650000000
1!
b111 %
1'
b111 +
#581660000000
0!
0'
#581670000000
1!
0$
b1000 %
1'
0*
b1000 +
#581680000000
0!
0'
#581690000000
1!
b1001 %
1'
b1001 +
#581700000000
0!
0'
#581710000000
1!
b0 %
1'
b0 +
#581720000000
0!
0'
#581730000000
1!
1$
b1 %
1'
1*
b1 +
#581740000000
0!
0'
#581750000000
1!
b10 %
1'
b10 +
#581760000000
0!
0'
#581770000000
1!
b11 %
1'
b11 +
#581780000000
0!
0'
#581790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#581800000000
0!
0'
#581810000000
1!
b101 %
1'
b101 +
#581820000000
0!
0'
#581830000000
1!
0$
b110 %
1'
0*
b110 +
#581840000000
0!
0'
#581850000000
1!
b111 %
1'
b111 +
#581860000000
0!
0'
#581870000000
1!
b1000 %
1'
b1000 +
#581880000000
0!
0'
#581890000000
1!
b1001 %
1'
b1001 +
#581900000000
0!
0'
#581910000000
1!
b0 %
1'
b0 +
#581920000000
0!
0'
#581930000000
1!
1$
b1 %
1'
1*
b1 +
#581940000000
0!
0'
#581950000000
1!
b10 %
1'
b10 +
#581960000000
0!
0'
#581970000000
1!
b11 %
1'
b11 +
#581980000000
0!
0'
#581990000000
1!
b100 %
1'
b100 +
#582000000000
1"
1(
#582010000000
0!
0"
b100 &
0'
0(
b100 ,
#582020000000
1!
b101 %
1'
b101 +
#582030000000
0!
0'
#582040000000
1!
b110 %
1'
b110 +
#582050000000
0!
0'
#582060000000
1!
b111 %
1'
b111 +
#582070000000
0!
0'
#582080000000
1!
0$
b1000 %
1'
0*
b1000 +
#582090000000
0!
0'
#582100000000
1!
b1001 %
1'
b1001 +
#582110000000
0!
0'
#582120000000
1!
b0 %
1'
b0 +
#582130000000
0!
0'
#582140000000
1!
1$
b1 %
1'
1*
b1 +
#582150000000
0!
0'
#582160000000
1!
b10 %
1'
b10 +
#582170000000
0!
0'
#582180000000
1!
b11 %
1'
b11 +
#582190000000
0!
0'
#582200000000
1!
b100 %
1'
b100 +
#582210000000
0!
0'
#582220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#582230000000
0!
0'
#582240000000
1!
0$
b110 %
1'
0*
b110 +
#582250000000
0!
0'
#582260000000
1!
b111 %
1'
b111 +
#582270000000
0!
0'
#582280000000
1!
b1000 %
1'
b1000 +
#582290000000
0!
0'
#582300000000
1!
b1001 %
1'
b1001 +
#582310000000
0!
0'
#582320000000
1!
b0 %
1'
b0 +
#582330000000
0!
0'
#582340000000
1!
1$
b1 %
1'
1*
b1 +
#582350000000
0!
0'
#582360000000
1!
b10 %
1'
b10 +
#582370000000
0!
0'
#582380000000
1!
b11 %
1'
b11 +
#582390000000
0!
0'
#582400000000
1!
b100 %
1'
b100 +
#582410000000
0!
0'
#582420000000
1!
b101 %
1'
b101 +
#582430000000
1"
1(
#582440000000
0!
0"
b100 &
0'
0(
b100 ,
#582450000000
1!
b110 %
1'
b110 +
#582460000000
0!
0'
#582470000000
1!
b111 %
1'
b111 +
#582480000000
0!
0'
#582490000000
1!
0$
b1000 %
1'
0*
b1000 +
#582500000000
0!
0'
#582510000000
1!
b1001 %
1'
b1001 +
#582520000000
0!
0'
#582530000000
1!
b0 %
1'
b0 +
#582540000000
0!
0'
#582550000000
1!
1$
b1 %
1'
1*
b1 +
#582560000000
0!
0'
#582570000000
1!
b10 %
1'
b10 +
#582580000000
0!
0'
#582590000000
1!
b11 %
1'
b11 +
#582600000000
0!
0'
#582610000000
1!
b100 %
1'
b100 +
#582620000000
0!
0'
#582630000000
1!
b101 %
1'
b101 +
#582640000000
0!
0'
#582650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#582660000000
0!
0'
#582670000000
1!
b111 %
1'
b111 +
#582680000000
0!
0'
#582690000000
1!
b1000 %
1'
b1000 +
#582700000000
0!
0'
#582710000000
1!
b1001 %
1'
b1001 +
#582720000000
0!
0'
#582730000000
1!
b0 %
1'
b0 +
#582740000000
0!
0'
#582750000000
1!
1$
b1 %
1'
1*
b1 +
#582760000000
0!
0'
#582770000000
1!
b10 %
1'
b10 +
#582780000000
0!
0'
#582790000000
1!
b11 %
1'
b11 +
#582800000000
0!
0'
#582810000000
1!
b100 %
1'
b100 +
#582820000000
0!
0'
#582830000000
1!
b101 %
1'
b101 +
#582840000000
0!
0'
#582850000000
1!
0$
b110 %
1'
0*
b110 +
#582860000000
1"
1(
#582870000000
0!
0"
b100 &
0'
0(
b100 ,
#582880000000
1!
1$
b111 %
1'
1*
b111 +
#582890000000
0!
0'
#582900000000
1!
0$
b1000 %
1'
0*
b1000 +
#582910000000
0!
0'
#582920000000
1!
b1001 %
1'
b1001 +
#582930000000
0!
0'
#582940000000
1!
b0 %
1'
b0 +
#582950000000
0!
0'
#582960000000
1!
1$
b1 %
1'
1*
b1 +
#582970000000
0!
0'
#582980000000
1!
b10 %
1'
b10 +
#582990000000
0!
0'
#583000000000
1!
b11 %
1'
b11 +
#583010000000
0!
0'
#583020000000
1!
b100 %
1'
b100 +
#583030000000
0!
0'
#583040000000
1!
b101 %
1'
b101 +
#583050000000
0!
0'
#583060000000
1!
b110 %
1'
b110 +
#583070000000
0!
0'
#583080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#583090000000
0!
0'
#583100000000
1!
b1000 %
1'
b1000 +
#583110000000
0!
0'
#583120000000
1!
b1001 %
1'
b1001 +
#583130000000
0!
0'
#583140000000
1!
b0 %
1'
b0 +
#583150000000
0!
0'
#583160000000
1!
1$
b1 %
1'
1*
b1 +
#583170000000
0!
0'
#583180000000
1!
b10 %
1'
b10 +
#583190000000
0!
0'
#583200000000
1!
b11 %
1'
b11 +
#583210000000
0!
0'
#583220000000
1!
b100 %
1'
b100 +
#583230000000
0!
0'
#583240000000
1!
b101 %
1'
b101 +
#583250000000
0!
0'
#583260000000
1!
0$
b110 %
1'
0*
b110 +
#583270000000
0!
0'
#583280000000
1!
b111 %
1'
b111 +
#583290000000
1"
1(
#583300000000
0!
0"
b100 &
0'
0(
b100 ,
#583310000000
1!
b1000 %
1'
b1000 +
#583320000000
0!
0'
#583330000000
1!
b1001 %
1'
b1001 +
#583340000000
0!
0'
#583350000000
1!
b0 %
1'
b0 +
#583360000000
0!
0'
#583370000000
1!
1$
b1 %
1'
1*
b1 +
#583380000000
0!
0'
#583390000000
1!
b10 %
1'
b10 +
#583400000000
0!
0'
#583410000000
1!
b11 %
1'
b11 +
#583420000000
0!
0'
#583430000000
1!
b100 %
1'
b100 +
#583440000000
0!
0'
#583450000000
1!
b101 %
1'
b101 +
#583460000000
0!
0'
#583470000000
1!
b110 %
1'
b110 +
#583480000000
0!
0'
#583490000000
1!
b111 %
1'
b111 +
#583500000000
0!
0'
#583510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#583520000000
0!
0'
#583530000000
1!
b1001 %
1'
b1001 +
#583540000000
0!
0'
#583550000000
1!
b0 %
1'
b0 +
#583560000000
0!
0'
#583570000000
1!
1$
b1 %
1'
1*
b1 +
#583580000000
0!
0'
#583590000000
1!
b10 %
1'
b10 +
#583600000000
0!
0'
#583610000000
1!
b11 %
1'
b11 +
#583620000000
0!
0'
#583630000000
1!
b100 %
1'
b100 +
#583640000000
0!
0'
#583650000000
1!
b101 %
1'
b101 +
#583660000000
0!
0'
#583670000000
1!
0$
b110 %
1'
0*
b110 +
#583680000000
0!
0'
#583690000000
1!
b111 %
1'
b111 +
#583700000000
0!
0'
#583710000000
1!
b1000 %
1'
b1000 +
#583720000000
1"
1(
#583730000000
0!
0"
b100 &
0'
0(
b100 ,
#583740000000
1!
b1001 %
1'
b1001 +
#583750000000
0!
0'
#583760000000
1!
b0 %
1'
b0 +
#583770000000
0!
0'
#583780000000
1!
1$
b1 %
1'
1*
b1 +
#583790000000
0!
0'
#583800000000
1!
b10 %
1'
b10 +
#583810000000
0!
0'
#583820000000
1!
b11 %
1'
b11 +
#583830000000
0!
0'
#583840000000
1!
b100 %
1'
b100 +
#583850000000
0!
0'
#583860000000
1!
b101 %
1'
b101 +
#583870000000
0!
0'
#583880000000
1!
b110 %
1'
b110 +
#583890000000
0!
0'
#583900000000
1!
b111 %
1'
b111 +
#583910000000
0!
0'
#583920000000
1!
0$
b1000 %
1'
0*
b1000 +
#583930000000
0!
0'
#583940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#583950000000
0!
0'
#583960000000
1!
b0 %
1'
b0 +
#583970000000
0!
0'
#583980000000
1!
1$
b1 %
1'
1*
b1 +
#583990000000
0!
0'
#584000000000
1!
b10 %
1'
b10 +
#584010000000
0!
0'
#584020000000
1!
b11 %
1'
b11 +
#584030000000
0!
0'
#584040000000
1!
b100 %
1'
b100 +
#584050000000
0!
0'
#584060000000
1!
b101 %
1'
b101 +
#584070000000
0!
0'
#584080000000
1!
0$
b110 %
1'
0*
b110 +
#584090000000
0!
0'
#584100000000
1!
b111 %
1'
b111 +
#584110000000
0!
0'
#584120000000
1!
b1000 %
1'
b1000 +
#584130000000
0!
0'
#584140000000
1!
b1001 %
1'
b1001 +
#584150000000
1"
1(
#584160000000
0!
0"
b100 &
0'
0(
b100 ,
#584170000000
1!
b0 %
1'
b0 +
#584180000000
0!
0'
#584190000000
1!
1$
b1 %
1'
1*
b1 +
#584200000000
0!
0'
#584210000000
1!
b10 %
1'
b10 +
#584220000000
0!
0'
#584230000000
1!
b11 %
1'
b11 +
#584240000000
0!
0'
#584250000000
1!
b100 %
1'
b100 +
#584260000000
0!
0'
#584270000000
1!
b101 %
1'
b101 +
#584280000000
0!
0'
#584290000000
1!
b110 %
1'
b110 +
#584300000000
0!
0'
#584310000000
1!
b111 %
1'
b111 +
#584320000000
0!
0'
#584330000000
1!
0$
b1000 %
1'
0*
b1000 +
#584340000000
0!
0'
#584350000000
1!
b1001 %
1'
b1001 +
#584360000000
0!
0'
#584370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#584380000000
0!
0'
#584390000000
1!
1$
b1 %
1'
1*
b1 +
#584400000000
0!
0'
#584410000000
1!
b10 %
1'
b10 +
#584420000000
0!
0'
#584430000000
1!
b11 %
1'
b11 +
#584440000000
0!
0'
#584450000000
1!
b100 %
1'
b100 +
#584460000000
0!
0'
#584470000000
1!
b101 %
1'
b101 +
#584480000000
0!
0'
#584490000000
1!
0$
b110 %
1'
0*
b110 +
#584500000000
0!
0'
#584510000000
1!
b111 %
1'
b111 +
#584520000000
0!
0'
#584530000000
1!
b1000 %
1'
b1000 +
#584540000000
0!
0'
#584550000000
1!
b1001 %
1'
b1001 +
#584560000000
0!
0'
#584570000000
1!
b0 %
1'
b0 +
#584580000000
1"
1(
#584590000000
0!
0"
b100 &
0'
0(
b100 ,
#584600000000
1!
1$
b1 %
1'
1*
b1 +
#584610000000
0!
0'
#584620000000
1!
b10 %
1'
b10 +
#584630000000
0!
0'
#584640000000
1!
b11 %
1'
b11 +
#584650000000
0!
0'
#584660000000
1!
b100 %
1'
b100 +
#584670000000
0!
0'
#584680000000
1!
b101 %
1'
b101 +
#584690000000
0!
0'
#584700000000
1!
b110 %
1'
b110 +
#584710000000
0!
0'
#584720000000
1!
b111 %
1'
b111 +
#584730000000
0!
0'
#584740000000
1!
0$
b1000 %
1'
0*
b1000 +
#584750000000
0!
0'
#584760000000
1!
b1001 %
1'
b1001 +
#584770000000
0!
0'
#584780000000
1!
b0 %
1'
b0 +
#584790000000
0!
0'
#584800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#584810000000
0!
0'
#584820000000
1!
b10 %
1'
b10 +
#584830000000
0!
0'
#584840000000
1!
b11 %
1'
b11 +
#584850000000
0!
0'
#584860000000
1!
b100 %
1'
b100 +
#584870000000
0!
0'
#584880000000
1!
b101 %
1'
b101 +
#584890000000
0!
0'
#584900000000
1!
0$
b110 %
1'
0*
b110 +
#584910000000
0!
0'
#584920000000
1!
b111 %
1'
b111 +
#584930000000
0!
0'
#584940000000
1!
b1000 %
1'
b1000 +
#584950000000
0!
0'
#584960000000
1!
b1001 %
1'
b1001 +
#584970000000
0!
0'
#584980000000
1!
b0 %
1'
b0 +
#584990000000
0!
0'
#585000000000
1!
1$
b1 %
1'
1*
b1 +
#585010000000
1"
1(
#585020000000
0!
0"
b100 &
0'
0(
b100 ,
#585030000000
1!
b10 %
1'
b10 +
#585040000000
0!
0'
#585050000000
1!
b11 %
1'
b11 +
#585060000000
0!
0'
#585070000000
1!
b100 %
1'
b100 +
#585080000000
0!
0'
#585090000000
1!
b101 %
1'
b101 +
#585100000000
0!
0'
#585110000000
1!
b110 %
1'
b110 +
#585120000000
0!
0'
#585130000000
1!
b111 %
1'
b111 +
#585140000000
0!
0'
#585150000000
1!
0$
b1000 %
1'
0*
b1000 +
#585160000000
0!
0'
#585170000000
1!
b1001 %
1'
b1001 +
#585180000000
0!
0'
#585190000000
1!
b0 %
1'
b0 +
#585200000000
0!
0'
#585210000000
1!
1$
b1 %
1'
1*
b1 +
#585220000000
0!
0'
#585230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#585240000000
0!
0'
#585250000000
1!
b11 %
1'
b11 +
#585260000000
0!
0'
#585270000000
1!
b100 %
1'
b100 +
#585280000000
0!
0'
#585290000000
1!
b101 %
1'
b101 +
#585300000000
0!
0'
#585310000000
1!
0$
b110 %
1'
0*
b110 +
#585320000000
0!
0'
#585330000000
1!
b111 %
1'
b111 +
#585340000000
0!
0'
#585350000000
1!
b1000 %
1'
b1000 +
#585360000000
0!
0'
#585370000000
1!
b1001 %
1'
b1001 +
#585380000000
0!
0'
#585390000000
1!
b0 %
1'
b0 +
#585400000000
0!
0'
#585410000000
1!
1$
b1 %
1'
1*
b1 +
#585420000000
0!
0'
#585430000000
1!
b10 %
1'
b10 +
#585440000000
1"
1(
#585450000000
0!
0"
b100 &
0'
0(
b100 ,
#585460000000
1!
b11 %
1'
b11 +
#585470000000
0!
0'
#585480000000
1!
b100 %
1'
b100 +
#585490000000
0!
0'
#585500000000
1!
b101 %
1'
b101 +
#585510000000
0!
0'
#585520000000
1!
b110 %
1'
b110 +
#585530000000
0!
0'
#585540000000
1!
b111 %
1'
b111 +
#585550000000
0!
0'
#585560000000
1!
0$
b1000 %
1'
0*
b1000 +
#585570000000
0!
0'
#585580000000
1!
b1001 %
1'
b1001 +
#585590000000
0!
0'
#585600000000
1!
b0 %
1'
b0 +
#585610000000
0!
0'
#585620000000
1!
1$
b1 %
1'
1*
b1 +
#585630000000
0!
0'
#585640000000
1!
b10 %
1'
b10 +
#585650000000
0!
0'
#585660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#585670000000
0!
0'
#585680000000
1!
b100 %
1'
b100 +
#585690000000
0!
0'
#585700000000
1!
b101 %
1'
b101 +
#585710000000
0!
0'
#585720000000
1!
0$
b110 %
1'
0*
b110 +
#585730000000
0!
0'
#585740000000
1!
b111 %
1'
b111 +
#585750000000
0!
0'
#585760000000
1!
b1000 %
1'
b1000 +
#585770000000
0!
0'
#585780000000
1!
b1001 %
1'
b1001 +
#585790000000
0!
0'
#585800000000
1!
b0 %
1'
b0 +
#585810000000
0!
0'
#585820000000
1!
1$
b1 %
1'
1*
b1 +
#585830000000
0!
0'
#585840000000
1!
b10 %
1'
b10 +
#585850000000
0!
0'
#585860000000
1!
b11 %
1'
b11 +
#585870000000
1"
1(
#585880000000
0!
0"
b100 &
0'
0(
b100 ,
#585890000000
1!
b100 %
1'
b100 +
#585900000000
0!
0'
#585910000000
1!
b101 %
1'
b101 +
#585920000000
0!
0'
#585930000000
1!
b110 %
1'
b110 +
#585940000000
0!
0'
#585950000000
1!
b111 %
1'
b111 +
#585960000000
0!
0'
#585970000000
1!
0$
b1000 %
1'
0*
b1000 +
#585980000000
0!
0'
#585990000000
1!
b1001 %
1'
b1001 +
#586000000000
0!
0'
#586010000000
1!
b0 %
1'
b0 +
#586020000000
0!
0'
#586030000000
1!
1$
b1 %
1'
1*
b1 +
#586040000000
0!
0'
#586050000000
1!
b10 %
1'
b10 +
#586060000000
0!
0'
#586070000000
1!
b11 %
1'
b11 +
#586080000000
0!
0'
#586090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#586100000000
0!
0'
#586110000000
1!
b101 %
1'
b101 +
#586120000000
0!
0'
#586130000000
1!
0$
b110 %
1'
0*
b110 +
#586140000000
0!
0'
#586150000000
1!
b111 %
1'
b111 +
#586160000000
0!
0'
#586170000000
1!
b1000 %
1'
b1000 +
#586180000000
0!
0'
#586190000000
1!
b1001 %
1'
b1001 +
#586200000000
0!
0'
#586210000000
1!
b0 %
1'
b0 +
#586220000000
0!
0'
#586230000000
1!
1$
b1 %
1'
1*
b1 +
#586240000000
0!
0'
#586250000000
1!
b10 %
1'
b10 +
#586260000000
0!
0'
#586270000000
1!
b11 %
1'
b11 +
#586280000000
0!
0'
#586290000000
1!
b100 %
1'
b100 +
#586300000000
1"
1(
#586310000000
0!
0"
b100 &
0'
0(
b100 ,
#586320000000
1!
b101 %
1'
b101 +
#586330000000
0!
0'
#586340000000
1!
b110 %
1'
b110 +
#586350000000
0!
0'
#586360000000
1!
b111 %
1'
b111 +
#586370000000
0!
0'
#586380000000
1!
0$
b1000 %
1'
0*
b1000 +
#586390000000
0!
0'
#586400000000
1!
b1001 %
1'
b1001 +
#586410000000
0!
0'
#586420000000
1!
b0 %
1'
b0 +
#586430000000
0!
0'
#586440000000
1!
1$
b1 %
1'
1*
b1 +
#586450000000
0!
0'
#586460000000
1!
b10 %
1'
b10 +
#586470000000
0!
0'
#586480000000
1!
b11 %
1'
b11 +
#586490000000
0!
0'
#586500000000
1!
b100 %
1'
b100 +
#586510000000
0!
0'
#586520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#586530000000
0!
0'
#586540000000
1!
0$
b110 %
1'
0*
b110 +
#586550000000
0!
0'
#586560000000
1!
b111 %
1'
b111 +
#586570000000
0!
0'
#586580000000
1!
b1000 %
1'
b1000 +
#586590000000
0!
0'
#586600000000
1!
b1001 %
1'
b1001 +
#586610000000
0!
0'
#586620000000
1!
b0 %
1'
b0 +
#586630000000
0!
0'
#586640000000
1!
1$
b1 %
1'
1*
b1 +
#586650000000
0!
0'
#586660000000
1!
b10 %
1'
b10 +
#586670000000
0!
0'
#586680000000
1!
b11 %
1'
b11 +
#586690000000
0!
0'
#586700000000
1!
b100 %
1'
b100 +
#586710000000
0!
0'
#586720000000
1!
b101 %
1'
b101 +
#586730000000
1"
1(
#586740000000
0!
0"
b100 &
0'
0(
b100 ,
#586750000000
1!
b110 %
1'
b110 +
#586760000000
0!
0'
#586770000000
1!
b111 %
1'
b111 +
#586780000000
0!
0'
#586790000000
1!
0$
b1000 %
1'
0*
b1000 +
#586800000000
0!
0'
#586810000000
1!
b1001 %
1'
b1001 +
#586820000000
0!
0'
#586830000000
1!
b0 %
1'
b0 +
#586840000000
0!
0'
#586850000000
1!
1$
b1 %
1'
1*
b1 +
#586860000000
0!
0'
#586870000000
1!
b10 %
1'
b10 +
#586880000000
0!
0'
#586890000000
1!
b11 %
1'
b11 +
#586900000000
0!
0'
#586910000000
1!
b100 %
1'
b100 +
#586920000000
0!
0'
#586930000000
1!
b101 %
1'
b101 +
#586940000000
0!
0'
#586950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#586960000000
0!
0'
#586970000000
1!
b111 %
1'
b111 +
#586980000000
0!
0'
#586990000000
1!
b1000 %
1'
b1000 +
#587000000000
0!
0'
#587010000000
1!
b1001 %
1'
b1001 +
#587020000000
0!
0'
#587030000000
1!
b0 %
1'
b0 +
#587040000000
0!
0'
#587050000000
1!
1$
b1 %
1'
1*
b1 +
#587060000000
0!
0'
#587070000000
1!
b10 %
1'
b10 +
#587080000000
0!
0'
#587090000000
1!
b11 %
1'
b11 +
#587100000000
0!
0'
#587110000000
1!
b100 %
1'
b100 +
#587120000000
0!
0'
#587130000000
1!
b101 %
1'
b101 +
#587140000000
0!
0'
#587150000000
1!
0$
b110 %
1'
0*
b110 +
#587160000000
1"
1(
#587170000000
0!
0"
b100 &
0'
0(
b100 ,
#587180000000
1!
1$
b111 %
1'
1*
b111 +
#587190000000
0!
0'
#587200000000
1!
0$
b1000 %
1'
0*
b1000 +
#587210000000
0!
0'
#587220000000
1!
b1001 %
1'
b1001 +
#587230000000
0!
0'
#587240000000
1!
b0 %
1'
b0 +
#587250000000
0!
0'
#587260000000
1!
1$
b1 %
1'
1*
b1 +
#587270000000
0!
0'
#587280000000
1!
b10 %
1'
b10 +
#587290000000
0!
0'
#587300000000
1!
b11 %
1'
b11 +
#587310000000
0!
0'
#587320000000
1!
b100 %
1'
b100 +
#587330000000
0!
0'
#587340000000
1!
b101 %
1'
b101 +
#587350000000
0!
0'
#587360000000
1!
b110 %
1'
b110 +
#587370000000
0!
0'
#587380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#587390000000
0!
0'
#587400000000
1!
b1000 %
1'
b1000 +
#587410000000
0!
0'
#587420000000
1!
b1001 %
1'
b1001 +
#587430000000
0!
0'
#587440000000
1!
b0 %
1'
b0 +
#587450000000
0!
0'
#587460000000
1!
1$
b1 %
1'
1*
b1 +
#587470000000
0!
0'
#587480000000
1!
b10 %
1'
b10 +
#587490000000
0!
0'
#587500000000
1!
b11 %
1'
b11 +
#587510000000
0!
0'
#587520000000
1!
b100 %
1'
b100 +
#587530000000
0!
0'
#587540000000
1!
b101 %
1'
b101 +
#587550000000
0!
0'
#587560000000
1!
0$
b110 %
1'
0*
b110 +
#587570000000
0!
0'
#587580000000
1!
b111 %
1'
b111 +
#587590000000
1"
1(
#587600000000
0!
0"
b100 &
0'
0(
b100 ,
#587610000000
1!
b1000 %
1'
b1000 +
#587620000000
0!
0'
#587630000000
1!
b1001 %
1'
b1001 +
#587640000000
0!
0'
#587650000000
1!
b0 %
1'
b0 +
#587660000000
0!
0'
#587670000000
1!
1$
b1 %
1'
1*
b1 +
#587680000000
0!
0'
#587690000000
1!
b10 %
1'
b10 +
#587700000000
0!
0'
#587710000000
1!
b11 %
1'
b11 +
#587720000000
0!
0'
#587730000000
1!
b100 %
1'
b100 +
#587740000000
0!
0'
#587750000000
1!
b101 %
1'
b101 +
#587760000000
0!
0'
#587770000000
1!
b110 %
1'
b110 +
#587780000000
0!
0'
#587790000000
1!
b111 %
1'
b111 +
#587800000000
0!
0'
#587810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#587820000000
0!
0'
#587830000000
1!
b1001 %
1'
b1001 +
#587840000000
0!
0'
#587850000000
1!
b0 %
1'
b0 +
#587860000000
0!
0'
#587870000000
1!
1$
b1 %
1'
1*
b1 +
#587880000000
0!
0'
#587890000000
1!
b10 %
1'
b10 +
#587900000000
0!
0'
#587910000000
1!
b11 %
1'
b11 +
#587920000000
0!
0'
#587930000000
1!
b100 %
1'
b100 +
#587940000000
0!
0'
#587950000000
1!
b101 %
1'
b101 +
#587960000000
0!
0'
#587970000000
1!
0$
b110 %
1'
0*
b110 +
#587980000000
0!
0'
#587990000000
1!
b111 %
1'
b111 +
#588000000000
0!
0'
#588010000000
1!
b1000 %
1'
b1000 +
#588020000000
1"
1(
#588030000000
0!
0"
b100 &
0'
0(
b100 ,
#588040000000
1!
b1001 %
1'
b1001 +
#588050000000
0!
0'
#588060000000
1!
b0 %
1'
b0 +
#588070000000
0!
0'
#588080000000
1!
1$
b1 %
1'
1*
b1 +
#588090000000
0!
0'
#588100000000
1!
b10 %
1'
b10 +
#588110000000
0!
0'
#588120000000
1!
b11 %
1'
b11 +
#588130000000
0!
0'
#588140000000
1!
b100 %
1'
b100 +
#588150000000
0!
0'
#588160000000
1!
b101 %
1'
b101 +
#588170000000
0!
0'
#588180000000
1!
b110 %
1'
b110 +
#588190000000
0!
0'
#588200000000
1!
b111 %
1'
b111 +
#588210000000
0!
0'
#588220000000
1!
0$
b1000 %
1'
0*
b1000 +
#588230000000
0!
0'
#588240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#588250000000
0!
0'
#588260000000
1!
b0 %
1'
b0 +
#588270000000
0!
0'
#588280000000
1!
1$
b1 %
1'
1*
b1 +
#588290000000
0!
0'
#588300000000
1!
b10 %
1'
b10 +
#588310000000
0!
0'
#588320000000
1!
b11 %
1'
b11 +
#588330000000
0!
0'
#588340000000
1!
b100 %
1'
b100 +
#588350000000
0!
0'
#588360000000
1!
b101 %
1'
b101 +
#588370000000
0!
0'
#588380000000
1!
0$
b110 %
1'
0*
b110 +
#588390000000
0!
0'
#588400000000
1!
b111 %
1'
b111 +
#588410000000
0!
0'
#588420000000
1!
b1000 %
1'
b1000 +
#588430000000
0!
0'
#588440000000
1!
b1001 %
1'
b1001 +
#588450000000
1"
1(
#588460000000
0!
0"
b100 &
0'
0(
b100 ,
#588470000000
1!
b0 %
1'
b0 +
#588480000000
0!
0'
#588490000000
1!
1$
b1 %
1'
1*
b1 +
#588500000000
0!
0'
#588510000000
1!
b10 %
1'
b10 +
#588520000000
0!
0'
#588530000000
1!
b11 %
1'
b11 +
#588540000000
0!
0'
#588550000000
1!
b100 %
1'
b100 +
#588560000000
0!
0'
#588570000000
1!
b101 %
1'
b101 +
#588580000000
0!
0'
#588590000000
1!
b110 %
1'
b110 +
#588600000000
0!
0'
#588610000000
1!
b111 %
1'
b111 +
#588620000000
0!
0'
#588630000000
1!
0$
b1000 %
1'
0*
b1000 +
#588640000000
0!
0'
#588650000000
1!
b1001 %
1'
b1001 +
#588660000000
0!
0'
#588670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#588680000000
0!
0'
#588690000000
1!
1$
b1 %
1'
1*
b1 +
#588700000000
0!
0'
#588710000000
1!
b10 %
1'
b10 +
#588720000000
0!
0'
#588730000000
1!
b11 %
1'
b11 +
#588740000000
0!
0'
#588750000000
1!
b100 %
1'
b100 +
#588760000000
0!
0'
#588770000000
1!
b101 %
1'
b101 +
#588780000000
0!
0'
#588790000000
1!
0$
b110 %
1'
0*
b110 +
#588800000000
0!
0'
#588810000000
1!
b111 %
1'
b111 +
#588820000000
0!
0'
#588830000000
1!
b1000 %
1'
b1000 +
#588840000000
0!
0'
#588850000000
1!
b1001 %
1'
b1001 +
#588860000000
0!
0'
#588870000000
1!
b0 %
1'
b0 +
#588880000000
1"
1(
#588890000000
0!
0"
b100 &
0'
0(
b100 ,
#588900000000
1!
1$
b1 %
1'
1*
b1 +
#588910000000
0!
0'
#588920000000
1!
b10 %
1'
b10 +
#588930000000
0!
0'
#588940000000
1!
b11 %
1'
b11 +
#588950000000
0!
0'
#588960000000
1!
b100 %
1'
b100 +
#588970000000
0!
0'
#588980000000
1!
b101 %
1'
b101 +
#588990000000
0!
0'
#589000000000
1!
b110 %
1'
b110 +
#589010000000
0!
0'
#589020000000
1!
b111 %
1'
b111 +
#589030000000
0!
0'
#589040000000
1!
0$
b1000 %
1'
0*
b1000 +
#589050000000
0!
0'
#589060000000
1!
b1001 %
1'
b1001 +
#589070000000
0!
0'
#589080000000
1!
b0 %
1'
b0 +
#589090000000
0!
0'
#589100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#589110000000
0!
0'
#589120000000
1!
b10 %
1'
b10 +
#589130000000
0!
0'
#589140000000
1!
b11 %
1'
b11 +
#589150000000
0!
0'
#589160000000
1!
b100 %
1'
b100 +
#589170000000
0!
0'
#589180000000
1!
b101 %
1'
b101 +
#589190000000
0!
0'
#589200000000
1!
0$
b110 %
1'
0*
b110 +
#589210000000
0!
0'
#589220000000
1!
b111 %
1'
b111 +
#589230000000
0!
0'
#589240000000
1!
b1000 %
1'
b1000 +
#589250000000
0!
0'
#589260000000
1!
b1001 %
1'
b1001 +
#589270000000
0!
0'
#589280000000
1!
b0 %
1'
b0 +
#589290000000
0!
0'
#589300000000
1!
1$
b1 %
1'
1*
b1 +
#589310000000
1"
1(
#589320000000
0!
0"
b100 &
0'
0(
b100 ,
#589330000000
1!
b10 %
1'
b10 +
#589340000000
0!
0'
#589350000000
1!
b11 %
1'
b11 +
#589360000000
0!
0'
#589370000000
1!
b100 %
1'
b100 +
#589380000000
0!
0'
#589390000000
1!
b101 %
1'
b101 +
#589400000000
0!
0'
#589410000000
1!
b110 %
1'
b110 +
#589420000000
0!
0'
#589430000000
1!
b111 %
1'
b111 +
#589440000000
0!
0'
#589450000000
1!
0$
b1000 %
1'
0*
b1000 +
#589460000000
0!
0'
#589470000000
1!
b1001 %
1'
b1001 +
#589480000000
0!
0'
#589490000000
1!
b0 %
1'
b0 +
#589500000000
0!
0'
#589510000000
1!
1$
b1 %
1'
1*
b1 +
#589520000000
0!
0'
#589530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#589540000000
0!
0'
#589550000000
1!
b11 %
1'
b11 +
#589560000000
0!
0'
#589570000000
1!
b100 %
1'
b100 +
#589580000000
0!
0'
#589590000000
1!
b101 %
1'
b101 +
#589600000000
0!
0'
#589610000000
1!
0$
b110 %
1'
0*
b110 +
#589620000000
0!
0'
#589630000000
1!
b111 %
1'
b111 +
#589640000000
0!
0'
#589650000000
1!
b1000 %
1'
b1000 +
#589660000000
0!
0'
#589670000000
1!
b1001 %
1'
b1001 +
#589680000000
0!
0'
#589690000000
1!
b0 %
1'
b0 +
#589700000000
0!
0'
#589710000000
1!
1$
b1 %
1'
1*
b1 +
#589720000000
0!
0'
#589730000000
1!
b10 %
1'
b10 +
#589740000000
1"
1(
#589750000000
0!
0"
b100 &
0'
0(
b100 ,
#589760000000
1!
b11 %
1'
b11 +
#589770000000
0!
0'
#589780000000
1!
b100 %
1'
b100 +
#589790000000
0!
0'
#589800000000
1!
b101 %
1'
b101 +
#589810000000
0!
0'
#589820000000
1!
b110 %
1'
b110 +
#589830000000
0!
0'
#589840000000
1!
b111 %
1'
b111 +
#589850000000
0!
0'
#589860000000
1!
0$
b1000 %
1'
0*
b1000 +
#589870000000
0!
0'
#589880000000
1!
b1001 %
1'
b1001 +
#589890000000
0!
0'
#589900000000
1!
b0 %
1'
b0 +
#589910000000
0!
0'
#589920000000
1!
1$
b1 %
1'
1*
b1 +
#589930000000
0!
0'
#589940000000
1!
b10 %
1'
b10 +
#589950000000
0!
0'
#589960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#589970000000
0!
0'
#589980000000
1!
b100 %
1'
b100 +
#589990000000
0!
0'
#590000000000
1!
b101 %
1'
b101 +
#590010000000
0!
0'
#590020000000
1!
0$
b110 %
1'
0*
b110 +
#590030000000
0!
0'
#590040000000
1!
b111 %
1'
b111 +
#590050000000
0!
0'
#590060000000
1!
b1000 %
1'
b1000 +
#590070000000
0!
0'
#590080000000
1!
b1001 %
1'
b1001 +
#590090000000
0!
0'
#590100000000
1!
b0 %
1'
b0 +
#590110000000
0!
0'
#590120000000
1!
1$
b1 %
1'
1*
b1 +
#590130000000
0!
0'
#590140000000
1!
b10 %
1'
b10 +
#590150000000
0!
0'
#590160000000
1!
b11 %
1'
b11 +
#590170000000
1"
1(
#590180000000
0!
0"
b100 &
0'
0(
b100 ,
#590190000000
1!
b100 %
1'
b100 +
#590200000000
0!
0'
#590210000000
1!
b101 %
1'
b101 +
#590220000000
0!
0'
#590230000000
1!
b110 %
1'
b110 +
#590240000000
0!
0'
#590250000000
1!
b111 %
1'
b111 +
#590260000000
0!
0'
#590270000000
1!
0$
b1000 %
1'
0*
b1000 +
#590280000000
0!
0'
#590290000000
1!
b1001 %
1'
b1001 +
#590300000000
0!
0'
#590310000000
1!
b0 %
1'
b0 +
#590320000000
0!
0'
#590330000000
1!
1$
b1 %
1'
1*
b1 +
#590340000000
0!
0'
#590350000000
1!
b10 %
1'
b10 +
#590360000000
0!
0'
#590370000000
1!
b11 %
1'
b11 +
#590380000000
0!
0'
#590390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#590400000000
0!
0'
#590410000000
1!
b101 %
1'
b101 +
#590420000000
0!
0'
#590430000000
1!
0$
b110 %
1'
0*
b110 +
#590440000000
0!
0'
#590450000000
1!
b111 %
1'
b111 +
#590460000000
0!
0'
#590470000000
1!
b1000 %
1'
b1000 +
#590480000000
0!
0'
#590490000000
1!
b1001 %
1'
b1001 +
#590500000000
0!
0'
#590510000000
1!
b0 %
1'
b0 +
#590520000000
0!
0'
#590530000000
1!
1$
b1 %
1'
1*
b1 +
#590540000000
0!
0'
#590550000000
1!
b10 %
1'
b10 +
#590560000000
0!
0'
#590570000000
1!
b11 %
1'
b11 +
#590580000000
0!
0'
#590590000000
1!
b100 %
1'
b100 +
#590600000000
1"
1(
#590610000000
0!
0"
b100 &
0'
0(
b100 ,
#590620000000
1!
b101 %
1'
b101 +
#590630000000
0!
0'
#590640000000
1!
b110 %
1'
b110 +
#590650000000
0!
0'
#590660000000
1!
b111 %
1'
b111 +
#590670000000
0!
0'
#590680000000
1!
0$
b1000 %
1'
0*
b1000 +
#590690000000
0!
0'
#590700000000
1!
b1001 %
1'
b1001 +
#590710000000
0!
0'
#590720000000
1!
b0 %
1'
b0 +
#590730000000
0!
0'
#590740000000
1!
1$
b1 %
1'
1*
b1 +
#590750000000
0!
0'
#590760000000
1!
b10 %
1'
b10 +
#590770000000
0!
0'
#590780000000
1!
b11 %
1'
b11 +
#590790000000
0!
0'
#590800000000
1!
b100 %
1'
b100 +
#590810000000
0!
0'
#590820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#590830000000
0!
0'
#590840000000
1!
0$
b110 %
1'
0*
b110 +
#590850000000
0!
0'
#590860000000
1!
b111 %
1'
b111 +
#590870000000
0!
0'
#590880000000
1!
b1000 %
1'
b1000 +
#590890000000
0!
0'
#590900000000
1!
b1001 %
1'
b1001 +
#590910000000
0!
0'
#590920000000
1!
b0 %
1'
b0 +
#590930000000
0!
0'
#590940000000
1!
1$
b1 %
1'
1*
b1 +
#590950000000
0!
0'
#590960000000
1!
b10 %
1'
b10 +
#590970000000
0!
0'
#590980000000
1!
b11 %
1'
b11 +
#590990000000
0!
0'
#591000000000
1!
b100 %
1'
b100 +
#591010000000
0!
0'
#591020000000
1!
b101 %
1'
b101 +
#591030000000
1"
1(
#591040000000
0!
0"
b100 &
0'
0(
b100 ,
#591050000000
1!
b110 %
1'
b110 +
#591060000000
0!
0'
#591070000000
1!
b111 %
1'
b111 +
#591080000000
0!
0'
#591090000000
1!
0$
b1000 %
1'
0*
b1000 +
#591100000000
0!
0'
#591110000000
1!
b1001 %
1'
b1001 +
#591120000000
0!
0'
#591130000000
1!
b0 %
1'
b0 +
#591140000000
0!
0'
#591150000000
1!
1$
b1 %
1'
1*
b1 +
#591160000000
0!
0'
#591170000000
1!
b10 %
1'
b10 +
#591180000000
0!
0'
#591190000000
1!
b11 %
1'
b11 +
#591200000000
0!
0'
#591210000000
1!
b100 %
1'
b100 +
#591220000000
0!
0'
#591230000000
1!
b101 %
1'
b101 +
#591240000000
0!
0'
#591250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#591260000000
0!
0'
#591270000000
1!
b111 %
1'
b111 +
#591280000000
0!
0'
#591290000000
1!
b1000 %
1'
b1000 +
#591300000000
0!
0'
#591310000000
1!
b1001 %
1'
b1001 +
#591320000000
0!
0'
#591330000000
1!
b0 %
1'
b0 +
#591340000000
0!
0'
#591350000000
1!
1$
b1 %
1'
1*
b1 +
#591360000000
0!
0'
#591370000000
1!
b10 %
1'
b10 +
#591380000000
0!
0'
#591390000000
1!
b11 %
1'
b11 +
#591400000000
0!
0'
#591410000000
1!
b100 %
1'
b100 +
#591420000000
0!
0'
#591430000000
1!
b101 %
1'
b101 +
#591440000000
0!
0'
#591450000000
1!
0$
b110 %
1'
0*
b110 +
#591460000000
1"
1(
#591470000000
0!
0"
b100 &
0'
0(
b100 ,
#591480000000
1!
1$
b111 %
1'
1*
b111 +
#591490000000
0!
0'
#591500000000
1!
0$
b1000 %
1'
0*
b1000 +
#591510000000
0!
0'
#591520000000
1!
b1001 %
1'
b1001 +
#591530000000
0!
0'
#591540000000
1!
b0 %
1'
b0 +
#591550000000
0!
0'
#591560000000
1!
1$
b1 %
1'
1*
b1 +
#591570000000
0!
0'
#591580000000
1!
b10 %
1'
b10 +
#591590000000
0!
0'
#591600000000
1!
b11 %
1'
b11 +
#591610000000
0!
0'
#591620000000
1!
b100 %
1'
b100 +
#591630000000
0!
0'
#591640000000
1!
b101 %
1'
b101 +
#591650000000
0!
0'
#591660000000
1!
b110 %
1'
b110 +
#591670000000
0!
0'
#591680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#591690000000
0!
0'
#591700000000
1!
b1000 %
1'
b1000 +
#591710000000
0!
0'
#591720000000
1!
b1001 %
1'
b1001 +
#591730000000
0!
0'
#591740000000
1!
b0 %
1'
b0 +
#591750000000
0!
0'
#591760000000
1!
1$
b1 %
1'
1*
b1 +
#591770000000
0!
0'
#591780000000
1!
b10 %
1'
b10 +
#591790000000
0!
0'
#591800000000
1!
b11 %
1'
b11 +
#591810000000
0!
0'
#591820000000
1!
b100 %
1'
b100 +
#591830000000
0!
0'
#591840000000
1!
b101 %
1'
b101 +
#591850000000
0!
0'
#591860000000
1!
0$
b110 %
1'
0*
b110 +
#591870000000
0!
0'
#591880000000
1!
b111 %
1'
b111 +
#591890000000
1"
1(
#591900000000
0!
0"
b100 &
0'
0(
b100 ,
#591910000000
1!
b1000 %
1'
b1000 +
#591920000000
0!
0'
#591930000000
1!
b1001 %
1'
b1001 +
#591940000000
0!
0'
#591950000000
1!
b0 %
1'
b0 +
#591960000000
0!
0'
#591970000000
1!
1$
b1 %
1'
1*
b1 +
#591980000000
0!
0'
#591990000000
1!
b10 %
1'
b10 +
#592000000000
0!
0'
#592010000000
1!
b11 %
1'
b11 +
#592020000000
0!
0'
#592030000000
1!
b100 %
1'
b100 +
#592040000000
0!
0'
#592050000000
1!
b101 %
1'
b101 +
#592060000000
0!
0'
#592070000000
1!
b110 %
1'
b110 +
#592080000000
0!
0'
#592090000000
1!
b111 %
1'
b111 +
#592100000000
0!
0'
#592110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#592120000000
0!
0'
#592130000000
1!
b1001 %
1'
b1001 +
#592140000000
0!
0'
#592150000000
1!
b0 %
1'
b0 +
#592160000000
0!
0'
#592170000000
1!
1$
b1 %
1'
1*
b1 +
#592180000000
0!
0'
#592190000000
1!
b10 %
1'
b10 +
#592200000000
0!
0'
#592210000000
1!
b11 %
1'
b11 +
#592220000000
0!
0'
#592230000000
1!
b100 %
1'
b100 +
#592240000000
0!
0'
#592250000000
1!
b101 %
1'
b101 +
#592260000000
0!
0'
#592270000000
1!
0$
b110 %
1'
0*
b110 +
#592280000000
0!
0'
#592290000000
1!
b111 %
1'
b111 +
#592300000000
0!
0'
#592310000000
1!
b1000 %
1'
b1000 +
#592320000000
1"
1(
#592330000000
0!
0"
b100 &
0'
0(
b100 ,
#592340000000
1!
b1001 %
1'
b1001 +
#592350000000
0!
0'
#592360000000
1!
b0 %
1'
b0 +
#592370000000
0!
0'
#592380000000
1!
1$
b1 %
1'
1*
b1 +
#592390000000
0!
0'
#592400000000
1!
b10 %
1'
b10 +
#592410000000
0!
0'
#592420000000
1!
b11 %
1'
b11 +
#592430000000
0!
0'
#592440000000
1!
b100 %
1'
b100 +
#592450000000
0!
0'
#592460000000
1!
b101 %
1'
b101 +
#592470000000
0!
0'
#592480000000
1!
b110 %
1'
b110 +
#592490000000
0!
0'
#592500000000
1!
b111 %
1'
b111 +
#592510000000
0!
0'
#592520000000
1!
0$
b1000 %
1'
0*
b1000 +
#592530000000
0!
0'
#592540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#592550000000
0!
0'
#592560000000
1!
b0 %
1'
b0 +
#592570000000
0!
0'
#592580000000
1!
1$
b1 %
1'
1*
b1 +
#592590000000
0!
0'
#592600000000
1!
b10 %
1'
b10 +
#592610000000
0!
0'
#592620000000
1!
b11 %
1'
b11 +
#592630000000
0!
0'
#592640000000
1!
b100 %
1'
b100 +
#592650000000
0!
0'
#592660000000
1!
b101 %
1'
b101 +
#592670000000
0!
0'
#592680000000
1!
0$
b110 %
1'
0*
b110 +
#592690000000
0!
0'
#592700000000
1!
b111 %
1'
b111 +
#592710000000
0!
0'
#592720000000
1!
b1000 %
1'
b1000 +
#592730000000
0!
0'
#592740000000
1!
b1001 %
1'
b1001 +
#592750000000
1"
1(
#592760000000
0!
0"
b100 &
0'
0(
b100 ,
#592770000000
1!
b0 %
1'
b0 +
#592780000000
0!
0'
#592790000000
1!
1$
b1 %
1'
1*
b1 +
#592800000000
0!
0'
#592810000000
1!
b10 %
1'
b10 +
#592820000000
0!
0'
#592830000000
1!
b11 %
1'
b11 +
#592840000000
0!
0'
#592850000000
1!
b100 %
1'
b100 +
#592860000000
0!
0'
#592870000000
1!
b101 %
1'
b101 +
#592880000000
0!
0'
#592890000000
1!
b110 %
1'
b110 +
#592900000000
0!
0'
#592910000000
1!
b111 %
1'
b111 +
#592920000000
0!
0'
#592930000000
1!
0$
b1000 %
1'
0*
b1000 +
#592940000000
0!
0'
#592950000000
1!
b1001 %
1'
b1001 +
#592960000000
0!
0'
#592970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#592980000000
0!
0'
#592990000000
1!
1$
b1 %
1'
1*
b1 +
#593000000000
0!
0'
#593010000000
1!
b10 %
1'
b10 +
#593020000000
0!
0'
#593030000000
1!
b11 %
1'
b11 +
#593040000000
0!
0'
#593050000000
1!
b100 %
1'
b100 +
#593060000000
0!
0'
#593070000000
1!
b101 %
1'
b101 +
#593080000000
0!
0'
#593090000000
1!
0$
b110 %
1'
0*
b110 +
#593100000000
0!
0'
#593110000000
1!
b111 %
1'
b111 +
#593120000000
0!
0'
#593130000000
1!
b1000 %
1'
b1000 +
#593140000000
0!
0'
#593150000000
1!
b1001 %
1'
b1001 +
#593160000000
0!
0'
#593170000000
1!
b0 %
1'
b0 +
#593180000000
1"
1(
#593190000000
0!
0"
b100 &
0'
0(
b100 ,
#593200000000
1!
1$
b1 %
1'
1*
b1 +
#593210000000
0!
0'
#593220000000
1!
b10 %
1'
b10 +
#593230000000
0!
0'
#593240000000
1!
b11 %
1'
b11 +
#593250000000
0!
0'
#593260000000
1!
b100 %
1'
b100 +
#593270000000
0!
0'
#593280000000
1!
b101 %
1'
b101 +
#593290000000
0!
0'
#593300000000
1!
b110 %
1'
b110 +
#593310000000
0!
0'
#593320000000
1!
b111 %
1'
b111 +
#593330000000
0!
0'
#593340000000
1!
0$
b1000 %
1'
0*
b1000 +
#593350000000
0!
0'
#593360000000
1!
b1001 %
1'
b1001 +
#593370000000
0!
0'
#593380000000
1!
b0 %
1'
b0 +
#593390000000
0!
0'
#593400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#593410000000
0!
0'
#593420000000
1!
b10 %
1'
b10 +
#593430000000
0!
0'
#593440000000
1!
b11 %
1'
b11 +
#593450000000
0!
0'
#593460000000
1!
b100 %
1'
b100 +
#593470000000
0!
0'
#593480000000
1!
b101 %
1'
b101 +
#593490000000
0!
0'
#593500000000
1!
0$
b110 %
1'
0*
b110 +
#593510000000
0!
0'
#593520000000
1!
b111 %
1'
b111 +
#593530000000
0!
0'
#593540000000
1!
b1000 %
1'
b1000 +
#593550000000
0!
0'
#593560000000
1!
b1001 %
1'
b1001 +
#593570000000
0!
0'
#593580000000
1!
b0 %
1'
b0 +
#593590000000
0!
0'
#593600000000
1!
1$
b1 %
1'
1*
b1 +
#593610000000
1"
1(
#593620000000
0!
0"
b100 &
0'
0(
b100 ,
#593630000000
1!
b10 %
1'
b10 +
#593640000000
0!
0'
#593650000000
1!
b11 %
1'
b11 +
#593660000000
0!
0'
#593670000000
1!
b100 %
1'
b100 +
#593680000000
0!
0'
#593690000000
1!
b101 %
1'
b101 +
#593700000000
0!
0'
#593710000000
1!
b110 %
1'
b110 +
#593720000000
0!
0'
#593730000000
1!
b111 %
1'
b111 +
#593740000000
0!
0'
#593750000000
1!
0$
b1000 %
1'
0*
b1000 +
#593760000000
0!
0'
#593770000000
1!
b1001 %
1'
b1001 +
#593780000000
0!
0'
#593790000000
1!
b0 %
1'
b0 +
#593800000000
0!
0'
#593810000000
1!
1$
b1 %
1'
1*
b1 +
#593820000000
0!
0'
#593830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#593840000000
0!
0'
#593850000000
1!
b11 %
1'
b11 +
#593860000000
0!
0'
#593870000000
1!
b100 %
1'
b100 +
#593880000000
0!
0'
#593890000000
1!
b101 %
1'
b101 +
#593900000000
0!
0'
#593910000000
1!
0$
b110 %
1'
0*
b110 +
#593920000000
0!
0'
#593930000000
1!
b111 %
1'
b111 +
#593940000000
0!
0'
#593950000000
1!
b1000 %
1'
b1000 +
#593960000000
0!
0'
#593970000000
1!
b1001 %
1'
b1001 +
#593980000000
0!
0'
#593990000000
1!
b0 %
1'
b0 +
#594000000000
0!
0'
#594010000000
1!
1$
b1 %
1'
1*
b1 +
#594020000000
0!
0'
#594030000000
1!
b10 %
1'
b10 +
#594040000000
1"
1(
#594050000000
0!
0"
b100 &
0'
0(
b100 ,
#594060000000
1!
b11 %
1'
b11 +
#594070000000
0!
0'
#594080000000
1!
b100 %
1'
b100 +
#594090000000
0!
0'
#594100000000
1!
b101 %
1'
b101 +
#594110000000
0!
0'
#594120000000
1!
b110 %
1'
b110 +
#594130000000
0!
0'
#594140000000
1!
b111 %
1'
b111 +
#594150000000
0!
0'
#594160000000
1!
0$
b1000 %
1'
0*
b1000 +
#594170000000
0!
0'
#594180000000
1!
b1001 %
1'
b1001 +
#594190000000
0!
0'
#594200000000
1!
b0 %
1'
b0 +
#594210000000
0!
0'
#594220000000
1!
1$
b1 %
1'
1*
b1 +
#594230000000
0!
0'
#594240000000
1!
b10 %
1'
b10 +
#594250000000
0!
0'
#594260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#594270000000
0!
0'
#594280000000
1!
b100 %
1'
b100 +
#594290000000
0!
0'
#594300000000
1!
b101 %
1'
b101 +
#594310000000
0!
0'
#594320000000
1!
0$
b110 %
1'
0*
b110 +
#594330000000
0!
0'
#594340000000
1!
b111 %
1'
b111 +
#594350000000
0!
0'
#594360000000
1!
b1000 %
1'
b1000 +
#594370000000
0!
0'
#594380000000
1!
b1001 %
1'
b1001 +
#594390000000
0!
0'
#594400000000
1!
b0 %
1'
b0 +
#594410000000
0!
0'
#594420000000
1!
1$
b1 %
1'
1*
b1 +
#594430000000
0!
0'
#594440000000
1!
b10 %
1'
b10 +
#594450000000
0!
0'
#594460000000
1!
b11 %
1'
b11 +
#594470000000
1"
1(
#594480000000
0!
0"
b100 &
0'
0(
b100 ,
#594490000000
1!
b100 %
1'
b100 +
#594500000000
0!
0'
#594510000000
1!
b101 %
1'
b101 +
#594520000000
0!
0'
#594530000000
1!
b110 %
1'
b110 +
#594540000000
0!
0'
#594550000000
1!
b111 %
1'
b111 +
#594560000000
0!
0'
#594570000000
1!
0$
b1000 %
1'
0*
b1000 +
#594580000000
0!
0'
#594590000000
1!
b1001 %
1'
b1001 +
#594600000000
0!
0'
#594610000000
1!
b0 %
1'
b0 +
#594620000000
0!
0'
#594630000000
1!
1$
b1 %
1'
1*
b1 +
#594640000000
0!
0'
#594650000000
1!
b10 %
1'
b10 +
#594660000000
0!
0'
#594670000000
1!
b11 %
1'
b11 +
#594680000000
0!
0'
#594690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#594700000000
0!
0'
#594710000000
1!
b101 %
1'
b101 +
#594720000000
0!
0'
#594730000000
1!
0$
b110 %
1'
0*
b110 +
#594740000000
0!
0'
#594750000000
1!
b111 %
1'
b111 +
#594760000000
0!
0'
#594770000000
1!
b1000 %
1'
b1000 +
#594780000000
0!
0'
#594790000000
1!
b1001 %
1'
b1001 +
#594800000000
0!
0'
#594810000000
1!
b0 %
1'
b0 +
#594820000000
0!
0'
#594830000000
1!
1$
b1 %
1'
1*
b1 +
#594840000000
0!
0'
#594850000000
1!
b10 %
1'
b10 +
#594860000000
0!
0'
#594870000000
1!
b11 %
1'
b11 +
#594880000000
0!
0'
#594890000000
1!
b100 %
1'
b100 +
#594900000000
1"
1(
#594910000000
0!
0"
b100 &
0'
0(
b100 ,
#594920000000
1!
b101 %
1'
b101 +
#594930000000
0!
0'
#594940000000
1!
b110 %
1'
b110 +
#594950000000
0!
0'
#594960000000
1!
b111 %
1'
b111 +
#594970000000
0!
0'
#594980000000
1!
0$
b1000 %
1'
0*
b1000 +
#594990000000
0!
0'
#595000000000
1!
b1001 %
1'
b1001 +
#595010000000
0!
0'
#595020000000
1!
b0 %
1'
b0 +
#595030000000
0!
0'
#595040000000
1!
1$
b1 %
1'
1*
b1 +
#595050000000
0!
0'
#595060000000
1!
b10 %
1'
b10 +
#595070000000
0!
0'
#595080000000
1!
b11 %
1'
b11 +
#595090000000
0!
0'
#595100000000
1!
b100 %
1'
b100 +
#595110000000
0!
0'
#595120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#595130000000
0!
0'
#595140000000
1!
0$
b110 %
1'
0*
b110 +
#595150000000
0!
0'
#595160000000
1!
b111 %
1'
b111 +
#595170000000
0!
0'
#595180000000
1!
b1000 %
1'
b1000 +
#595190000000
0!
0'
#595200000000
1!
b1001 %
1'
b1001 +
#595210000000
0!
0'
#595220000000
1!
b0 %
1'
b0 +
#595230000000
0!
0'
#595240000000
1!
1$
b1 %
1'
1*
b1 +
#595250000000
0!
0'
#595260000000
1!
b10 %
1'
b10 +
#595270000000
0!
0'
#595280000000
1!
b11 %
1'
b11 +
#595290000000
0!
0'
#595300000000
1!
b100 %
1'
b100 +
#595310000000
0!
0'
#595320000000
1!
b101 %
1'
b101 +
#595330000000
1"
1(
#595340000000
0!
0"
b100 &
0'
0(
b100 ,
#595350000000
1!
b110 %
1'
b110 +
#595360000000
0!
0'
#595370000000
1!
b111 %
1'
b111 +
#595380000000
0!
0'
#595390000000
1!
0$
b1000 %
1'
0*
b1000 +
#595400000000
0!
0'
#595410000000
1!
b1001 %
1'
b1001 +
#595420000000
0!
0'
#595430000000
1!
b0 %
1'
b0 +
#595440000000
0!
0'
#595450000000
1!
1$
b1 %
1'
1*
b1 +
#595460000000
0!
0'
#595470000000
1!
b10 %
1'
b10 +
#595480000000
0!
0'
#595490000000
1!
b11 %
1'
b11 +
#595500000000
0!
0'
#595510000000
1!
b100 %
1'
b100 +
#595520000000
0!
0'
#595530000000
1!
b101 %
1'
b101 +
#595540000000
0!
0'
#595550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#595560000000
0!
0'
#595570000000
1!
b111 %
1'
b111 +
#595580000000
0!
0'
#595590000000
1!
b1000 %
1'
b1000 +
#595600000000
0!
0'
#595610000000
1!
b1001 %
1'
b1001 +
#595620000000
0!
0'
#595630000000
1!
b0 %
1'
b0 +
#595640000000
0!
0'
#595650000000
1!
1$
b1 %
1'
1*
b1 +
#595660000000
0!
0'
#595670000000
1!
b10 %
1'
b10 +
#595680000000
0!
0'
#595690000000
1!
b11 %
1'
b11 +
#595700000000
0!
0'
#595710000000
1!
b100 %
1'
b100 +
#595720000000
0!
0'
#595730000000
1!
b101 %
1'
b101 +
#595740000000
0!
0'
#595750000000
1!
0$
b110 %
1'
0*
b110 +
#595760000000
1"
1(
#595770000000
0!
0"
b100 &
0'
0(
b100 ,
#595780000000
1!
1$
b111 %
1'
1*
b111 +
#595790000000
0!
0'
#595800000000
1!
0$
b1000 %
1'
0*
b1000 +
#595810000000
0!
0'
#595820000000
1!
b1001 %
1'
b1001 +
#595830000000
0!
0'
#595840000000
1!
b0 %
1'
b0 +
#595850000000
0!
0'
#595860000000
1!
1$
b1 %
1'
1*
b1 +
#595870000000
0!
0'
#595880000000
1!
b10 %
1'
b10 +
#595890000000
0!
0'
#595900000000
1!
b11 %
1'
b11 +
#595910000000
0!
0'
#595920000000
1!
b100 %
1'
b100 +
#595930000000
0!
0'
#595940000000
1!
b101 %
1'
b101 +
#595950000000
0!
0'
#595960000000
1!
b110 %
1'
b110 +
#595970000000
0!
0'
#595980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#595990000000
0!
0'
#596000000000
1!
b1000 %
1'
b1000 +
#596010000000
0!
0'
#596020000000
1!
b1001 %
1'
b1001 +
#596030000000
0!
0'
#596040000000
1!
b0 %
1'
b0 +
#596050000000
0!
0'
#596060000000
1!
1$
b1 %
1'
1*
b1 +
#596070000000
0!
0'
#596080000000
1!
b10 %
1'
b10 +
#596090000000
0!
0'
#596100000000
1!
b11 %
1'
b11 +
#596110000000
0!
0'
#596120000000
1!
b100 %
1'
b100 +
#596130000000
0!
0'
#596140000000
1!
b101 %
1'
b101 +
#596150000000
0!
0'
#596160000000
1!
0$
b110 %
1'
0*
b110 +
#596170000000
0!
0'
#596180000000
1!
b111 %
1'
b111 +
#596190000000
1"
1(
#596200000000
0!
0"
b100 &
0'
0(
b100 ,
#596210000000
1!
b1000 %
1'
b1000 +
#596220000000
0!
0'
#596230000000
1!
b1001 %
1'
b1001 +
#596240000000
0!
0'
#596250000000
1!
b0 %
1'
b0 +
#596260000000
0!
0'
#596270000000
1!
1$
b1 %
1'
1*
b1 +
#596280000000
0!
0'
#596290000000
1!
b10 %
1'
b10 +
#596300000000
0!
0'
#596310000000
1!
b11 %
1'
b11 +
#596320000000
0!
0'
#596330000000
1!
b100 %
1'
b100 +
#596340000000
0!
0'
#596350000000
1!
b101 %
1'
b101 +
#596360000000
0!
0'
#596370000000
1!
b110 %
1'
b110 +
#596380000000
0!
0'
#596390000000
1!
b111 %
1'
b111 +
#596400000000
0!
0'
#596410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#596420000000
0!
0'
#596430000000
1!
b1001 %
1'
b1001 +
#596440000000
0!
0'
#596450000000
1!
b0 %
1'
b0 +
#596460000000
0!
0'
#596470000000
1!
1$
b1 %
1'
1*
b1 +
#596480000000
0!
0'
#596490000000
1!
b10 %
1'
b10 +
#596500000000
0!
0'
#596510000000
1!
b11 %
1'
b11 +
#596520000000
0!
0'
#596530000000
1!
b100 %
1'
b100 +
#596540000000
0!
0'
#596550000000
1!
b101 %
1'
b101 +
#596560000000
0!
0'
#596570000000
1!
0$
b110 %
1'
0*
b110 +
#596580000000
0!
0'
#596590000000
1!
b111 %
1'
b111 +
#596600000000
0!
0'
#596610000000
1!
b1000 %
1'
b1000 +
#596620000000
1"
1(
#596630000000
0!
0"
b100 &
0'
0(
b100 ,
#596640000000
1!
b1001 %
1'
b1001 +
#596650000000
0!
0'
#596660000000
1!
b0 %
1'
b0 +
#596670000000
0!
0'
#596680000000
1!
1$
b1 %
1'
1*
b1 +
#596690000000
0!
0'
#596700000000
1!
b10 %
1'
b10 +
#596710000000
0!
0'
#596720000000
1!
b11 %
1'
b11 +
#596730000000
0!
0'
#596740000000
1!
b100 %
1'
b100 +
#596750000000
0!
0'
#596760000000
1!
b101 %
1'
b101 +
#596770000000
0!
0'
#596780000000
1!
b110 %
1'
b110 +
#596790000000
0!
0'
#596800000000
1!
b111 %
1'
b111 +
#596810000000
0!
0'
#596820000000
1!
0$
b1000 %
1'
0*
b1000 +
#596830000000
0!
0'
#596840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#596850000000
0!
0'
#596860000000
1!
b0 %
1'
b0 +
#596870000000
0!
0'
#596880000000
1!
1$
b1 %
1'
1*
b1 +
#596890000000
0!
0'
#596900000000
1!
b10 %
1'
b10 +
#596910000000
0!
0'
#596920000000
1!
b11 %
1'
b11 +
#596930000000
0!
0'
#596940000000
1!
b100 %
1'
b100 +
#596950000000
0!
0'
#596960000000
1!
b101 %
1'
b101 +
#596970000000
0!
0'
#596980000000
1!
0$
b110 %
1'
0*
b110 +
#596990000000
0!
0'
#597000000000
1!
b111 %
1'
b111 +
#597010000000
0!
0'
#597020000000
1!
b1000 %
1'
b1000 +
#597030000000
0!
0'
#597040000000
1!
b1001 %
1'
b1001 +
#597050000000
1"
1(
#597060000000
0!
0"
b100 &
0'
0(
b100 ,
#597070000000
1!
b0 %
1'
b0 +
#597080000000
0!
0'
#597090000000
1!
1$
b1 %
1'
1*
b1 +
#597100000000
0!
0'
#597110000000
1!
b10 %
1'
b10 +
#597120000000
0!
0'
#597130000000
1!
b11 %
1'
b11 +
#597140000000
0!
0'
#597150000000
1!
b100 %
1'
b100 +
#597160000000
0!
0'
#597170000000
1!
b101 %
1'
b101 +
#597180000000
0!
0'
#597190000000
1!
b110 %
1'
b110 +
#597200000000
0!
0'
#597210000000
1!
b111 %
1'
b111 +
#597220000000
0!
0'
#597230000000
1!
0$
b1000 %
1'
0*
b1000 +
#597240000000
0!
0'
#597250000000
1!
b1001 %
1'
b1001 +
#597260000000
0!
0'
#597270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#597280000000
0!
0'
#597290000000
1!
1$
b1 %
1'
1*
b1 +
#597300000000
0!
0'
#597310000000
1!
b10 %
1'
b10 +
#597320000000
0!
0'
#597330000000
1!
b11 %
1'
b11 +
#597340000000
0!
0'
#597350000000
1!
b100 %
1'
b100 +
#597360000000
0!
0'
#597370000000
1!
b101 %
1'
b101 +
#597380000000
0!
0'
#597390000000
1!
0$
b110 %
1'
0*
b110 +
#597400000000
0!
0'
#597410000000
1!
b111 %
1'
b111 +
#597420000000
0!
0'
#597430000000
1!
b1000 %
1'
b1000 +
#597440000000
0!
0'
#597450000000
1!
b1001 %
1'
b1001 +
#597460000000
0!
0'
#597470000000
1!
b0 %
1'
b0 +
#597480000000
1"
1(
#597490000000
0!
0"
b100 &
0'
0(
b100 ,
#597500000000
1!
1$
b1 %
1'
1*
b1 +
#597510000000
0!
0'
#597520000000
1!
b10 %
1'
b10 +
#597530000000
0!
0'
#597540000000
1!
b11 %
1'
b11 +
#597550000000
0!
0'
#597560000000
1!
b100 %
1'
b100 +
#597570000000
0!
0'
#597580000000
1!
b101 %
1'
b101 +
#597590000000
0!
0'
#597600000000
1!
b110 %
1'
b110 +
#597610000000
0!
0'
#597620000000
1!
b111 %
1'
b111 +
#597630000000
0!
0'
#597640000000
1!
0$
b1000 %
1'
0*
b1000 +
#597650000000
0!
0'
#597660000000
1!
b1001 %
1'
b1001 +
#597670000000
0!
0'
#597680000000
1!
b0 %
1'
b0 +
#597690000000
0!
0'
#597700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#597710000000
0!
0'
#597720000000
1!
b10 %
1'
b10 +
#597730000000
0!
0'
#597740000000
1!
b11 %
1'
b11 +
#597750000000
0!
0'
#597760000000
1!
b100 %
1'
b100 +
#597770000000
0!
0'
#597780000000
1!
b101 %
1'
b101 +
#597790000000
0!
0'
#597800000000
1!
0$
b110 %
1'
0*
b110 +
#597810000000
0!
0'
#597820000000
1!
b111 %
1'
b111 +
#597830000000
0!
0'
#597840000000
1!
b1000 %
1'
b1000 +
#597850000000
0!
0'
#597860000000
1!
b1001 %
1'
b1001 +
#597870000000
0!
0'
#597880000000
1!
b0 %
1'
b0 +
#597890000000
0!
0'
#597900000000
1!
1$
b1 %
1'
1*
b1 +
#597910000000
1"
1(
#597920000000
0!
0"
b100 &
0'
0(
b100 ,
#597930000000
1!
b10 %
1'
b10 +
#597940000000
0!
0'
#597950000000
1!
b11 %
1'
b11 +
#597960000000
0!
0'
#597970000000
1!
b100 %
1'
b100 +
#597980000000
0!
0'
#597990000000
1!
b101 %
1'
b101 +
#598000000000
0!
0'
#598010000000
1!
b110 %
1'
b110 +
#598020000000
0!
0'
#598030000000
1!
b111 %
1'
b111 +
#598040000000
0!
0'
#598050000000
1!
0$
b1000 %
1'
0*
b1000 +
#598060000000
0!
0'
#598070000000
1!
b1001 %
1'
b1001 +
#598080000000
0!
0'
#598090000000
1!
b0 %
1'
b0 +
#598100000000
0!
0'
#598110000000
1!
1$
b1 %
1'
1*
b1 +
#598120000000
0!
0'
#598130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#598140000000
0!
0'
#598150000000
1!
b11 %
1'
b11 +
#598160000000
0!
0'
#598170000000
1!
b100 %
1'
b100 +
#598180000000
0!
0'
#598190000000
1!
b101 %
1'
b101 +
#598200000000
0!
0'
#598210000000
1!
0$
b110 %
1'
0*
b110 +
#598220000000
0!
0'
#598230000000
1!
b111 %
1'
b111 +
#598240000000
0!
0'
#598250000000
1!
b1000 %
1'
b1000 +
#598260000000
0!
0'
#598270000000
1!
b1001 %
1'
b1001 +
#598280000000
0!
0'
#598290000000
1!
b0 %
1'
b0 +
#598300000000
0!
0'
#598310000000
1!
1$
b1 %
1'
1*
b1 +
#598320000000
0!
0'
#598330000000
1!
b10 %
1'
b10 +
#598340000000
1"
1(
#598350000000
0!
0"
b100 &
0'
0(
b100 ,
#598360000000
1!
b11 %
1'
b11 +
#598370000000
0!
0'
#598380000000
1!
b100 %
1'
b100 +
#598390000000
0!
0'
#598400000000
1!
b101 %
1'
b101 +
#598410000000
0!
0'
#598420000000
1!
b110 %
1'
b110 +
#598430000000
0!
0'
#598440000000
1!
b111 %
1'
b111 +
#598450000000
0!
0'
#598460000000
1!
0$
b1000 %
1'
0*
b1000 +
#598470000000
0!
0'
#598480000000
1!
b1001 %
1'
b1001 +
#598490000000
0!
0'
#598500000000
1!
b0 %
1'
b0 +
#598510000000
0!
0'
#598520000000
1!
1$
b1 %
1'
1*
b1 +
#598530000000
0!
0'
#598540000000
1!
b10 %
1'
b10 +
#598550000000
0!
0'
#598560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#598570000000
0!
0'
#598580000000
1!
b100 %
1'
b100 +
#598590000000
0!
0'
#598600000000
1!
b101 %
1'
b101 +
#598610000000
0!
0'
#598620000000
1!
0$
b110 %
1'
0*
b110 +
#598630000000
0!
0'
#598640000000
1!
b111 %
1'
b111 +
#598650000000
0!
0'
#598660000000
1!
b1000 %
1'
b1000 +
#598670000000
0!
0'
#598680000000
1!
b1001 %
1'
b1001 +
#598690000000
0!
0'
#598700000000
1!
b0 %
1'
b0 +
#598710000000
0!
0'
#598720000000
1!
1$
b1 %
1'
1*
b1 +
#598730000000
0!
0'
#598740000000
1!
b10 %
1'
b10 +
#598750000000
0!
0'
#598760000000
1!
b11 %
1'
b11 +
#598770000000
1"
1(
#598780000000
0!
0"
b100 &
0'
0(
b100 ,
#598790000000
1!
b100 %
1'
b100 +
#598800000000
0!
0'
#598810000000
1!
b101 %
1'
b101 +
#598820000000
0!
0'
#598830000000
1!
b110 %
1'
b110 +
#598840000000
0!
0'
#598850000000
1!
b111 %
1'
b111 +
#598860000000
0!
0'
#598870000000
1!
0$
b1000 %
1'
0*
b1000 +
#598880000000
0!
0'
#598890000000
1!
b1001 %
1'
b1001 +
#598900000000
0!
0'
#598910000000
1!
b0 %
1'
b0 +
#598920000000
0!
0'
#598930000000
1!
1$
b1 %
1'
1*
b1 +
#598940000000
0!
0'
#598950000000
1!
b10 %
1'
b10 +
#598960000000
0!
0'
#598970000000
1!
b11 %
1'
b11 +
#598980000000
0!
0'
#598990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#599000000000
0!
0'
#599010000000
1!
b101 %
1'
b101 +
#599020000000
0!
0'
#599030000000
1!
0$
b110 %
1'
0*
b110 +
#599040000000
0!
0'
#599050000000
1!
b111 %
1'
b111 +
#599060000000
0!
0'
#599070000000
1!
b1000 %
1'
b1000 +
#599080000000
0!
0'
#599090000000
1!
b1001 %
1'
b1001 +
#599100000000
0!
0'
#599110000000
1!
b0 %
1'
b0 +
#599120000000
0!
0'
#599130000000
1!
1$
b1 %
1'
1*
b1 +
#599140000000
0!
0'
#599150000000
1!
b10 %
1'
b10 +
#599160000000
0!
0'
#599170000000
1!
b11 %
1'
b11 +
#599180000000
0!
0'
#599190000000
1!
b100 %
1'
b100 +
#599200000000
1"
1(
#599210000000
0!
0"
b100 &
0'
0(
b100 ,
#599220000000
1!
b101 %
1'
b101 +
#599230000000
0!
0'
#599240000000
1!
b110 %
1'
b110 +
#599250000000
0!
0'
#599260000000
1!
b111 %
1'
b111 +
#599270000000
0!
0'
#599280000000
1!
0$
b1000 %
1'
0*
b1000 +
#599290000000
0!
0'
#599300000000
1!
b1001 %
1'
b1001 +
#599310000000
0!
0'
#599320000000
1!
b0 %
1'
b0 +
#599330000000
0!
0'
#599340000000
1!
1$
b1 %
1'
1*
b1 +
#599350000000
0!
0'
#599360000000
1!
b10 %
1'
b10 +
#599370000000
0!
0'
#599380000000
1!
b11 %
1'
b11 +
#599390000000
0!
0'
#599400000000
1!
b100 %
1'
b100 +
#599410000000
0!
0'
#599420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#599430000000
0!
0'
#599440000000
1!
0$
b110 %
1'
0*
b110 +
#599450000000
0!
0'
#599460000000
1!
b111 %
1'
b111 +
#599470000000
0!
0'
#599480000000
1!
b1000 %
1'
b1000 +
#599490000000
0!
0'
#599500000000
1!
b1001 %
1'
b1001 +
#599510000000
0!
0'
#599520000000
1!
b0 %
1'
b0 +
#599530000000
0!
0'
#599540000000
1!
1$
b1 %
1'
1*
b1 +
#599550000000
0!
0'
#599560000000
1!
b10 %
1'
b10 +
#599570000000
0!
0'
#599580000000
1!
b11 %
1'
b11 +
#599590000000
0!
0'
#599600000000
1!
b100 %
1'
b100 +
#599610000000
0!
0'
#599620000000
1!
b101 %
1'
b101 +
#599630000000
1"
1(
#599640000000
0!
0"
b100 &
0'
0(
b100 ,
#599650000000
1!
b110 %
1'
b110 +
#599660000000
0!
0'
#599670000000
1!
b111 %
1'
b111 +
#599680000000
0!
0'
#599690000000
1!
0$
b1000 %
1'
0*
b1000 +
#599700000000
0!
0'
#599710000000
1!
b1001 %
1'
b1001 +
#599720000000
0!
0'
#599730000000
1!
b0 %
1'
b0 +
#599740000000
0!
0'
#599750000000
1!
1$
b1 %
1'
1*
b1 +
#599760000000
0!
0'
#599770000000
1!
b10 %
1'
b10 +
#599780000000
0!
0'
#599790000000
1!
b11 %
1'
b11 +
#599800000000
0!
0'
#599810000000
1!
b100 %
1'
b100 +
#599820000000
0!
0'
#599830000000
1!
b101 %
1'
b101 +
#599840000000
0!
0'
#599850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#599860000000
0!
0'
#599870000000
1!
b111 %
1'
b111 +
#599880000000
0!
0'
#599890000000
1!
b1000 %
1'
b1000 +
#599900000000
0!
0'
#599910000000
1!
b1001 %
1'
b1001 +
#599920000000
0!
0'
#599930000000
1!
b0 %
1'
b0 +
#599940000000
0!
0'
#599950000000
1!
1$
b1 %
1'
1*
b1 +
#599960000000
0!
0'
#599970000000
1!
b10 %
1'
b10 +
#599980000000
0!
0'
#599990000000
1!
b11 %
1'
b11 +
#600000000000
0!
0'
#600010000000
1!
b100 %
1'
b100 +
#600020000000
0!
0'
#600030000000
1!
b101 %
1'
b101 +
#600040000000
0!
0'
#600050000000
1!
0$
b110 %
1'
0*
b110 +
#600060000000
1"
1(
#600070000000
0!
0"
b100 &
0'
0(
b100 ,
#600080000000
1!
1$
b111 %
1'
1*
b111 +
#600090000000
0!
0'
#600100000000
1!
0$
b1000 %
1'
0*
b1000 +
#600110000000
0!
0'
#600120000000
1!
b1001 %
1'
b1001 +
#600130000000
0!
0'
#600140000000
1!
b0 %
1'
b0 +
#600150000000
0!
0'
#600160000000
1!
1$
b1 %
1'
1*
b1 +
#600170000000
0!
0'
#600180000000
1!
b10 %
1'
b10 +
#600190000000
0!
0'
#600200000000
1!
b11 %
1'
b11 +
#600210000000
0!
0'
#600220000000
1!
b100 %
1'
b100 +
#600230000000
0!
0'
#600240000000
1!
b101 %
1'
b101 +
#600250000000
0!
0'
#600260000000
1!
b110 %
1'
b110 +
#600270000000
0!
0'
#600280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#600290000000
0!
0'
#600300000000
1!
b1000 %
1'
b1000 +
#600310000000
0!
0'
#600320000000
1!
b1001 %
1'
b1001 +
#600330000000
0!
0'
#600340000000
1!
b0 %
1'
b0 +
#600350000000
0!
0'
#600360000000
1!
1$
b1 %
1'
1*
b1 +
#600370000000
0!
0'
#600380000000
1!
b10 %
1'
b10 +
#600390000000
0!
0'
#600400000000
1!
b11 %
1'
b11 +
#600410000000
0!
0'
#600420000000
1!
b100 %
1'
b100 +
#600430000000
0!
0'
#600440000000
1!
b101 %
1'
b101 +
#600450000000
0!
0'
#600460000000
1!
0$
b110 %
1'
0*
b110 +
#600470000000
0!
0'
#600480000000
1!
b111 %
1'
b111 +
#600490000000
1"
1(
#600500000000
0!
0"
b100 &
0'
0(
b100 ,
#600510000000
1!
b1000 %
1'
b1000 +
#600520000000
0!
0'
#600530000000
1!
b1001 %
1'
b1001 +
#600540000000
0!
0'
#600550000000
1!
b0 %
1'
b0 +
#600560000000
0!
0'
#600570000000
1!
1$
b1 %
1'
1*
b1 +
#600580000000
0!
0'
#600590000000
1!
b10 %
1'
b10 +
#600600000000
0!
0'
#600610000000
1!
b11 %
1'
b11 +
#600620000000
0!
0'
#600630000000
1!
b100 %
1'
b100 +
#600640000000
0!
0'
#600650000000
1!
b101 %
1'
b101 +
#600660000000
0!
0'
#600670000000
1!
b110 %
1'
b110 +
#600680000000
0!
0'
#600690000000
1!
b111 %
1'
b111 +
#600700000000
0!
0'
#600710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#600720000000
0!
0'
#600730000000
1!
b1001 %
1'
b1001 +
#600740000000
0!
0'
#600750000000
1!
b0 %
1'
b0 +
#600760000000
0!
0'
#600770000000
1!
1$
b1 %
1'
1*
b1 +
#600780000000
0!
0'
#600790000000
1!
b10 %
1'
b10 +
#600800000000
0!
0'
#600810000000
1!
b11 %
1'
b11 +
#600820000000
0!
0'
#600830000000
1!
b100 %
1'
b100 +
#600840000000
0!
0'
#600850000000
1!
b101 %
1'
b101 +
#600860000000
0!
0'
#600870000000
1!
0$
b110 %
1'
0*
b110 +
#600880000000
0!
0'
#600890000000
1!
b111 %
1'
b111 +
#600900000000
0!
0'
#600910000000
1!
b1000 %
1'
b1000 +
#600920000000
1"
1(
#600930000000
0!
0"
b100 &
0'
0(
b100 ,
#600940000000
1!
b1001 %
1'
b1001 +
#600950000000
0!
0'
#600960000000
1!
b0 %
1'
b0 +
#600970000000
0!
0'
#600980000000
1!
1$
b1 %
1'
1*
b1 +
#600990000000
0!
0'
#601000000000
1!
b10 %
1'
b10 +
#601010000000
0!
0'
#601020000000
1!
b11 %
1'
b11 +
#601030000000
0!
0'
#601040000000
1!
b100 %
1'
b100 +
#601050000000
0!
0'
#601060000000
1!
b101 %
1'
b101 +
#601070000000
0!
0'
#601080000000
1!
b110 %
1'
b110 +
#601090000000
0!
0'
#601100000000
1!
b111 %
1'
b111 +
#601110000000
0!
0'
#601120000000
1!
0$
b1000 %
1'
0*
b1000 +
#601130000000
0!
0'
#601140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#601150000000
0!
0'
#601160000000
1!
b0 %
1'
b0 +
#601170000000
0!
0'
#601180000000
1!
1$
b1 %
1'
1*
b1 +
#601190000000
0!
0'
#601200000000
1!
b10 %
1'
b10 +
#601210000000
0!
0'
#601220000000
1!
b11 %
1'
b11 +
#601230000000
0!
0'
#601240000000
1!
b100 %
1'
b100 +
#601250000000
0!
0'
#601260000000
1!
b101 %
1'
b101 +
#601270000000
0!
0'
#601280000000
1!
0$
b110 %
1'
0*
b110 +
#601290000000
0!
0'
#601300000000
1!
b111 %
1'
b111 +
#601310000000
0!
0'
#601320000000
1!
b1000 %
1'
b1000 +
#601330000000
0!
0'
#601340000000
1!
b1001 %
1'
b1001 +
#601350000000
1"
1(
#601360000000
0!
0"
b100 &
0'
0(
b100 ,
#601370000000
1!
b0 %
1'
b0 +
#601380000000
0!
0'
#601390000000
1!
1$
b1 %
1'
1*
b1 +
#601400000000
0!
0'
#601410000000
1!
b10 %
1'
b10 +
#601420000000
0!
0'
#601430000000
1!
b11 %
1'
b11 +
#601440000000
0!
0'
#601450000000
1!
b100 %
1'
b100 +
#601460000000
0!
0'
#601470000000
1!
b101 %
1'
b101 +
#601480000000
0!
0'
#601490000000
1!
b110 %
1'
b110 +
#601500000000
0!
0'
#601510000000
1!
b111 %
1'
b111 +
#601520000000
0!
0'
#601530000000
1!
0$
b1000 %
1'
0*
b1000 +
#601540000000
0!
0'
#601550000000
1!
b1001 %
1'
b1001 +
#601560000000
0!
0'
#601570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#601580000000
0!
0'
#601590000000
1!
1$
b1 %
1'
1*
b1 +
#601600000000
0!
0'
#601610000000
1!
b10 %
1'
b10 +
#601620000000
0!
0'
#601630000000
1!
b11 %
1'
b11 +
#601640000000
0!
0'
#601650000000
1!
b100 %
1'
b100 +
#601660000000
0!
0'
#601670000000
1!
b101 %
1'
b101 +
#601680000000
0!
0'
#601690000000
1!
0$
b110 %
1'
0*
b110 +
#601700000000
0!
0'
#601710000000
1!
b111 %
1'
b111 +
#601720000000
0!
0'
#601730000000
1!
b1000 %
1'
b1000 +
#601740000000
0!
0'
#601750000000
1!
b1001 %
1'
b1001 +
#601760000000
0!
0'
#601770000000
1!
b0 %
1'
b0 +
#601780000000
1"
1(
#601790000000
0!
0"
b100 &
0'
0(
b100 ,
#601800000000
1!
1$
b1 %
1'
1*
b1 +
#601810000000
0!
0'
#601820000000
1!
b10 %
1'
b10 +
#601830000000
0!
0'
#601840000000
1!
b11 %
1'
b11 +
#601850000000
0!
0'
#601860000000
1!
b100 %
1'
b100 +
#601870000000
0!
0'
#601880000000
1!
b101 %
1'
b101 +
#601890000000
0!
0'
#601900000000
1!
b110 %
1'
b110 +
#601910000000
0!
0'
#601920000000
1!
b111 %
1'
b111 +
#601930000000
0!
0'
#601940000000
1!
0$
b1000 %
1'
0*
b1000 +
#601950000000
0!
0'
#601960000000
1!
b1001 %
1'
b1001 +
#601970000000
0!
0'
#601980000000
1!
b0 %
1'
b0 +
#601990000000
0!
0'
#602000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#602010000000
0!
0'
#602020000000
1!
b10 %
1'
b10 +
#602030000000
0!
0'
#602040000000
1!
b11 %
1'
b11 +
#602050000000
0!
0'
#602060000000
1!
b100 %
1'
b100 +
#602070000000
0!
0'
#602080000000
1!
b101 %
1'
b101 +
#602090000000
0!
0'
#602100000000
1!
0$
b110 %
1'
0*
b110 +
#602110000000
0!
0'
#602120000000
1!
b111 %
1'
b111 +
#602130000000
0!
0'
#602140000000
1!
b1000 %
1'
b1000 +
#602150000000
0!
0'
#602160000000
1!
b1001 %
1'
b1001 +
#602170000000
0!
0'
#602180000000
1!
b0 %
1'
b0 +
#602190000000
0!
0'
#602200000000
1!
1$
b1 %
1'
1*
b1 +
#602210000000
1"
1(
#602220000000
0!
0"
b100 &
0'
0(
b100 ,
#602230000000
1!
b10 %
1'
b10 +
#602240000000
0!
0'
#602250000000
1!
b11 %
1'
b11 +
#602260000000
0!
0'
#602270000000
1!
b100 %
1'
b100 +
#602280000000
0!
0'
#602290000000
1!
b101 %
1'
b101 +
#602300000000
0!
0'
#602310000000
1!
b110 %
1'
b110 +
#602320000000
0!
0'
#602330000000
1!
b111 %
1'
b111 +
#602340000000
0!
0'
#602350000000
1!
0$
b1000 %
1'
0*
b1000 +
#602360000000
0!
0'
#602370000000
1!
b1001 %
1'
b1001 +
#602380000000
0!
0'
#602390000000
1!
b0 %
1'
b0 +
#602400000000
0!
0'
#602410000000
1!
1$
b1 %
1'
1*
b1 +
#602420000000
0!
0'
#602430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#602440000000
0!
0'
#602450000000
1!
b11 %
1'
b11 +
#602460000000
0!
0'
#602470000000
1!
b100 %
1'
b100 +
#602480000000
0!
0'
#602490000000
1!
b101 %
1'
b101 +
#602500000000
0!
0'
#602510000000
1!
0$
b110 %
1'
0*
b110 +
#602520000000
0!
0'
#602530000000
1!
b111 %
1'
b111 +
#602540000000
0!
0'
#602550000000
1!
b1000 %
1'
b1000 +
#602560000000
0!
0'
#602570000000
1!
b1001 %
1'
b1001 +
#602580000000
0!
0'
#602590000000
1!
b0 %
1'
b0 +
#602600000000
0!
0'
#602610000000
1!
1$
b1 %
1'
1*
b1 +
#602620000000
0!
0'
#602630000000
1!
b10 %
1'
b10 +
#602640000000
1"
1(
#602650000000
0!
0"
b100 &
0'
0(
b100 ,
#602660000000
1!
b11 %
1'
b11 +
#602670000000
0!
0'
#602680000000
1!
b100 %
1'
b100 +
#602690000000
0!
0'
#602700000000
1!
b101 %
1'
b101 +
#602710000000
0!
0'
#602720000000
1!
b110 %
1'
b110 +
#602730000000
0!
0'
#602740000000
1!
b111 %
1'
b111 +
#602750000000
0!
0'
#602760000000
1!
0$
b1000 %
1'
0*
b1000 +
#602770000000
0!
0'
#602780000000
1!
b1001 %
1'
b1001 +
#602790000000
0!
0'
#602800000000
1!
b0 %
1'
b0 +
#602810000000
0!
0'
#602820000000
1!
1$
b1 %
1'
1*
b1 +
#602830000000
0!
0'
#602840000000
1!
b10 %
1'
b10 +
#602850000000
0!
0'
#602860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#602870000000
0!
0'
#602880000000
1!
b100 %
1'
b100 +
#602890000000
0!
0'
#602900000000
1!
b101 %
1'
b101 +
#602910000000
0!
0'
#602920000000
1!
0$
b110 %
1'
0*
b110 +
#602930000000
0!
0'
#602940000000
1!
b111 %
1'
b111 +
#602950000000
0!
0'
#602960000000
1!
b1000 %
1'
b1000 +
#602970000000
0!
0'
#602980000000
1!
b1001 %
1'
b1001 +
#602990000000
0!
0'
#603000000000
1!
b0 %
1'
b0 +
#603010000000
0!
0'
#603020000000
1!
1$
b1 %
1'
1*
b1 +
#603030000000
0!
0'
#603040000000
1!
b10 %
1'
b10 +
#603050000000
0!
0'
#603060000000
1!
b11 %
1'
b11 +
#603070000000
1"
1(
#603080000000
0!
0"
b100 &
0'
0(
b100 ,
#603090000000
1!
b100 %
1'
b100 +
#603100000000
0!
0'
#603110000000
1!
b101 %
1'
b101 +
#603120000000
0!
0'
#603130000000
1!
b110 %
1'
b110 +
#603140000000
0!
0'
#603150000000
1!
b111 %
1'
b111 +
#603160000000
0!
0'
#603170000000
1!
0$
b1000 %
1'
0*
b1000 +
#603180000000
0!
0'
#603190000000
1!
b1001 %
1'
b1001 +
#603200000000
0!
0'
#603210000000
1!
b0 %
1'
b0 +
#603220000000
0!
0'
#603230000000
1!
1$
b1 %
1'
1*
b1 +
#603240000000
0!
0'
#603250000000
1!
b10 %
1'
b10 +
#603260000000
0!
0'
#603270000000
1!
b11 %
1'
b11 +
#603280000000
0!
0'
#603290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#603300000000
0!
0'
#603310000000
1!
b101 %
1'
b101 +
#603320000000
0!
0'
#603330000000
1!
0$
b110 %
1'
0*
b110 +
#603340000000
0!
0'
#603350000000
1!
b111 %
1'
b111 +
#603360000000
0!
0'
#603370000000
1!
b1000 %
1'
b1000 +
#603380000000
0!
0'
#603390000000
1!
b1001 %
1'
b1001 +
#603400000000
0!
0'
#603410000000
1!
b0 %
1'
b0 +
#603420000000
0!
0'
#603430000000
1!
1$
b1 %
1'
1*
b1 +
#603440000000
0!
0'
#603450000000
1!
b10 %
1'
b10 +
#603460000000
0!
0'
#603470000000
1!
b11 %
1'
b11 +
#603480000000
0!
0'
#603490000000
1!
b100 %
1'
b100 +
#603500000000
1"
1(
#603510000000
0!
0"
b100 &
0'
0(
b100 ,
#603520000000
1!
b101 %
1'
b101 +
#603530000000
0!
0'
#603540000000
1!
b110 %
1'
b110 +
#603550000000
0!
0'
#603560000000
1!
b111 %
1'
b111 +
#603570000000
0!
0'
#603580000000
1!
0$
b1000 %
1'
0*
b1000 +
#603590000000
0!
0'
#603600000000
1!
b1001 %
1'
b1001 +
#603610000000
0!
0'
#603620000000
1!
b0 %
1'
b0 +
#603630000000
0!
0'
#603640000000
1!
1$
b1 %
1'
1*
b1 +
#603650000000
0!
0'
#603660000000
1!
b10 %
1'
b10 +
#603670000000
0!
0'
#603680000000
1!
b11 %
1'
b11 +
#603690000000
0!
0'
#603700000000
1!
b100 %
1'
b100 +
#603710000000
0!
0'
#603720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#603730000000
0!
0'
#603740000000
1!
0$
b110 %
1'
0*
b110 +
#603750000000
0!
0'
#603760000000
1!
b111 %
1'
b111 +
#603770000000
0!
0'
#603780000000
1!
b1000 %
1'
b1000 +
#603790000000
0!
0'
#603800000000
1!
b1001 %
1'
b1001 +
#603810000000
0!
0'
#603820000000
1!
b0 %
1'
b0 +
#603830000000
0!
0'
#603840000000
1!
1$
b1 %
1'
1*
b1 +
#603850000000
0!
0'
#603860000000
1!
b10 %
1'
b10 +
#603870000000
0!
0'
#603880000000
1!
b11 %
1'
b11 +
#603890000000
0!
0'
#603900000000
1!
b100 %
1'
b100 +
#603910000000
0!
0'
#603920000000
1!
b101 %
1'
b101 +
#603930000000
1"
1(
#603940000000
0!
0"
b100 &
0'
0(
b100 ,
#603950000000
1!
b110 %
1'
b110 +
#603960000000
0!
0'
#603970000000
1!
b111 %
1'
b111 +
#603980000000
0!
0'
#603990000000
1!
0$
b1000 %
1'
0*
b1000 +
#604000000000
0!
0'
#604010000000
1!
b1001 %
1'
b1001 +
#604020000000
0!
0'
#604030000000
1!
b0 %
1'
b0 +
#604040000000
0!
0'
#604050000000
1!
1$
b1 %
1'
1*
b1 +
#604060000000
0!
0'
#604070000000
1!
b10 %
1'
b10 +
#604080000000
0!
0'
#604090000000
1!
b11 %
1'
b11 +
#604100000000
0!
0'
#604110000000
1!
b100 %
1'
b100 +
#604120000000
0!
0'
#604130000000
1!
b101 %
1'
b101 +
#604140000000
0!
0'
#604150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#604160000000
0!
0'
#604170000000
1!
b111 %
1'
b111 +
#604180000000
0!
0'
#604190000000
1!
b1000 %
1'
b1000 +
#604200000000
0!
0'
#604210000000
1!
b1001 %
1'
b1001 +
#604220000000
0!
0'
#604230000000
1!
b0 %
1'
b0 +
#604240000000
0!
0'
#604250000000
1!
1$
b1 %
1'
1*
b1 +
#604260000000
0!
0'
#604270000000
1!
b10 %
1'
b10 +
#604280000000
0!
0'
#604290000000
1!
b11 %
1'
b11 +
#604300000000
0!
0'
#604310000000
1!
b100 %
1'
b100 +
#604320000000
0!
0'
#604330000000
1!
b101 %
1'
b101 +
#604340000000
0!
0'
#604350000000
1!
0$
b110 %
1'
0*
b110 +
#604360000000
1"
1(
#604370000000
0!
0"
b100 &
0'
0(
b100 ,
#604380000000
1!
1$
b111 %
1'
1*
b111 +
#604390000000
0!
0'
#604400000000
1!
0$
b1000 %
1'
0*
b1000 +
#604410000000
0!
0'
#604420000000
1!
b1001 %
1'
b1001 +
#604430000000
0!
0'
#604440000000
1!
b0 %
1'
b0 +
#604450000000
0!
0'
#604460000000
1!
1$
b1 %
1'
1*
b1 +
#604470000000
0!
0'
#604480000000
1!
b10 %
1'
b10 +
#604490000000
0!
0'
#604500000000
1!
b11 %
1'
b11 +
#604510000000
0!
0'
#604520000000
1!
b100 %
1'
b100 +
#604530000000
0!
0'
#604540000000
1!
b101 %
1'
b101 +
#604550000000
0!
0'
#604560000000
1!
b110 %
1'
b110 +
#604570000000
0!
0'
#604580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#604590000000
0!
0'
#604600000000
1!
b1000 %
1'
b1000 +
#604610000000
0!
0'
#604620000000
1!
b1001 %
1'
b1001 +
#604630000000
0!
0'
#604640000000
1!
b0 %
1'
b0 +
#604650000000
0!
0'
#604660000000
1!
1$
b1 %
1'
1*
b1 +
#604670000000
0!
0'
#604680000000
1!
b10 %
1'
b10 +
#604690000000
0!
0'
#604700000000
1!
b11 %
1'
b11 +
#604710000000
0!
0'
#604720000000
1!
b100 %
1'
b100 +
#604730000000
0!
0'
#604740000000
1!
b101 %
1'
b101 +
#604750000000
0!
0'
#604760000000
1!
0$
b110 %
1'
0*
b110 +
#604770000000
0!
0'
#604780000000
1!
b111 %
1'
b111 +
#604790000000
1"
1(
#604800000000
0!
0"
b100 &
0'
0(
b100 ,
#604810000000
1!
b1000 %
1'
b1000 +
#604820000000
0!
0'
#604830000000
1!
b1001 %
1'
b1001 +
#604840000000
0!
0'
#604850000000
1!
b0 %
1'
b0 +
#604860000000
0!
0'
#604870000000
1!
1$
b1 %
1'
1*
b1 +
#604880000000
0!
0'
#604890000000
1!
b10 %
1'
b10 +
#604900000000
0!
0'
#604910000000
1!
b11 %
1'
b11 +
#604920000000
0!
0'
#604930000000
1!
b100 %
1'
b100 +
#604940000000
0!
0'
#604950000000
1!
b101 %
1'
b101 +
#604960000000
0!
0'
#604970000000
1!
b110 %
1'
b110 +
#604980000000
0!
0'
#604990000000
1!
b111 %
1'
b111 +
#605000000000
0!
0'
#605010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#605020000000
0!
0'
#605030000000
1!
b1001 %
1'
b1001 +
#605040000000
0!
0'
#605050000000
1!
b0 %
1'
b0 +
#605060000000
0!
0'
#605070000000
1!
1$
b1 %
1'
1*
b1 +
#605080000000
0!
0'
#605090000000
1!
b10 %
1'
b10 +
#605100000000
0!
0'
#605110000000
1!
b11 %
1'
b11 +
#605120000000
0!
0'
#605130000000
1!
b100 %
1'
b100 +
#605140000000
0!
0'
#605150000000
1!
b101 %
1'
b101 +
#605160000000
0!
0'
#605170000000
1!
0$
b110 %
1'
0*
b110 +
#605180000000
0!
0'
#605190000000
1!
b111 %
1'
b111 +
#605200000000
0!
0'
#605210000000
1!
b1000 %
1'
b1000 +
#605220000000
1"
1(
#605230000000
0!
0"
b100 &
0'
0(
b100 ,
#605240000000
1!
b1001 %
1'
b1001 +
#605250000000
0!
0'
#605260000000
1!
b0 %
1'
b0 +
#605270000000
0!
0'
#605280000000
1!
1$
b1 %
1'
1*
b1 +
#605290000000
0!
0'
#605300000000
1!
b10 %
1'
b10 +
#605310000000
0!
0'
#605320000000
1!
b11 %
1'
b11 +
#605330000000
0!
0'
#605340000000
1!
b100 %
1'
b100 +
#605350000000
0!
0'
#605360000000
1!
b101 %
1'
b101 +
#605370000000
0!
0'
#605380000000
1!
b110 %
1'
b110 +
#605390000000
0!
0'
#605400000000
1!
b111 %
1'
b111 +
#605410000000
0!
0'
#605420000000
1!
0$
b1000 %
1'
0*
b1000 +
#605430000000
0!
0'
#605440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#605450000000
0!
0'
#605460000000
1!
b0 %
1'
b0 +
#605470000000
0!
0'
#605480000000
1!
1$
b1 %
1'
1*
b1 +
#605490000000
0!
0'
#605500000000
1!
b10 %
1'
b10 +
#605510000000
0!
0'
#605520000000
1!
b11 %
1'
b11 +
#605530000000
0!
0'
#605540000000
1!
b100 %
1'
b100 +
#605550000000
0!
0'
#605560000000
1!
b101 %
1'
b101 +
#605570000000
0!
0'
#605580000000
1!
0$
b110 %
1'
0*
b110 +
#605590000000
0!
0'
#605600000000
1!
b111 %
1'
b111 +
#605610000000
0!
0'
#605620000000
1!
b1000 %
1'
b1000 +
#605630000000
0!
0'
#605640000000
1!
b1001 %
1'
b1001 +
#605650000000
1"
1(
#605660000000
0!
0"
b100 &
0'
0(
b100 ,
#605670000000
1!
b0 %
1'
b0 +
#605680000000
0!
0'
#605690000000
1!
1$
b1 %
1'
1*
b1 +
#605700000000
0!
0'
#605710000000
1!
b10 %
1'
b10 +
#605720000000
0!
0'
#605730000000
1!
b11 %
1'
b11 +
#605740000000
0!
0'
#605750000000
1!
b100 %
1'
b100 +
#605760000000
0!
0'
#605770000000
1!
b101 %
1'
b101 +
#605780000000
0!
0'
#605790000000
1!
b110 %
1'
b110 +
#605800000000
0!
0'
#605810000000
1!
b111 %
1'
b111 +
#605820000000
0!
0'
#605830000000
1!
0$
b1000 %
1'
0*
b1000 +
#605840000000
0!
0'
#605850000000
1!
b1001 %
1'
b1001 +
#605860000000
0!
0'
#605870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#605880000000
0!
0'
#605890000000
1!
1$
b1 %
1'
1*
b1 +
#605900000000
0!
0'
#605910000000
1!
b10 %
1'
b10 +
#605920000000
0!
0'
#605930000000
1!
b11 %
1'
b11 +
#605940000000
0!
0'
#605950000000
1!
b100 %
1'
b100 +
#605960000000
0!
0'
#605970000000
1!
b101 %
1'
b101 +
#605980000000
0!
0'
#605990000000
1!
0$
b110 %
1'
0*
b110 +
#606000000000
0!
0'
#606010000000
1!
b111 %
1'
b111 +
#606020000000
0!
0'
#606030000000
1!
b1000 %
1'
b1000 +
#606040000000
0!
0'
#606050000000
1!
b1001 %
1'
b1001 +
#606060000000
0!
0'
#606070000000
1!
b0 %
1'
b0 +
#606080000000
1"
1(
#606090000000
0!
0"
b100 &
0'
0(
b100 ,
#606100000000
1!
1$
b1 %
1'
1*
b1 +
#606110000000
0!
0'
#606120000000
1!
b10 %
1'
b10 +
#606130000000
0!
0'
#606140000000
1!
b11 %
1'
b11 +
#606150000000
0!
0'
#606160000000
1!
b100 %
1'
b100 +
#606170000000
0!
0'
#606180000000
1!
b101 %
1'
b101 +
#606190000000
0!
0'
#606200000000
1!
b110 %
1'
b110 +
#606210000000
0!
0'
#606220000000
1!
b111 %
1'
b111 +
#606230000000
0!
0'
#606240000000
1!
0$
b1000 %
1'
0*
b1000 +
#606250000000
0!
0'
#606260000000
1!
b1001 %
1'
b1001 +
#606270000000
0!
0'
#606280000000
1!
b0 %
1'
b0 +
#606290000000
0!
0'
#606300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#606310000000
0!
0'
#606320000000
1!
b10 %
1'
b10 +
#606330000000
0!
0'
#606340000000
1!
b11 %
1'
b11 +
#606350000000
0!
0'
#606360000000
1!
b100 %
1'
b100 +
#606370000000
0!
0'
#606380000000
1!
b101 %
1'
b101 +
#606390000000
0!
0'
#606400000000
1!
0$
b110 %
1'
0*
b110 +
#606410000000
0!
0'
#606420000000
1!
b111 %
1'
b111 +
#606430000000
0!
0'
#606440000000
1!
b1000 %
1'
b1000 +
#606450000000
0!
0'
#606460000000
1!
b1001 %
1'
b1001 +
#606470000000
0!
0'
#606480000000
1!
b0 %
1'
b0 +
#606490000000
0!
0'
#606500000000
1!
1$
b1 %
1'
1*
b1 +
#606510000000
1"
1(
#606520000000
0!
0"
b100 &
0'
0(
b100 ,
#606530000000
1!
b10 %
1'
b10 +
#606540000000
0!
0'
#606550000000
1!
b11 %
1'
b11 +
#606560000000
0!
0'
#606570000000
1!
b100 %
1'
b100 +
#606580000000
0!
0'
#606590000000
1!
b101 %
1'
b101 +
#606600000000
0!
0'
#606610000000
1!
b110 %
1'
b110 +
#606620000000
0!
0'
#606630000000
1!
b111 %
1'
b111 +
#606640000000
0!
0'
#606650000000
1!
0$
b1000 %
1'
0*
b1000 +
#606660000000
0!
0'
#606670000000
1!
b1001 %
1'
b1001 +
#606680000000
0!
0'
#606690000000
1!
b0 %
1'
b0 +
#606700000000
0!
0'
#606710000000
1!
1$
b1 %
1'
1*
b1 +
#606720000000
0!
0'
#606730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#606740000000
0!
0'
#606750000000
1!
b11 %
1'
b11 +
#606760000000
0!
0'
#606770000000
1!
b100 %
1'
b100 +
#606780000000
0!
0'
#606790000000
1!
b101 %
1'
b101 +
#606800000000
0!
0'
#606810000000
1!
0$
b110 %
1'
0*
b110 +
#606820000000
0!
0'
#606830000000
1!
b111 %
1'
b111 +
#606840000000
0!
0'
#606850000000
1!
b1000 %
1'
b1000 +
#606860000000
0!
0'
#606870000000
1!
b1001 %
1'
b1001 +
#606880000000
0!
0'
#606890000000
1!
b0 %
1'
b0 +
#606900000000
0!
0'
#606910000000
1!
1$
b1 %
1'
1*
b1 +
#606920000000
0!
0'
#606930000000
1!
b10 %
1'
b10 +
#606940000000
1"
1(
#606950000000
0!
0"
b100 &
0'
0(
b100 ,
#606960000000
1!
b11 %
1'
b11 +
#606970000000
0!
0'
#606980000000
1!
b100 %
1'
b100 +
#606990000000
0!
0'
#607000000000
1!
b101 %
1'
b101 +
#607010000000
0!
0'
#607020000000
1!
b110 %
1'
b110 +
#607030000000
0!
0'
#607040000000
1!
b111 %
1'
b111 +
#607050000000
0!
0'
#607060000000
1!
0$
b1000 %
1'
0*
b1000 +
#607070000000
0!
0'
#607080000000
1!
b1001 %
1'
b1001 +
#607090000000
0!
0'
#607100000000
1!
b0 %
1'
b0 +
#607110000000
0!
0'
#607120000000
1!
1$
b1 %
1'
1*
b1 +
#607130000000
0!
0'
#607140000000
1!
b10 %
1'
b10 +
#607150000000
0!
0'
#607160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#607170000000
0!
0'
#607180000000
1!
b100 %
1'
b100 +
#607190000000
0!
0'
#607200000000
1!
b101 %
1'
b101 +
#607210000000
0!
0'
#607220000000
1!
0$
b110 %
1'
0*
b110 +
#607230000000
0!
0'
#607240000000
1!
b111 %
1'
b111 +
#607250000000
0!
0'
#607260000000
1!
b1000 %
1'
b1000 +
#607270000000
0!
0'
#607280000000
1!
b1001 %
1'
b1001 +
#607290000000
0!
0'
#607300000000
1!
b0 %
1'
b0 +
#607310000000
0!
0'
#607320000000
1!
1$
b1 %
1'
1*
b1 +
#607330000000
0!
0'
#607340000000
1!
b10 %
1'
b10 +
#607350000000
0!
0'
#607360000000
1!
b11 %
1'
b11 +
#607370000000
1"
1(
#607380000000
0!
0"
b100 &
0'
0(
b100 ,
#607390000000
1!
b100 %
1'
b100 +
#607400000000
0!
0'
#607410000000
1!
b101 %
1'
b101 +
#607420000000
0!
0'
#607430000000
1!
b110 %
1'
b110 +
#607440000000
0!
0'
#607450000000
1!
b111 %
1'
b111 +
#607460000000
0!
0'
#607470000000
1!
0$
b1000 %
1'
0*
b1000 +
#607480000000
0!
0'
#607490000000
1!
b1001 %
1'
b1001 +
#607500000000
0!
0'
#607510000000
1!
b0 %
1'
b0 +
#607520000000
0!
0'
#607530000000
1!
1$
b1 %
1'
1*
b1 +
#607540000000
0!
0'
#607550000000
1!
b10 %
1'
b10 +
#607560000000
0!
0'
#607570000000
1!
b11 %
1'
b11 +
#607580000000
0!
0'
#607590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#607600000000
0!
0'
#607610000000
1!
b101 %
1'
b101 +
#607620000000
0!
0'
#607630000000
1!
0$
b110 %
1'
0*
b110 +
#607640000000
0!
0'
#607650000000
1!
b111 %
1'
b111 +
#607660000000
0!
0'
#607670000000
1!
b1000 %
1'
b1000 +
#607680000000
0!
0'
#607690000000
1!
b1001 %
1'
b1001 +
#607700000000
0!
0'
#607710000000
1!
b0 %
1'
b0 +
#607720000000
0!
0'
#607730000000
1!
1$
b1 %
1'
1*
b1 +
#607740000000
0!
0'
#607750000000
1!
b10 %
1'
b10 +
#607760000000
0!
0'
#607770000000
1!
b11 %
1'
b11 +
#607780000000
0!
0'
#607790000000
1!
b100 %
1'
b100 +
#607800000000
1"
1(
#607810000000
0!
0"
b100 &
0'
0(
b100 ,
#607820000000
1!
b101 %
1'
b101 +
#607830000000
0!
0'
#607840000000
1!
b110 %
1'
b110 +
#607850000000
0!
0'
#607860000000
1!
b111 %
1'
b111 +
#607870000000
0!
0'
#607880000000
1!
0$
b1000 %
1'
0*
b1000 +
#607890000000
0!
0'
#607900000000
1!
b1001 %
1'
b1001 +
#607910000000
0!
0'
#607920000000
1!
b0 %
1'
b0 +
#607930000000
0!
0'
#607940000000
1!
1$
b1 %
1'
1*
b1 +
#607950000000
0!
0'
#607960000000
1!
b10 %
1'
b10 +
#607970000000
0!
0'
#607980000000
1!
b11 %
1'
b11 +
#607990000000
0!
0'
#608000000000
1!
b100 %
1'
b100 +
#608010000000
0!
0'
#608020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#608030000000
0!
0'
#608040000000
1!
0$
b110 %
1'
0*
b110 +
#608050000000
0!
0'
#608060000000
1!
b111 %
1'
b111 +
#608070000000
0!
0'
#608080000000
1!
b1000 %
1'
b1000 +
#608090000000
0!
0'
#608100000000
1!
b1001 %
1'
b1001 +
#608110000000
0!
0'
#608120000000
1!
b0 %
1'
b0 +
#608130000000
0!
0'
#608140000000
1!
1$
b1 %
1'
1*
b1 +
#608150000000
0!
0'
#608160000000
1!
b10 %
1'
b10 +
#608170000000
0!
0'
#608180000000
1!
b11 %
1'
b11 +
#608190000000
0!
0'
#608200000000
1!
b100 %
1'
b100 +
#608210000000
0!
0'
#608220000000
1!
b101 %
1'
b101 +
#608230000000
1"
1(
#608240000000
0!
0"
b100 &
0'
0(
b100 ,
#608250000000
1!
b110 %
1'
b110 +
#608260000000
0!
0'
#608270000000
1!
b111 %
1'
b111 +
#608280000000
0!
0'
#608290000000
1!
0$
b1000 %
1'
0*
b1000 +
#608300000000
0!
0'
#608310000000
1!
b1001 %
1'
b1001 +
#608320000000
0!
0'
#608330000000
1!
b0 %
1'
b0 +
#608340000000
0!
0'
#608350000000
1!
1$
b1 %
1'
1*
b1 +
#608360000000
0!
0'
#608370000000
1!
b10 %
1'
b10 +
#608380000000
0!
0'
#608390000000
1!
b11 %
1'
b11 +
#608400000000
0!
0'
#608410000000
1!
b100 %
1'
b100 +
#608420000000
0!
0'
#608430000000
1!
b101 %
1'
b101 +
#608440000000
0!
0'
#608450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#608460000000
0!
0'
#608470000000
1!
b111 %
1'
b111 +
#608480000000
0!
0'
#608490000000
1!
b1000 %
1'
b1000 +
#608500000000
0!
0'
#608510000000
1!
b1001 %
1'
b1001 +
#608520000000
0!
0'
#608530000000
1!
b0 %
1'
b0 +
#608540000000
0!
0'
#608550000000
1!
1$
b1 %
1'
1*
b1 +
#608560000000
0!
0'
#608570000000
1!
b10 %
1'
b10 +
#608580000000
0!
0'
#608590000000
1!
b11 %
1'
b11 +
#608600000000
0!
0'
#608610000000
1!
b100 %
1'
b100 +
#608620000000
0!
0'
#608630000000
1!
b101 %
1'
b101 +
#608640000000
0!
0'
#608650000000
1!
0$
b110 %
1'
0*
b110 +
#608660000000
1"
1(
#608670000000
0!
0"
b100 &
0'
0(
b100 ,
#608680000000
1!
1$
b111 %
1'
1*
b111 +
#608690000000
0!
0'
#608700000000
1!
0$
b1000 %
1'
0*
b1000 +
#608710000000
0!
0'
#608720000000
1!
b1001 %
1'
b1001 +
#608730000000
0!
0'
#608740000000
1!
b0 %
1'
b0 +
#608750000000
0!
0'
#608760000000
1!
1$
b1 %
1'
1*
b1 +
#608770000000
0!
0'
#608780000000
1!
b10 %
1'
b10 +
#608790000000
0!
0'
#608800000000
1!
b11 %
1'
b11 +
#608810000000
0!
0'
#608820000000
1!
b100 %
1'
b100 +
#608830000000
0!
0'
#608840000000
1!
b101 %
1'
b101 +
#608850000000
0!
0'
#608860000000
1!
b110 %
1'
b110 +
#608870000000
0!
0'
#608880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#608890000000
0!
0'
#608900000000
1!
b1000 %
1'
b1000 +
#608910000000
0!
0'
#608920000000
1!
b1001 %
1'
b1001 +
#608930000000
0!
0'
#608940000000
1!
b0 %
1'
b0 +
#608950000000
0!
0'
#608960000000
1!
1$
b1 %
1'
1*
b1 +
#608970000000
0!
0'
#608980000000
1!
b10 %
1'
b10 +
#608990000000
0!
0'
#609000000000
1!
b11 %
1'
b11 +
#609010000000
0!
0'
#609020000000
1!
b100 %
1'
b100 +
#609030000000
0!
0'
#609040000000
1!
b101 %
1'
b101 +
#609050000000
0!
0'
#609060000000
1!
0$
b110 %
1'
0*
b110 +
#609070000000
0!
0'
#609080000000
1!
b111 %
1'
b111 +
#609090000000
1"
1(
#609100000000
0!
0"
b100 &
0'
0(
b100 ,
#609110000000
1!
b1000 %
1'
b1000 +
#609120000000
0!
0'
#609130000000
1!
b1001 %
1'
b1001 +
#609140000000
0!
0'
#609150000000
1!
b0 %
1'
b0 +
#609160000000
0!
0'
#609170000000
1!
1$
b1 %
1'
1*
b1 +
#609180000000
0!
0'
#609190000000
1!
b10 %
1'
b10 +
#609200000000
0!
0'
#609210000000
1!
b11 %
1'
b11 +
#609220000000
0!
0'
#609230000000
1!
b100 %
1'
b100 +
#609240000000
0!
0'
#609250000000
1!
b101 %
1'
b101 +
#609260000000
0!
0'
#609270000000
1!
b110 %
1'
b110 +
#609280000000
0!
0'
#609290000000
1!
b111 %
1'
b111 +
#609300000000
0!
0'
#609310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#609320000000
0!
0'
#609330000000
1!
b1001 %
1'
b1001 +
#609340000000
0!
0'
#609350000000
1!
b0 %
1'
b0 +
#609360000000
0!
0'
#609370000000
1!
1$
b1 %
1'
1*
b1 +
#609380000000
0!
0'
#609390000000
1!
b10 %
1'
b10 +
#609400000000
0!
0'
#609410000000
1!
b11 %
1'
b11 +
#609420000000
0!
0'
#609430000000
1!
b100 %
1'
b100 +
#609440000000
0!
0'
#609450000000
1!
b101 %
1'
b101 +
#609460000000
0!
0'
#609470000000
1!
0$
b110 %
1'
0*
b110 +
#609480000000
0!
0'
#609490000000
1!
b111 %
1'
b111 +
#609500000000
0!
0'
#609510000000
1!
b1000 %
1'
b1000 +
#609520000000
1"
1(
#609530000000
0!
0"
b100 &
0'
0(
b100 ,
#609540000000
1!
b1001 %
1'
b1001 +
#609550000000
0!
0'
#609560000000
1!
b0 %
1'
b0 +
#609570000000
0!
0'
#609580000000
1!
1$
b1 %
1'
1*
b1 +
#609590000000
0!
0'
#609600000000
1!
b10 %
1'
b10 +
#609610000000
0!
0'
#609620000000
1!
b11 %
1'
b11 +
#609630000000
0!
0'
#609640000000
1!
b100 %
1'
b100 +
#609650000000
0!
0'
#609660000000
1!
b101 %
1'
b101 +
#609670000000
0!
0'
#609680000000
1!
b110 %
1'
b110 +
#609690000000
0!
0'
#609700000000
1!
b111 %
1'
b111 +
#609710000000
0!
0'
#609720000000
1!
0$
b1000 %
1'
0*
b1000 +
#609730000000
0!
0'
#609740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#609750000000
0!
0'
#609760000000
1!
b0 %
1'
b0 +
#609770000000
0!
0'
#609780000000
1!
1$
b1 %
1'
1*
b1 +
#609790000000
0!
0'
#609800000000
1!
b10 %
1'
b10 +
#609810000000
0!
0'
#609820000000
1!
b11 %
1'
b11 +
#609830000000
0!
0'
#609840000000
1!
b100 %
1'
b100 +
#609850000000
0!
0'
#609860000000
1!
b101 %
1'
b101 +
#609870000000
0!
0'
#609880000000
1!
0$
b110 %
1'
0*
b110 +
#609890000000
0!
0'
#609900000000
1!
b111 %
1'
b111 +
#609910000000
0!
0'
#609920000000
1!
b1000 %
1'
b1000 +
#609930000000
0!
0'
#609940000000
1!
b1001 %
1'
b1001 +
#609950000000
1"
1(
#609960000000
0!
0"
b100 &
0'
0(
b100 ,
#609970000000
1!
b0 %
1'
b0 +
#609980000000
0!
0'
#609990000000
1!
1$
b1 %
1'
1*
b1 +
#610000000000
0!
0'
#610010000000
1!
b10 %
1'
b10 +
#610020000000
0!
0'
#610030000000
1!
b11 %
1'
b11 +
#610040000000
0!
0'
#610050000000
1!
b100 %
1'
b100 +
#610060000000
0!
0'
#610070000000
1!
b101 %
1'
b101 +
#610080000000
0!
0'
#610090000000
1!
b110 %
1'
b110 +
#610100000000
0!
0'
#610110000000
1!
b111 %
1'
b111 +
#610120000000
0!
0'
#610130000000
1!
0$
b1000 %
1'
0*
b1000 +
#610140000000
0!
0'
#610150000000
1!
b1001 %
1'
b1001 +
#610160000000
0!
0'
#610170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#610180000000
0!
0'
#610190000000
1!
1$
b1 %
1'
1*
b1 +
#610200000000
0!
0'
#610210000000
1!
b10 %
1'
b10 +
#610220000000
0!
0'
#610230000000
1!
b11 %
1'
b11 +
#610240000000
0!
0'
#610250000000
1!
b100 %
1'
b100 +
#610260000000
0!
0'
#610270000000
1!
b101 %
1'
b101 +
#610280000000
0!
0'
#610290000000
1!
0$
b110 %
1'
0*
b110 +
#610300000000
0!
0'
#610310000000
1!
b111 %
1'
b111 +
#610320000000
0!
0'
#610330000000
1!
b1000 %
1'
b1000 +
#610340000000
0!
0'
#610350000000
1!
b1001 %
1'
b1001 +
#610360000000
0!
0'
#610370000000
1!
b0 %
1'
b0 +
#610380000000
1"
1(
#610390000000
0!
0"
b100 &
0'
0(
b100 ,
#610400000000
1!
1$
b1 %
1'
1*
b1 +
#610410000000
0!
0'
#610420000000
1!
b10 %
1'
b10 +
#610430000000
0!
0'
#610440000000
1!
b11 %
1'
b11 +
#610450000000
0!
0'
#610460000000
1!
b100 %
1'
b100 +
#610470000000
0!
0'
#610480000000
1!
b101 %
1'
b101 +
#610490000000
0!
0'
#610500000000
1!
b110 %
1'
b110 +
#610510000000
0!
0'
#610520000000
1!
b111 %
1'
b111 +
#610530000000
0!
0'
#610540000000
1!
0$
b1000 %
1'
0*
b1000 +
#610550000000
0!
0'
#610560000000
1!
b1001 %
1'
b1001 +
#610570000000
0!
0'
#610580000000
1!
b0 %
1'
b0 +
#610590000000
0!
0'
#610600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#610610000000
0!
0'
#610620000000
1!
b10 %
1'
b10 +
#610630000000
0!
0'
#610640000000
1!
b11 %
1'
b11 +
#610650000000
0!
0'
#610660000000
1!
b100 %
1'
b100 +
#610670000000
0!
0'
#610680000000
1!
b101 %
1'
b101 +
#610690000000
0!
0'
#610700000000
1!
0$
b110 %
1'
0*
b110 +
#610710000000
0!
0'
#610720000000
1!
b111 %
1'
b111 +
#610730000000
0!
0'
#610740000000
1!
b1000 %
1'
b1000 +
#610750000000
0!
0'
#610760000000
1!
b1001 %
1'
b1001 +
#610770000000
0!
0'
#610780000000
1!
b0 %
1'
b0 +
#610790000000
0!
0'
#610800000000
1!
1$
b1 %
1'
1*
b1 +
#610810000000
1"
1(
#610820000000
0!
0"
b100 &
0'
0(
b100 ,
#610830000000
1!
b10 %
1'
b10 +
#610840000000
0!
0'
#610850000000
1!
b11 %
1'
b11 +
#610860000000
0!
0'
#610870000000
1!
b100 %
1'
b100 +
#610880000000
0!
0'
#610890000000
1!
b101 %
1'
b101 +
#610900000000
0!
0'
#610910000000
1!
b110 %
1'
b110 +
#610920000000
0!
0'
#610930000000
1!
b111 %
1'
b111 +
#610940000000
0!
0'
#610950000000
1!
0$
b1000 %
1'
0*
b1000 +
#610960000000
0!
0'
#610970000000
1!
b1001 %
1'
b1001 +
#610980000000
0!
0'
#610990000000
1!
b0 %
1'
b0 +
#611000000000
0!
0'
#611010000000
1!
1$
b1 %
1'
1*
b1 +
#611020000000
0!
0'
#611030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#611040000000
0!
0'
#611050000000
1!
b11 %
1'
b11 +
#611060000000
0!
0'
#611070000000
1!
b100 %
1'
b100 +
#611080000000
0!
0'
#611090000000
1!
b101 %
1'
b101 +
#611100000000
0!
0'
#611110000000
1!
0$
b110 %
1'
0*
b110 +
#611120000000
0!
0'
#611130000000
1!
b111 %
1'
b111 +
#611140000000
0!
0'
#611150000000
1!
b1000 %
1'
b1000 +
#611160000000
0!
0'
#611170000000
1!
b1001 %
1'
b1001 +
#611180000000
0!
0'
#611190000000
1!
b0 %
1'
b0 +
#611200000000
0!
0'
#611210000000
1!
1$
b1 %
1'
1*
b1 +
#611220000000
0!
0'
#611230000000
1!
b10 %
1'
b10 +
#611240000000
1"
1(
#611250000000
0!
0"
b100 &
0'
0(
b100 ,
#611260000000
1!
b11 %
1'
b11 +
#611270000000
0!
0'
#611280000000
1!
b100 %
1'
b100 +
#611290000000
0!
0'
#611300000000
1!
b101 %
1'
b101 +
#611310000000
0!
0'
#611320000000
1!
b110 %
1'
b110 +
#611330000000
0!
0'
#611340000000
1!
b111 %
1'
b111 +
#611350000000
0!
0'
#611360000000
1!
0$
b1000 %
1'
0*
b1000 +
#611370000000
0!
0'
#611380000000
1!
b1001 %
1'
b1001 +
#611390000000
0!
0'
#611400000000
1!
b0 %
1'
b0 +
#611410000000
0!
0'
#611420000000
1!
1$
b1 %
1'
1*
b1 +
#611430000000
0!
0'
#611440000000
1!
b10 %
1'
b10 +
#611450000000
0!
0'
#611460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#611470000000
0!
0'
#611480000000
1!
b100 %
1'
b100 +
#611490000000
0!
0'
#611500000000
1!
b101 %
1'
b101 +
#611510000000
0!
0'
#611520000000
1!
0$
b110 %
1'
0*
b110 +
#611530000000
0!
0'
#611540000000
1!
b111 %
1'
b111 +
#611550000000
0!
0'
#611560000000
1!
b1000 %
1'
b1000 +
#611570000000
0!
0'
#611580000000
1!
b1001 %
1'
b1001 +
#611590000000
0!
0'
#611600000000
1!
b0 %
1'
b0 +
#611610000000
0!
0'
#611620000000
1!
1$
b1 %
1'
1*
b1 +
#611630000000
0!
0'
#611640000000
1!
b10 %
1'
b10 +
#611650000000
0!
0'
#611660000000
1!
b11 %
1'
b11 +
#611670000000
1"
1(
#611680000000
0!
0"
b100 &
0'
0(
b100 ,
#611690000000
1!
b100 %
1'
b100 +
#611700000000
0!
0'
#611710000000
1!
b101 %
1'
b101 +
#611720000000
0!
0'
#611730000000
1!
b110 %
1'
b110 +
#611740000000
0!
0'
#611750000000
1!
b111 %
1'
b111 +
#611760000000
0!
0'
#611770000000
1!
0$
b1000 %
1'
0*
b1000 +
#611780000000
0!
0'
#611790000000
1!
b1001 %
1'
b1001 +
#611800000000
0!
0'
#611810000000
1!
b0 %
1'
b0 +
#611820000000
0!
0'
#611830000000
1!
1$
b1 %
1'
1*
b1 +
#611840000000
0!
0'
#611850000000
1!
b10 %
1'
b10 +
#611860000000
0!
0'
#611870000000
1!
b11 %
1'
b11 +
#611880000000
0!
0'
#611890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#611900000000
0!
0'
#611910000000
1!
b101 %
1'
b101 +
#611920000000
0!
0'
#611930000000
1!
0$
b110 %
1'
0*
b110 +
#611940000000
0!
0'
#611950000000
1!
b111 %
1'
b111 +
#611960000000
0!
0'
#611970000000
1!
b1000 %
1'
b1000 +
#611980000000
0!
0'
#611990000000
1!
b1001 %
1'
b1001 +
#612000000000
0!
0'
#612010000000
1!
b0 %
1'
b0 +
#612020000000
0!
0'
#612030000000
1!
1$
b1 %
1'
1*
b1 +
#612040000000
0!
0'
#612050000000
1!
b10 %
1'
b10 +
#612060000000
0!
0'
#612070000000
1!
b11 %
1'
b11 +
#612080000000
0!
0'
#612090000000
1!
b100 %
1'
b100 +
#612100000000
1"
1(
#612110000000
0!
0"
b100 &
0'
0(
b100 ,
#612120000000
1!
b101 %
1'
b101 +
#612130000000
0!
0'
#612140000000
1!
b110 %
1'
b110 +
#612150000000
0!
0'
#612160000000
1!
b111 %
1'
b111 +
#612170000000
0!
0'
#612180000000
1!
0$
b1000 %
1'
0*
b1000 +
#612190000000
0!
0'
#612200000000
1!
b1001 %
1'
b1001 +
#612210000000
0!
0'
#612220000000
1!
b0 %
1'
b0 +
#612230000000
0!
0'
#612240000000
1!
1$
b1 %
1'
1*
b1 +
#612250000000
0!
0'
#612260000000
1!
b10 %
1'
b10 +
#612270000000
0!
0'
#612280000000
1!
b11 %
1'
b11 +
#612290000000
0!
0'
#612300000000
1!
b100 %
1'
b100 +
#612310000000
0!
0'
#612320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#612330000000
0!
0'
#612340000000
1!
0$
b110 %
1'
0*
b110 +
#612350000000
0!
0'
#612360000000
1!
b111 %
1'
b111 +
#612370000000
0!
0'
#612380000000
1!
b1000 %
1'
b1000 +
#612390000000
0!
0'
#612400000000
1!
b1001 %
1'
b1001 +
#612410000000
0!
0'
#612420000000
1!
b0 %
1'
b0 +
#612430000000
0!
0'
#612440000000
1!
1$
b1 %
1'
1*
b1 +
#612450000000
0!
0'
#612460000000
1!
b10 %
1'
b10 +
#612470000000
0!
0'
#612480000000
1!
b11 %
1'
b11 +
#612490000000
0!
0'
#612500000000
1!
b100 %
1'
b100 +
#612510000000
0!
0'
#612520000000
1!
b101 %
1'
b101 +
#612530000000
1"
1(
#612540000000
0!
0"
b100 &
0'
0(
b100 ,
#612550000000
1!
b110 %
1'
b110 +
#612560000000
0!
0'
#612570000000
1!
b111 %
1'
b111 +
#612580000000
0!
0'
#612590000000
1!
0$
b1000 %
1'
0*
b1000 +
#612600000000
0!
0'
#612610000000
1!
b1001 %
1'
b1001 +
#612620000000
0!
0'
#612630000000
1!
b0 %
1'
b0 +
#612640000000
0!
0'
#612650000000
1!
1$
b1 %
1'
1*
b1 +
#612660000000
0!
0'
#612670000000
1!
b10 %
1'
b10 +
#612680000000
0!
0'
#612690000000
1!
b11 %
1'
b11 +
#612700000000
0!
0'
#612710000000
1!
b100 %
1'
b100 +
#612720000000
0!
0'
#612730000000
1!
b101 %
1'
b101 +
#612740000000
0!
0'
#612750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#612760000000
0!
0'
#612770000000
1!
b111 %
1'
b111 +
#612780000000
0!
0'
#612790000000
1!
b1000 %
1'
b1000 +
#612800000000
0!
0'
#612810000000
1!
b1001 %
1'
b1001 +
#612820000000
0!
0'
#612830000000
1!
b0 %
1'
b0 +
#612840000000
0!
0'
#612850000000
1!
1$
b1 %
1'
1*
b1 +
#612860000000
0!
0'
#612870000000
1!
b10 %
1'
b10 +
#612880000000
0!
0'
#612890000000
1!
b11 %
1'
b11 +
#612900000000
0!
0'
#612910000000
1!
b100 %
1'
b100 +
#612920000000
0!
0'
#612930000000
1!
b101 %
1'
b101 +
#612940000000
0!
0'
#612950000000
1!
0$
b110 %
1'
0*
b110 +
#612960000000
1"
1(
#612970000000
0!
0"
b100 &
0'
0(
b100 ,
#612980000000
1!
1$
b111 %
1'
1*
b111 +
#612990000000
0!
0'
#613000000000
1!
0$
b1000 %
1'
0*
b1000 +
#613010000000
0!
0'
#613020000000
1!
b1001 %
1'
b1001 +
#613030000000
0!
0'
#613040000000
1!
b0 %
1'
b0 +
#613050000000
0!
0'
#613060000000
1!
1$
b1 %
1'
1*
b1 +
#613070000000
0!
0'
#613080000000
1!
b10 %
1'
b10 +
#613090000000
0!
0'
#613100000000
1!
b11 %
1'
b11 +
#613110000000
0!
0'
#613120000000
1!
b100 %
1'
b100 +
#613130000000
0!
0'
#613140000000
1!
b101 %
1'
b101 +
#613150000000
0!
0'
#613160000000
1!
b110 %
1'
b110 +
#613170000000
0!
0'
#613180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#613190000000
0!
0'
#613200000000
1!
b1000 %
1'
b1000 +
#613210000000
0!
0'
#613220000000
1!
b1001 %
1'
b1001 +
#613230000000
0!
0'
#613240000000
1!
b0 %
1'
b0 +
#613250000000
0!
0'
#613260000000
1!
1$
b1 %
1'
1*
b1 +
#613270000000
0!
0'
#613280000000
1!
b10 %
1'
b10 +
#613290000000
0!
0'
#613300000000
1!
b11 %
1'
b11 +
#613310000000
0!
0'
#613320000000
1!
b100 %
1'
b100 +
#613330000000
0!
0'
#613340000000
1!
b101 %
1'
b101 +
#613350000000
0!
0'
#613360000000
1!
0$
b110 %
1'
0*
b110 +
#613370000000
0!
0'
#613380000000
1!
b111 %
1'
b111 +
#613390000000
1"
1(
#613400000000
0!
0"
b100 &
0'
0(
b100 ,
#613410000000
1!
b1000 %
1'
b1000 +
#613420000000
0!
0'
#613430000000
1!
b1001 %
1'
b1001 +
#613440000000
0!
0'
#613450000000
1!
b0 %
1'
b0 +
#613460000000
0!
0'
#613470000000
1!
1$
b1 %
1'
1*
b1 +
#613480000000
0!
0'
#613490000000
1!
b10 %
1'
b10 +
#613500000000
0!
0'
#613510000000
1!
b11 %
1'
b11 +
#613520000000
0!
0'
#613530000000
1!
b100 %
1'
b100 +
#613540000000
0!
0'
#613550000000
1!
b101 %
1'
b101 +
#613560000000
0!
0'
#613570000000
1!
b110 %
1'
b110 +
#613580000000
0!
0'
#613590000000
1!
b111 %
1'
b111 +
#613600000000
0!
0'
#613610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#613620000000
0!
0'
#613630000000
1!
b1001 %
1'
b1001 +
#613640000000
0!
0'
#613650000000
1!
b0 %
1'
b0 +
#613660000000
0!
0'
#613670000000
1!
1$
b1 %
1'
1*
b1 +
#613680000000
0!
0'
#613690000000
1!
b10 %
1'
b10 +
#613700000000
0!
0'
#613710000000
1!
b11 %
1'
b11 +
#613720000000
0!
0'
#613730000000
1!
b100 %
1'
b100 +
#613740000000
0!
0'
#613750000000
1!
b101 %
1'
b101 +
#613760000000
0!
0'
#613770000000
1!
0$
b110 %
1'
0*
b110 +
#613780000000
0!
0'
#613790000000
1!
b111 %
1'
b111 +
#613800000000
0!
0'
#613810000000
1!
b1000 %
1'
b1000 +
#613820000000
1"
1(
#613830000000
0!
0"
b100 &
0'
0(
b100 ,
#613840000000
1!
b1001 %
1'
b1001 +
#613850000000
0!
0'
#613860000000
1!
b0 %
1'
b0 +
#613870000000
0!
0'
#613880000000
1!
1$
b1 %
1'
1*
b1 +
#613890000000
0!
0'
#613900000000
1!
b10 %
1'
b10 +
#613910000000
0!
0'
#613920000000
1!
b11 %
1'
b11 +
#613930000000
0!
0'
#613940000000
1!
b100 %
1'
b100 +
#613950000000
0!
0'
#613960000000
1!
b101 %
1'
b101 +
#613970000000
0!
0'
#613980000000
1!
b110 %
1'
b110 +
#613990000000
0!
0'
#614000000000
1!
b111 %
1'
b111 +
#614010000000
0!
0'
#614020000000
1!
0$
b1000 %
1'
0*
b1000 +
#614030000000
0!
0'
#614040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#614050000000
0!
0'
#614060000000
1!
b0 %
1'
b0 +
#614070000000
0!
0'
#614080000000
1!
1$
b1 %
1'
1*
b1 +
#614090000000
0!
0'
#614100000000
1!
b10 %
1'
b10 +
#614110000000
0!
0'
#614120000000
1!
b11 %
1'
b11 +
#614130000000
0!
0'
#614140000000
1!
b100 %
1'
b100 +
#614150000000
0!
0'
#614160000000
1!
b101 %
1'
b101 +
#614170000000
0!
0'
#614180000000
1!
0$
b110 %
1'
0*
b110 +
#614190000000
0!
0'
#614200000000
1!
b111 %
1'
b111 +
#614210000000
0!
0'
#614220000000
1!
b1000 %
1'
b1000 +
#614230000000
0!
0'
#614240000000
1!
b1001 %
1'
b1001 +
#614250000000
1"
1(
#614260000000
0!
0"
b100 &
0'
0(
b100 ,
#614270000000
1!
b0 %
1'
b0 +
#614280000000
0!
0'
#614290000000
1!
1$
b1 %
1'
1*
b1 +
#614300000000
0!
0'
#614310000000
1!
b10 %
1'
b10 +
#614320000000
0!
0'
#614330000000
1!
b11 %
1'
b11 +
#614340000000
0!
0'
#614350000000
1!
b100 %
1'
b100 +
#614360000000
0!
0'
#614370000000
1!
b101 %
1'
b101 +
#614380000000
0!
0'
#614390000000
1!
b110 %
1'
b110 +
#614400000000
0!
0'
#614410000000
1!
b111 %
1'
b111 +
#614420000000
0!
0'
#614430000000
1!
0$
b1000 %
1'
0*
b1000 +
#614440000000
0!
0'
#614450000000
1!
b1001 %
1'
b1001 +
#614460000000
0!
0'
#614470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#614480000000
0!
0'
#614490000000
1!
1$
b1 %
1'
1*
b1 +
#614500000000
0!
0'
#614510000000
1!
b10 %
1'
b10 +
#614520000000
0!
0'
#614530000000
1!
b11 %
1'
b11 +
#614540000000
0!
0'
#614550000000
1!
b100 %
1'
b100 +
#614560000000
0!
0'
#614570000000
1!
b101 %
1'
b101 +
#614580000000
0!
0'
#614590000000
1!
0$
b110 %
1'
0*
b110 +
#614600000000
0!
0'
#614610000000
1!
b111 %
1'
b111 +
#614620000000
0!
0'
#614630000000
1!
b1000 %
1'
b1000 +
#614640000000
0!
0'
#614650000000
1!
b1001 %
1'
b1001 +
#614660000000
0!
0'
#614670000000
1!
b0 %
1'
b0 +
#614680000000
1"
1(
#614690000000
0!
0"
b100 &
0'
0(
b100 ,
#614700000000
1!
1$
b1 %
1'
1*
b1 +
#614710000000
0!
0'
#614720000000
1!
b10 %
1'
b10 +
#614730000000
0!
0'
#614740000000
1!
b11 %
1'
b11 +
#614750000000
0!
0'
#614760000000
1!
b100 %
1'
b100 +
#614770000000
0!
0'
#614780000000
1!
b101 %
1'
b101 +
#614790000000
0!
0'
#614800000000
1!
b110 %
1'
b110 +
#614810000000
0!
0'
#614820000000
1!
b111 %
1'
b111 +
#614830000000
0!
0'
#614840000000
1!
0$
b1000 %
1'
0*
b1000 +
#614850000000
0!
0'
#614860000000
1!
b1001 %
1'
b1001 +
#614870000000
0!
0'
#614880000000
1!
b0 %
1'
b0 +
#614890000000
0!
0'
#614900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#614910000000
0!
0'
#614920000000
1!
b10 %
1'
b10 +
#614930000000
0!
0'
#614940000000
1!
b11 %
1'
b11 +
#614950000000
0!
0'
#614960000000
1!
b100 %
1'
b100 +
#614970000000
0!
0'
#614980000000
1!
b101 %
1'
b101 +
#614990000000
0!
0'
#615000000000
1!
0$
b110 %
1'
0*
b110 +
#615010000000
0!
0'
#615020000000
1!
b111 %
1'
b111 +
#615030000000
0!
0'
#615040000000
1!
b1000 %
1'
b1000 +
#615050000000
0!
0'
#615060000000
1!
b1001 %
1'
b1001 +
#615070000000
0!
0'
#615080000000
1!
b0 %
1'
b0 +
#615090000000
0!
0'
#615100000000
1!
1$
b1 %
1'
1*
b1 +
#615110000000
1"
1(
#615120000000
0!
0"
b100 &
0'
0(
b100 ,
#615130000000
1!
b10 %
1'
b10 +
#615140000000
0!
0'
#615150000000
1!
b11 %
1'
b11 +
#615160000000
0!
0'
#615170000000
1!
b100 %
1'
b100 +
#615180000000
0!
0'
#615190000000
1!
b101 %
1'
b101 +
#615200000000
0!
0'
#615210000000
1!
b110 %
1'
b110 +
#615220000000
0!
0'
#615230000000
1!
b111 %
1'
b111 +
#615240000000
0!
0'
#615250000000
1!
0$
b1000 %
1'
0*
b1000 +
#615260000000
0!
0'
#615270000000
1!
b1001 %
1'
b1001 +
#615280000000
0!
0'
#615290000000
1!
b0 %
1'
b0 +
#615300000000
0!
0'
#615310000000
1!
1$
b1 %
1'
1*
b1 +
#615320000000
0!
0'
#615330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#615340000000
0!
0'
#615350000000
1!
b11 %
1'
b11 +
#615360000000
0!
0'
#615370000000
1!
b100 %
1'
b100 +
#615380000000
0!
0'
#615390000000
1!
b101 %
1'
b101 +
#615400000000
0!
0'
#615410000000
1!
0$
b110 %
1'
0*
b110 +
#615420000000
0!
0'
#615430000000
1!
b111 %
1'
b111 +
#615440000000
0!
0'
#615450000000
1!
b1000 %
1'
b1000 +
#615460000000
0!
0'
#615470000000
1!
b1001 %
1'
b1001 +
#615480000000
0!
0'
#615490000000
1!
b0 %
1'
b0 +
#615500000000
0!
0'
#615510000000
1!
1$
b1 %
1'
1*
b1 +
#615520000000
0!
0'
#615530000000
1!
b10 %
1'
b10 +
#615540000000
1"
1(
#615550000000
0!
0"
b100 &
0'
0(
b100 ,
#615560000000
1!
b11 %
1'
b11 +
#615570000000
0!
0'
#615580000000
1!
b100 %
1'
b100 +
#615590000000
0!
0'
#615600000000
1!
b101 %
1'
b101 +
#615610000000
0!
0'
#615620000000
1!
b110 %
1'
b110 +
#615630000000
0!
0'
#615640000000
1!
b111 %
1'
b111 +
#615650000000
0!
0'
#615660000000
1!
0$
b1000 %
1'
0*
b1000 +
#615670000000
0!
0'
#615680000000
1!
b1001 %
1'
b1001 +
#615690000000
0!
0'
#615700000000
1!
b0 %
1'
b0 +
#615710000000
0!
0'
#615720000000
1!
1$
b1 %
1'
1*
b1 +
#615730000000
0!
0'
#615740000000
1!
b10 %
1'
b10 +
#615750000000
0!
0'
#615760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#615770000000
0!
0'
#615780000000
1!
b100 %
1'
b100 +
#615790000000
0!
0'
#615800000000
1!
b101 %
1'
b101 +
#615810000000
0!
0'
#615820000000
1!
0$
b110 %
1'
0*
b110 +
#615830000000
0!
0'
#615840000000
1!
b111 %
1'
b111 +
#615850000000
0!
0'
#615860000000
1!
b1000 %
1'
b1000 +
#615870000000
0!
0'
#615880000000
1!
b1001 %
1'
b1001 +
#615890000000
0!
0'
#615900000000
1!
b0 %
1'
b0 +
#615910000000
0!
0'
#615920000000
1!
1$
b1 %
1'
1*
b1 +
#615930000000
0!
0'
#615940000000
1!
b10 %
1'
b10 +
#615950000000
0!
0'
#615960000000
1!
b11 %
1'
b11 +
#615970000000
1"
1(
#615980000000
0!
0"
b100 &
0'
0(
b100 ,
#615990000000
1!
b100 %
1'
b100 +
#616000000000
0!
0'
#616010000000
1!
b101 %
1'
b101 +
#616020000000
0!
0'
#616030000000
1!
b110 %
1'
b110 +
#616040000000
0!
0'
#616050000000
1!
b111 %
1'
b111 +
#616060000000
0!
0'
#616070000000
1!
0$
b1000 %
1'
0*
b1000 +
#616080000000
0!
0'
#616090000000
1!
b1001 %
1'
b1001 +
#616100000000
0!
0'
#616110000000
1!
b0 %
1'
b0 +
#616120000000
0!
0'
#616130000000
1!
1$
b1 %
1'
1*
b1 +
#616140000000
0!
0'
#616150000000
1!
b10 %
1'
b10 +
#616160000000
0!
0'
#616170000000
1!
b11 %
1'
b11 +
#616180000000
0!
0'
#616190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#616200000000
0!
0'
#616210000000
1!
b101 %
1'
b101 +
#616220000000
0!
0'
#616230000000
1!
0$
b110 %
1'
0*
b110 +
#616240000000
0!
0'
#616250000000
1!
b111 %
1'
b111 +
#616260000000
0!
0'
#616270000000
1!
b1000 %
1'
b1000 +
#616280000000
0!
0'
#616290000000
1!
b1001 %
1'
b1001 +
#616300000000
0!
0'
#616310000000
1!
b0 %
1'
b0 +
#616320000000
0!
0'
#616330000000
1!
1$
b1 %
1'
1*
b1 +
#616340000000
0!
0'
#616350000000
1!
b10 %
1'
b10 +
#616360000000
0!
0'
#616370000000
1!
b11 %
1'
b11 +
#616380000000
0!
0'
#616390000000
1!
b100 %
1'
b100 +
#616400000000
1"
1(
#616410000000
0!
0"
b100 &
0'
0(
b100 ,
#616420000000
1!
b101 %
1'
b101 +
#616430000000
0!
0'
#616440000000
1!
b110 %
1'
b110 +
#616450000000
0!
0'
#616460000000
1!
b111 %
1'
b111 +
#616470000000
0!
0'
#616480000000
1!
0$
b1000 %
1'
0*
b1000 +
#616490000000
0!
0'
#616500000000
1!
b1001 %
1'
b1001 +
#616510000000
0!
0'
#616520000000
1!
b0 %
1'
b0 +
#616530000000
0!
0'
#616540000000
1!
1$
b1 %
1'
1*
b1 +
#616550000000
0!
0'
#616560000000
1!
b10 %
1'
b10 +
#616570000000
0!
0'
#616580000000
1!
b11 %
1'
b11 +
#616590000000
0!
0'
#616600000000
1!
b100 %
1'
b100 +
#616610000000
0!
0'
#616620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#616630000000
0!
0'
#616640000000
1!
0$
b110 %
1'
0*
b110 +
#616650000000
0!
0'
#616660000000
1!
b111 %
1'
b111 +
#616670000000
0!
0'
#616680000000
1!
b1000 %
1'
b1000 +
#616690000000
0!
0'
#616700000000
1!
b1001 %
1'
b1001 +
#616710000000
0!
0'
#616720000000
1!
b0 %
1'
b0 +
#616730000000
0!
0'
#616740000000
1!
1$
b1 %
1'
1*
b1 +
#616750000000
0!
0'
#616760000000
1!
b10 %
1'
b10 +
#616770000000
0!
0'
#616780000000
1!
b11 %
1'
b11 +
#616790000000
0!
0'
#616800000000
1!
b100 %
1'
b100 +
#616810000000
0!
0'
#616820000000
1!
b101 %
1'
b101 +
#616830000000
1"
1(
#616840000000
0!
0"
b100 &
0'
0(
b100 ,
#616850000000
1!
b110 %
1'
b110 +
#616860000000
0!
0'
#616870000000
1!
b111 %
1'
b111 +
#616880000000
0!
0'
#616890000000
1!
0$
b1000 %
1'
0*
b1000 +
#616900000000
0!
0'
#616910000000
1!
b1001 %
1'
b1001 +
#616920000000
0!
0'
#616930000000
1!
b0 %
1'
b0 +
#616940000000
0!
0'
#616950000000
1!
1$
b1 %
1'
1*
b1 +
#616960000000
0!
0'
#616970000000
1!
b10 %
1'
b10 +
#616980000000
0!
0'
#616990000000
1!
b11 %
1'
b11 +
#617000000000
0!
0'
#617010000000
1!
b100 %
1'
b100 +
#617020000000
0!
0'
#617030000000
1!
b101 %
1'
b101 +
#617040000000
0!
0'
#617050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#617060000000
0!
0'
#617070000000
1!
b111 %
1'
b111 +
#617080000000
0!
0'
#617090000000
1!
b1000 %
1'
b1000 +
#617100000000
0!
0'
#617110000000
1!
b1001 %
1'
b1001 +
#617120000000
0!
0'
#617130000000
1!
b0 %
1'
b0 +
#617140000000
0!
0'
#617150000000
1!
1$
b1 %
1'
1*
b1 +
#617160000000
0!
0'
#617170000000
1!
b10 %
1'
b10 +
#617180000000
0!
0'
#617190000000
1!
b11 %
1'
b11 +
#617200000000
0!
0'
#617210000000
1!
b100 %
1'
b100 +
#617220000000
0!
0'
#617230000000
1!
b101 %
1'
b101 +
#617240000000
0!
0'
#617250000000
1!
0$
b110 %
1'
0*
b110 +
#617260000000
1"
1(
#617270000000
0!
0"
b100 &
0'
0(
b100 ,
#617280000000
1!
1$
b111 %
1'
1*
b111 +
#617290000000
0!
0'
#617300000000
1!
0$
b1000 %
1'
0*
b1000 +
#617310000000
0!
0'
#617320000000
1!
b1001 %
1'
b1001 +
#617330000000
0!
0'
#617340000000
1!
b0 %
1'
b0 +
#617350000000
0!
0'
#617360000000
1!
1$
b1 %
1'
1*
b1 +
#617370000000
0!
0'
#617380000000
1!
b10 %
1'
b10 +
#617390000000
0!
0'
#617400000000
1!
b11 %
1'
b11 +
#617410000000
0!
0'
#617420000000
1!
b100 %
1'
b100 +
#617430000000
0!
0'
#617440000000
1!
b101 %
1'
b101 +
#617450000000
0!
0'
#617460000000
1!
b110 %
1'
b110 +
#617470000000
0!
0'
#617480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#617490000000
0!
0'
#617500000000
1!
b1000 %
1'
b1000 +
#617510000000
0!
0'
#617520000000
1!
b1001 %
1'
b1001 +
#617530000000
0!
0'
#617540000000
1!
b0 %
1'
b0 +
#617550000000
0!
0'
#617560000000
1!
1$
b1 %
1'
1*
b1 +
#617570000000
0!
0'
#617580000000
1!
b10 %
1'
b10 +
#617590000000
0!
0'
#617600000000
1!
b11 %
1'
b11 +
#617610000000
0!
0'
#617620000000
1!
b100 %
1'
b100 +
#617630000000
0!
0'
#617640000000
1!
b101 %
1'
b101 +
#617650000000
0!
0'
#617660000000
1!
0$
b110 %
1'
0*
b110 +
#617670000000
0!
0'
#617680000000
1!
b111 %
1'
b111 +
#617690000000
1"
1(
#617700000000
0!
0"
b100 &
0'
0(
b100 ,
#617710000000
1!
b1000 %
1'
b1000 +
#617720000000
0!
0'
#617730000000
1!
b1001 %
1'
b1001 +
#617740000000
0!
0'
#617750000000
1!
b0 %
1'
b0 +
#617760000000
0!
0'
#617770000000
1!
1$
b1 %
1'
1*
b1 +
#617780000000
0!
0'
#617790000000
1!
b10 %
1'
b10 +
#617800000000
0!
0'
#617810000000
1!
b11 %
1'
b11 +
#617820000000
0!
0'
#617830000000
1!
b100 %
1'
b100 +
#617840000000
0!
0'
#617850000000
1!
b101 %
1'
b101 +
#617860000000
0!
0'
#617870000000
1!
b110 %
1'
b110 +
#617880000000
0!
0'
#617890000000
1!
b111 %
1'
b111 +
#617900000000
0!
0'
#617910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#617920000000
0!
0'
#617930000000
1!
b1001 %
1'
b1001 +
#617940000000
0!
0'
#617950000000
1!
b0 %
1'
b0 +
#617960000000
0!
0'
#617970000000
1!
1$
b1 %
1'
1*
b1 +
#617980000000
0!
0'
#617990000000
1!
b10 %
1'
b10 +
#618000000000
0!
0'
#618010000000
1!
b11 %
1'
b11 +
#618020000000
0!
0'
#618030000000
1!
b100 %
1'
b100 +
#618040000000
0!
0'
#618050000000
1!
b101 %
1'
b101 +
#618060000000
0!
0'
#618070000000
1!
0$
b110 %
1'
0*
b110 +
#618080000000
0!
0'
#618090000000
1!
b111 %
1'
b111 +
#618100000000
0!
0'
#618110000000
1!
b1000 %
1'
b1000 +
#618120000000
1"
1(
#618130000000
0!
0"
b100 &
0'
0(
b100 ,
#618140000000
1!
b1001 %
1'
b1001 +
#618150000000
0!
0'
#618160000000
1!
b0 %
1'
b0 +
#618170000000
0!
0'
#618180000000
1!
1$
b1 %
1'
1*
b1 +
#618190000000
0!
0'
#618200000000
1!
b10 %
1'
b10 +
#618210000000
0!
0'
#618220000000
1!
b11 %
1'
b11 +
#618230000000
0!
0'
#618240000000
1!
b100 %
1'
b100 +
#618250000000
0!
0'
#618260000000
1!
b101 %
1'
b101 +
#618270000000
0!
0'
#618280000000
1!
b110 %
1'
b110 +
#618290000000
0!
0'
#618300000000
1!
b111 %
1'
b111 +
#618310000000
0!
0'
#618320000000
1!
0$
b1000 %
1'
0*
b1000 +
#618330000000
0!
0'
#618340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#618350000000
0!
0'
#618360000000
1!
b0 %
1'
b0 +
#618370000000
0!
0'
#618380000000
1!
1$
b1 %
1'
1*
b1 +
#618390000000
0!
0'
#618400000000
1!
b10 %
1'
b10 +
#618410000000
0!
0'
#618420000000
1!
b11 %
1'
b11 +
#618430000000
0!
0'
#618440000000
1!
b100 %
1'
b100 +
#618450000000
0!
0'
#618460000000
1!
b101 %
1'
b101 +
#618470000000
0!
0'
#618480000000
1!
0$
b110 %
1'
0*
b110 +
#618490000000
0!
0'
#618500000000
1!
b111 %
1'
b111 +
#618510000000
0!
0'
#618520000000
1!
b1000 %
1'
b1000 +
#618530000000
0!
0'
#618540000000
1!
b1001 %
1'
b1001 +
#618550000000
1"
1(
#618560000000
0!
0"
b100 &
0'
0(
b100 ,
#618570000000
1!
b0 %
1'
b0 +
#618580000000
0!
0'
#618590000000
1!
1$
b1 %
1'
1*
b1 +
#618600000000
0!
0'
#618610000000
1!
b10 %
1'
b10 +
#618620000000
0!
0'
#618630000000
1!
b11 %
1'
b11 +
#618640000000
0!
0'
#618650000000
1!
b100 %
1'
b100 +
#618660000000
0!
0'
#618670000000
1!
b101 %
1'
b101 +
#618680000000
0!
0'
#618690000000
1!
b110 %
1'
b110 +
#618700000000
0!
0'
#618710000000
1!
b111 %
1'
b111 +
#618720000000
0!
0'
#618730000000
1!
0$
b1000 %
1'
0*
b1000 +
#618740000000
0!
0'
#618750000000
1!
b1001 %
1'
b1001 +
#618760000000
0!
0'
#618770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#618780000000
0!
0'
#618790000000
1!
1$
b1 %
1'
1*
b1 +
#618800000000
0!
0'
#618810000000
1!
b10 %
1'
b10 +
#618820000000
0!
0'
#618830000000
1!
b11 %
1'
b11 +
#618840000000
0!
0'
#618850000000
1!
b100 %
1'
b100 +
#618860000000
0!
0'
#618870000000
1!
b101 %
1'
b101 +
#618880000000
0!
0'
#618890000000
1!
0$
b110 %
1'
0*
b110 +
#618900000000
0!
0'
#618910000000
1!
b111 %
1'
b111 +
#618920000000
0!
0'
#618930000000
1!
b1000 %
1'
b1000 +
#618940000000
0!
0'
#618950000000
1!
b1001 %
1'
b1001 +
#618960000000
0!
0'
#618970000000
1!
b0 %
1'
b0 +
#618980000000
1"
1(
#618990000000
0!
0"
b100 &
0'
0(
b100 ,
#619000000000
1!
1$
b1 %
1'
1*
b1 +
#619010000000
0!
0'
#619020000000
1!
b10 %
1'
b10 +
#619030000000
0!
0'
#619040000000
1!
b11 %
1'
b11 +
#619050000000
0!
0'
#619060000000
1!
b100 %
1'
b100 +
#619070000000
0!
0'
#619080000000
1!
b101 %
1'
b101 +
#619090000000
0!
0'
#619100000000
1!
b110 %
1'
b110 +
#619110000000
0!
0'
#619120000000
1!
b111 %
1'
b111 +
#619130000000
0!
0'
#619140000000
1!
0$
b1000 %
1'
0*
b1000 +
#619150000000
0!
0'
#619160000000
1!
b1001 %
1'
b1001 +
#619170000000
0!
0'
#619180000000
1!
b0 %
1'
b0 +
#619190000000
0!
0'
#619200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#619210000000
0!
0'
#619220000000
1!
b10 %
1'
b10 +
#619230000000
0!
0'
#619240000000
1!
b11 %
1'
b11 +
#619250000000
0!
0'
#619260000000
1!
b100 %
1'
b100 +
#619270000000
0!
0'
#619280000000
1!
b101 %
1'
b101 +
#619290000000
0!
0'
#619300000000
1!
0$
b110 %
1'
0*
b110 +
#619310000000
0!
0'
#619320000000
1!
b111 %
1'
b111 +
#619330000000
0!
0'
#619340000000
1!
b1000 %
1'
b1000 +
#619350000000
0!
0'
#619360000000
1!
b1001 %
1'
b1001 +
#619370000000
0!
0'
#619380000000
1!
b0 %
1'
b0 +
#619390000000
0!
0'
#619400000000
1!
1$
b1 %
1'
1*
b1 +
#619410000000
1"
1(
#619420000000
0!
0"
b100 &
0'
0(
b100 ,
#619430000000
1!
b10 %
1'
b10 +
#619440000000
0!
0'
#619450000000
1!
b11 %
1'
b11 +
#619460000000
0!
0'
#619470000000
1!
b100 %
1'
b100 +
#619480000000
0!
0'
#619490000000
1!
b101 %
1'
b101 +
#619500000000
0!
0'
#619510000000
1!
b110 %
1'
b110 +
#619520000000
0!
0'
#619530000000
1!
b111 %
1'
b111 +
#619540000000
0!
0'
#619550000000
1!
0$
b1000 %
1'
0*
b1000 +
#619560000000
0!
0'
#619570000000
1!
b1001 %
1'
b1001 +
#619580000000
0!
0'
#619590000000
1!
b0 %
1'
b0 +
#619600000000
0!
0'
#619610000000
1!
1$
b1 %
1'
1*
b1 +
#619620000000
0!
0'
#619630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#619640000000
0!
0'
#619650000000
1!
b11 %
1'
b11 +
#619660000000
0!
0'
#619670000000
1!
b100 %
1'
b100 +
#619680000000
0!
0'
#619690000000
1!
b101 %
1'
b101 +
#619700000000
0!
0'
#619710000000
1!
0$
b110 %
1'
0*
b110 +
#619720000000
0!
0'
#619730000000
1!
b111 %
1'
b111 +
#619740000000
0!
0'
#619750000000
1!
b1000 %
1'
b1000 +
#619760000000
0!
0'
#619770000000
1!
b1001 %
1'
b1001 +
#619780000000
0!
0'
#619790000000
1!
b0 %
1'
b0 +
#619800000000
0!
0'
#619810000000
1!
1$
b1 %
1'
1*
b1 +
#619820000000
0!
0'
#619830000000
1!
b10 %
1'
b10 +
#619840000000
1"
1(
#619850000000
0!
0"
b100 &
0'
0(
b100 ,
#619860000000
1!
b11 %
1'
b11 +
#619870000000
0!
0'
#619880000000
1!
b100 %
1'
b100 +
#619890000000
0!
0'
#619900000000
1!
b101 %
1'
b101 +
#619910000000
0!
0'
#619920000000
1!
b110 %
1'
b110 +
#619930000000
0!
0'
#619940000000
1!
b111 %
1'
b111 +
#619950000000
0!
0'
#619960000000
1!
0$
b1000 %
1'
0*
b1000 +
#619970000000
0!
0'
#619980000000
1!
b1001 %
1'
b1001 +
#619990000000
0!
0'
#620000000000
1!
b0 %
1'
b0 +
#620010000000
0!
0'
#620020000000
1!
1$
b1 %
1'
1*
b1 +
#620030000000
0!
0'
#620040000000
1!
b10 %
1'
b10 +
#620050000000
0!
0'
#620060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#620070000000
0!
0'
#620080000000
1!
b100 %
1'
b100 +
#620090000000
0!
0'
#620100000000
1!
b101 %
1'
b101 +
#620110000000
0!
0'
#620120000000
1!
0$
b110 %
1'
0*
b110 +
#620130000000
0!
0'
#620140000000
1!
b111 %
1'
b111 +
#620150000000
0!
0'
#620160000000
1!
b1000 %
1'
b1000 +
#620170000000
0!
0'
#620180000000
1!
b1001 %
1'
b1001 +
#620190000000
0!
0'
#620200000000
1!
b0 %
1'
b0 +
#620210000000
0!
0'
#620220000000
1!
1$
b1 %
1'
1*
b1 +
#620230000000
0!
0'
#620240000000
1!
b10 %
1'
b10 +
#620250000000
0!
0'
#620260000000
1!
b11 %
1'
b11 +
#620270000000
1"
1(
#620280000000
0!
0"
b100 &
0'
0(
b100 ,
#620290000000
1!
b100 %
1'
b100 +
#620300000000
0!
0'
#620310000000
1!
b101 %
1'
b101 +
#620320000000
0!
0'
#620330000000
1!
b110 %
1'
b110 +
#620340000000
0!
0'
#620350000000
1!
b111 %
1'
b111 +
#620360000000
0!
0'
#620370000000
1!
0$
b1000 %
1'
0*
b1000 +
#620380000000
0!
0'
#620390000000
1!
b1001 %
1'
b1001 +
#620400000000
0!
0'
#620410000000
1!
b0 %
1'
b0 +
#620420000000
0!
0'
#620430000000
1!
1$
b1 %
1'
1*
b1 +
#620440000000
0!
0'
#620450000000
1!
b10 %
1'
b10 +
#620460000000
0!
0'
#620470000000
1!
b11 %
1'
b11 +
#620480000000
0!
0'
#620490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#620500000000
0!
0'
#620510000000
1!
b101 %
1'
b101 +
#620520000000
0!
0'
#620530000000
1!
0$
b110 %
1'
0*
b110 +
#620540000000
0!
0'
#620550000000
1!
b111 %
1'
b111 +
#620560000000
0!
0'
#620570000000
1!
b1000 %
1'
b1000 +
#620580000000
0!
0'
#620590000000
1!
b1001 %
1'
b1001 +
#620600000000
0!
0'
#620610000000
1!
b0 %
1'
b0 +
#620620000000
0!
0'
#620630000000
1!
1$
b1 %
1'
1*
b1 +
#620640000000
0!
0'
#620650000000
1!
b10 %
1'
b10 +
#620660000000
0!
0'
#620670000000
1!
b11 %
1'
b11 +
#620680000000
0!
0'
#620690000000
1!
b100 %
1'
b100 +
#620700000000
1"
1(
#620710000000
0!
0"
b100 &
0'
0(
b100 ,
#620720000000
1!
b101 %
1'
b101 +
#620730000000
0!
0'
#620740000000
1!
b110 %
1'
b110 +
#620750000000
0!
0'
#620760000000
1!
b111 %
1'
b111 +
#620770000000
0!
0'
#620780000000
1!
0$
b1000 %
1'
0*
b1000 +
#620790000000
0!
0'
#620800000000
1!
b1001 %
1'
b1001 +
#620810000000
0!
0'
#620820000000
1!
b0 %
1'
b0 +
#620830000000
0!
0'
#620840000000
1!
1$
b1 %
1'
1*
b1 +
#620850000000
0!
0'
#620860000000
1!
b10 %
1'
b10 +
#620870000000
0!
0'
#620880000000
1!
b11 %
1'
b11 +
#620890000000
0!
0'
#620900000000
1!
b100 %
1'
b100 +
#620910000000
0!
0'
#620920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#620930000000
0!
0'
#620940000000
1!
0$
b110 %
1'
0*
b110 +
#620950000000
0!
0'
#620960000000
1!
b111 %
1'
b111 +
#620970000000
0!
0'
#620980000000
1!
b1000 %
1'
b1000 +
#620990000000
0!
0'
#621000000000
1!
b1001 %
1'
b1001 +
#621010000000
0!
0'
#621020000000
1!
b0 %
1'
b0 +
#621030000000
0!
0'
#621040000000
1!
1$
b1 %
1'
1*
b1 +
#621050000000
0!
0'
#621060000000
1!
b10 %
1'
b10 +
#621070000000
0!
0'
#621080000000
1!
b11 %
1'
b11 +
#621090000000
0!
0'
#621100000000
1!
b100 %
1'
b100 +
#621110000000
0!
0'
#621120000000
1!
b101 %
1'
b101 +
#621130000000
1"
1(
#621140000000
0!
0"
b100 &
0'
0(
b100 ,
#621150000000
1!
b110 %
1'
b110 +
#621160000000
0!
0'
#621170000000
1!
b111 %
1'
b111 +
#621180000000
0!
0'
#621190000000
1!
0$
b1000 %
1'
0*
b1000 +
#621200000000
0!
0'
#621210000000
1!
b1001 %
1'
b1001 +
#621220000000
0!
0'
#621230000000
1!
b0 %
1'
b0 +
#621240000000
0!
0'
#621250000000
1!
1$
b1 %
1'
1*
b1 +
#621260000000
0!
0'
#621270000000
1!
b10 %
1'
b10 +
#621280000000
0!
0'
#621290000000
1!
b11 %
1'
b11 +
#621300000000
0!
0'
#621310000000
1!
b100 %
1'
b100 +
#621320000000
0!
0'
#621330000000
1!
b101 %
1'
b101 +
#621340000000
0!
0'
#621350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#621360000000
0!
0'
#621370000000
1!
b111 %
1'
b111 +
#621380000000
0!
0'
#621390000000
1!
b1000 %
1'
b1000 +
#621400000000
0!
0'
#621410000000
1!
b1001 %
1'
b1001 +
#621420000000
0!
0'
#621430000000
1!
b0 %
1'
b0 +
#621440000000
0!
0'
#621450000000
1!
1$
b1 %
1'
1*
b1 +
#621460000000
0!
0'
#621470000000
1!
b10 %
1'
b10 +
#621480000000
0!
0'
#621490000000
1!
b11 %
1'
b11 +
#621500000000
0!
0'
#621510000000
1!
b100 %
1'
b100 +
#621520000000
0!
0'
#621530000000
1!
b101 %
1'
b101 +
#621540000000
0!
0'
#621550000000
1!
0$
b110 %
1'
0*
b110 +
#621560000000
1"
1(
#621570000000
0!
0"
b100 &
0'
0(
b100 ,
#621580000000
1!
1$
b111 %
1'
1*
b111 +
#621590000000
0!
0'
#621600000000
1!
0$
b1000 %
1'
0*
b1000 +
#621610000000
0!
0'
#621620000000
1!
b1001 %
1'
b1001 +
#621630000000
0!
0'
#621640000000
1!
b0 %
1'
b0 +
#621650000000
0!
0'
#621660000000
1!
1$
b1 %
1'
1*
b1 +
#621670000000
0!
0'
#621680000000
1!
b10 %
1'
b10 +
#621690000000
0!
0'
#621700000000
1!
b11 %
1'
b11 +
#621710000000
0!
0'
#621720000000
1!
b100 %
1'
b100 +
#621730000000
0!
0'
#621740000000
1!
b101 %
1'
b101 +
#621750000000
0!
0'
#621760000000
1!
b110 %
1'
b110 +
#621770000000
0!
0'
#621780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#621790000000
0!
0'
#621800000000
1!
b1000 %
1'
b1000 +
#621810000000
0!
0'
#621820000000
1!
b1001 %
1'
b1001 +
#621830000000
0!
0'
#621840000000
1!
b0 %
1'
b0 +
#621850000000
0!
0'
#621860000000
1!
1$
b1 %
1'
1*
b1 +
#621870000000
0!
0'
#621880000000
1!
b10 %
1'
b10 +
#621890000000
0!
0'
#621900000000
1!
b11 %
1'
b11 +
#621910000000
0!
0'
#621920000000
1!
b100 %
1'
b100 +
#621930000000
0!
0'
#621940000000
1!
b101 %
1'
b101 +
#621950000000
0!
0'
#621960000000
1!
0$
b110 %
1'
0*
b110 +
#621970000000
0!
0'
#621980000000
1!
b111 %
1'
b111 +
#621990000000
1"
1(
#622000000000
0!
0"
b100 &
0'
0(
b100 ,
#622010000000
1!
b1000 %
1'
b1000 +
#622020000000
0!
0'
#622030000000
1!
b1001 %
1'
b1001 +
#622040000000
0!
0'
#622050000000
1!
b0 %
1'
b0 +
#622060000000
0!
0'
#622070000000
1!
1$
b1 %
1'
1*
b1 +
#622080000000
0!
0'
#622090000000
1!
b10 %
1'
b10 +
#622100000000
0!
0'
#622110000000
1!
b11 %
1'
b11 +
#622120000000
0!
0'
#622130000000
1!
b100 %
1'
b100 +
#622140000000
0!
0'
#622150000000
1!
b101 %
1'
b101 +
#622160000000
0!
0'
#622170000000
1!
b110 %
1'
b110 +
#622180000000
0!
0'
#622190000000
1!
b111 %
1'
b111 +
#622200000000
0!
0'
#622210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#622220000000
0!
0'
#622230000000
1!
b1001 %
1'
b1001 +
#622240000000
0!
0'
#622250000000
1!
b0 %
1'
b0 +
#622260000000
0!
0'
#622270000000
1!
1$
b1 %
1'
1*
b1 +
#622280000000
0!
0'
#622290000000
1!
b10 %
1'
b10 +
#622300000000
0!
0'
#622310000000
1!
b11 %
1'
b11 +
#622320000000
0!
0'
#622330000000
1!
b100 %
1'
b100 +
#622340000000
0!
0'
#622350000000
1!
b101 %
1'
b101 +
#622360000000
0!
0'
#622370000000
1!
0$
b110 %
1'
0*
b110 +
#622380000000
0!
0'
#622390000000
1!
b111 %
1'
b111 +
#622400000000
0!
0'
#622410000000
1!
b1000 %
1'
b1000 +
#622420000000
1"
1(
#622430000000
0!
0"
b100 &
0'
0(
b100 ,
#622440000000
1!
b1001 %
1'
b1001 +
#622450000000
0!
0'
#622460000000
1!
b0 %
1'
b0 +
#622470000000
0!
0'
#622480000000
1!
1$
b1 %
1'
1*
b1 +
#622490000000
0!
0'
#622500000000
1!
b10 %
1'
b10 +
#622510000000
0!
0'
#622520000000
1!
b11 %
1'
b11 +
#622530000000
0!
0'
#622540000000
1!
b100 %
1'
b100 +
#622550000000
0!
0'
#622560000000
1!
b101 %
1'
b101 +
#622570000000
0!
0'
#622580000000
1!
b110 %
1'
b110 +
#622590000000
0!
0'
#622600000000
1!
b111 %
1'
b111 +
#622610000000
0!
0'
#622620000000
1!
0$
b1000 %
1'
0*
b1000 +
#622630000000
0!
0'
#622640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#622650000000
0!
0'
#622660000000
1!
b0 %
1'
b0 +
#622670000000
0!
0'
#622680000000
1!
1$
b1 %
1'
1*
b1 +
#622690000000
0!
0'
#622700000000
1!
b10 %
1'
b10 +
#622710000000
0!
0'
#622720000000
1!
b11 %
1'
b11 +
#622730000000
0!
0'
#622740000000
1!
b100 %
1'
b100 +
#622750000000
0!
0'
#622760000000
1!
b101 %
1'
b101 +
#622770000000
0!
0'
#622780000000
1!
0$
b110 %
1'
0*
b110 +
#622790000000
0!
0'
#622800000000
1!
b111 %
1'
b111 +
#622810000000
0!
0'
#622820000000
1!
b1000 %
1'
b1000 +
#622830000000
0!
0'
#622840000000
1!
b1001 %
1'
b1001 +
#622850000000
1"
1(
#622860000000
0!
0"
b100 &
0'
0(
b100 ,
#622870000000
1!
b0 %
1'
b0 +
#622880000000
0!
0'
#622890000000
1!
1$
b1 %
1'
1*
b1 +
#622900000000
0!
0'
#622910000000
1!
b10 %
1'
b10 +
#622920000000
0!
0'
#622930000000
1!
b11 %
1'
b11 +
#622940000000
0!
0'
#622950000000
1!
b100 %
1'
b100 +
#622960000000
0!
0'
#622970000000
1!
b101 %
1'
b101 +
#622980000000
0!
0'
#622990000000
1!
b110 %
1'
b110 +
#623000000000
0!
0'
#623010000000
1!
b111 %
1'
b111 +
#623020000000
0!
0'
#623030000000
1!
0$
b1000 %
1'
0*
b1000 +
#623040000000
0!
0'
#623050000000
1!
b1001 %
1'
b1001 +
#623060000000
0!
0'
#623070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#623080000000
0!
0'
#623090000000
1!
1$
b1 %
1'
1*
b1 +
#623100000000
0!
0'
#623110000000
1!
b10 %
1'
b10 +
#623120000000
0!
0'
#623130000000
1!
b11 %
1'
b11 +
#623140000000
0!
0'
#623150000000
1!
b100 %
1'
b100 +
#623160000000
0!
0'
#623170000000
1!
b101 %
1'
b101 +
#623180000000
0!
0'
#623190000000
1!
0$
b110 %
1'
0*
b110 +
#623200000000
0!
0'
#623210000000
1!
b111 %
1'
b111 +
#623220000000
0!
0'
#623230000000
1!
b1000 %
1'
b1000 +
#623240000000
0!
0'
#623250000000
1!
b1001 %
1'
b1001 +
#623260000000
0!
0'
#623270000000
1!
b0 %
1'
b0 +
#623280000000
1"
1(
#623290000000
0!
0"
b100 &
0'
0(
b100 ,
#623300000000
1!
1$
b1 %
1'
1*
b1 +
#623310000000
0!
0'
#623320000000
1!
b10 %
1'
b10 +
#623330000000
0!
0'
#623340000000
1!
b11 %
1'
b11 +
#623350000000
0!
0'
#623360000000
1!
b100 %
1'
b100 +
#623370000000
0!
0'
#623380000000
1!
b101 %
1'
b101 +
#623390000000
0!
0'
#623400000000
1!
b110 %
1'
b110 +
#623410000000
0!
0'
#623420000000
1!
b111 %
1'
b111 +
#623430000000
0!
0'
#623440000000
1!
0$
b1000 %
1'
0*
b1000 +
#623450000000
0!
0'
#623460000000
1!
b1001 %
1'
b1001 +
#623470000000
0!
0'
#623480000000
1!
b0 %
1'
b0 +
#623490000000
0!
0'
#623500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#623510000000
0!
0'
#623520000000
1!
b10 %
1'
b10 +
#623530000000
0!
0'
#623540000000
1!
b11 %
1'
b11 +
#623550000000
0!
0'
#623560000000
1!
b100 %
1'
b100 +
#623570000000
0!
0'
#623580000000
1!
b101 %
1'
b101 +
#623590000000
0!
0'
#623600000000
1!
0$
b110 %
1'
0*
b110 +
#623610000000
0!
0'
#623620000000
1!
b111 %
1'
b111 +
#623630000000
0!
0'
#623640000000
1!
b1000 %
1'
b1000 +
#623650000000
0!
0'
#623660000000
1!
b1001 %
1'
b1001 +
#623670000000
0!
0'
#623680000000
1!
b0 %
1'
b0 +
#623690000000
0!
0'
#623700000000
1!
1$
b1 %
1'
1*
b1 +
#623710000000
1"
1(
#623720000000
0!
0"
b100 &
0'
0(
b100 ,
#623730000000
1!
b10 %
1'
b10 +
#623740000000
0!
0'
#623750000000
1!
b11 %
1'
b11 +
#623760000000
0!
0'
#623770000000
1!
b100 %
1'
b100 +
#623780000000
0!
0'
#623790000000
1!
b101 %
1'
b101 +
#623800000000
0!
0'
#623810000000
1!
b110 %
1'
b110 +
#623820000000
0!
0'
#623830000000
1!
b111 %
1'
b111 +
#623840000000
0!
0'
#623850000000
1!
0$
b1000 %
1'
0*
b1000 +
#623860000000
0!
0'
#623870000000
1!
b1001 %
1'
b1001 +
#623880000000
0!
0'
#623890000000
1!
b0 %
1'
b0 +
#623900000000
0!
0'
#623910000000
1!
1$
b1 %
1'
1*
b1 +
#623920000000
0!
0'
#623930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#623940000000
0!
0'
#623950000000
1!
b11 %
1'
b11 +
#623960000000
0!
0'
#623970000000
1!
b100 %
1'
b100 +
#623980000000
0!
0'
#623990000000
1!
b101 %
1'
b101 +
#624000000000
0!
0'
#624010000000
1!
0$
b110 %
1'
0*
b110 +
#624020000000
0!
0'
#624030000000
1!
b111 %
1'
b111 +
#624040000000
0!
0'
#624050000000
1!
b1000 %
1'
b1000 +
#624060000000
0!
0'
#624070000000
1!
b1001 %
1'
b1001 +
#624080000000
0!
0'
#624090000000
1!
b0 %
1'
b0 +
#624100000000
0!
0'
#624110000000
1!
1$
b1 %
1'
1*
b1 +
#624120000000
0!
0'
#624130000000
1!
b10 %
1'
b10 +
#624140000000
1"
1(
#624150000000
0!
0"
b100 &
0'
0(
b100 ,
#624160000000
1!
b11 %
1'
b11 +
#624170000000
0!
0'
#624180000000
1!
b100 %
1'
b100 +
#624190000000
0!
0'
#624200000000
1!
b101 %
1'
b101 +
#624210000000
0!
0'
#624220000000
1!
b110 %
1'
b110 +
#624230000000
0!
0'
#624240000000
1!
b111 %
1'
b111 +
#624250000000
0!
0'
#624260000000
1!
0$
b1000 %
1'
0*
b1000 +
#624270000000
0!
0'
#624280000000
1!
b1001 %
1'
b1001 +
#624290000000
0!
0'
#624300000000
1!
b0 %
1'
b0 +
#624310000000
0!
0'
#624320000000
1!
1$
b1 %
1'
1*
b1 +
#624330000000
0!
0'
#624340000000
1!
b10 %
1'
b10 +
#624350000000
0!
0'
#624360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#624370000000
0!
0'
#624380000000
1!
b100 %
1'
b100 +
#624390000000
0!
0'
#624400000000
1!
b101 %
1'
b101 +
#624410000000
0!
0'
#624420000000
1!
0$
b110 %
1'
0*
b110 +
#624430000000
0!
0'
#624440000000
1!
b111 %
1'
b111 +
#624450000000
0!
0'
#624460000000
1!
b1000 %
1'
b1000 +
#624470000000
0!
0'
#624480000000
1!
b1001 %
1'
b1001 +
#624490000000
0!
0'
#624500000000
1!
b0 %
1'
b0 +
#624510000000
0!
0'
#624520000000
1!
1$
b1 %
1'
1*
b1 +
#624530000000
0!
0'
#624540000000
1!
b10 %
1'
b10 +
#624550000000
0!
0'
#624560000000
1!
b11 %
1'
b11 +
#624570000000
1"
1(
#624580000000
0!
0"
b100 &
0'
0(
b100 ,
#624590000000
1!
b100 %
1'
b100 +
#624600000000
0!
0'
#624610000000
1!
b101 %
1'
b101 +
#624620000000
0!
0'
#624630000000
1!
b110 %
1'
b110 +
#624640000000
0!
0'
#624650000000
1!
b111 %
1'
b111 +
#624660000000
0!
0'
#624670000000
1!
0$
b1000 %
1'
0*
b1000 +
#624680000000
0!
0'
#624690000000
1!
b1001 %
1'
b1001 +
#624700000000
0!
0'
#624710000000
1!
b0 %
1'
b0 +
#624720000000
0!
0'
#624730000000
1!
1$
b1 %
1'
1*
b1 +
#624740000000
0!
0'
#624750000000
1!
b10 %
1'
b10 +
#624760000000
0!
0'
#624770000000
1!
b11 %
1'
b11 +
#624780000000
0!
0'
#624790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#624800000000
0!
0'
#624810000000
1!
b101 %
1'
b101 +
#624820000000
0!
0'
#624830000000
1!
0$
b110 %
1'
0*
b110 +
#624840000000
0!
0'
#624850000000
1!
b111 %
1'
b111 +
#624860000000
0!
0'
#624870000000
1!
b1000 %
1'
b1000 +
#624880000000
0!
0'
#624890000000
1!
b1001 %
1'
b1001 +
#624900000000
0!
0'
#624910000000
1!
b0 %
1'
b0 +
#624920000000
0!
0'
#624930000000
1!
1$
b1 %
1'
1*
b1 +
#624940000000
0!
0'
#624950000000
1!
b10 %
1'
b10 +
#624960000000
0!
0'
#624970000000
1!
b11 %
1'
b11 +
#624980000000
0!
0'
#624990000000
1!
b100 %
1'
b100 +
#625000000000
1"
1(
#625010000000
0!
0"
b100 &
0'
0(
b100 ,
#625020000000
1!
b101 %
1'
b101 +
#625030000000
0!
0'
#625040000000
1!
b110 %
1'
b110 +
#625050000000
0!
0'
#625060000000
1!
b111 %
1'
b111 +
#625070000000
0!
0'
#625080000000
1!
0$
b1000 %
1'
0*
b1000 +
#625090000000
0!
0'
#625100000000
1!
b1001 %
1'
b1001 +
#625110000000
0!
0'
#625120000000
1!
b0 %
1'
b0 +
#625130000000
0!
0'
#625140000000
1!
1$
b1 %
1'
1*
b1 +
#625150000000
0!
0'
#625160000000
1!
b10 %
1'
b10 +
#625170000000
0!
0'
#625180000000
1!
b11 %
1'
b11 +
#625190000000
0!
0'
#625200000000
1!
b100 %
1'
b100 +
#625210000000
0!
0'
#625220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#625230000000
0!
0'
#625240000000
1!
0$
b110 %
1'
0*
b110 +
#625250000000
0!
0'
#625260000000
1!
b111 %
1'
b111 +
#625270000000
0!
0'
#625280000000
1!
b1000 %
1'
b1000 +
#625290000000
0!
0'
#625300000000
1!
b1001 %
1'
b1001 +
#625310000000
0!
0'
#625320000000
1!
b0 %
1'
b0 +
#625330000000
0!
0'
#625340000000
1!
1$
b1 %
1'
1*
b1 +
#625350000000
0!
0'
#625360000000
1!
b10 %
1'
b10 +
#625370000000
0!
0'
#625380000000
1!
b11 %
1'
b11 +
#625390000000
0!
0'
#625400000000
1!
b100 %
1'
b100 +
#625410000000
0!
0'
#625420000000
1!
b101 %
1'
b101 +
#625430000000
1"
1(
#625440000000
0!
0"
b100 &
0'
0(
b100 ,
#625450000000
1!
b110 %
1'
b110 +
#625460000000
0!
0'
#625470000000
1!
b111 %
1'
b111 +
#625480000000
0!
0'
#625490000000
1!
0$
b1000 %
1'
0*
b1000 +
#625500000000
0!
0'
#625510000000
1!
b1001 %
1'
b1001 +
#625520000000
0!
0'
#625530000000
1!
b0 %
1'
b0 +
#625540000000
0!
0'
#625550000000
1!
1$
b1 %
1'
1*
b1 +
#625560000000
0!
0'
#625570000000
1!
b10 %
1'
b10 +
#625580000000
0!
0'
#625590000000
1!
b11 %
1'
b11 +
#625600000000
0!
0'
#625610000000
1!
b100 %
1'
b100 +
#625620000000
0!
0'
#625630000000
1!
b101 %
1'
b101 +
#625640000000
0!
0'
#625650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#625660000000
0!
0'
#625670000000
1!
b111 %
1'
b111 +
#625680000000
0!
0'
#625690000000
1!
b1000 %
1'
b1000 +
#625700000000
0!
0'
#625710000000
1!
b1001 %
1'
b1001 +
#625720000000
0!
0'
#625730000000
1!
b0 %
1'
b0 +
#625740000000
0!
0'
#625750000000
1!
1$
b1 %
1'
1*
b1 +
#625760000000
0!
0'
#625770000000
1!
b10 %
1'
b10 +
#625780000000
0!
0'
#625790000000
1!
b11 %
1'
b11 +
#625800000000
0!
0'
#625810000000
1!
b100 %
1'
b100 +
#625820000000
0!
0'
#625830000000
1!
b101 %
1'
b101 +
#625840000000
0!
0'
#625850000000
1!
0$
b110 %
1'
0*
b110 +
#625860000000
1"
1(
#625870000000
0!
0"
b100 &
0'
0(
b100 ,
#625880000000
1!
1$
b111 %
1'
1*
b111 +
#625890000000
0!
0'
#625900000000
1!
0$
b1000 %
1'
0*
b1000 +
#625910000000
0!
0'
#625920000000
1!
b1001 %
1'
b1001 +
#625930000000
0!
0'
#625940000000
1!
b0 %
1'
b0 +
#625950000000
0!
0'
#625960000000
1!
1$
b1 %
1'
1*
b1 +
#625970000000
0!
0'
#625980000000
1!
b10 %
1'
b10 +
#625990000000
0!
0'
#626000000000
1!
b11 %
1'
b11 +
#626010000000
0!
0'
#626020000000
1!
b100 %
1'
b100 +
#626030000000
0!
0'
#626040000000
1!
b101 %
1'
b101 +
#626050000000
0!
0'
#626060000000
1!
b110 %
1'
b110 +
#626070000000
0!
0'
#626080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#626090000000
0!
0'
#626100000000
1!
b1000 %
1'
b1000 +
#626110000000
0!
0'
#626120000000
1!
b1001 %
1'
b1001 +
#626130000000
0!
0'
#626140000000
1!
b0 %
1'
b0 +
#626150000000
0!
0'
#626160000000
1!
1$
b1 %
1'
1*
b1 +
#626170000000
0!
0'
#626180000000
1!
b10 %
1'
b10 +
#626190000000
0!
0'
#626200000000
1!
b11 %
1'
b11 +
#626210000000
0!
0'
#626220000000
1!
b100 %
1'
b100 +
#626230000000
0!
0'
#626240000000
1!
b101 %
1'
b101 +
#626250000000
0!
0'
#626260000000
1!
0$
b110 %
1'
0*
b110 +
#626270000000
0!
0'
#626280000000
1!
b111 %
1'
b111 +
#626290000000
1"
1(
#626300000000
0!
0"
b100 &
0'
0(
b100 ,
#626310000000
1!
b1000 %
1'
b1000 +
#626320000000
0!
0'
#626330000000
1!
b1001 %
1'
b1001 +
#626340000000
0!
0'
#626350000000
1!
b0 %
1'
b0 +
#626360000000
0!
0'
#626370000000
1!
1$
b1 %
1'
1*
b1 +
#626380000000
0!
0'
#626390000000
1!
b10 %
1'
b10 +
#626400000000
0!
0'
#626410000000
1!
b11 %
1'
b11 +
#626420000000
0!
0'
#626430000000
1!
b100 %
1'
b100 +
#626440000000
0!
0'
#626450000000
1!
b101 %
1'
b101 +
#626460000000
0!
0'
#626470000000
1!
b110 %
1'
b110 +
#626480000000
0!
0'
#626490000000
1!
b111 %
1'
b111 +
#626500000000
0!
0'
#626510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#626520000000
0!
0'
#626530000000
1!
b1001 %
1'
b1001 +
#626540000000
0!
0'
#626550000000
1!
b0 %
1'
b0 +
#626560000000
0!
0'
#626570000000
1!
1$
b1 %
1'
1*
b1 +
#626580000000
0!
0'
#626590000000
1!
b10 %
1'
b10 +
#626600000000
0!
0'
#626610000000
1!
b11 %
1'
b11 +
#626620000000
0!
0'
#626630000000
1!
b100 %
1'
b100 +
#626640000000
0!
0'
#626650000000
1!
b101 %
1'
b101 +
#626660000000
0!
0'
#626670000000
1!
0$
b110 %
1'
0*
b110 +
#626680000000
0!
0'
#626690000000
1!
b111 %
1'
b111 +
#626700000000
0!
0'
#626710000000
1!
b1000 %
1'
b1000 +
#626720000000
1"
1(
#626730000000
0!
0"
b100 &
0'
0(
b100 ,
#626740000000
1!
b1001 %
1'
b1001 +
#626750000000
0!
0'
#626760000000
1!
b0 %
1'
b0 +
#626770000000
0!
0'
#626780000000
1!
1$
b1 %
1'
1*
b1 +
#626790000000
0!
0'
#626800000000
1!
b10 %
1'
b10 +
#626810000000
0!
0'
#626820000000
1!
b11 %
1'
b11 +
#626830000000
0!
0'
#626840000000
1!
b100 %
1'
b100 +
#626850000000
0!
0'
#626860000000
1!
b101 %
1'
b101 +
#626870000000
0!
0'
#626880000000
1!
b110 %
1'
b110 +
#626890000000
0!
0'
#626900000000
1!
b111 %
1'
b111 +
#626910000000
0!
0'
#626920000000
1!
0$
b1000 %
1'
0*
b1000 +
#626930000000
0!
0'
#626940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#626950000000
0!
0'
#626960000000
1!
b0 %
1'
b0 +
#626970000000
0!
0'
#626980000000
1!
1$
b1 %
1'
1*
b1 +
#626990000000
0!
0'
#627000000000
1!
b10 %
1'
b10 +
#627010000000
0!
0'
#627020000000
1!
b11 %
1'
b11 +
#627030000000
0!
0'
#627040000000
1!
b100 %
1'
b100 +
#627050000000
0!
0'
#627060000000
1!
b101 %
1'
b101 +
#627070000000
0!
0'
#627080000000
1!
0$
b110 %
1'
0*
b110 +
#627090000000
0!
0'
#627100000000
1!
b111 %
1'
b111 +
#627110000000
0!
0'
#627120000000
1!
b1000 %
1'
b1000 +
#627130000000
0!
0'
#627140000000
1!
b1001 %
1'
b1001 +
#627150000000
1"
1(
#627160000000
0!
0"
b100 &
0'
0(
b100 ,
#627170000000
1!
b0 %
1'
b0 +
#627180000000
0!
0'
#627190000000
1!
1$
b1 %
1'
1*
b1 +
#627200000000
0!
0'
#627210000000
1!
b10 %
1'
b10 +
#627220000000
0!
0'
#627230000000
1!
b11 %
1'
b11 +
#627240000000
0!
0'
#627250000000
1!
b100 %
1'
b100 +
#627260000000
0!
0'
#627270000000
1!
b101 %
1'
b101 +
#627280000000
0!
0'
#627290000000
1!
b110 %
1'
b110 +
#627300000000
0!
0'
#627310000000
1!
b111 %
1'
b111 +
#627320000000
0!
0'
#627330000000
1!
0$
b1000 %
1'
0*
b1000 +
#627340000000
0!
0'
#627350000000
1!
b1001 %
1'
b1001 +
#627360000000
0!
0'
#627370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#627380000000
0!
0'
#627390000000
1!
1$
b1 %
1'
1*
b1 +
#627400000000
0!
0'
#627410000000
1!
b10 %
1'
b10 +
#627420000000
0!
0'
#627430000000
1!
b11 %
1'
b11 +
#627440000000
0!
0'
#627450000000
1!
b100 %
1'
b100 +
#627460000000
0!
0'
#627470000000
1!
b101 %
1'
b101 +
#627480000000
0!
0'
#627490000000
1!
0$
b110 %
1'
0*
b110 +
#627500000000
0!
0'
#627510000000
1!
b111 %
1'
b111 +
#627520000000
0!
0'
#627530000000
1!
b1000 %
1'
b1000 +
#627540000000
0!
0'
#627550000000
1!
b1001 %
1'
b1001 +
#627560000000
0!
0'
#627570000000
1!
b0 %
1'
b0 +
#627580000000
1"
1(
#627590000000
0!
0"
b100 &
0'
0(
b100 ,
#627600000000
1!
1$
b1 %
1'
1*
b1 +
#627610000000
0!
0'
#627620000000
1!
b10 %
1'
b10 +
#627630000000
0!
0'
#627640000000
1!
b11 %
1'
b11 +
#627650000000
0!
0'
#627660000000
1!
b100 %
1'
b100 +
#627670000000
0!
0'
#627680000000
1!
b101 %
1'
b101 +
#627690000000
0!
0'
#627700000000
1!
b110 %
1'
b110 +
#627710000000
0!
0'
#627720000000
1!
b111 %
1'
b111 +
#627730000000
0!
0'
#627740000000
1!
0$
b1000 %
1'
0*
b1000 +
#627750000000
0!
0'
#627760000000
1!
b1001 %
1'
b1001 +
#627770000000
0!
0'
#627780000000
1!
b0 %
1'
b0 +
#627790000000
0!
0'
#627800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#627810000000
0!
0'
#627820000000
1!
b10 %
1'
b10 +
#627830000000
0!
0'
#627840000000
1!
b11 %
1'
b11 +
#627850000000
0!
0'
#627860000000
1!
b100 %
1'
b100 +
#627870000000
0!
0'
#627880000000
1!
b101 %
1'
b101 +
#627890000000
0!
0'
#627900000000
1!
0$
b110 %
1'
0*
b110 +
#627910000000
0!
0'
#627920000000
1!
b111 %
1'
b111 +
#627930000000
0!
0'
#627940000000
1!
b1000 %
1'
b1000 +
#627950000000
0!
0'
#627960000000
1!
b1001 %
1'
b1001 +
#627970000000
0!
0'
#627980000000
1!
b0 %
1'
b0 +
#627990000000
0!
0'
#628000000000
1!
1$
b1 %
1'
1*
b1 +
#628010000000
1"
1(
#628020000000
0!
0"
b100 &
0'
0(
b100 ,
#628030000000
1!
b10 %
1'
b10 +
#628040000000
0!
0'
#628050000000
1!
b11 %
1'
b11 +
#628060000000
0!
0'
#628070000000
1!
b100 %
1'
b100 +
#628080000000
0!
0'
#628090000000
1!
b101 %
1'
b101 +
#628100000000
0!
0'
#628110000000
1!
b110 %
1'
b110 +
#628120000000
0!
0'
#628130000000
1!
b111 %
1'
b111 +
#628140000000
0!
0'
#628150000000
1!
0$
b1000 %
1'
0*
b1000 +
#628160000000
0!
0'
#628170000000
1!
b1001 %
1'
b1001 +
#628180000000
0!
0'
#628190000000
1!
b0 %
1'
b0 +
#628200000000
0!
0'
#628210000000
1!
1$
b1 %
1'
1*
b1 +
#628220000000
0!
0'
#628230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#628240000000
0!
0'
#628250000000
1!
b11 %
1'
b11 +
#628260000000
0!
0'
#628270000000
1!
b100 %
1'
b100 +
#628280000000
0!
0'
#628290000000
1!
b101 %
1'
b101 +
#628300000000
0!
0'
#628310000000
1!
0$
b110 %
1'
0*
b110 +
#628320000000
0!
0'
#628330000000
1!
b111 %
1'
b111 +
#628340000000
0!
0'
#628350000000
1!
b1000 %
1'
b1000 +
#628360000000
0!
0'
#628370000000
1!
b1001 %
1'
b1001 +
#628380000000
0!
0'
#628390000000
1!
b0 %
1'
b0 +
#628400000000
0!
0'
#628410000000
1!
1$
b1 %
1'
1*
b1 +
#628420000000
0!
0'
#628430000000
1!
b10 %
1'
b10 +
#628440000000
1"
1(
#628450000000
0!
0"
b100 &
0'
0(
b100 ,
#628460000000
1!
b11 %
1'
b11 +
#628470000000
0!
0'
#628480000000
1!
b100 %
1'
b100 +
#628490000000
0!
0'
#628500000000
1!
b101 %
1'
b101 +
#628510000000
0!
0'
#628520000000
1!
b110 %
1'
b110 +
#628530000000
0!
0'
#628540000000
1!
b111 %
1'
b111 +
#628550000000
0!
0'
#628560000000
1!
0$
b1000 %
1'
0*
b1000 +
#628570000000
0!
0'
#628580000000
1!
b1001 %
1'
b1001 +
#628590000000
0!
0'
#628600000000
1!
b0 %
1'
b0 +
#628610000000
0!
0'
#628620000000
1!
1$
b1 %
1'
1*
b1 +
#628630000000
0!
0'
#628640000000
1!
b10 %
1'
b10 +
#628650000000
0!
0'
#628660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#628670000000
0!
0'
#628680000000
1!
b100 %
1'
b100 +
#628690000000
0!
0'
#628700000000
1!
b101 %
1'
b101 +
#628710000000
0!
0'
#628720000000
1!
0$
b110 %
1'
0*
b110 +
#628730000000
0!
0'
#628740000000
1!
b111 %
1'
b111 +
#628750000000
0!
0'
#628760000000
1!
b1000 %
1'
b1000 +
#628770000000
0!
0'
#628780000000
1!
b1001 %
1'
b1001 +
#628790000000
0!
0'
#628800000000
1!
b0 %
1'
b0 +
#628810000000
0!
0'
#628820000000
1!
1$
b1 %
1'
1*
b1 +
#628830000000
0!
0'
#628840000000
1!
b10 %
1'
b10 +
#628850000000
0!
0'
#628860000000
1!
b11 %
1'
b11 +
#628870000000
1"
1(
#628880000000
0!
0"
b100 &
0'
0(
b100 ,
#628890000000
1!
b100 %
1'
b100 +
#628900000000
0!
0'
#628910000000
1!
b101 %
1'
b101 +
#628920000000
0!
0'
#628930000000
1!
b110 %
1'
b110 +
#628940000000
0!
0'
#628950000000
1!
b111 %
1'
b111 +
#628960000000
0!
0'
#628970000000
1!
0$
b1000 %
1'
0*
b1000 +
#628980000000
0!
0'
#628990000000
1!
b1001 %
1'
b1001 +
#629000000000
0!
0'
#629010000000
1!
b0 %
1'
b0 +
#629020000000
0!
0'
#629030000000
1!
1$
b1 %
1'
1*
b1 +
#629040000000
0!
0'
#629050000000
1!
b10 %
1'
b10 +
#629060000000
0!
0'
#629070000000
1!
b11 %
1'
b11 +
#629080000000
0!
0'
#629090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#629100000000
0!
0'
#629110000000
1!
b101 %
1'
b101 +
#629120000000
0!
0'
#629130000000
1!
0$
b110 %
1'
0*
b110 +
#629140000000
0!
0'
#629150000000
1!
b111 %
1'
b111 +
#629160000000
0!
0'
#629170000000
1!
b1000 %
1'
b1000 +
#629180000000
0!
0'
#629190000000
1!
b1001 %
1'
b1001 +
#629200000000
0!
0'
#629210000000
1!
b0 %
1'
b0 +
#629220000000
0!
0'
#629230000000
1!
1$
b1 %
1'
1*
b1 +
#629240000000
0!
0'
#629250000000
1!
b10 %
1'
b10 +
#629260000000
0!
0'
#629270000000
1!
b11 %
1'
b11 +
#629280000000
0!
0'
#629290000000
1!
b100 %
1'
b100 +
#629300000000
1"
1(
#629310000000
0!
0"
b100 &
0'
0(
b100 ,
#629320000000
1!
b101 %
1'
b101 +
#629330000000
0!
0'
#629340000000
1!
b110 %
1'
b110 +
#629350000000
0!
0'
#629360000000
1!
b111 %
1'
b111 +
#629370000000
0!
0'
#629380000000
1!
0$
b1000 %
1'
0*
b1000 +
#629390000000
0!
0'
#629400000000
1!
b1001 %
1'
b1001 +
#629410000000
0!
0'
#629420000000
1!
b0 %
1'
b0 +
#629430000000
0!
0'
#629440000000
1!
1$
b1 %
1'
1*
b1 +
#629450000000
0!
0'
#629460000000
1!
b10 %
1'
b10 +
#629470000000
0!
0'
#629480000000
1!
b11 %
1'
b11 +
#629490000000
0!
0'
#629500000000
1!
b100 %
1'
b100 +
#629510000000
0!
0'
#629520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#629530000000
0!
0'
#629540000000
1!
0$
b110 %
1'
0*
b110 +
#629550000000
0!
0'
#629560000000
1!
b111 %
1'
b111 +
#629570000000
0!
0'
#629580000000
1!
b1000 %
1'
b1000 +
#629590000000
0!
0'
#629600000000
1!
b1001 %
1'
b1001 +
#629610000000
0!
0'
#629620000000
1!
b0 %
1'
b0 +
#629630000000
0!
0'
#629640000000
1!
1$
b1 %
1'
1*
b1 +
#629650000000
0!
0'
#629660000000
1!
b10 %
1'
b10 +
#629670000000
0!
0'
#629680000000
1!
b11 %
1'
b11 +
#629690000000
0!
0'
#629700000000
1!
b100 %
1'
b100 +
#629710000000
0!
0'
#629720000000
1!
b101 %
1'
b101 +
#629730000000
1"
1(
#629740000000
0!
0"
b100 &
0'
0(
b100 ,
#629750000000
1!
b110 %
1'
b110 +
#629760000000
0!
0'
#629770000000
1!
b111 %
1'
b111 +
#629780000000
0!
0'
#629790000000
1!
0$
b1000 %
1'
0*
b1000 +
#629800000000
0!
0'
#629810000000
1!
b1001 %
1'
b1001 +
#629820000000
0!
0'
#629830000000
1!
b0 %
1'
b0 +
#629840000000
0!
0'
#629850000000
1!
1$
b1 %
1'
1*
b1 +
#629860000000
0!
0'
#629870000000
1!
b10 %
1'
b10 +
#629880000000
0!
0'
#629890000000
1!
b11 %
1'
b11 +
#629900000000
0!
0'
#629910000000
1!
b100 %
1'
b100 +
#629920000000
0!
0'
#629930000000
1!
b101 %
1'
b101 +
#629940000000
0!
0'
#629950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#629960000000
0!
0'
#629970000000
1!
b111 %
1'
b111 +
#629980000000
0!
0'
#629990000000
1!
b1000 %
1'
b1000 +
#630000000000
0!
0'
#630010000000
1!
b1001 %
1'
b1001 +
#630020000000
0!
0'
#630030000000
1!
b0 %
1'
b0 +
#630040000000
0!
0'
#630050000000
1!
1$
b1 %
1'
1*
b1 +
#630060000000
0!
0'
#630070000000
1!
b10 %
1'
b10 +
#630080000000
0!
0'
#630090000000
1!
b11 %
1'
b11 +
#630100000000
0!
0'
#630110000000
1!
b100 %
1'
b100 +
#630120000000
0!
0'
#630130000000
1!
b101 %
1'
b101 +
#630140000000
0!
0'
#630150000000
1!
0$
b110 %
1'
0*
b110 +
#630160000000
1"
1(
#630170000000
0!
0"
b100 &
0'
0(
b100 ,
#630180000000
1!
1$
b111 %
1'
1*
b111 +
#630190000000
0!
0'
#630200000000
1!
0$
b1000 %
1'
0*
b1000 +
#630210000000
0!
0'
#630220000000
1!
b1001 %
1'
b1001 +
#630230000000
0!
0'
#630240000000
1!
b0 %
1'
b0 +
#630250000000
0!
0'
#630260000000
1!
1$
b1 %
1'
1*
b1 +
#630270000000
0!
0'
#630280000000
1!
b10 %
1'
b10 +
#630290000000
0!
0'
#630300000000
1!
b11 %
1'
b11 +
#630310000000
0!
0'
#630320000000
1!
b100 %
1'
b100 +
#630330000000
0!
0'
#630340000000
1!
b101 %
1'
b101 +
#630350000000
0!
0'
#630360000000
1!
b110 %
1'
b110 +
#630370000000
0!
0'
#630380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#630390000000
0!
0'
#630400000000
1!
b1000 %
1'
b1000 +
#630410000000
0!
0'
#630420000000
1!
b1001 %
1'
b1001 +
#630430000000
0!
0'
#630440000000
1!
b0 %
1'
b0 +
#630450000000
0!
0'
#630460000000
1!
1$
b1 %
1'
1*
b1 +
#630470000000
0!
0'
#630480000000
1!
b10 %
1'
b10 +
#630490000000
0!
0'
#630500000000
1!
b11 %
1'
b11 +
#630510000000
0!
0'
#630520000000
1!
b100 %
1'
b100 +
#630530000000
0!
0'
#630540000000
1!
b101 %
1'
b101 +
#630550000000
0!
0'
#630560000000
1!
0$
b110 %
1'
0*
b110 +
#630570000000
0!
0'
#630580000000
1!
b111 %
1'
b111 +
#630590000000
1"
1(
#630600000000
0!
0"
b100 &
0'
0(
b100 ,
#630610000000
1!
b1000 %
1'
b1000 +
#630620000000
0!
0'
#630630000000
1!
b1001 %
1'
b1001 +
#630640000000
0!
0'
#630650000000
1!
b0 %
1'
b0 +
#630660000000
0!
0'
#630670000000
1!
1$
b1 %
1'
1*
b1 +
#630680000000
0!
0'
#630690000000
1!
b10 %
1'
b10 +
#630700000000
0!
0'
#630710000000
1!
b11 %
1'
b11 +
#630720000000
0!
0'
#630730000000
1!
b100 %
1'
b100 +
#630740000000
0!
0'
#630750000000
1!
b101 %
1'
b101 +
#630760000000
0!
0'
#630770000000
1!
b110 %
1'
b110 +
#630780000000
0!
0'
#630790000000
1!
b111 %
1'
b111 +
#630800000000
0!
0'
#630810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#630820000000
0!
0'
#630830000000
1!
b1001 %
1'
b1001 +
#630840000000
0!
0'
#630850000000
1!
b0 %
1'
b0 +
#630860000000
0!
0'
#630870000000
1!
1$
b1 %
1'
1*
b1 +
#630880000000
0!
0'
#630890000000
1!
b10 %
1'
b10 +
#630900000000
0!
0'
#630910000000
1!
b11 %
1'
b11 +
#630920000000
0!
0'
#630930000000
1!
b100 %
1'
b100 +
#630940000000
0!
0'
#630950000000
1!
b101 %
1'
b101 +
#630960000000
0!
0'
#630970000000
1!
0$
b110 %
1'
0*
b110 +
#630980000000
0!
0'
#630990000000
1!
b111 %
1'
b111 +
#631000000000
0!
0'
#631010000000
1!
b1000 %
1'
b1000 +
#631020000000
1"
1(
#631030000000
0!
0"
b100 &
0'
0(
b100 ,
#631040000000
1!
b1001 %
1'
b1001 +
#631050000000
0!
0'
#631060000000
1!
b0 %
1'
b0 +
#631070000000
0!
0'
#631080000000
1!
1$
b1 %
1'
1*
b1 +
#631090000000
0!
0'
#631100000000
1!
b10 %
1'
b10 +
#631110000000
0!
0'
#631120000000
1!
b11 %
1'
b11 +
#631130000000
0!
0'
#631140000000
1!
b100 %
1'
b100 +
#631150000000
0!
0'
#631160000000
1!
b101 %
1'
b101 +
#631170000000
0!
0'
#631180000000
1!
b110 %
1'
b110 +
#631190000000
0!
0'
#631200000000
1!
b111 %
1'
b111 +
#631210000000
0!
0'
#631220000000
1!
0$
b1000 %
1'
0*
b1000 +
#631230000000
0!
0'
#631240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#631250000000
0!
0'
#631260000000
1!
b0 %
1'
b0 +
#631270000000
0!
0'
#631280000000
1!
1$
b1 %
1'
1*
b1 +
#631290000000
0!
0'
#631300000000
1!
b10 %
1'
b10 +
#631310000000
0!
0'
#631320000000
1!
b11 %
1'
b11 +
#631330000000
0!
0'
#631340000000
1!
b100 %
1'
b100 +
#631350000000
0!
0'
#631360000000
1!
b101 %
1'
b101 +
#631370000000
0!
0'
#631380000000
1!
0$
b110 %
1'
0*
b110 +
#631390000000
0!
0'
#631400000000
1!
b111 %
1'
b111 +
#631410000000
0!
0'
#631420000000
1!
b1000 %
1'
b1000 +
#631430000000
0!
0'
#631440000000
1!
b1001 %
1'
b1001 +
#631450000000
1"
1(
#631460000000
0!
0"
b100 &
0'
0(
b100 ,
#631470000000
1!
b0 %
1'
b0 +
#631480000000
0!
0'
#631490000000
1!
1$
b1 %
1'
1*
b1 +
#631500000000
0!
0'
#631510000000
1!
b10 %
1'
b10 +
#631520000000
0!
0'
#631530000000
1!
b11 %
1'
b11 +
#631540000000
0!
0'
#631550000000
1!
b100 %
1'
b100 +
#631560000000
0!
0'
#631570000000
1!
b101 %
1'
b101 +
#631580000000
0!
0'
#631590000000
1!
b110 %
1'
b110 +
#631600000000
0!
0'
#631610000000
1!
b111 %
1'
b111 +
#631620000000
0!
0'
#631630000000
1!
0$
b1000 %
1'
0*
b1000 +
#631640000000
0!
0'
#631650000000
1!
b1001 %
1'
b1001 +
#631660000000
0!
0'
#631670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#631680000000
0!
0'
#631690000000
1!
1$
b1 %
1'
1*
b1 +
#631700000000
0!
0'
#631710000000
1!
b10 %
1'
b10 +
#631720000000
0!
0'
#631730000000
1!
b11 %
1'
b11 +
#631740000000
0!
0'
#631750000000
1!
b100 %
1'
b100 +
#631760000000
0!
0'
#631770000000
1!
b101 %
1'
b101 +
#631780000000
0!
0'
#631790000000
1!
0$
b110 %
1'
0*
b110 +
#631800000000
0!
0'
#631810000000
1!
b111 %
1'
b111 +
#631820000000
0!
0'
#631830000000
1!
b1000 %
1'
b1000 +
#631840000000
0!
0'
#631850000000
1!
b1001 %
1'
b1001 +
#631860000000
0!
0'
#631870000000
1!
b0 %
1'
b0 +
#631880000000
1"
1(
#631890000000
0!
0"
b100 &
0'
0(
b100 ,
#631900000000
1!
1$
b1 %
1'
1*
b1 +
#631910000000
0!
0'
#631920000000
1!
b10 %
1'
b10 +
#631930000000
0!
0'
#631940000000
1!
b11 %
1'
b11 +
#631950000000
0!
0'
#631960000000
1!
b100 %
1'
b100 +
#631970000000
0!
0'
#631980000000
1!
b101 %
1'
b101 +
#631990000000
0!
0'
#632000000000
1!
b110 %
1'
b110 +
#632010000000
0!
0'
#632020000000
1!
b111 %
1'
b111 +
#632030000000
0!
0'
#632040000000
1!
0$
b1000 %
1'
0*
b1000 +
#632050000000
0!
0'
#632060000000
1!
b1001 %
1'
b1001 +
#632070000000
0!
0'
#632080000000
1!
b0 %
1'
b0 +
#632090000000
0!
0'
#632100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#632110000000
0!
0'
#632120000000
1!
b10 %
1'
b10 +
#632130000000
0!
0'
#632140000000
1!
b11 %
1'
b11 +
#632150000000
0!
0'
#632160000000
1!
b100 %
1'
b100 +
#632170000000
0!
0'
#632180000000
1!
b101 %
1'
b101 +
#632190000000
0!
0'
#632200000000
1!
0$
b110 %
1'
0*
b110 +
#632210000000
0!
0'
#632220000000
1!
b111 %
1'
b111 +
#632230000000
0!
0'
#632240000000
1!
b1000 %
1'
b1000 +
#632250000000
0!
0'
#632260000000
1!
b1001 %
1'
b1001 +
#632270000000
0!
0'
#632280000000
1!
b0 %
1'
b0 +
#632290000000
0!
0'
#632300000000
1!
1$
b1 %
1'
1*
b1 +
#632310000000
1"
1(
#632320000000
0!
0"
b100 &
0'
0(
b100 ,
#632330000000
1!
b10 %
1'
b10 +
#632340000000
0!
0'
#632350000000
1!
b11 %
1'
b11 +
#632360000000
0!
0'
#632370000000
1!
b100 %
1'
b100 +
#632380000000
0!
0'
#632390000000
1!
b101 %
1'
b101 +
#632400000000
0!
0'
#632410000000
1!
b110 %
1'
b110 +
#632420000000
0!
0'
#632430000000
1!
b111 %
1'
b111 +
#632440000000
0!
0'
#632450000000
1!
0$
b1000 %
1'
0*
b1000 +
#632460000000
0!
0'
#632470000000
1!
b1001 %
1'
b1001 +
#632480000000
0!
0'
#632490000000
1!
b0 %
1'
b0 +
#632500000000
0!
0'
#632510000000
1!
1$
b1 %
1'
1*
b1 +
#632520000000
0!
0'
#632530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#632540000000
0!
0'
#632550000000
1!
b11 %
1'
b11 +
#632560000000
0!
0'
#632570000000
1!
b100 %
1'
b100 +
#632580000000
0!
0'
#632590000000
1!
b101 %
1'
b101 +
#632600000000
0!
0'
#632610000000
1!
0$
b110 %
1'
0*
b110 +
#632620000000
0!
0'
#632630000000
1!
b111 %
1'
b111 +
#632640000000
0!
0'
#632650000000
1!
b1000 %
1'
b1000 +
#632660000000
0!
0'
#632670000000
1!
b1001 %
1'
b1001 +
#632680000000
0!
0'
#632690000000
1!
b0 %
1'
b0 +
#632700000000
0!
0'
#632710000000
1!
1$
b1 %
1'
1*
b1 +
#632720000000
0!
0'
#632730000000
1!
b10 %
1'
b10 +
#632740000000
1"
1(
#632750000000
0!
0"
b100 &
0'
0(
b100 ,
#632760000000
1!
b11 %
1'
b11 +
#632770000000
0!
0'
#632780000000
1!
b100 %
1'
b100 +
#632790000000
0!
0'
#632800000000
1!
b101 %
1'
b101 +
#632810000000
0!
0'
#632820000000
1!
b110 %
1'
b110 +
#632830000000
0!
0'
#632840000000
1!
b111 %
1'
b111 +
#632850000000
0!
0'
#632860000000
1!
0$
b1000 %
1'
0*
b1000 +
#632870000000
0!
0'
#632880000000
1!
b1001 %
1'
b1001 +
#632890000000
0!
0'
#632900000000
1!
b0 %
1'
b0 +
#632910000000
0!
0'
#632920000000
1!
1$
b1 %
1'
1*
b1 +
#632930000000
0!
0'
#632940000000
1!
b10 %
1'
b10 +
#632950000000
0!
0'
#632960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#632970000000
0!
0'
#632980000000
1!
b100 %
1'
b100 +
#632990000000
0!
0'
#633000000000
1!
b101 %
1'
b101 +
#633010000000
0!
0'
#633020000000
1!
0$
b110 %
1'
0*
b110 +
#633030000000
0!
0'
#633040000000
1!
b111 %
1'
b111 +
#633050000000
0!
0'
#633060000000
1!
b1000 %
1'
b1000 +
#633070000000
0!
0'
#633080000000
1!
b1001 %
1'
b1001 +
#633090000000
0!
0'
#633100000000
1!
b0 %
1'
b0 +
#633110000000
0!
0'
#633120000000
1!
1$
b1 %
1'
1*
b1 +
#633130000000
0!
0'
#633140000000
1!
b10 %
1'
b10 +
#633150000000
0!
0'
#633160000000
1!
b11 %
1'
b11 +
#633170000000
1"
1(
#633180000000
0!
0"
b100 &
0'
0(
b100 ,
#633190000000
1!
b100 %
1'
b100 +
#633200000000
0!
0'
#633210000000
1!
b101 %
1'
b101 +
#633220000000
0!
0'
#633230000000
1!
b110 %
1'
b110 +
#633240000000
0!
0'
#633250000000
1!
b111 %
1'
b111 +
#633260000000
0!
0'
#633270000000
1!
0$
b1000 %
1'
0*
b1000 +
#633280000000
0!
0'
#633290000000
1!
b1001 %
1'
b1001 +
#633300000000
0!
0'
#633310000000
1!
b0 %
1'
b0 +
#633320000000
0!
0'
#633330000000
1!
1$
b1 %
1'
1*
b1 +
#633340000000
0!
0'
#633350000000
1!
b10 %
1'
b10 +
#633360000000
0!
0'
#633370000000
1!
b11 %
1'
b11 +
#633380000000
0!
0'
#633390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#633400000000
0!
0'
#633410000000
1!
b101 %
1'
b101 +
#633420000000
0!
0'
#633430000000
1!
0$
b110 %
1'
0*
b110 +
#633440000000
0!
0'
#633450000000
1!
b111 %
1'
b111 +
#633460000000
0!
0'
#633470000000
1!
b1000 %
1'
b1000 +
#633480000000
0!
0'
#633490000000
1!
b1001 %
1'
b1001 +
#633500000000
0!
0'
#633510000000
1!
b0 %
1'
b0 +
#633520000000
0!
0'
#633530000000
1!
1$
b1 %
1'
1*
b1 +
#633540000000
0!
0'
#633550000000
1!
b10 %
1'
b10 +
#633560000000
0!
0'
#633570000000
1!
b11 %
1'
b11 +
#633580000000
0!
0'
#633590000000
1!
b100 %
1'
b100 +
#633600000000
1"
1(
#633610000000
0!
0"
b100 &
0'
0(
b100 ,
#633620000000
1!
b101 %
1'
b101 +
#633630000000
0!
0'
#633640000000
1!
b110 %
1'
b110 +
#633650000000
0!
0'
#633660000000
1!
b111 %
1'
b111 +
#633670000000
0!
0'
#633680000000
1!
0$
b1000 %
1'
0*
b1000 +
#633690000000
0!
0'
#633700000000
1!
b1001 %
1'
b1001 +
#633710000000
0!
0'
#633720000000
1!
b0 %
1'
b0 +
#633730000000
0!
0'
#633740000000
1!
1$
b1 %
1'
1*
b1 +
#633750000000
0!
0'
#633760000000
1!
b10 %
1'
b10 +
#633770000000
0!
0'
#633780000000
1!
b11 %
1'
b11 +
#633790000000
0!
0'
#633800000000
1!
b100 %
1'
b100 +
#633810000000
0!
0'
#633820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#633830000000
0!
0'
#633840000000
1!
0$
b110 %
1'
0*
b110 +
#633850000000
0!
0'
#633860000000
1!
b111 %
1'
b111 +
#633870000000
0!
0'
#633880000000
1!
b1000 %
1'
b1000 +
#633890000000
0!
0'
#633900000000
1!
b1001 %
1'
b1001 +
#633910000000
0!
0'
#633920000000
1!
b0 %
1'
b0 +
#633930000000
0!
0'
#633940000000
1!
1$
b1 %
1'
1*
b1 +
#633950000000
0!
0'
#633960000000
1!
b10 %
1'
b10 +
#633970000000
0!
0'
#633980000000
1!
b11 %
1'
b11 +
#633990000000
0!
0'
#634000000000
1!
b100 %
1'
b100 +
#634010000000
0!
0'
#634020000000
1!
b101 %
1'
b101 +
#634030000000
1"
1(
#634040000000
0!
0"
b100 &
0'
0(
b100 ,
#634050000000
1!
b110 %
1'
b110 +
#634060000000
0!
0'
#634070000000
1!
b111 %
1'
b111 +
#634080000000
0!
0'
#634090000000
1!
0$
b1000 %
1'
0*
b1000 +
#634100000000
0!
0'
#634110000000
1!
b1001 %
1'
b1001 +
#634120000000
0!
0'
#634130000000
1!
b0 %
1'
b0 +
#634140000000
0!
0'
#634150000000
1!
1$
b1 %
1'
1*
b1 +
#634160000000
0!
0'
#634170000000
1!
b10 %
1'
b10 +
#634180000000
0!
0'
#634190000000
1!
b11 %
1'
b11 +
#634200000000
0!
0'
#634210000000
1!
b100 %
1'
b100 +
#634220000000
0!
0'
#634230000000
1!
b101 %
1'
b101 +
#634240000000
0!
0'
#634250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#634260000000
0!
0'
#634270000000
1!
b111 %
1'
b111 +
#634280000000
0!
0'
#634290000000
1!
b1000 %
1'
b1000 +
#634300000000
0!
0'
#634310000000
1!
b1001 %
1'
b1001 +
#634320000000
0!
0'
#634330000000
1!
b0 %
1'
b0 +
#634340000000
0!
0'
#634350000000
1!
1$
b1 %
1'
1*
b1 +
#634360000000
0!
0'
#634370000000
1!
b10 %
1'
b10 +
#634380000000
0!
0'
#634390000000
1!
b11 %
1'
b11 +
#634400000000
0!
0'
#634410000000
1!
b100 %
1'
b100 +
#634420000000
0!
0'
#634430000000
1!
b101 %
1'
b101 +
#634440000000
0!
0'
#634450000000
1!
0$
b110 %
1'
0*
b110 +
#634460000000
1"
1(
#634470000000
0!
0"
b100 &
0'
0(
b100 ,
#634480000000
1!
1$
b111 %
1'
1*
b111 +
#634490000000
0!
0'
#634500000000
1!
0$
b1000 %
1'
0*
b1000 +
#634510000000
0!
0'
#634520000000
1!
b1001 %
1'
b1001 +
#634530000000
0!
0'
#634540000000
1!
b0 %
1'
b0 +
#634550000000
0!
0'
#634560000000
1!
1$
b1 %
1'
1*
b1 +
#634570000000
0!
0'
#634580000000
1!
b10 %
1'
b10 +
#634590000000
0!
0'
#634600000000
1!
b11 %
1'
b11 +
#634610000000
0!
0'
#634620000000
1!
b100 %
1'
b100 +
#634630000000
0!
0'
#634640000000
1!
b101 %
1'
b101 +
#634650000000
0!
0'
#634660000000
1!
b110 %
1'
b110 +
#634670000000
0!
0'
#634680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#634690000000
0!
0'
#634700000000
1!
b1000 %
1'
b1000 +
#634710000000
0!
0'
#634720000000
1!
b1001 %
1'
b1001 +
#634730000000
0!
0'
#634740000000
1!
b0 %
1'
b0 +
#634750000000
0!
0'
#634760000000
1!
1$
b1 %
1'
1*
b1 +
#634770000000
0!
0'
#634780000000
1!
b10 %
1'
b10 +
#634790000000
0!
0'
#634800000000
1!
b11 %
1'
b11 +
#634810000000
0!
0'
#634820000000
1!
b100 %
1'
b100 +
#634830000000
0!
0'
#634840000000
1!
b101 %
1'
b101 +
#634850000000
0!
0'
#634860000000
1!
0$
b110 %
1'
0*
b110 +
#634870000000
0!
0'
#634880000000
1!
b111 %
1'
b111 +
#634890000000
1"
1(
#634900000000
0!
0"
b100 &
0'
0(
b100 ,
#634910000000
1!
b1000 %
1'
b1000 +
#634920000000
0!
0'
#634930000000
1!
b1001 %
1'
b1001 +
#634940000000
0!
0'
#634950000000
1!
b0 %
1'
b0 +
#634960000000
0!
0'
#634970000000
1!
1$
b1 %
1'
1*
b1 +
#634980000000
0!
0'
#634990000000
1!
b10 %
1'
b10 +
#635000000000
0!
0'
#635010000000
1!
b11 %
1'
b11 +
#635020000000
0!
0'
#635030000000
1!
b100 %
1'
b100 +
#635040000000
0!
0'
#635050000000
1!
b101 %
1'
b101 +
#635060000000
0!
0'
#635070000000
1!
b110 %
1'
b110 +
#635080000000
0!
0'
#635090000000
1!
b111 %
1'
b111 +
#635100000000
0!
0'
#635110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#635120000000
0!
0'
#635130000000
1!
b1001 %
1'
b1001 +
#635140000000
0!
0'
#635150000000
1!
b0 %
1'
b0 +
#635160000000
0!
0'
#635170000000
1!
1$
b1 %
1'
1*
b1 +
#635180000000
0!
0'
#635190000000
1!
b10 %
1'
b10 +
#635200000000
0!
0'
#635210000000
1!
b11 %
1'
b11 +
#635220000000
0!
0'
#635230000000
1!
b100 %
1'
b100 +
#635240000000
0!
0'
#635250000000
1!
b101 %
1'
b101 +
#635260000000
0!
0'
#635270000000
1!
0$
b110 %
1'
0*
b110 +
#635280000000
0!
0'
#635290000000
1!
b111 %
1'
b111 +
#635300000000
0!
0'
#635310000000
1!
b1000 %
1'
b1000 +
#635320000000
1"
1(
#635330000000
0!
0"
b100 &
0'
0(
b100 ,
#635340000000
1!
b1001 %
1'
b1001 +
#635350000000
0!
0'
#635360000000
1!
b0 %
1'
b0 +
#635370000000
0!
0'
#635380000000
1!
1$
b1 %
1'
1*
b1 +
#635390000000
0!
0'
#635400000000
1!
b10 %
1'
b10 +
#635410000000
0!
0'
#635420000000
1!
b11 %
1'
b11 +
#635430000000
0!
0'
#635440000000
1!
b100 %
1'
b100 +
#635450000000
0!
0'
#635460000000
1!
b101 %
1'
b101 +
#635470000000
0!
0'
#635480000000
1!
b110 %
1'
b110 +
#635490000000
0!
0'
#635500000000
1!
b111 %
1'
b111 +
#635510000000
0!
0'
#635520000000
1!
0$
b1000 %
1'
0*
b1000 +
#635530000000
0!
0'
#635540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#635550000000
0!
0'
#635560000000
1!
b0 %
1'
b0 +
#635570000000
0!
0'
#635580000000
1!
1$
b1 %
1'
1*
b1 +
#635590000000
0!
0'
#635600000000
1!
b10 %
1'
b10 +
#635610000000
0!
0'
#635620000000
1!
b11 %
1'
b11 +
#635630000000
0!
0'
#635640000000
1!
b100 %
1'
b100 +
#635650000000
0!
0'
#635660000000
1!
b101 %
1'
b101 +
#635670000000
0!
0'
#635680000000
1!
0$
b110 %
1'
0*
b110 +
#635690000000
0!
0'
#635700000000
1!
b111 %
1'
b111 +
#635710000000
0!
0'
#635720000000
1!
b1000 %
1'
b1000 +
#635730000000
0!
0'
#635740000000
1!
b1001 %
1'
b1001 +
#635750000000
1"
1(
#635760000000
0!
0"
b100 &
0'
0(
b100 ,
#635770000000
1!
b0 %
1'
b0 +
#635780000000
0!
0'
#635790000000
1!
1$
b1 %
1'
1*
b1 +
#635800000000
0!
0'
#635810000000
1!
b10 %
1'
b10 +
#635820000000
0!
0'
#635830000000
1!
b11 %
1'
b11 +
#635840000000
0!
0'
#635850000000
1!
b100 %
1'
b100 +
#635860000000
0!
0'
#635870000000
1!
b101 %
1'
b101 +
#635880000000
0!
0'
#635890000000
1!
b110 %
1'
b110 +
#635900000000
0!
0'
#635910000000
1!
b111 %
1'
b111 +
#635920000000
0!
0'
#635930000000
1!
0$
b1000 %
1'
0*
b1000 +
#635940000000
0!
0'
#635950000000
1!
b1001 %
1'
b1001 +
#635960000000
0!
0'
#635970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#635980000000
0!
0'
#635990000000
1!
1$
b1 %
1'
1*
b1 +
#636000000000
0!
0'
#636010000000
1!
b10 %
1'
b10 +
#636020000000
0!
0'
#636030000000
1!
b11 %
1'
b11 +
#636040000000
0!
0'
#636050000000
1!
b100 %
1'
b100 +
#636060000000
0!
0'
#636070000000
1!
b101 %
1'
b101 +
#636080000000
0!
0'
#636090000000
1!
0$
b110 %
1'
0*
b110 +
#636100000000
0!
0'
#636110000000
1!
b111 %
1'
b111 +
#636120000000
0!
0'
#636130000000
1!
b1000 %
1'
b1000 +
#636140000000
0!
0'
#636150000000
1!
b1001 %
1'
b1001 +
#636160000000
0!
0'
#636170000000
1!
b0 %
1'
b0 +
#636180000000
1"
1(
#636190000000
0!
0"
b100 &
0'
0(
b100 ,
#636200000000
1!
1$
b1 %
1'
1*
b1 +
#636210000000
0!
0'
#636220000000
1!
b10 %
1'
b10 +
#636230000000
0!
0'
#636240000000
1!
b11 %
1'
b11 +
#636250000000
0!
0'
#636260000000
1!
b100 %
1'
b100 +
#636270000000
0!
0'
#636280000000
1!
b101 %
1'
b101 +
#636290000000
0!
0'
#636300000000
1!
b110 %
1'
b110 +
#636310000000
0!
0'
#636320000000
1!
b111 %
1'
b111 +
#636330000000
0!
0'
#636340000000
1!
0$
b1000 %
1'
0*
b1000 +
#636350000000
0!
0'
#636360000000
1!
b1001 %
1'
b1001 +
#636370000000
0!
0'
#636380000000
1!
b0 %
1'
b0 +
#636390000000
0!
0'
#636400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#636410000000
0!
0'
#636420000000
1!
b10 %
1'
b10 +
#636430000000
0!
0'
#636440000000
1!
b11 %
1'
b11 +
#636450000000
0!
0'
#636460000000
1!
b100 %
1'
b100 +
#636470000000
0!
0'
#636480000000
1!
b101 %
1'
b101 +
#636490000000
0!
0'
#636500000000
1!
0$
b110 %
1'
0*
b110 +
#636510000000
0!
0'
#636520000000
1!
b111 %
1'
b111 +
#636530000000
0!
0'
#636540000000
1!
b1000 %
1'
b1000 +
#636550000000
0!
0'
#636560000000
1!
b1001 %
1'
b1001 +
#636570000000
0!
0'
#636580000000
1!
b0 %
1'
b0 +
#636590000000
0!
0'
#636600000000
1!
1$
b1 %
1'
1*
b1 +
#636610000000
1"
1(
#636620000000
0!
0"
b100 &
0'
0(
b100 ,
#636630000000
1!
b10 %
1'
b10 +
#636640000000
0!
0'
#636650000000
1!
b11 %
1'
b11 +
#636660000000
0!
0'
#636670000000
1!
b100 %
1'
b100 +
#636680000000
0!
0'
#636690000000
1!
b101 %
1'
b101 +
#636700000000
0!
0'
#636710000000
1!
b110 %
1'
b110 +
#636720000000
0!
0'
#636730000000
1!
b111 %
1'
b111 +
#636740000000
0!
0'
#636750000000
1!
0$
b1000 %
1'
0*
b1000 +
#636760000000
0!
0'
#636770000000
1!
b1001 %
1'
b1001 +
#636780000000
0!
0'
#636790000000
1!
b0 %
1'
b0 +
#636800000000
0!
0'
#636810000000
1!
1$
b1 %
1'
1*
b1 +
#636820000000
0!
0'
#636830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#636840000000
0!
0'
#636850000000
1!
b11 %
1'
b11 +
#636860000000
0!
0'
#636870000000
1!
b100 %
1'
b100 +
#636880000000
0!
0'
#636890000000
1!
b101 %
1'
b101 +
#636900000000
0!
0'
#636910000000
1!
0$
b110 %
1'
0*
b110 +
#636920000000
0!
0'
#636930000000
1!
b111 %
1'
b111 +
#636940000000
0!
0'
#636950000000
1!
b1000 %
1'
b1000 +
#636960000000
0!
0'
#636970000000
1!
b1001 %
1'
b1001 +
#636980000000
0!
0'
#636990000000
1!
b0 %
1'
b0 +
#637000000000
0!
0'
#637010000000
1!
1$
b1 %
1'
1*
b1 +
#637020000000
0!
0'
#637030000000
1!
b10 %
1'
b10 +
#637040000000
1"
1(
#637050000000
0!
0"
b100 &
0'
0(
b100 ,
#637060000000
1!
b11 %
1'
b11 +
#637070000000
0!
0'
#637080000000
1!
b100 %
1'
b100 +
#637090000000
0!
0'
#637100000000
1!
b101 %
1'
b101 +
#637110000000
0!
0'
#637120000000
1!
b110 %
1'
b110 +
#637130000000
0!
0'
#637140000000
1!
b111 %
1'
b111 +
#637150000000
0!
0'
#637160000000
1!
0$
b1000 %
1'
0*
b1000 +
#637170000000
0!
0'
#637180000000
1!
b1001 %
1'
b1001 +
#637190000000
0!
0'
#637200000000
1!
b0 %
1'
b0 +
#637210000000
0!
0'
#637220000000
1!
1$
b1 %
1'
1*
b1 +
#637230000000
0!
0'
#637240000000
1!
b10 %
1'
b10 +
#637250000000
0!
0'
#637260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#637270000000
0!
0'
#637280000000
1!
b100 %
1'
b100 +
#637290000000
0!
0'
#637300000000
1!
b101 %
1'
b101 +
#637310000000
0!
0'
#637320000000
1!
0$
b110 %
1'
0*
b110 +
#637330000000
0!
0'
#637340000000
1!
b111 %
1'
b111 +
#637350000000
0!
0'
#637360000000
1!
b1000 %
1'
b1000 +
#637370000000
0!
0'
#637380000000
1!
b1001 %
1'
b1001 +
#637390000000
0!
0'
#637400000000
1!
b0 %
1'
b0 +
#637410000000
0!
0'
#637420000000
1!
1$
b1 %
1'
1*
b1 +
#637430000000
0!
0'
#637440000000
1!
b10 %
1'
b10 +
#637450000000
0!
0'
#637460000000
1!
b11 %
1'
b11 +
#637470000000
1"
1(
#637480000000
0!
0"
b100 &
0'
0(
b100 ,
#637490000000
1!
b100 %
1'
b100 +
#637500000000
0!
0'
#637510000000
1!
b101 %
1'
b101 +
#637520000000
0!
0'
#637530000000
1!
b110 %
1'
b110 +
#637540000000
0!
0'
#637550000000
1!
b111 %
1'
b111 +
#637560000000
0!
0'
#637570000000
1!
0$
b1000 %
1'
0*
b1000 +
#637580000000
0!
0'
#637590000000
1!
b1001 %
1'
b1001 +
#637600000000
0!
0'
#637610000000
1!
b0 %
1'
b0 +
#637620000000
0!
0'
#637630000000
1!
1$
b1 %
1'
1*
b1 +
#637640000000
0!
0'
#637650000000
1!
b10 %
1'
b10 +
#637660000000
0!
0'
#637670000000
1!
b11 %
1'
b11 +
#637680000000
0!
0'
#637690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#637700000000
0!
0'
#637710000000
1!
b101 %
1'
b101 +
#637720000000
0!
0'
#637730000000
1!
0$
b110 %
1'
0*
b110 +
#637740000000
0!
0'
#637750000000
1!
b111 %
1'
b111 +
#637760000000
0!
0'
#637770000000
1!
b1000 %
1'
b1000 +
#637780000000
0!
0'
#637790000000
1!
b1001 %
1'
b1001 +
#637800000000
0!
0'
#637810000000
1!
b0 %
1'
b0 +
#637820000000
0!
0'
#637830000000
1!
1$
b1 %
1'
1*
b1 +
#637840000000
0!
0'
#637850000000
1!
b10 %
1'
b10 +
#637860000000
0!
0'
#637870000000
1!
b11 %
1'
b11 +
#637880000000
0!
0'
#637890000000
1!
b100 %
1'
b100 +
#637900000000
1"
1(
#637910000000
0!
0"
b100 &
0'
0(
b100 ,
#637920000000
1!
b101 %
1'
b101 +
#637930000000
0!
0'
#637940000000
1!
b110 %
1'
b110 +
#637950000000
0!
0'
#637960000000
1!
b111 %
1'
b111 +
#637970000000
0!
0'
#637980000000
1!
0$
b1000 %
1'
0*
b1000 +
#637990000000
0!
0'
#638000000000
1!
b1001 %
1'
b1001 +
#638010000000
0!
0'
#638020000000
1!
b0 %
1'
b0 +
#638030000000
0!
0'
#638040000000
1!
1$
b1 %
1'
1*
b1 +
#638050000000
0!
0'
#638060000000
1!
b10 %
1'
b10 +
#638070000000
0!
0'
#638080000000
1!
b11 %
1'
b11 +
#638090000000
0!
0'
#638100000000
1!
b100 %
1'
b100 +
#638110000000
0!
0'
#638120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#638130000000
0!
0'
#638140000000
1!
0$
b110 %
1'
0*
b110 +
#638150000000
0!
0'
#638160000000
1!
b111 %
1'
b111 +
#638170000000
0!
0'
#638180000000
1!
b1000 %
1'
b1000 +
#638190000000
0!
0'
#638200000000
1!
b1001 %
1'
b1001 +
#638210000000
0!
0'
#638220000000
1!
b0 %
1'
b0 +
#638230000000
0!
0'
#638240000000
1!
1$
b1 %
1'
1*
b1 +
#638250000000
0!
0'
#638260000000
1!
b10 %
1'
b10 +
#638270000000
0!
0'
#638280000000
1!
b11 %
1'
b11 +
#638290000000
0!
0'
#638300000000
1!
b100 %
1'
b100 +
#638310000000
0!
0'
#638320000000
1!
b101 %
1'
b101 +
#638330000000
1"
1(
#638340000000
0!
0"
b100 &
0'
0(
b100 ,
#638350000000
1!
b110 %
1'
b110 +
#638360000000
0!
0'
#638370000000
1!
b111 %
1'
b111 +
#638380000000
0!
0'
#638390000000
1!
0$
b1000 %
1'
0*
b1000 +
#638400000000
0!
0'
#638410000000
1!
b1001 %
1'
b1001 +
#638420000000
0!
0'
#638430000000
1!
b0 %
1'
b0 +
#638440000000
0!
0'
#638450000000
1!
1$
b1 %
1'
1*
b1 +
#638460000000
0!
0'
#638470000000
1!
b10 %
1'
b10 +
#638480000000
0!
0'
#638490000000
1!
b11 %
1'
b11 +
#638500000000
0!
0'
#638510000000
1!
b100 %
1'
b100 +
#638520000000
0!
0'
#638530000000
1!
b101 %
1'
b101 +
#638540000000
0!
0'
#638550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#638560000000
0!
0'
#638570000000
1!
b111 %
1'
b111 +
#638580000000
0!
0'
#638590000000
1!
b1000 %
1'
b1000 +
#638600000000
0!
0'
#638610000000
1!
b1001 %
1'
b1001 +
#638620000000
0!
0'
#638630000000
1!
b0 %
1'
b0 +
#638640000000
0!
0'
#638650000000
1!
1$
b1 %
1'
1*
b1 +
#638660000000
0!
0'
#638670000000
1!
b10 %
1'
b10 +
#638680000000
0!
0'
#638690000000
1!
b11 %
1'
b11 +
#638700000000
0!
0'
#638710000000
1!
b100 %
1'
b100 +
#638720000000
0!
0'
#638730000000
1!
b101 %
1'
b101 +
#638740000000
0!
0'
#638750000000
1!
0$
b110 %
1'
0*
b110 +
#638760000000
1"
1(
#638770000000
0!
0"
b100 &
0'
0(
b100 ,
#638780000000
1!
1$
b111 %
1'
1*
b111 +
#638790000000
0!
0'
#638800000000
1!
0$
b1000 %
1'
0*
b1000 +
#638810000000
0!
0'
#638820000000
1!
b1001 %
1'
b1001 +
#638830000000
0!
0'
#638840000000
1!
b0 %
1'
b0 +
#638850000000
0!
0'
#638860000000
1!
1$
b1 %
1'
1*
b1 +
#638870000000
0!
0'
#638880000000
1!
b10 %
1'
b10 +
#638890000000
0!
0'
#638900000000
1!
b11 %
1'
b11 +
#638910000000
0!
0'
#638920000000
1!
b100 %
1'
b100 +
#638930000000
0!
0'
#638940000000
1!
b101 %
1'
b101 +
#638950000000
0!
0'
#638960000000
1!
b110 %
1'
b110 +
#638970000000
0!
0'
#638980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#638990000000
0!
0'
#639000000000
1!
b1000 %
1'
b1000 +
#639010000000
0!
0'
#639020000000
1!
b1001 %
1'
b1001 +
#639030000000
0!
0'
#639040000000
1!
b0 %
1'
b0 +
#639050000000
0!
0'
#639060000000
1!
1$
b1 %
1'
1*
b1 +
#639070000000
0!
0'
#639080000000
1!
b10 %
1'
b10 +
#639090000000
0!
0'
#639100000000
1!
b11 %
1'
b11 +
#639110000000
0!
0'
#639120000000
1!
b100 %
1'
b100 +
#639130000000
0!
0'
#639140000000
1!
b101 %
1'
b101 +
#639150000000
0!
0'
#639160000000
1!
0$
b110 %
1'
0*
b110 +
#639170000000
0!
0'
#639180000000
1!
b111 %
1'
b111 +
#639190000000
1"
1(
#639200000000
0!
0"
b100 &
0'
0(
b100 ,
#639210000000
1!
b1000 %
1'
b1000 +
#639220000000
0!
0'
#639230000000
1!
b1001 %
1'
b1001 +
#639240000000
0!
0'
#639250000000
1!
b0 %
1'
b0 +
#639260000000
0!
0'
#639270000000
1!
1$
b1 %
1'
1*
b1 +
#639280000000
0!
0'
#639290000000
1!
b10 %
1'
b10 +
#639300000000
0!
0'
#639310000000
1!
b11 %
1'
b11 +
#639320000000
0!
0'
#639330000000
1!
b100 %
1'
b100 +
#639340000000
0!
0'
#639350000000
1!
b101 %
1'
b101 +
#639360000000
0!
0'
#639370000000
1!
b110 %
1'
b110 +
#639380000000
0!
0'
#639390000000
1!
b111 %
1'
b111 +
#639400000000
0!
0'
#639410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#639420000000
0!
0'
#639430000000
1!
b1001 %
1'
b1001 +
#639440000000
0!
0'
#639450000000
1!
b0 %
1'
b0 +
#639460000000
0!
0'
#639470000000
1!
1$
b1 %
1'
1*
b1 +
#639480000000
0!
0'
#639490000000
1!
b10 %
1'
b10 +
#639500000000
0!
0'
#639510000000
1!
b11 %
1'
b11 +
#639520000000
0!
0'
#639530000000
1!
b100 %
1'
b100 +
#639540000000
0!
0'
#639550000000
1!
b101 %
1'
b101 +
#639560000000
0!
0'
#639570000000
1!
0$
b110 %
1'
0*
b110 +
#639580000000
0!
0'
#639590000000
1!
b111 %
1'
b111 +
#639600000000
0!
0'
#639610000000
1!
b1000 %
1'
b1000 +
#639620000000
1"
1(
#639630000000
0!
0"
b100 &
0'
0(
b100 ,
#639640000000
1!
b1001 %
1'
b1001 +
#639650000000
0!
0'
#639660000000
1!
b0 %
1'
b0 +
#639670000000
0!
0'
#639680000000
1!
1$
b1 %
1'
1*
b1 +
#639690000000
0!
0'
#639700000000
1!
b10 %
1'
b10 +
#639710000000
0!
0'
#639720000000
1!
b11 %
1'
b11 +
#639730000000
0!
0'
#639740000000
1!
b100 %
1'
b100 +
#639750000000
0!
0'
#639760000000
1!
b101 %
1'
b101 +
#639770000000
0!
0'
#639780000000
1!
b110 %
1'
b110 +
#639790000000
0!
0'
#639800000000
1!
b111 %
1'
b111 +
#639810000000
0!
0'
#639820000000
1!
0$
b1000 %
1'
0*
b1000 +
#639830000000
0!
0'
#639840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#639850000000
0!
0'
#639860000000
1!
b0 %
1'
b0 +
#639870000000
0!
0'
#639880000000
1!
1$
b1 %
1'
1*
b1 +
#639890000000
0!
0'
#639900000000
1!
b10 %
1'
b10 +
#639910000000
0!
0'
#639920000000
1!
b11 %
1'
b11 +
#639930000000
0!
0'
#639940000000
1!
b100 %
1'
b100 +
#639950000000
0!
0'
#639960000000
1!
b101 %
1'
b101 +
#639970000000
0!
0'
#639980000000
1!
0$
b110 %
1'
0*
b110 +
#639990000000
0!
0'
#640000000000
1!
b111 %
1'
b111 +
#640010000000
0!
0'
#640020000000
1!
b1000 %
1'
b1000 +
#640030000000
0!
0'
#640040000000
1!
b1001 %
1'
b1001 +
#640050000000
1"
1(
#640060000000
0!
0"
b100 &
0'
0(
b100 ,
#640070000000
1!
b0 %
1'
b0 +
#640080000000
0!
0'
#640090000000
1!
1$
b1 %
1'
1*
b1 +
#640100000000
0!
0'
#640110000000
1!
b10 %
1'
b10 +
#640120000000
0!
0'
#640130000000
1!
b11 %
1'
b11 +
#640140000000
0!
0'
#640150000000
1!
b100 %
1'
b100 +
#640160000000
0!
0'
#640170000000
1!
b101 %
1'
b101 +
#640180000000
0!
0'
#640190000000
1!
b110 %
1'
b110 +
#640200000000
0!
0'
#640210000000
1!
b111 %
1'
b111 +
#640220000000
0!
0'
#640230000000
1!
0$
b1000 %
1'
0*
b1000 +
#640240000000
0!
0'
#640250000000
1!
b1001 %
1'
b1001 +
#640260000000
0!
0'
#640270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#640280000000
0!
0'
#640290000000
1!
1$
b1 %
1'
1*
b1 +
#640300000000
0!
0'
#640310000000
1!
b10 %
1'
b10 +
#640320000000
0!
0'
#640330000000
1!
b11 %
1'
b11 +
#640340000000
0!
0'
#640350000000
1!
b100 %
1'
b100 +
#640360000000
0!
0'
#640370000000
1!
b101 %
1'
b101 +
#640380000000
0!
0'
#640390000000
1!
0$
b110 %
1'
0*
b110 +
#640400000000
0!
0'
#640410000000
1!
b111 %
1'
b111 +
#640420000000
0!
0'
#640430000000
1!
b1000 %
1'
b1000 +
#640440000000
0!
0'
#640450000000
1!
b1001 %
1'
b1001 +
#640460000000
0!
0'
#640470000000
1!
b0 %
1'
b0 +
#640480000000
1"
1(
#640490000000
0!
0"
b100 &
0'
0(
b100 ,
#640500000000
1!
1$
b1 %
1'
1*
b1 +
#640510000000
0!
0'
#640520000000
1!
b10 %
1'
b10 +
#640530000000
0!
0'
#640540000000
1!
b11 %
1'
b11 +
#640550000000
0!
0'
#640560000000
1!
b100 %
1'
b100 +
#640570000000
0!
0'
#640580000000
1!
b101 %
1'
b101 +
#640590000000
0!
0'
#640600000000
1!
b110 %
1'
b110 +
#640610000000
0!
0'
#640620000000
1!
b111 %
1'
b111 +
#640630000000
0!
0'
#640640000000
1!
0$
b1000 %
1'
0*
b1000 +
#640650000000
0!
0'
#640660000000
1!
b1001 %
1'
b1001 +
#640670000000
0!
0'
#640680000000
1!
b0 %
1'
b0 +
#640690000000
0!
0'
#640700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#640710000000
0!
0'
#640720000000
1!
b10 %
1'
b10 +
#640730000000
0!
0'
#640740000000
1!
b11 %
1'
b11 +
#640750000000
0!
0'
#640760000000
1!
b100 %
1'
b100 +
#640770000000
0!
0'
#640780000000
1!
b101 %
1'
b101 +
#640790000000
0!
0'
#640800000000
1!
0$
b110 %
1'
0*
b110 +
#640810000000
0!
0'
#640820000000
1!
b111 %
1'
b111 +
#640830000000
0!
0'
#640840000000
1!
b1000 %
1'
b1000 +
#640850000000
0!
0'
#640860000000
1!
b1001 %
1'
b1001 +
#640870000000
0!
0'
#640880000000
1!
b0 %
1'
b0 +
#640890000000
0!
0'
#640900000000
1!
1$
b1 %
1'
1*
b1 +
#640910000000
1"
1(
#640920000000
0!
0"
b100 &
0'
0(
b100 ,
#640930000000
1!
b10 %
1'
b10 +
#640940000000
0!
0'
#640950000000
1!
b11 %
1'
b11 +
#640960000000
0!
0'
#640970000000
1!
b100 %
1'
b100 +
#640980000000
0!
0'
#640990000000
1!
b101 %
1'
b101 +
#641000000000
0!
0'
#641010000000
1!
b110 %
1'
b110 +
#641020000000
0!
0'
#641030000000
1!
b111 %
1'
b111 +
#641040000000
0!
0'
#641050000000
1!
0$
b1000 %
1'
0*
b1000 +
#641060000000
0!
0'
#641070000000
1!
b1001 %
1'
b1001 +
#641080000000
0!
0'
#641090000000
1!
b0 %
1'
b0 +
#641100000000
0!
0'
#641110000000
1!
1$
b1 %
1'
1*
b1 +
#641120000000
0!
0'
#641130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#641140000000
0!
0'
#641150000000
1!
b11 %
1'
b11 +
#641160000000
0!
0'
#641170000000
1!
b100 %
1'
b100 +
#641180000000
0!
0'
#641190000000
1!
b101 %
1'
b101 +
#641200000000
0!
0'
#641210000000
1!
0$
b110 %
1'
0*
b110 +
#641220000000
0!
0'
#641230000000
1!
b111 %
1'
b111 +
#641240000000
0!
0'
#641250000000
1!
b1000 %
1'
b1000 +
#641260000000
0!
0'
#641270000000
1!
b1001 %
1'
b1001 +
#641280000000
0!
0'
#641290000000
1!
b0 %
1'
b0 +
#641300000000
0!
0'
#641310000000
1!
1$
b1 %
1'
1*
b1 +
#641320000000
0!
0'
#641330000000
1!
b10 %
1'
b10 +
#641340000000
1"
1(
#641350000000
0!
0"
b100 &
0'
0(
b100 ,
#641360000000
1!
b11 %
1'
b11 +
#641370000000
0!
0'
#641380000000
1!
b100 %
1'
b100 +
#641390000000
0!
0'
#641400000000
1!
b101 %
1'
b101 +
#641410000000
0!
0'
#641420000000
1!
b110 %
1'
b110 +
#641430000000
0!
0'
#641440000000
1!
b111 %
1'
b111 +
#641450000000
0!
0'
#641460000000
1!
0$
b1000 %
1'
0*
b1000 +
#641470000000
0!
0'
#641480000000
1!
b1001 %
1'
b1001 +
#641490000000
0!
0'
#641500000000
1!
b0 %
1'
b0 +
#641510000000
0!
0'
#641520000000
1!
1$
b1 %
1'
1*
b1 +
#641530000000
0!
0'
#641540000000
1!
b10 %
1'
b10 +
#641550000000
0!
0'
#641560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#641570000000
0!
0'
#641580000000
1!
b100 %
1'
b100 +
#641590000000
0!
0'
#641600000000
1!
b101 %
1'
b101 +
#641610000000
0!
0'
#641620000000
1!
0$
b110 %
1'
0*
b110 +
#641630000000
0!
0'
#641640000000
1!
b111 %
1'
b111 +
#641650000000
0!
0'
#641660000000
1!
b1000 %
1'
b1000 +
#641670000000
0!
0'
#641680000000
1!
b1001 %
1'
b1001 +
#641690000000
0!
0'
#641700000000
1!
b0 %
1'
b0 +
#641710000000
0!
0'
#641720000000
1!
1$
b1 %
1'
1*
b1 +
#641730000000
0!
0'
#641740000000
1!
b10 %
1'
b10 +
#641750000000
0!
0'
#641760000000
1!
b11 %
1'
b11 +
#641770000000
1"
1(
#641780000000
0!
0"
b100 &
0'
0(
b100 ,
#641790000000
1!
b100 %
1'
b100 +
#641800000000
0!
0'
#641810000000
1!
b101 %
1'
b101 +
#641820000000
0!
0'
#641830000000
1!
b110 %
1'
b110 +
#641840000000
0!
0'
#641850000000
1!
b111 %
1'
b111 +
#641860000000
0!
0'
#641870000000
1!
0$
b1000 %
1'
0*
b1000 +
#641880000000
0!
0'
#641890000000
1!
b1001 %
1'
b1001 +
#641900000000
0!
0'
#641910000000
1!
b0 %
1'
b0 +
#641920000000
0!
0'
#641930000000
1!
1$
b1 %
1'
1*
b1 +
#641940000000
0!
0'
#641950000000
1!
b10 %
1'
b10 +
#641960000000
0!
0'
#641970000000
1!
b11 %
1'
b11 +
#641980000000
0!
0'
#641990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#642000000000
0!
0'
#642010000000
1!
b101 %
1'
b101 +
#642020000000
0!
0'
#642030000000
1!
0$
b110 %
1'
0*
b110 +
#642040000000
0!
0'
#642050000000
1!
b111 %
1'
b111 +
#642060000000
0!
0'
#642070000000
1!
b1000 %
1'
b1000 +
#642080000000
0!
0'
#642090000000
1!
b1001 %
1'
b1001 +
#642100000000
0!
0'
#642110000000
1!
b0 %
1'
b0 +
#642120000000
0!
0'
#642130000000
1!
1$
b1 %
1'
1*
b1 +
#642140000000
0!
0'
#642150000000
1!
b10 %
1'
b10 +
#642160000000
0!
0'
#642170000000
1!
b11 %
1'
b11 +
#642180000000
0!
0'
#642190000000
1!
b100 %
1'
b100 +
#642200000000
1"
1(
#642210000000
0!
0"
b100 &
0'
0(
b100 ,
#642220000000
1!
b101 %
1'
b101 +
#642230000000
0!
0'
#642240000000
1!
b110 %
1'
b110 +
#642250000000
0!
0'
#642260000000
1!
b111 %
1'
b111 +
#642270000000
0!
0'
#642280000000
1!
0$
b1000 %
1'
0*
b1000 +
#642290000000
0!
0'
#642300000000
1!
b1001 %
1'
b1001 +
#642310000000
0!
0'
#642320000000
1!
b0 %
1'
b0 +
#642330000000
0!
0'
#642340000000
1!
1$
b1 %
1'
1*
b1 +
#642350000000
0!
0'
#642360000000
1!
b10 %
1'
b10 +
#642370000000
0!
0'
#642380000000
1!
b11 %
1'
b11 +
#642390000000
0!
0'
#642400000000
1!
b100 %
1'
b100 +
#642410000000
0!
0'
#642420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#642430000000
0!
0'
#642440000000
1!
0$
b110 %
1'
0*
b110 +
#642450000000
0!
0'
#642460000000
1!
b111 %
1'
b111 +
#642470000000
0!
0'
#642480000000
1!
b1000 %
1'
b1000 +
#642490000000
0!
0'
#642500000000
1!
b1001 %
1'
b1001 +
#642510000000
0!
0'
#642520000000
1!
b0 %
1'
b0 +
#642530000000
0!
0'
#642540000000
1!
1$
b1 %
1'
1*
b1 +
#642550000000
0!
0'
#642560000000
1!
b10 %
1'
b10 +
#642570000000
0!
0'
#642580000000
1!
b11 %
1'
b11 +
#642590000000
0!
0'
#642600000000
1!
b100 %
1'
b100 +
#642610000000
0!
0'
#642620000000
1!
b101 %
1'
b101 +
#642630000000
1"
1(
#642640000000
0!
0"
b100 &
0'
0(
b100 ,
#642650000000
1!
b110 %
1'
b110 +
#642660000000
0!
0'
#642670000000
1!
b111 %
1'
b111 +
#642680000000
0!
0'
#642690000000
1!
0$
b1000 %
1'
0*
b1000 +
#642700000000
0!
0'
#642710000000
1!
b1001 %
1'
b1001 +
#642720000000
0!
0'
#642730000000
1!
b0 %
1'
b0 +
#642740000000
0!
0'
#642750000000
1!
1$
b1 %
1'
1*
b1 +
#642760000000
0!
0'
#642770000000
1!
b10 %
1'
b10 +
#642780000000
0!
0'
#642790000000
1!
b11 %
1'
b11 +
#642800000000
0!
0'
#642810000000
1!
b100 %
1'
b100 +
#642820000000
0!
0'
#642830000000
1!
b101 %
1'
b101 +
#642840000000
0!
0'
#642850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#642860000000
0!
0'
#642870000000
1!
b111 %
1'
b111 +
#642880000000
0!
0'
#642890000000
1!
b1000 %
1'
b1000 +
#642900000000
0!
0'
#642910000000
1!
b1001 %
1'
b1001 +
#642920000000
0!
0'
#642930000000
1!
b0 %
1'
b0 +
#642940000000
0!
0'
#642950000000
1!
1$
b1 %
1'
1*
b1 +
#642960000000
0!
0'
#642970000000
1!
b10 %
1'
b10 +
#642980000000
0!
0'
#642990000000
1!
b11 %
1'
b11 +
#643000000000
0!
0'
#643010000000
1!
b100 %
1'
b100 +
#643020000000
0!
0'
#643030000000
1!
b101 %
1'
b101 +
#643040000000
0!
0'
#643050000000
1!
0$
b110 %
1'
0*
b110 +
#643060000000
1"
1(
#643070000000
0!
0"
b100 &
0'
0(
b100 ,
#643080000000
1!
1$
b111 %
1'
1*
b111 +
#643090000000
0!
0'
#643100000000
1!
0$
b1000 %
1'
0*
b1000 +
#643110000000
0!
0'
#643120000000
1!
b1001 %
1'
b1001 +
#643130000000
0!
0'
#643140000000
1!
b0 %
1'
b0 +
#643150000000
0!
0'
#643160000000
1!
1$
b1 %
1'
1*
b1 +
#643170000000
0!
0'
#643180000000
1!
b10 %
1'
b10 +
#643190000000
0!
0'
#643200000000
1!
b11 %
1'
b11 +
#643210000000
0!
0'
#643220000000
1!
b100 %
1'
b100 +
#643230000000
0!
0'
#643240000000
1!
b101 %
1'
b101 +
#643250000000
0!
0'
#643260000000
1!
b110 %
1'
b110 +
#643270000000
0!
0'
#643280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#643290000000
0!
0'
#643300000000
1!
b1000 %
1'
b1000 +
#643310000000
0!
0'
#643320000000
1!
b1001 %
1'
b1001 +
#643330000000
0!
0'
#643340000000
1!
b0 %
1'
b0 +
#643350000000
0!
0'
#643360000000
1!
1$
b1 %
1'
1*
b1 +
#643370000000
0!
0'
#643380000000
1!
b10 %
1'
b10 +
#643390000000
0!
0'
#643400000000
1!
b11 %
1'
b11 +
#643410000000
0!
0'
#643420000000
1!
b100 %
1'
b100 +
#643430000000
0!
0'
#643440000000
1!
b101 %
1'
b101 +
#643450000000
0!
0'
#643460000000
1!
0$
b110 %
1'
0*
b110 +
#643470000000
0!
0'
#643480000000
1!
b111 %
1'
b111 +
#643490000000
1"
1(
#643500000000
0!
0"
b100 &
0'
0(
b100 ,
#643510000000
1!
b1000 %
1'
b1000 +
#643520000000
0!
0'
#643530000000
1!
b1001 %
1'
b1001 +
#643540000000
0!
0'
#643550000000
1!
b0 %
1'
b0 +
#643560000000
0!
0'
#643570000000
1!
1$
b1 %
1'
1*
b1 +
#643580000000
0!
0'
#643590000000
1!
b10 %
1'
b10 +
#643600000000
0!
0'
#643610000000
1!
b11 %
1'
b11 +
#643620000000
0!
0'
#643630000000
1!
b100 %
1'
b100 +
#643640000000
0!
0'
#643650000000
1!
b101 %
1'
b101 +
#643660000000
0!
0'
#643670000000
1!
b110 %
1'
b110 +
#643680000000
0!
0'
#643690000000
1!
b111 %
1'
b111 +
#643700000000
0!
0'
#643710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#643720000000
0!
0'
#643730000000
1!
b1001 %
1'
b1001 +
#643740000000
0!
0'
#643750000000
1!
b0 %
1'
b0 +
#643760000000
0!
0'
#643770000000
1!
1$
b1 %
1'
1*
b1 +
#643780000000
0!
0'
#643790000000
1!
b10 %
1'
b10 +
#643800000000
0!
0'
#643810000000
1!
b11 %
1'
b11 +
#643820000000
0!
0'
#643830000000
1!
b100 %
1'
b100 +
#643840000000
0!
0'
#643850000000
1!
b101 %
1'
b101 +
#643860000000
0!
0'
#643870000000
1!
0$
b110 %
1'
0*
b110 +
#643880000000
0!
0'
#643890000000
1!
b111 %
1'
b111 +
#643900000000
0!
0'
#643910000000
1!
b1000 %
1'
b1000 +
#643920000000
1"
1(
#643930000000
0!
0"
b100 &
0'
0(
b100 ,
#643940000000
1!
b1001 %
1'
b1001 +
#643950000000
0!
0'
#643960000000
1!
b0 %
1'
b0 +
#643970000000
0!
0'
#643980000000
1!
1$
b1 %
1'
1*
b1 +
#643990000000
0!
0'
#644000000000
1!
b10 %
1'
b10 +
#644010000000
0!
0'
#644020000000
1!
b11 %
1'
b11 +
#644030000000
0!
0'
#644040000000
1!
b100 %
1'
b100 +
#644050000000
0!
0'
#644060000000
1!
b101 %
1'
b101 +
#644070000000
0!
0'
#644080000000
1!
b110 %
1'
b110 +
#644090000000
0!
0'
#644100000000
1!
b111 %
1'
b111 +
#644110000000
0!
0'
#644120000000
1!
0$
b1000 %
1'
0*
b1000 +
#644130000000
0!
0'
#644140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#644150000000
0!
0'
#644160000000
1!
b0 %
1'
b0 +
#644170000000
0!
0'
#644180000000
1!
1$
b1 %
1'
1*
b1 +
#644190000000
0!
0'
#644200000000
1!
b10 %
1'
b10 +
#644210000000
0!
0'
#644220000000
1!
b11 %
1'
b11 +
#644230000000
0!
0'
#644240000000
1!
b100 %
1'
b100 +
#644250000000
0!
0'
#644260000000
1!
b101 %
1'
b101 +
#644270000000
0!
0'
#644280000000
1!
0$
b110 %
1'
0*
b110 +
#644290000000
0!
0'
#644300000000
1!
b111 %
1'
b111 +
#644310000000
0!
0'
#644320000000
1!
b1000 %
1'
b1000 +
#644330000000
0!
0'
#644340000000
1!
b1001 %
1'
b1001 +
#644350000000
1"
1(
#644360000000
0!
0"
b100 &
0'
0(
b100 ,
#644370000000
1!
b0 %
1'
b0 +
#644380000000
0!
0'
#644390000000
1!
1$
b1 %
1'
1*
b1 +
#644400000000
0!
0'
#644410000000
1!
b10 %
1'
b10 +
#644420000000
0!
0'
#644430000000
1!
b11 %
1'
b11 +
#644440000000
0!
0'
#644450000000
1!
b100 %
1'
b100 +
#644460000000
0!
0'
#644470000000
1!
b101 %
1'
b101 +
#644480000000
0!
0'
#644490000000
1!
b110 %
1'
b110 +
#644500000000
0!
0'
#644510000000
1!
b111 %
1'
b111 +
#644520000000
0!
0'
#644530000000
1!
0$
b1000 %
1'
0*
b1000 +
#644540000000
0!
0'
#644550000000
1!
b1001 %
1'
b1001 +
#644560000000
0!
0'
#644570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#644580000000
0!
0'
#644590000000
1!
1$
b1 %
1'
1*
b1 +
#644600000000
0!
0'
#644610000000
1!
b10 %
1'
b10 +
#644620000000
0!
0'
#644630000000
1!
b11 %
1'
b11 +
#644640000000
0!
0'
#644650000000
1!
b100 %
1'
b100 +
#644660000000
0!
0'
#644670000000
1!
b101 %
1'
b101 +
#644680000000
0!
0'
#644690000000
1!
0$
b110 %
1'
0*
b110 +
#644700000000
0!
0'
#644710000000
1!
b111 %
1'
b111 +
#644720000000
0!
0'
#644730000000
1!
b1000 %
1'
b1000 +
#644740000000
0!
0'
#644750000000
1!
b1001 %
1'
b1001 +
#644760000000
0!
0'
#644770000000
1!
b0 %
1'
b0 +
#644780000000
1"
1(
#644790000000
0!
0"
b100 &
0'
0(
b100 ,
#644800000000
1!
1$
b1 %
1'
1*
b1 +
#644810000000
0!
0'
#644820000000
1!
b10 %
1'
b10 +
#644830000000
0!
0'
#644840000000
1!
b11 %
1'
b11 +
#644850000000
0!
0'
#644860000000
1!
b100 %
1'
b100 +
#644870000000
0!
0'
#644880000000
1!
b101 %
1'
b101 +
#644890000000
0!
0'
#644900000000
1!
b110 %
1'
b110 +
#644910000000
0!
0'
#644920000000
1!
b111 %
1'
b111 +
#644930000000
0!
0'
#644940000000
1!
0$
b1000 %
1'
0*
b1000 +
#644950000000
0!
0'
#644960000000
1!
b1001 %
1'
b1001 +
#644970000000
0!
0'
#644980000000
1!
b0 %
1'
b0 +
#644990000000
0!
0'
#645000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#645010000000
0!
0'
#645020000000
1!
b10 %
1'
b10 +
#645030000000
0!
0'
#645040000000
1!
b11 %
1'
b11 +
#645050000000
0!
0'
#645060000000
1!
b100 %
1'
b100 +
#645070000000
0!
0'
#645080000000
1!
b101 %
1'
b101 +
#645090000000
0!
0'
#645100000000
1!
0$
b110 %
1'
0*
b110 +
#645110000000
0!
0'
#645120000000
1!
b111 %
1'
b111 +
#645130000000
0!
0'
#645140000000
1!
b1000 %
1'
b1000 +
#645150000000
0!
0'
#645160000000
1!
b1001 %
1'
b1001 +
#645170000000
0!
0'
#645180000000
1!
b0 %
1'
b0 +
#645190000000
0!
0'
#645200000000
1!
1$
b1 %
1'
1*
b1 +
#645210000000
1"
1(
#645220000000
0!
0"
b100 &
0'
0(
b100 ,
#645230000000
1!
b10 %
1'
b10 +
#645240000000
0!
0'
#645250000000
1!
b11 %
1'
b11 +
#645260000000
0!
0'
#645270000000
1!
b100 %
1'
b100 +
#645280000000
0!
0'
#645290000000
1!
b101 %
1'
b101 +
#645300000000
0!
0'
#645310000000
1!
b110 %
1'
b110 +
#645320000000
0!
0'
#645330000000
1!
b111 %
1'
b111 +
#645340000000
0!
0'
#645350000000
1!
0$
b1000 %
1'
0*
b1000 +
#645360000000
0!
0'
#645370000000
1!
b1001 %
1'
b1001 +
#645380000000
0!
0'
#645390000000
1!
b0 %
1'
b0 +
#645400000000
0!
0'
#645410000000
1!
1$
b1 %
1'
1*
b1 +
#645420000000
0!
0'
#645430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#645440000000
0!
0'
#645450000000
1!
b11 %
1'
b11 +
#645460000000
0!
0'
#645470000000
1!
b100 %
1'
b100 +
#645480000000
0!
0'
#645490000000
1!
b101 %
1'
b101 +
#645500000000
0!
0'
#645510000000
1!
0$
b110 %
1'
0*
b110 +
#645520000000
0!
0'
#645530000000
1!
b111 %
1'
b111 +
#645540000000
0!
0'
#645550000000
1!
b1000 %
1'
b1000 +
#645560000000
0!
0'
#645570000000
1!
b1001 %
1'
b1001 +
#645580000000
0!
0'
#645590000000
1!
b0 %
1'
b0 +
#645600000000
0!
0'
#645610000000
1!
1$
b1 %
1'
1*
b1 +
#645620000000
0!
0'
#645630000000
1!
b10 %
1'
b10 +
#645640000000
1"
1(
#645650000000
0!
0"
b100 &
0'
0(
b100 ,
#645660000000
1!
b11 %
1'
b11 +
#645670000000
0!
0'
#645680000000
1!
b100 %
1'
b100 +
#645690000000
0!
0'
#645700000000
1!
b101 %
1'
b101 +
#645710000000
0!
0'
#645720000000
1!
b110 %
1'
b110 +
#645730000000
0!
0'
#645740000000
1!
b111 %
1'
b111 +
#645750000000
0!
0'
#645760000000
1!
0$
b1000 %
1'
0*
b1000 +
#645770000000
0!
0'
#645780000000
1!
b1001 %
1'
b1001 +
#645790000000
0!
0'
#645800000000
1!
b0 %
1'
b0 +
#645810000000
0!
0'
#645820000000
1!
1$
b1 %
1'
1*
b1 +
#645830000000
0!
0'
#645840000000
1!
b10 %
1'
b10 +
#645850000000
0!
0'
#645860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#645870000000
0!
0'
#645880000000
1!
b100 %
1'
b100 +
#645890000000
0!
0'
#645900000000
1!
b101 %
1'
b101 +
#645910000000
0!
0'
#645920000000
1!
0$
b110 %
1'
0*
b110 +
#645930000000
0!
0'
#645940000000
1!
b111 %
1'
b111 +
#645950000000
0!
0'
#645960000000
1!
b1000 %
1'
b1000 +
#645970000000
0!
0'
#645980000000
1!
b1001 %
1'
b1001 +
#645990000000
0!
0'
#646000000000
1!
b0 %
1'
b0 +
#646010000000
0!
0'
#646020000000
1!
1$
b1 %
1'
1*
b1 +
#646030000000
0!
0'
#646040000000
1!
b10 %
1'
b10 +
#646050000000
0!
0'
#646060000000
1!
b11 %
1'
b11 +
#646070000000
1"
1(
#646080000000
0!
0"
b100 &
0'
0(
b100 ,
#646090000000
1!
b100 %
1'
b100 +
#646100000000
0!
0'
#646110000000
1!
b101 %
1'
b101 +
#646120000000
0!
0'
#646130000000
1!
b110 %
1'
b110 +
#646140000000
0!
0'
#646150000000
1!
b111 %
1'
b111 +
#646160000000
0!
0'
#646170000000
1!
0$
b1000 %
1'
0*
b1000 +
#646180000000
0!
0'
#646190000000
1!
b1001 %
1'
b1001 +
#646200000000
0!
0'
#646210000000
1!
b0 %
1'
b0 +
#646220000000
0!
0'
#646230000000
1!
1$
b1 %
1'
1*
b1 +
#646240000000
0!
0'
#646250000000
1!
b10 %
1'
b10 +
#646260000000
0!
0'
#646270000000
1!
b11 %
1'
b11 +
#646280000000
0!
0'
#646290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#646300000000
0!
0'
#646310000000
1!
b101 %
1'
b101 +
#646320000000
0!
0'
#646330000000
1!
0$
b110 %
1'
0*
b110 +
#646340000000
0!
0'
#646350000000
1!
b111 %
1'
b111 +
#646360000000
0!
0'
#646370000000
1!
b1000 %
1'
b1000 +
#646380000000
0!
0'
#646390000000
1!
b1001 %
1'
b1001 +
#646400000000
0!
0'
#646410000000
1!
b0 %
1'
b0 +
#646420000000
0!
0'
#646430000000
1!
1$
b1 %
1'
1*
b1 +
#646440000000
0!
0'
#646450000000
1!
b10 %
1'
b10 +
#646460000000
0!
0'
#646470000000
1!
b11 %
1'
b11 +
#646480000000
0!
0'
#646490000000
1!
b100 %
1'
b100 +
#646500000000
1"
1(
#646510000000
0!
0"
b100 &
0'
0(
b100 ,
#646520000000
1!
b101 %
1'
b101 +
#646530000000
0!
0'
#646540000000
1!
b110 %
1'
b110 +
#646550000000
0!
0'
#646560000000
1!
b111 %
1'
b111 +
#646570000000
0!
0'
#646580000000
1!
0$
b1000 %
1'
0*
b1000 +
#646590000000
0!
0'
#646600000000
1!
b1001 %
1'
b1001 +
#646610000000
0!
0'
#646620000000
1!
b0 %
1'
b0 +
#646630000000
0!
0'
#646640000000
1!
1$
b1 %
1'
1*
b1 +
#646650000000
0!
0'
#646660000000
1!
b10 %
1'
b10 +
#646670000000
0!
0'
#646680000000
1!
b11 %
1'
b11 +
#646690000000
0!
0'
#646700000000
1!
b100 %
1'
b100 +
#646710000000
0!
0'
#646720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#646730000000
0!
0'
#646740000000
1!
0$
b110 %
1'
0*
b110 +
#646750000000
0!
0'
#646760000000
1!
b111 %
1'
b111 +
#646770000000
0!
0'
#646780000000
1!
b1000 %
1'
b1000 +
#646790000000
0!
0'
#646800000000
1!
b1001 %
1'
b1001 +
#646810000000
0!
0'
#646820000000
1!
b0 %
1'
b0 +
#646830000000
0!
0'
#646840000000
1!
1$
b1 %
1'
1*
b1 +
#646850000000
0!
0'
#646860000000
1!
b10 %
1'
b10 +
#646870000000
0!
0'
#646880000000
1!
b11 %
1'
b11 +
#646890000000
0!
0'
#646900000000
1!
b100 %
1'
b100 +
#646910000000
0!
0'
#646920000000
1!
b101 %
1'
b101 +
#646930000000
1"
1(
#646940000000
0!
0"
b100 &
0'
0(
b100 ,
#646950000000
1!
b110 %
1'
b110 +
#646960000000
0!
0'
#646970000000
1!
b111 %
1'
b111 +
#646980000000
0!
0'
#646990000000
1!
0$
b1000 %
1'
0*
b1000 +
#647000000000
0!
0'
#647010000000
1!
b1001 %
1'
b1001 +
#647020000000
0!
0'
#647030000000
1!
b0 %
1'
b0 +
#647040000000
0!
0'
#647050000000
1!
1$
b1 %
1'
1*
b1 +
#647060000000
0!
0'
#647070000000
1!
b10 %
1'
b10 +
#647080000000
0!
0'
#647090000000
1!
b11 %
1'
b11 +
#647100000000
0!
0'
#647110000000
1!
b100 %
1'
b100 +
#647120000000
0!
0'
#647130000000
1!
b101 %
1'
b101 +
#647140000000
0!
0'
#647150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#647160000000
0!
0'
#647170000000
1!
b111 %
1'
b111 +
#647180000000
0!
0'
#647190000000
1!
b1000 %
1'
b1000 +
#647200000000
0!
0'
#647210000000
1!
b1001 %
1'
b1001 +
#647220000000
0!
0'
#647230000000
1!
b0 %
1'
b0 +
#647240000000
0!
0'
#647250000000
1!
1$
b1 %
1'
1*
b1 +
#647260000000
0!
0'
#647270000000
1!
b10 %
1'
b10 +
#647280000000
0!
0'
#647290000000
1!
b11 %
1'
b11 +
#647300000000
0!
0'
#647310000000
1!
b100 %
1'
b100 +
#647320000000
0!
0'
#647330000000
1!
b101 %
1'
b101 +
#647340000000
0!
0'
#647350000000
1!
0$
b110 %
1'
0*
b110 +
#647360000000
1"
1(
#647370000000
0!
0"
b100 &
0'
0(
b100 ,
#647380000000
1!
1$
b111 %
1'
1*
b111 +
#647390000000
0!
0'
#647400000000
1!
0$
b1000 %
1'
0*
b1000 +
#647410000000
0!
0'
#647420000000
1!
b1001 %
1'
b1001 +
#647430000000
0!
0'
#647440000000
1!
b0 %
1'
b0 +
#647450000000
0!
0'
#647460000000
1!
1$
b1 %
1'
1*
b1 +
#647470000000
0!
0'
#647480000000
1!
b10 %
1'
b10 +
#647490000000
0!
0'
#647500000000
1!
b11 %
1'
b11 +
#647510000000
0!
0'
#647520000000
1!
b100 %
1'
b100 +
#647530000000
0!
0'
#647540000000
1!
b101 %
1'
b101 +
#647550000000
0!
0'
#647560000000
1!
b110 %
1'
b110 +
#647570000000
0!
0'
#647580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#647590000000
0!
0'
#647600000000
1!
b1000 %
1'
b1000 +
#647610000000
0!
0'
#647620000000
1!
b1001 %
1'
b1001 +
#647630000000
0!
0'
#647640000000
1!
b0 %
1'
b0 +
#647650000000
0!
0'
#647660000000
1!
1$
b1 %
1'
1*
b1 +
#647670000000
0!
0'
#647680000000
1!
b10 %
1'
b10 +
#647690000000
0!
0'
#647700000000
1!
b11 %
1'
b11 +
#647710000000
0!
0'
#647720000000
1!
b100 %
1'
b100 +
#647730000000
0!
0'
#647740000000
1!
b101 %
1'
b101 +
#647750000000
0!
0'
#647760000000
1!
0$
b110 %
1'
0*
b110 +
#647770000000
0!
0'
#647780000000
1!
b111 %
1'
b111 +
#647790000000
1"
1(
#647800000000
0!
0"
b100 &
0'
0(
b100 ,
#647810000000
1!
b1000 %
1'
b1000 +
#647820000000
0!
0'
#647830000000
1!
b1001 %
1'
b1001 +
#647840000000
0!
0'
#647850000000
1!
b0 %
1'
b0 +
#647860000000
0!
0'
#647870000000
1!
1$
b1 %
1'
1*
b1 +
#647880000000
0!
0'
#647890000000
1!
b10 %
1'
b10 +
#647900000000
0!
0'
#647910000000
1!
b11 %
1'
b11 +
#647920000000
0!
0'
#647930000000
1!
b100 %
1'
b100 +
#647940000000
0!
0'
#647950000000
1!
b101 %
1'
b101 +
#647960000000
0!
0'
#647970000000
1!
b110 %
1'
b110 +
#647980000000
0!
0'
#647990000000
1!
b111 %
1'
b111 +
#648000000000
0!
0'
#648010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#648020000000
0!
0'
#648030000000
1!
b1001 %
1'
b1001 +
#648040000000
0!
0'
#648050000000
1!
b0 %
1'
b0 +
#648060000000
0!
0'
#648070000000
1!
1$
b1 %
1'
1*
b1 +
#648080000000
0!
0'
#648090000000
1!
b10 %
1'
b10 +
#648100000000
0!
0'
#648110000000
1!
b11 %
1'
b11 +
#648120000000
0!
0'
#648130000000
1!
b100 %
1'
b100 +
#648140000000
0!
0'
#648150000000
1!
b101 %
1'
b101 +
#648160000000
0!
0'
#648170000000
1!
0$
b110 %
1'
0*
b110 +
#648180000000
0!
0'
#648190000000
1!
b111 %
1'
b111 +
#648200000000
0!
0'
#648210000000
1!
b1000 %
1'
b1000 +
#648220000000
1"
1(
#648230000000
0!
0"
b100 &
0'
0(
b100 ,
#648240000000
1!
b1001 %
1'
b1001 +
#648250000000
0!
0'
#648260000000
1!
b0 %
1'
b0 +
#648270000000
0!
0'
#648280000000
1!
1$
b1 %
1'
1*
b1 +
#648290000000
0!
0'
#648300000000
1!
b10 %
1'
b10 +
#648310000000
0!
0'
#648320000000
1!
b11 %
1'
b11 +
#648330000000
0!
0'
#648340000000
1!
b100 %
1'
b100 +
#648350000000
0!
0'
#648360000000
1!
b101 %
1'
b101 +
#648370000000
0!
0'
#648380000000
1!
b110 %
1'
b110 +
#648390000000
0!
0'
#648400000000
1!
b111 %
1'
b111 +
#648410000000
0!
0'
#648420000000
1!
0$
b1000 %
1'
0*
b1000 +
#648430000000
0!
0'
#648440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#648450000000
0!
0'
#648460000000
1!
b0 %
1'
b0 +
#648470000000
0!
0'
#648480000000
1!
1$
b1 %
1'
1*
b1 +
#648490000000
0!
0'
#648500000000
1!
b10 %
1'
b10 +
#648510000000
0!
0'
#648520000000
1!
b11 %
1'
b11 +
#648530000000
0!
0'
#648540000000
1!
b100 %
1'
b100 +
#648550000000
0!
0'
#648560000000
1!
b101 %
1'
b101 +
#648570000000
0!
0'
#648580000000
1!
0$
b110 %
1'
0*
b110 +
#648590000000
0!
0'
#648600000000
1!
b111 %
1'
b111 +
#648610000000
0!
0'
#648620000000
1!
b1000 %
1'
b1000 +
#648630000000
0!
0'
#648640000000
1!
b1001 %
1'
b1001 +
#648650000000
1"
1(
#648660000000
0!
0"
b100 &
0'
0(
b100 ,
#648670000000
1!
b0 %
1'
b0 +
#648680000000
0!
0'
#648690000000
1!
1$
b1 %
1'
1*
b1 +
#648700000000
0!
0'
#648710000000
1!
b10 %
1'
b10 +
#648720000000
0!
0'
#648730000000
1!
b11 %
1'
b11 +
#648740000000
0!
0'
#648750000000
1!
b100 %
1'
b100 +
#648760000000
0!
0'
#648770000000
1!
b101 %
1'
b101 +
#648780000000
0!
0'
#648790000000
1!
b110 %
1'
b110 +
#648800000000
0!
0'
#648810000000
1!
b111 %
1'
b111 +
#648820000000
0!
0'
#648830000000
1!
0$
b1000 %
1'
0*
b1000 +
#648840000000
0!
0'
#648850000000
1!
b1001 %
1'
b1001 +
#648860000000
0!
0'
#648870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#648880000000
0!
0'
#648890000000
1!
1$
b1 %
1'
1*
b1 +
#648900000000
0!
0'
#648910000000
1!
b10 %
1'
b10 +
#648920000000
0!
0'
#648930000000
1!
b11 %
1'
b11 +
#648940000000
0!
0'
#648950000000
1!
b100 %
1'
b100 +
#648960000000
0!
0'
#648970000000
1!
b101 %
1'
b101 +
#648980000000
0!
0'
#648990000000
1!
0$
b110 %
1'
0*
b110 +
#649000000000
0!
0'
#649010000000
1!
b111 %
1'
b111 +
#649020000000
0!
0'
#649030000000
1!
b1000 %
1'
b1000 +
#649040000000
0!
0'
#649050000000
1!
b1001 %
1'
b1001 +
#649060000000
0!
0'
#649070000000
1!
b0 %
1'
b0 +
#649080000000
1"
1(
#649090000000
0!
0"
b100 &
0'
0(
b100 ,
#649100000000
1!
1$
b1 %
1'
1*
b1 +
#649110000000
0!
0'
#649120000000
1!
b10 %
1'
b10 +
#649130000000
0!
0'
#649140000000
1!
b11 %
1'
b11 +
#649150000000
0!
0'
#649160000000
1!
b100 %
1'
b100 +
#649170000000
0!
0'
#649180000000
1!
b101 %
1'
b101 +
#649190000000
0!
0'
#649200000000
1!
b110 %
1'
b110 +
#649210000000
0!
0'
#649220000000
1!
b111 %
1'
b111 +
#649230000000
0!
0'
#649240000000
1!
0$
b1000 %
1'
0*
b1000 +
#649250000000
0!
0'
#649260000000
1!
b1001 %
1'
b1001 +
#649270000000
0!
0'
#649280000000
1!
b0 %
1'
b0 +
#649290000000
0!
0'
#649300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#649310000000
0!
0'
#649320000000
1!
b10 %
1'
b10 +
#649330000000
0!
0'
#649340000000
1!
b11 %
1'
b11 +
#649350000000
0!
0'
#649360000000
1!
b100 %
1'
b100 +
#649370000000
0!
0'
#649380000000
1!
b101 %
1'
b101 +
#649390000000
0!
0'
#649400000000
1!
0$
b110 %
1'
0*
b110 +
#649410000000
0!
0'
#649420000000
1!
b111 %
1'
b111 +
#649430000000
0!
0'
#649440000000
1!
b1000 %
1'
b1000 +
#649450000000
0!
0'
#649460000000
1!
b1001 %
1'
b1001 +
#649470000000
0!
0'
#649480000000
1!
b0 %
1'
b0 +
#649490000000
0!
0'
#649500000000
1!
1$
b1 %
1'
1*
b1 +
#649510000000
1"
1(
#649520000000
0!
0"
b100 &
0'
0(
b100 ,
#649530000000
1!
b10 %
1'
b10 +
#649540000000
0!
0'
#649550000000
1!
b11 %
1'
b11 +
#649560000000
0!
0'
#649570000000
1!
b100 %
1'
b100 +
#649580000000
0!
0'
#649590000000
1!
b101 %
1'
b101 +
#649600000000
0!
0'
#649610000000
1!
b110 %
1'
b110 +
#649620000000
0!
0'
#649630000000
1!
b111 %
1'
b111 +
#649640000000
0!
0'
#649650000000
1!
0$
b1000 %
1'
0*
b1000 +
#649660000000
0!
0'
#649670000000
1!
b1001 %
1'
b1001 +
#649680000000
0!
0'
#649690000000
1!
b0 %
1'
b0 +
#649700000000
0!
0'
#649710000000
1!
1$
b1 %
1'
1*
b1 +
#649720000000
0!
0'
#649730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#649740000000
0!
0'
#649750000000
1!
b11 %
1'
b11 +
#649760000000
0!
0'
#649770000000
1!
b100 %
1'
b100 +
#649780000000
0!
0'
#649790000000
1!
b101 %
1'
b101 +
#649800000000
0!
0'
#649810000000
1!
0$
b110 %
1'
0*
b110 +
#649820000000
0!
0'
#649830000000
1!
b111 %
1'
b111 +
#649840000000
0!
0'
#649850000000
1!
b1000 %
1'
b1000 +
#649860000000
0!
0'
#649870000000
1!
b1001 %
1'
b1001 +
#649880000000
0!
0'
#649890000000
1!
b0 %
1'
b0 +
#649900000000
0!
0'
#649910000000
1!
1$
b1 %
1'
1*
b1 +
#649920000000
0!
0'
#649930000000
1!
b10 %
1'
b10 +
#649940000000
1"
1(
#649950000000
0!
0"
b100 &
0'
0(
b100 ,
#649960000000
1!
b11 %
1'
b11 +
#649970000000
0!
0'
#649980000000
1!
b100 %
1'
b100 +
#649990000000
0!
0'
#650000000000
1!
b101 %
1'
b101 +
#650010000000
0!
0'
#650020000000
1!
b110 %
1'
b110 +
#650030000000
0!
0'
#650040000000
1!
b111 %
1'
b111 +
#650050000000
0!
0'
#650060000000
1!
0$
b1000 %
1'
0*
b1000 +
#650070000000
0!
0'
#650080000000
1!
b1001 %
1'
b1001 +
#650090000000
0!
0'
#650100000000
1!
b0 %
1'
b0 +
#650110000000
0!
0'
#650120000000
1!
1$
b1 %
1'
1*
b1 +
#650130000000
0!
0'
#650140000000
1!
b10 %
1'
b10 +
#650150000000
0!
0'
#650160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#650170000000
0!
0'
#650180000000
1!
b100 %
1'
b100 +
#650190000000
0!
0'
#650200000000
1!
b101 %
1'
b101 +
#650210000000
0!
0'
#650220000000
1!
0$
b110 %
1'
0*
b110 +
#650230000000
0!
0'
#650240000000
1!
b111 %
1'
b111 +
#650250000000
0!
0'
#650260000000
1!
b1000 %
1'
b1000 +
#650270000000
0!
0'
#650280000000
1!
b1001 %
1'
b1001 +
#650290000000
0!
0'
#650300000000
1!
b0 %
1'
b0 +
#650310000000
0!
0'
#650320000000
1!
1$
b1 %
1'
1*
b1 +
#650330000000
0!
0'
#650340000000
1!
b10 %
1'
b10 +
#650350000000
0!
0'
#650360000000
1!
b11 %
1'
b11 +
#650370000000
1"
1(
#650380000000
0!
0"
b100 &
0'
0(
b100 ,
#650390000000
1!
b100 %
1'
b100 +
#650400000000
0!
0'
#650410000000
1!
b101 %
1'
b101 +
#650420000000
0!
0'
#650430000000
1!
b110 %
1'
b110 +
#650440000000
0!
0'
#650450000000
1!
b111 %
1'
b111 +
#650460000000
0!
0'
#650470000000
1!
0$
b1000 %
1'
0*
b1000 +
#650480000000
0!
0'
#650490000000
1!
b1001 %
1'
b1001 +
#650500000000
0!
0'
#650510000000
1!
b0 %
1'
b0 +
#650520000000
0!
0'
#650530000000
1!
1$
b1 %
1'
1*
b1 +
#650540000000
0!
0'
#650550000000
1!
b10 %
1'
b10 +
#650560000000
0!
0'
#650570000000
1!
b11 %
1'
b11 +
#650580000000
0!
0'
#650590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#650600000000
0!
0'
#650610000000
1!
b101 %
1'
b101 +
#650620000000
0!
0'
#650630000000
1!
0$
b110 %
1'
0*
b110 +
#650640000000
0!
0'
#650650000000
1!
b111 %
1'
b111 +
#650660000000
0!
0'
#650670000000
1!
b1000 %
1'
b1000 +
#650680000000
0!
0'
#650690000000
1!
b1001 %
1'
b1001 +
#650700000000
0!
0'
#650710000000
1!
b0 %
1'
b0 +
#650720000000
0!
0'
#650730000000
1!
1$
b1 %
1'
1*
b1 +
#650740000000
0!
0'
#650750000000
1!
b10 %
1'
b10 +
#650760000000
0!
0'
#650770000000
1!
b11 %
1'
b11 +
#650780000000
0!
0'
#650790000000
1!
b100 %
1'
b100 +
#650800000000
1"
1(
#650810000000
0!
0"
b100 &
0'
0(
b100 ,
#650820000000
1!
b101 %
1'
b101 +
#650830000000
0!
0'
#650840000000
1!
b110 %
1'
b110 +
#650850000000
0!
0'
#650860000000
1!
b111 %
1'
b111 +
#650870000000
0!
0'
#650880000000
1!
0$
b1000 %
1'
0*
b1000 +
#650890000000
0!
0'
#650900000000
1!
b1001 %
1'
b1001 +
#650910000000
0!
0'
#650920000000
1!
b0 %
1'
b0 +
#650930000000
0!
0'
#650940000000
1!
1$
b1 %
1'
1*
b1 +
#650950000000
0!
0'
#650960000000
1!
b10 %
1'
b10 +
#650970000000
0!
0'
#650980000000
1!
b11 %
1'
b11 +
#650990000000
0!
0'
#651000000000
1!
b100 %
1'
b100 +
#651010000000
0!
0'
#651020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#651030000000
0!
0'
#651040000000
1!
0$
b110 %
1'
0*
b110 +
#651050000000
0!
0'
#651060000000
1!
b111 %
1'
b111 +
#651070000000
0!
0'
#651080000000
1!
b1000 %
1'
b1000 +
#651090000000
0!
0'
#651100000000
1!
b1001 %
1'
b1001 +
#651110000000
0!
0'
#651120000000
1!
b0 %
1'
b0 +
#651130000000
0!
0'
#651140000000
1!
1$
b1 %
1'
1*
b1 +
#651150000000
0!
0'
#651160000000
1!
b10 %
1'
b10 +
#651170000000
0!
0'
#651180000000
1!
b11 %
1'
b11 +
#651190000000
0!
0'
#651200000000
1!
b100 %
1'
b100 +
#651210000000
0!
0'
#651220000000
1!
b101 %
1'
b101 +
#651230000000
1"
1(
#651240000000
0!
0"
b100 &
0'
0(
b100 ,
#651250000000
1!
b110 %
1'
b110 +
#651260000000
0!
0'
#651270000000
1!
b111 %
1'
b111 +
#651280000000
0!
0'
#651290000000
1!
0$
b1000 %
1'
0*
b1000 +
#651300000000
0!
0'
#651310000000
1!
b1001 %
1'
b1001 +
#651320000000
0!
0'
#651330000000
1!
b0 %
1'
b0 +
#651340000000
0!
0'
#651350000000
1!
1$
b1 %
1'
1*
b1 +
#651360000000
0!
0'
#651370000000
1!
b10 %
1'
b10 +
#651380000000
0!
0'
#651390000000
1!
b11 %
1'
b11 +
#651400000000
0!
0'
#651410000000
1!
b100 %
1'
b100 +
#651420000000
0!
0'
#651430000000
1!
b101 %
1'
b101 +
#651440000000
0!
0'
#651450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#651460000000
0!
0'
#651470000000
1!
b111 %
1'
b111 +
#651480000000
0!
0'
#651490000000
1!
b1000 %
1'
b1000 +
#651500000000
0!
0'
#651510000000
1!
b1001 %
1'
b1001 +
#651520000000
0!
0'
#651530000000
1!
b0 %
1'
b0 +
#651540000000
0!
0'
#651550000000
1!
1$
b1 %
1'
1*
b1 +
#651560000000
0!
0'
#651570000000
1!
b10 %
1'
b10 +
#651580000000
0!
0'
#651590000000
1!
b11 %
1'
b11 +
#651600000000
0!
0'
#651610000000
1!
b100 %
1'
b100 +
#651620000000
0!
0'
#651630000000
1!
b101 %
1'
b101 +
#651640000000
0!
0'
#651650000000
1!
0$
b110 %
1'
0*
b110 +
#651660000000
1"
1(
#651670000000
0!
0"
b100 &
0'
0(
b100 ,
#651680000000
1!
1$
b111 %
1'
1*
b111 +
#651690000000
0!
0'
#651700000000
1!
0$
b1000 %
1'
0*
b1000 +
#651710000000
0!
0'
#651720000000
1!
b1001 %
1'
b1001 +
#651730000000
0!
0'
#651740000000
1!
b0 %
1'
b0 +
#651750000000
0!
0'
#651760000000
1!
1$
b1 %
1'
1*
b1 +
#651770000000
0!
0'
#651780000000
1!
b10 %
1'
b10 +
#651790000000
0!
0'
#651800000000
1!
b11 %
1'
b11 +
#651810000000
0!
0'
#651820000000
1!
b100 %
1'
b100 +
#651830000000
0!
0'
#651840000000
1!
b101 %
1'
b101 +
#651850000000
0!
0'
#651860000000
1!
b110 %
1'
b110 +
#651870000000
0!
0'
#651880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#651890000000
0!
0'
#651900000000
1!
b1000 %
1'
b1000 +
#651910000000
0!
0'
#651920000000
1!
b1001 %
1'
b1001 +
#651930000000
0!
0'
#651940000000
1!
b0 %
1'
b0 +
#651950000000
0!
0'
#651960000000
1!
1$
b1 %
1'
1*
b1 +
#651970000000
0!
0'
#651980000000
1!
b10 %
1'
b10 +
#651990000000
0!
0'
#652000000000
1!
b11 %
1'
b11 +
#652010000000
0!
0'
#652020000000
1!
b100 %
1'
b100 +
#652030000000
0!
0'
#652040000000
1!
b101 %
1'
b101 +
#652050000000
0!
0'
#652060000000
1!
0$
b110 %
1'
0*
b110 +
#652070000000
0!
0'
#652080000000
1!
b111 %
1'
b111 +
#652090000000
1"
1(
#652100000000
0!
0"
b100 &
0'
0(
b100 ,
#652110000000
1!
b1000 %
1'
b1000 +
#652120000000
0!
0'
#652130000000
1!
b1001 %
1'
b1001 +
#652140000000
0!
0'
#652150000000
1!
b0 %
1'
b0 +
#652160000000
0!
0'
#652170000000
1!
1$
b1 %
1'
1*
b1 +
#652180000000
0!
0'
#652190000000
1!
b10 %
1'
b10 +
#652200000000
0!
0'
#652210000000
1!
b11 %
1'
b11 +
#652220000000
0!
0'
#652230000000
1!
b100 %
1'
b100 +
#652240000000
0!
0'
#652250000000
1!
b101 %
1'
b101 +
#652260000000
0!
0'
#652270000000
1!
b110 %
1'
b110 +
#652280000000
0!
0'
#652290000000
1!
b111 %
1'
b111 +
#652300000000
0!
0'
#652310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#652320000000
0!
0'
#652330000000
1!
b1001 %
1'
b1001 +
#652340000000
0!
0'
#652350000000
1!
b0 %
1'
b0 +
#652360000000
0!
0'
#652370000000
1!
1$
b1 %
1'
1*
b1 +
#652380000000
0!
0'
#652390000000
1!
b10 %
1'
b10 +
#652400000000
0!
0'
#652410000000
1!
b11 %
1'
b11 +
#652420000000
0!
0'
#652430000000
1!
b100 %
1'
b100 +
#652440000000
0!
0'
#652450000000
1!
b101 %
1'
b101 +
#652460000000
0!
0'
#652470000000
1!
0$
b110 %
1'
0*
b110 +
#652480000000
0!
0'
#652490000000
1!
b111 %
1'
b111 +
#652500000000
0!
0'
#652510000000
1!
b1000 %
1'
b1000 +
#652520000000
1"
1(
#652530000000
0!
0"
b100 &
0'
0(
b100 ,
#652540000000
1!
b1001 %
1'
b1001 +
#652550000000
0!
0'
#652560000000
1!
b0 %
1'
b0 +
#652570000000
0!
0'
#652580000000
1!
1$
b1 %
1'
1*
b1 +
#652590000000
0!
0'
#652600000000
1!
b10 %
1'
b10 +
#652610000000
0!
0'
#652620000000
1!
b11 %
1'
b11 +
#652630000000
0!
0'
#652640000000
1!
b100 %
1'
b100 +
#652650000000
0!
0'
#652660000000
1!
b101 %
1'
b101 +
#652670000000
0!
0'
#652680000000
1!
b110 %
1'
b110 +
#652690000000
0!
0'
#652700000000
1!
b111 %
1'
b111 +
#652710000000
0!
0'
#652720000000
1!
0$
b1000 %
1'
0*
b1000 +
#652730000000
0!
0'
#652740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#652750000000
0!
0'
#652760000000
1!
b0 %
1'
b0 +
#652770000000
0!
0'
#652780000000
1!
1$
b1 %
1'
1*
b1 +
#652790000000
0!
0'
#652800000000
1!
b10 %
1'
b10 +
#652810000000
0!
0'
#652820000000
1!
b11 %
1'
b11 +
#652830000000
0!
0'
#652840000000
1!
b100 %
1'
b100 +
#652850000000
0!
0'
#652860000000
1!
b101 %
1'
b101 +
#652870000000
0!
0'
#652880000000
1!
0$
b110 %
1'
0*
b110 +
#652890000000
0!
0'
#652900000000
1!
b111 %
1'
b111 +
#652910000000
0!
0'
#652920000000
1!
b1000 %
1'
b1000 +
#652930000000
0!
0'
#652940000000
1!
b1001 %
1'
b1001 +
#652950000000
1"
1(
#652960000000
0!
0"
b100 &
0'
0(
b100 ,
#652970000000
1!
b0 %
1'
b0 +
#652980000000
0!
0'
#652990000000
1!
1$
b1 %
1'
1*
b1 +
#653000000000
0!
0'
#653010000000
1!
b10 %
1'
b10 +
#653020000000
0!
0'
#653030000000
1!
b11 %
1'
b11 +
#653040000000
0!
0'
#653050000000
1!
b100 %
1'
b100 +
#653060000000
0!
0'
#653070000000
1!
b101 %
1'
b101 +
#653080000000
0!
0'
#653090000000
1!
b110 %
1'
b110 +
#653100000000
0!
0'
#653110000000
1!
b111 %
1'
b111 +
#653120000000
0!
0'
#653130000000
1!
0$
b1000 %
1'
0*
b1000 +
#653140000000
0!
0'
#653150000000
1!
b1001 %
1'
b1001 +
#653160000000
0!
0'
#653170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#653180000000
0!
0'
#653190000000
1!
1$
b1 %
1'
1*
b1 +
#653200000000
0!
0'
#653210000000
1!
b10 %
1'
b10 +
#653220000000
0!
0'
#653230000000
1!
b11 %
1'
b11 +
#653240000000
0!
0'
#653250000000
1!
b100 %
1'
b100 +
#653260000000
0!
0'
#653270000000
1!
b101 %
1'
b101 +
#653280000000
0!
0'
#653290000000
1!
0$
b110 %
1'
0*
b110 +
#653300000000
0!
0'
#653310000000
1!
b111 %
1'
b111 +
#653320000000
0!
0'
#653330000000
1!
b1000 %
1'
b1000 +
#653340000000
0!
0'
#653350000000
1!
b1001 %
1'
b1001 +
#653360000000
0!
0'
#653370000000
1!
b0 %
1'
b0 +
#653380000000
1"
1(
#653390000000
0!
0"
b100 &
0'
0(
b100 ,
#653400000000
1!
1$
b1 %
1'
1*
b1 +
#653410000000
0!
0'
#653420000000
1!
b10 %
1'
b10 +
#653430000000
0!
0'
#653440000000
1!
b11 %
1'
b11 +
#653450000000
0!
0'
#653460000000
1!
b100 %
1'
b100 +
#653470000000
0!
0'
#653480000000
1!
b101 %
1'
b101 +
#653490000000
0!
0'
#653500000000
1!
b110 %
1'
b110 +
#653510000000
0!
0'
#653520000000
1!
b111 %
1'
b111 +
#653530000000
0!
0'
#653540000000
1!
0$
b1000 %
1'
0*
b1000 +
#653550000000
0!
0'
#653560000000
1!
b1001 %
1'
b1001 +
#653570000000
0!
0'
#653580000000
1!
b0 %
1'
b0 +
#653590000000
0!
0'
#653600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#653610000000
0!
0'
#653620000000
1!
b10 %
1'
b10 +
#653630000000
0!
0'
#653640000000
1!
b11 %
1'
b11 +
#653650000000
0!
0'
#653660000000
1!
b100 %
1'
b100 +
#653670000000
0!
0'
#653680000000
1!
b101 %
1'
b101 +
#653690000000
0!
0'
#653700000000
1!
0$
b110 %
1'
0*
b110 +
#653710000000
0!
0'
#653720000000
1!
b111 %
1'
b111 +
#653730000000
0!
0'
#653740000000
1!
b1000 %
1'
b1000 +
#653750000000
0!
0'
#653760000000
1!
b1001 %
1'
b1001 +
#653770000000
0!
0'
#653780000000
1!
b0 %
1'
b0 +
#653790000000
0!
0'
#653800000000
1!
1$
b1 %
1'
1*
b1 +
#653810000000
1"
1(
#653820000000
0!
0"
b100 &
0'
0(
b100 ,
#653830000000
1!
b10 %
1'
b10 +
#653840000000
0!
0'
#653850000000
1!
b11 %
1'
b11 +
#653860000000
0!
0'
#653870000000
1!
b100 %
1'
b100 +
#653880000000
0!
0'
#653890000000
1!
b101 %
1'
b101 +
#653900000000
0!
0'
#653910000000
1!
b110 %
1'
b110 +
#653920000000
0!
0'
#653930000000
1!
b111 %
1'
b111 +
#653940000000
0!
0'
#653950000000
1!
0$
b1000 %
1'
0*
b1000 +
#653960000000
0!
0'
#653970000000
1!
b1001 %
1'
b1001 +
#653980000000
0!
0'
#653990000000
1!
b0 %
1'
b0 +
#654000000000
0!
0'
#654010000000
1!
1$
b1 %
1'
1*
b1 +
#654020000000
0!
0'
#654030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#654040000000
0!
0'
#654050000000
1!
b11 %
1'
b11 +
#654060000000
0!
0'
#654070000000
1!
b100 %
1'
b100 +
#654080000000
0!
0'
#654090000000
1!
b101 %
1'
b101 +
#654100000000
0!
0'
#654110000000
1!
0$
b110 %
1'
0*
b110 +
#654120000000
0!
0'
#654130000000
1!
b111 %
1'
b111 +
#654140000000
0!
0'
#654150000000
1!
b1000 %
1'
b1000 +
#654160000000
0!
0'
#654170000000
1!
b1001 %
1'
b1001 +
#654180000000
0!
0'
#654190000000
1!
b0 %
1'
b0 +
#654200000000
0!
0'
#654210000000
1!
1$
b1 %
1'
1*
b1 +
#654220000000
0!
0'
#654230000000
1!
b10 %
1'
b10 +
#654240000000
1"
1(
#654250000000
0!
0"
b100 &
0'
0(
b100 ,
#654260000000
1!
b11 %
1'
b11 +
#654270000000
0!
0'
#654280000000
1!
b100 %
1'
b100 +
#654290000000
0!
0'
#654300000000
1!
b101 %
1'
b101 +
#654310000000
0!
0'
#654320000000
1!
b110 %
1'
b110 +
#654330000000
0!
0'
#654340000000
1!
b111 %
1'
b111 +
#654350000000
0!
0'
#654360000000
1!
0$
b1000 %
1'
0*
b1000 +
#654370000000
0!
0'
#654380000000
1!
b1001 %
1'
b1001 +
#654390000000
0!
0'
#654400000000
1!
b0 %
1'
b0 +
#654410000000
0!
0'
#654420000000
1!
1$
b1 %
1'
1*
b1 +
#654430000000
0!
0'
#654440000000
1!
b10 %
1'
b10 +
#654450000000
0!
0'
#654460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#654470000000
0!
0'
#654480000000
1!
b100 %
1'
b100 +
#654490000000
0!
0'
#654500000000
1!
b101 %
1'
b101 +
#654510000000
0!
0'
#654520000000
1!
0$
b110 %
1'
0*
b110 +
#654530000000
0!
0'
#654540000000
1!
b111 %
1'
b111 +
#654550000000
0!
0'
#654560000000
1!
b1000 %
1'
b1000 +
#654570000000
0!
0'
#654580000000
1!
b1001 %
1'
b1001 +
#654590000000
0!
0'
#654600000000
1!
b0 %
1'
b0 +
#654610000000
0!
0'
#654620000000
1!
1$
b1 %
1'
1*
b1 +
#654630000000
0!
0'
#654640000000
1!
b10 %
1'
b10 +
#654650000000
0!
0'
#654660000000
1!
b11 %
1'
b11 +
#654670000000
1"
1(
#654680000000
0!
0"
b100 &
0'
0(
b100 ,
#654690000000
1!
b100 %
1'
b100 +
#654700000000
0!
0'
#654710000000
1!
b101 %
1'
b101 +
#654720000000
0!
0'
#654730000000
1!
b110 %
1'
b110 +
#654740000000
0!
0'
#654750000000
1!
b111 %
1'
b111 +
#654760000000
0!
0'
#654770000000
1!
0$
b1000 %
1'
0*
b1000 +
#654780000000
0!
0'
#654790000000
1!
b1001 %
1'
b1001 +
#654800000000
0!
0'
#654810000000
1!
b0 %
1'
b0 +
#654820000000
0!
0'
#654830000000
1!
1$
b1 %
1'
1*
b1 +
#654840000000
0!
0'
#654850000000
1!
b10 %
1'
b10 +
#654860000000
0!
0'
#654870000000
1!
b11 %
1'
b11 +
#654880000000
0!
0'
#654890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#654900000000
0!
0'
#654910000000
1!
b101 %
1'
b101 +
#654920000000
0!
0'
#654930000000
1!
0$
b110 %
1'
0*
b110 +
#654940000000
0!
0'
#654950000000
1!
b111 %
1'
b111 +
#654960000000
0!
0'
#654970000000
1!
b1000 %
1'
b1000 +
#654980000000
0!
0'
#654990000000
1!
b1001 %
1'
b1001 +
#655000000000
0!
0'
#655010000000
1!
b0 %
1'
b0 +
#655020000000
0!
0'
#655030000000
1!
1$
b1 %
1'
1*
b1 +
#655040000000
0!
0'
#655050000000
1!
b10 %
1'
b10 +
#655060000000
0!
0'
#655070000000
1!
b11 %
1'
b11 +
#655080000000
0!
0'
#655090000000
1!
b100 %
1'
b100 +
#655100000000
1"
1(
#655110000000
0!
0"
b100 &
0'
0(
b100 ,
#655120000000
1!
b101 %
1'
b101 +
#655130000000
0!
0'
#655140000000
1!
b110 %
1'
b110 +
#655150000000
0!
0'
#655160000000
1!
b111 %
1'
b111 +
#655170000000
0!
0'
#655180000000
1!
0$
b1000 %
1'
0*
b1000 +
#655190000000
0!
0'
#655200000000
1!
b1001 %
1'
b1001 +
#655210000000
0!
0'
#655220000000
1!
b0 %
1'
b0 +
#655230000000
0!
0'
#655240000000
1!
1$
b1 %
1'
1*
b1 +
#655250000000
0!
0'
#655260000000
1!
b10 %
1'
b10 +
#655270000000
0!
0'
#655280000000
1!
b11 %
1'
b11 +
#655290000000
0!
0'
#655300000000
1!
b100 %
1'
b100 +
#655310000000
0!
0'
#655320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#655330000000
0!
0'
#655340000000
1!
0$
b110 %
1'
0*
b110 +
#655350000000
0!
0'
#655360000000
1!
b111 %
1'
b111 +
#655370000000
0!
0'
#655380000000
1!
b1000 %
1'
b1000 +
#655390000000
0!
0'
#655400000000
1!
b1001 %
1'
b1001 +
#655410000000
0!
0'
#655420000000
1!
b0 %
1'
b0 +
#655430000000
0!
0'
#655440000000
1!
1$
b1 %
1'
1*
b1 +
#655450000000
0!
0'
#655460000000
1!
b10 %
1'
b10 +
#655470000000
0!
0'
#655480000000
1!
b11 %
1'
b11 +
#655490000000
0!
0'
#655500000000
1!
b100 %
1'
b100 +
#655510000000
0!
0'
#655520000000
1!
b101 %
1'
b101 +
#655530000000
1"
1(
#655540000000
0!
0"
b100 &
0'
0(
b100 ,
#655550000000
1!
b110 %
1'
b110 +
#655560000000
0!
0'
#655570000000
1!
b111 %
1'
b111 +
#655580000000
0!
0'
#655590000000
1!
0$
b1000 %
1'
0*
b1000 +
#655600000000
0!
0'
#655610000000
1!
b1001 %
1'
b1001 +
#655620000000
0!
0'
#655630000000
1!
b0 %
1'
b0 +
#655640000000
0!
0'
#655650000000
1!
1$
b1 %
1'
1*
b1 +
#655660000000
0!
0'
#655670000000
1!
b10 %
1'
b10 +
#655680000000
0!
0'
#655690000000
1!
b11 %
1'
b11 +
#655700000000
0!
0'
#655710000000
1!
b100 %
1'
b100 +
#655720000000
0!
0'
#655730000000
1!
b101 %
1'
b101 +
#655740000000
0!
0'
#655750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#655760000000
0!
0'
#655770000000
1!
b111 %
1'
b111 +
#655780000000
0!
0'
#655790000000
1!
b1000 %
1'
b1000 +
#655800000000
0!
0'
#655810000000
1!
b1001 %
1'
b1001 +
#655820000000
0!
0'
#655830000000
1!
b0 %
1'
b0 +
#655840000000
0!
0'
#655850000000
1!
1$
b1 %
1'
1*
b1 +
#655860000000
0!
0'
#655870000000
1!
b10 %
1'
b10 +
#655880000000
0!
0'
#655890000000
1!
b11 %
1'
b11 +
#655900000000
0!
0'
#655910000000
1!
b100 %
1'
b100 +
#655920000000
0!
0'
#655930000000
1!
b101 %
1'
b101 +
#655940000000
0!
0'
#655950000000
1!
0$
b110 %
1'
0*
b110 +
#655960000000
1"
1(
#655970000000
0!
0"
b100 &
0'
0(
b100 ,
#655980000000
1!
1$
b111 %
1'
1*
b111 +
#655990000000
0!
0'
#656000000000
1!
0$
b1000 %
1'
0*
b1000 +
#656010000000
0!
0'
#656020000000
1!
b1001 %
1'
b1001 +
#656030000000
0!
0'
#656040000000
1!
b0 %
1'
b0 +
#656050000000
0!
0'
#656060000000
1!
1$
b1 %
1'
1*
b1 +
#656070000000
0!
0'
#656080000000
1!
b10 %
1'
b10 +
#656090000000
0!
0'
#656100000000
1!
b11 %
1'
b11 +
#656110000000
0!
0'
#656120000000
1!
b100 %
1'
b100 +
#656130000000
0!
0'
#656140000000
1!
b101 %
1'
b101 +
#656150000000
0!
0'
#656160000000
1!
b110 %
1'
b110 +
#656170000000
0!
0'
#656180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#656190000000
0!
0'
#656200000000
1!
b1000 %
1'
b1000 +
#656210000000
0!
0'
#656220000000
1!
b1001 %
1'
b1001 +
#656230000000
0!
0'
#656240000000
1!
b0 %
1'
b0 +
#656250000000
0!
0'
#656260000000
1!
1$
b1 %
1'
1*
b1 +
#656270000000
0!
0'
#656280000000
1!
b10 %
1'
b10 +
#656290000000
0!
0'
#656300000000
1!
b11 %
1'
b11 +
#656310000000
0!
0'
#656320000000
1!
b100 %
1'
b100 +
#656330000000
0!
0'
#656340000000
1!
b101 %
1'
b101 +
#656350000000
0!
0'
#656360000000
1!
0$
b110 %
1'
0*
b110 +
#656370000000
0!
0'
#656380000000
1!
b111 %
1'
b111 +
#656390000000
1"
1(
#656400000000
0!
0"
b100 &
0'
0(
b100 ,
#656410000000
1!
b1000 %
1'
b1000 +
#656420000000
0!
0'
#656430000000
1!
b1001 %
1'
b1001 +
#656440000000
0!
0'
#656450000000
1!
b0 %
1'
b0 +
#656460000000
0!
0'
#656470000000
1!
1$
b1 %
1'
1*
b1 +
#656480000000
0!
0'
#656490000000
1!
b10 %
1'
b10 +
#656500000000
0!
0'
#656510000000
1!
b11 %
1'
b11 +
#656520000000
0!
0'
#656530000000
1!
b100 %
1'
b100 +
#656540000000
0!
0'
#656550000000
1!
b101 %
1'
b101 +
#656560000000
0!
0'
#656570000000
1!
b110 %
1'
b110 +
#656580000000
0!
0'
#656590000000
1!
b111 %
1'
b111 +
#656600000000
0!
0'
#656610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#656620000000
0!
0'
#656630000000
1!
b1001 %
1'
b1001 +
#656640000000
0!
0'
#656650000000
1!
b0 %
1'
b0 +
#656660000000
0!
0'
#656670000000
1!
1$
b1 %
1'
1*
b1 +
#656680000000
0!
0'
#656690000000
1!
b10 %
1'
b10 +
#656700000000
0!
0'
#656710000000
1!
b11 %
1'
b11 +
#656720000000
0!
0'
#656730000000
1!
b100 %
1'
b100 +
#656740000000
0!
0'
#656750000000
1!
b101 %
1'
b101 +
#656760000000
0!
0'
#656770000000
1!
0$
b110 %
1'
0*
b110 +
#656780000000
0!
0'
#656790000000
1!
b111 %
1'
b111 +
#656800000000
0!
0'
#656810000000
1!
b1000 %
1'
b1000 +
#656820000000
1"
1(
#656830000000
0!
0"
b100 &
0'
0(
b100 ,
#656840000000
1!
b1001 %
1'
b1001 +
#656850000000
0!
0'
#656860000000
1!
b0 %
1'
b0 +
#656870000000
0!
0'
#656880000000
1!
1$
b1 %
1'
1*
b1 +
#656890000000
0!
0'
#656900000000
1!
b10 %
1'
b10 +
#656910000000
0!
0'
#656920000000
1!
b11 %
1'
b11 +
#656930000000
0!
0'
#656940000000
1!
b100 %
1'
b100 +
#656950000000
0!
0'
#656960000000
1!
b101 %
1'
b101 +
#656970000000
0!
0'
#656980000000
1!
b110 %
1'
b110 +
#656990000000
0!
0'
#657000000000
1!
b111 %
1'
b111 +
#657010000000
0!
0'
#657020000000
1!
0$
b1000 %
1'
0*
b1000 +
#657030000000
0!
0'
#657040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#657050000000
0!
0'
#657060000000
1!
b0 %
1'
b0 +
#657070000000
0!
0'
#657080000000
1!
1$
b1 %
1'
1*
b1 +
#657090000000
0!
0'
#657100000000
1!
b10 %
1'
b10 +
#657110000000
0!
0'
#657120000000
1!
b11 %
1'
b11 +
#657130000000
0!
0'
#657140000000
1!
b100 %
1'
b100 +
#657150000000
0!
0'
#657160000000
1!
b101 %
1'
b101 +
#657170000000
0!
0'
#657180000000
1!
0$
b110 %
1'
0*
b110 +
#657190000000
0!
0'
#657200000000
1!
b111 %
1'
b111 +
#657210000000
0!
0'
#657220000000
1!
b1000 %
1'
b1000 +
#657230000000
0!
0'
#657240000000
1!
b1001 %
1'
b1001 +
#657250000000
1"
1(
#657260000000
0!
0"
b100 &
0'
0(
b100 ,
#657270000000
1!
b0 %
1'
b0 +
#657280000000
0!
0'
#657290000000
1!
1$
b1 %
1'
1*
b1 +
#657300000000
0!
0'
#657310000000
1!
b10 %
1'
b10 +
#657320000000
0!
0'
#657330000000
1!
b11 %
1'
b11 +
#657340000000
0!
0'
#657350000000
1!
b100 %
1'
b100 +
#657360000000
0!
0'
#657370000000
1!
b101 %
1'
b101 +
#657380000000
0!
0'
#657390000000
1!
b110 %
1'
b110 +
#657400000000
0!
0'
#657410000000
1!
b111 %
1'
b111 +
#657420000000
0!
0'
#657430000000
1!
0$
b1000 %
1'
0*
b1000 +
#657440000000
0!
0'
#657450000000
1!
b1001 %
1'
b1001 +
#657460000000
0!
0'
#657470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#657480000000
0!
0'
#657490000000
1!
1$
b1 %
1'
1*
b1 +
#657500000000
0!
0'
#657510000000
1!
b10 %
1'
b10 +
#657520000000
0!
0'
#657530000000
1!
b11 %
1'
b11 +
#657540000000
0!
0'
#657550000000
1!
b100 %
1'
b100 +
#657560000000
0!
0'
#657570000000
1!
b101 %
1'
b101 +
#657580000000
0!
0'
#657590000000
1!
0$
b110 %
1'
0*
b110 +
#657600000000
0!
0'
#657610000000
1!
b111 %
1'
b111 +
#657620000000
0!
0'
#657630000000
1!
b1000 %
1'
b1000 +
#657640000000
0!
0'
#657650000000
1!
b1001 %
1'
b1001 +
#657660000000
0!
0'
#657670000000
1!
b0 %
1'
b0 +
#657680000000
1"
1(
#657690000000
0!
0"
b100 &
0'
0(
b100 ,
#657700000000
1!
1$
b1 %
1'
1*
b1 +
#657710000000
0!
0'
#657720000000
1!
b10 %
1'
b10 +
#657730000000
0!
0'
#657740000000
1!
b11 %
1'
b11 +
#657750000000
0!
0'
#657760000000
1!
b100 %
1'
b100 +
#657770000000
0!
0'
#657780000000
1!
b101 %
1'
b101 +
#657790000000
0!
0'
#657800000000
1!
b110 %
1'
b110 +
#657810000000
0!
0'
#657820000000
1!
b111 %
1'
b111 +
#657830000000
0!
0'
#657840000000
1!
0$
b1000 %
1'
0*
b1000 +
#657850000000
0!
0'
#657860000000
1!
b1001 %
1'
b1001 +
#657870000000
0!
0'
#657880000000
1!
b0 %
1'
b0 +
#657890000000
0!
0'
#657900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#657910000000
0!
0'
#657920000000
1!
b10 %
1'
b10 +
#657930000000
0!
0'
#657940000000
1!
b11 %
1'
b11 +
#657950000000
0!
0'
#657960000000
1!
b100 %
1'
b100 +
#657970000000
0!
0'
#657980000000
1!
b101 %
1'
b101 +
#657990000000
0!
0'
#658000000000
1!
0$
b110 %
1'
0*
b110 +
#658010000000
0!
0'
#658020000000
1!
b111 %
1'
b111 +
#658030000000
0!
0'
#658040000000
1!
b1000 %
1'
b1000 +
#658050000000
0!
0'
#658060000000
1!
b1001 %
1'
b1001 +
#658070000000
0!
0'
#658080000000
1!
b0 %
1'
b0 +
#658090000000
0!
0'
#658100000000
1!
1$
b1 %
1'
1*
b1 +
#658110000000
1"
1(
#658120000000
0!
0"
b100 &
0'
0(
b100 ,
#658130000000
1!
b10 %
1'
b10 +
#658140000000
0!
0'
#658150000000
1!
b11 %
1'
b11 +
#658160000000
0!
0'
#658170000000
1!
b100 %
1'
b100 +
#658180000000
0!
0'
#658190000000
1!
b101 %
1'
b101 +
#658200000000
0!
0'
#658210000000
1!
b110 %
1'
b110 +
#658220000000
0!
0'
#658230000000
1!
b111 %
1'
b111 +
#658240000000
0!
0'
#658250000000
1!
0$
b1000 %
1'
0*
b1000 +
#658260000000
0!
0'
#658270000000
1!
b1001 %
1'
b1001 +
#658280000000
0!
0'
#658290000000
1!
b0 %
1'
b0 +
#658300000000
0!
0'
#658310000000
1!
1$
b1 %
1'
1*
b1 +
#658320000000
0!
0'
#658330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#658340000000
0!
0'
#658350000000
1!
b11 %
1'
b11 +
#658360000000
0!
0'
#658370000000
1!
b100 %
1'
b100 +
#658380000000
0!
0'
#658390000000
1!
b101 %
1'
b101 +
#658400000000
0!
0'
#658410000000
1!
0$
b110 %
1'
0*
b110 +
#658420000000
0!
0'
#658430000000
1!
b111 %
1'
b111 +
#658440000000
0!
0'
#658450000000
1!
b1000 %
1'
b1000 +
#658460000000
0!
0'
#658470000000
1!
b1001 %
1'
b1001 +
#658480000000
0!
0'
#658490000000
1!
b0 %
1'
b0 +
#658500000000
0!
0'
#658510000000
1!
1$
b1 %
1'
1*
b1 +
#658520000000
0!
0'
#658530000000
1!
b10 %
1'
b10 +
#658540000000
1"
1(
#658550000000
0!
0"
b100 &
0'
0(
b100 ,
#658560000000
1!
b11 %
1'
b11 +
#658570000000
0!
0'
#658580000000
1!
b100 %
1'
b100 +
#658590000000
0!
0'
#658600000000
1!
b101 %
1'
b101 +
#658610000000
0!
0'
#658620000000
1!
b110 %
1'
b110 +
#658630000000
0!
0'
#658640000000
1!
b111 %
1'
b111 +
#658650000000
0!
0'
#658660000000
1!
0$
b1000 %
1'
0*
b1000 +
#658670000000
0!
0'
#658680000000
1!
b1001 %
1'
b1001 +
#658690000000
0!
0'
#658700000000
1!
b0 %
1'
b0 +
#658710000000
0!
0'
#658720000000
1!
1$
b1 %
1'
1*
b1 +
#658730000000
0!
0'
#658740000000
1!
b10 %
1'
b10 +
#658750000000
0!
0'
#658760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#658770000000
0!
0'
#658780000000
1!
b100 %
1'
b100 +
#658790000000
0!
0'
#658800000000
1!
b101 %
1'
b101 +
#658810000000
0!
0'
#658820000000
1!
0$
b110 %
1'
0*
b110 +
#658830000000
0!
0'
#658840000000
1!
b111 %
1'
b111 +
#658850000000
0!
0'
#658860000000
1!
b1000 %
1'
b1000 +
#658870000000
0!
0'
#658880000000
1!
b1001 %
1'
b1001 +
#658890000000
0!
0'
#658900000000
1!
b0 %
1'
b0 +
#658910000000
0!
0'
#658920000000
1!
1$
b1 %
1'
1*
b1 +
#658930000000
0!
0'
#658940000000
1!
b10 %
1'
b10 +
#658950000000
0!
0'
#658960000000
1!
b11 %
1'
b11 +
#658970000000
1"
1(
#658980000000
0!
0"
b100 &
0'
0(
b100 ,
#658990000000
1!
b100 %
1'
b100 +
#659000000000
0!
0'
#659010000000
1!
b101 %
1'
b101 +
#659020000000
0!
0'
#659030000000
1!
b110 %
1'
b110 +
#659040000000
0!
0'
#659050000000
1!
b111 %
1'
b111 +
#659060000000
0!
0'
#659070000000
1!
0$
b1000 %
1'
0*
b1000 +
#659080000000
0!
0'
#659090000000
1!
b1001 %
1'
b1001 +
#659100000000
0!
0'
#659110000000
1!
b0 %
1'
b0 +
#659120000000
0!
0'
#659130000000
1!
1$
b1 %
1'
1*
b1 +
#659140000000
0!
0'
#659150000000
1!
b10 %
1'
b10 +
#659160000000
0!
0'
#659170000000
1!
b11 %
1'
b11 +
#659180000000
0!
0'
#659190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#659200000000
0!
0'
#659210000000
1!
b101 %
1'
b101 +
#659220000000
0!
0'
#659230000000
1!
0$
b110 %
1'
0*
b110 +
#659240000000
0!
0'
#659250000000
1!
b111 %
1'
b111 +
#659260000000
0!
0'
#659270000000
1!
b1000 %
1'
b1000 +
#659280000000
0!
0'
#659290000000
1!
b1001 %
1'
b1001 +
#659300000000
0!
0'
#659310000000
1!
b0 %
1'
b0 +
#659320000000
0!
0'
#659330000000
1!
1$
b1 %
1'
1*
b1 +
#659340000000
0!
0'
#659350000000
1!
b10 %
1'
b10 +
#659360000000
0!
0'
#659370000000
1!
b11 %
1'
b11 +
#659380000000
0!
0'
#659390000000
1!
b100 %
1'
b100 +
#659400000000
1"
1(
#659410000000
0!
0"
b100 &
0'
0(
b100 ,
#659420000000
1!
b101 %
1'
b101 +
#659430000000
0!
0'
#659440000000
1!
b110 %
1'
b110 +
#659450000000
0!
0'
#659460000000
1!
b111 %
1'
b111 +
#659470000000
0!
0'
#659480000000
1!
0$
b1000 %
1'
0*
b1000 +
#659490000000
0!
0'
#659500000000
1!
b1001 %
1'
b1001 +
#659510000000
0!
0'
#659520000000
1!
b0 %
1'
b0 +
#659530000000
0!
0'
#659540000000
1!
1$
b1 %
1'
1*
b1 +
#659550000000
0!
0'
#659560000000
1!
b10 %
1'
b10 +
#659570000000
0!
0'
#659580000000
1!
b11 %
1'
b11 +
#659590000000
0!
0'
#659600000000
1!
b100 %
1'
b100 +
#659610000000
0!
0'
#659620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#659630000000
0!
0'
#659640000000
1!
0$
b110 %
1'
0*
b110 +
#659650000000
0!
0'
#659660000000
1!
b111 %
1'
b111 +
#659670000000
0!
0'
#659680000000
1!
b1000 %
1'
b1000 +
#659690000000
0!
0'
#659700000000
1!
b1001 %
1'
b1001 +
#659710000000
0!
0'
#659720000000
1!
b0 %
1'
b0 +
#659730000000
0!
0'
#659740000000
1!
1$
b1 %
1'
1*
b1 +
#659750000000
0!
0'
#659760000000
1!
b10 %
1'
b10 +
#659770000000
0!
0'
#659780000000
1!
b11 %
1'
b11 +
#659790000000
0!
0'
#659800000000
1!
b100 %
1'
b100 +
#659810000000
0!
0'
#659820000000
1!
b101 %
1'
b101 +
#659830000000
1"
1(
#659840000000
0!
0"
b100 &
0'
0(
b100 ,
#659850000000
1!
b110 %
1'
b110 +
#659860000000
0!
0'
#659870000000
1!
b111 %
1'
b111 +
#659880000000
0!
0'
#659890000000
1!
0$
b1000 %
1'
0*
b1000 +
#659900000000
0!
0'
#659910000000
1!
b1001 %
1'
b1001 +
#659920000000
0!
0'
#659930000000
1!
b0 %
1'
b0 +
#659940000000
0!
0'
#659950000000
1!
1$
b1 %
1'
1*
b1 +
#659960000000
0!
0'
#659970000000
1!
b10 %
1'
b10 +
#659980000000
0!
0'
#659990000000
1!
b11 %
1'
b11 +
#660000000000
0!
0'
#660010000000
1!
b100 %
1'
b100 +
#660020000000
0!
0'
#660030000000
1!
b101 %
1'
b101 +
#660040000000
0!
0'
#660050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#660060000000
0!
0'
#660070000000
1!
b111 %
1'
b111 +
#660080000000
0!
0'
#660090000000
1!
b1000 %
1'
b1000 +
#660100000000
0!
0'
#660110000000
1!
b1001 %
1'
b1001 +
#660120000000
0!
0'
#660130000000
1!
b0 %
1'
b0 +
#660140000000
0!
0'
#660150000000
1!
1$
b1 %
1'
1*
b1 +
#660160000000
0!
0'
#660170000000
1!
b10 %
1'
b10 +
#660180000000
0!
0'
#660190000000
1!
b11 %
1'
b11 +
#660200000000
0!
0'
#660210000000
1!
b100 %
1'
b100 +
#660220000000
0!
0'
#660230000000
1!
b101 %
1'
b101 +
#660240000000
0!
0'
#660250000000
1!
0$
b110 %
1'
0*
b110 +
#660260000000
1"
1(
#660270000000
0!
0"
b100 &
0'
0(
b100 ,
#660280000000
1!
1$
b111 %
1'
1*
b111 +
#660290000000
0!
0'
#660300000000
1!
0$
b1000 %
1'
0*
b1000 +
#660310000000
0!
0'
#660320000000
1!
b1001 %
1'
b1001 +
#660330000000
0!
0'
#660340000000
1!
b0 %
1'
b0 +
#660350000000
0!
0'
#660360000000
1!
1$
b1 %
1'
1*
b1 +
#660370000000
0!
0'
#660380000000
1!
b10 %
1'
b10 +
#660390000000
0!
0'
#660400000000
1!
b11 %
1'
b11 +
#660410000000
0!
0'
#660420000000
1!
b100 %
1'
b100 +
#660430000000
0!
0'
#660440000000
1!
b101 %
1'
b101 +
#660450000000
0!
0'
#660460000000
1!
b110 %
1'
b110 +
#660470000000
0!
0'
#660480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#660490000000
0!
0'
#660500000000
1!
b1000 %
1'
b1000 +
#660510000000
0!
0'
#660520000000
1!
b1001 %
1'
b1001 +
#660530000000
0!
0'
#660540000000
1!
b0 %
1'
b0 +
#660550000000
0!
0'
#660560000000
1!
1$
b1 %
1'
1*
b1 +
#660570000000
0!
0'
#660580000000
1!
b10 %
1'
b10 +
#660590000000
0!
0'
#660600000000
1!
b11 %
1'
b11 +
#660610000000
0!
0'
#660620000000
1!
b100 %
1'
b100 +
#660630000000
0!
0'
#660640000000
1!
b101 %
1'
b101 +
#660650000000
0!
0'
#660660000000
1!
0$
b110 %
1'
0*
b110 +
#660670000000
0!
0'
#660680000000
1!
b111 %
1'
b111 +
#660690000000
1"
1(
#660700000000
0!
0"
b100 &
0'
0(
b100 ,
#660710000000
1!
b1000 %
1'
b1000 +
#660720000000
0!
0'
#660730000000
1!
b1001 %
1'
b1001 +
#660740000000
0!
0'
#660750000000
1!
b0 %
1'
b0 +
#660760000000
0!
0'
#660770000000
1!
1$
b1 %
1'
1*
b1 +
#660780000000
0!
0'
#660790000000
1!
b10 %
1'
b10 +
#660800000000
0!
0'
#660810000000
1!
b11 %
1'
b11 +
#660820000000
0!
0'
#660830000000
1!
b100 %
1'
b100 +
#660840000000
0!
0'
#660850000000
1!
b101 %
1'
b101 +
#660860000000
0!
0'
#660870000000
1!
b110 %
1'
b110 +
#660880000000
0!
0'
#660890000000
1!
b111 %
1'
b111 +
#660900000000
0!
0'
#660910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#660920000000
0!
0'
#660930000000
1!
b1001 %
1'
b1001 +
#660940000000
0!
0'
#660950000000
1!
b0 %
1'
b0 +
#660960000000
0!
0'
#660970000000
1!
1$
b1 %
1'
1*
b1 +
#660980000000
0!
0'
#660990000000
1!
b10 %
1'
b10 +
#661000000000
0!
0'
#661010000000
1!
b11 %
1'
b11 +
#661020000000
0!
0'
#661030000000
1!
b100 %
1'
b100 +
#661040000000
0!
0'
#661050000000
1!
b101 %
1'
b101 +
#661060000000
0!
0'
#661070000000
1!
0$
b110 %
1'
0*
b110 +
#661080000000
0!
0'
#661090000000
1!
b111 %
1'
b111 +
#661100000000
0!
0'
#661110000000
1!
b1000 %
1'
b1000 +
#661120000000
1"
1(
#661130000000
0!
0"
b100 &
0'
0(
b100 ,
#661140000000
1!
b1001 %
1'
b1001 +
#661150000000
0!
0'
#661160000000
1!
b0 %
1'
b0 +
#661170000000
0!
0'
#661180000000
1!
1$
b1 %
1'
1*
b1 +
#661190000000
0!
0'
#661200000000
1!
b10 %
1'
b10 +
#661210000000
0!
0'
#661220000000
1!
b11 %
1'
b11 +
#661230000000
0!
0'
#661240000000
1!
b100 %
1'
b100 +
#661250000000
0!
0'
#661260000000
1!
b101 %
1'
b101 +
#661270000000
0!
0'
#661280000000
1!
b110 %
1'
b110 +
#661290000000
0!
0'
#661300000000
1!
b111 %
1'
b111 +
#661310000000
0!
0'
#661320000000
1!
0$
b1000 %
1'
0*
b1000 +
#661330000000
0!
0'
#661340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#661350000000
0!
0'
#661360000000
1!
b0 %
1'
b0 +
#661370000000
0!
0'
#661380000000
1!
1$
b1 %
1'
1*
b1 +
#661390000000
0!
0'
#661400000000
1!
b10 %
1'
b10 +
#661410000000
0!
0'
#661420000000
1!
b11 %
1'
b11 +
#661430000000
0!
0'
#661440000000
1!
b100 %
1'
b100 +
#661450000000
0!
0'
#661460000000
1!
b101 %
1'
b101 +
#661470000000
0!
0'
#661480000000
1!
0$
b110 %
1'
0*
b110 +
#661490000000
0!
0'
#661500000000
1!
b111 %
1'
b111 +
#661510000000
0!
0'
#661520000000
1!
b1000 %
1'
b1000 +
#661530000000
0!
0'
#661540000000
1!
b1001 %
1'
b1001 +
#661550000000
1"
1(
#661560000000
0!
0"
b100 &
0'
0(
b100 ,
#661570000000
1!
b0 %
1'
b0 +
#661580000000
0!
0'
#661590000000
1!
1$
b1 %
1'
1*
b1 +
#661600000000
0!
0'
#661610000000
1!
b10 %
1'
b10 +
#661620000000
0!
0'
#661630000000
1!
b11 %
1'
b11 +
#661640000000
0!
0'
#661650000000
1!
b100 %
1'
b100 +
#661660000000
0!
0'
#661670000000
1!
b101 %
1'
b101 +
#661680000000
0!
0'
#661690000000
1!
b110 %
1'
b110 +
#661700000000
0!
0'
#661710000000
1!
b111 %
1'
b111 +
#661720000000
0!
0'
#661730000000
1!
0$
b1000 %
1'
0*
b1000 +
#661740000000
0!
0'
#661750000000
1!
b1001 %
1'
b1001 +
#661760000000
0!
0'
#661770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#661780000000
0!
0'
#661790000000
1!
1$
b1 %
1'
1*
b1 +
#661800000000
0!
0'
#661810000000
1!
b10 %
1'
b10 +
#661820000000
0!
0'
#661830000000
1!
b11 %
1'
b11 +
#661840000000
0!
0'
#661850000000
1!
b100 %
1'
b100 +
#661860000000
0!
0'
#661870000000
1!
b101 %
1'
b101 +
#661880000000
0!
0'
#661890000000
1!
0$
b110 %
1'
0*
b110 +
#661900000000
0!
0'
#661910000000
1!
b111 %
1'
b111 +
#661920000000
0!
0'
#661930000000
1!
b1000 %
1'
b1000 +
#661940000000
0!
0'
#661950000000
1!
b1001 %
1'
b1001 +
#661960000000
0!
0'
#661970000000
1!
b0 %
1'
b0 +
#661980000000
1"
1(
#661990000000
0!
0"
b100 &
0'
0(
b100 ,
#662000000000
1!
1$
b1 %
1'
1*
b1 +
#662010000000
0!
0'
#662020000000
1!
b10 %
1'
b10 +
#662030000000
0!
0'
#662040000000
1!
b11 %
1'
b11 +
#662050000000
0!
0'
#662060000000
1!
b100 %
1'
b100 +
#662070000000
0!
0'
#662080000000
1!
b101 %
1'
b101 +
#662090000000
0!
0'
#662100000000
1!
b110 %
1'
b110 +
#662110000000
0!
0'
#662120000000
1!
b111 %
1'
b111 +
#662130000000
0!
0'
#662140000000
1!
0$
b1000 %
1'
0*
b1000 +
#662150000000
0!
0'
#662160000000
1!
b1001 %
1'
b1001 +
#662170000000
0!
0'
#662180000000
1!
b0 %
1'
b0 +
#662190000000
0!
0'
#662200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#662210000000
0!
0'
#662220000000
1!
b10 %
1'
b10 +
#662230000000
0!
0'
#662240000000
1!
b11 %
1'
b11 +
#662250000000
0!
0'
#662260000000
1!
b100 %
1'
b100 +
#662270000000
0!
0'
#662280000000
1!
b101 %
1'
b101 +
#662290000000
0!
0'
#662300000000
1!
0$
b110 %
1'
0*
b110 +
#662310000000
0!
0'
#662320000000
1!
b111 %
1'
b111 +
#662330000000
0!
0'
#662340000000
1!
b1000 %
1'
b1000 +
#662350000000
0!
0'
#662360000000
1!
b1001 %
1'
b1001 +
#662370000000
0!
0'
#662380000000
1!
b0 %
1'
b0 +
#662390000000
0!
0'
#662400000000
1!
1$
b1 %
1'
1*
b1 +
#662410000000
1"
1(
#662420000000
0!
0"
b100 &
0'
0(
b100 ,
#662430000000
1!
b10 %
1'
b10 +
#662440000000
0!
0'
#662450000000
1!
b11 %
1'
b11 +
#662460000000
0!
0'
#662470000000
1!
b100 %
1'
b100 +
#662480000000
0!
0'
#662490000000
1!
b101 %
1'
b101 +
#662500000000
0!
0'
#662510000000
1!
b110 %
1'
b110 +
#662520000000
0!
0'
#662530000000
1!
b111 %
1'
b111 +
#662540000000
0!
0'
#662550000000
1!
0$
b1000 %
1'
0*
b1000 +
#662560000000
0!
0'
#662570000000
1!
b1001 %
1'
b1001 +
#662580000000
0!
0'
#662590000000
1!
b0 %
1'
b0 +
#662600000000
0!
0'
#662610000000
1!
1$
b1 %
1'
1*
b1 +
#662620000000
0!
0'
#662630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#662640000000
0!
0'
#662650000000
1!
b11 %
1'
b11 +
#662660000000
0!
0'
#662670000000
1!
b100 %
1'
b100 +
#662680000000
0!
0'
#662690000000
1!
b101 %
1'
b101 +
#662700000000
0!
0'
#662710000000
1!
0$
b110 %
1'
0*
b110 +
#662720000000
0!
0'
#662730000000
1!
b111 %
1'
b111 +
#662740000000
0!
0'
#662750000000
1!
b1000 %
1'
b1000 +
#662760000000
0!
0'
#662770000000
1!
b1001 %
1'
b1001 +
#662780000000
0!
0'
#662790000000
1!
b0 %
1'
b0 +
#662800000000
0!
0'
#662810000000
1!
1$
b1 %
1'
1*
b1 +
#662820000000
0!
0'
#662830000000
1!
b10 %
1'
b10 +
#662840000000
1"
1(
#662850000000
0!
0"
b100 &
0'
0(
b100 ,
#662860000000
1!
b11 %
1'
b11 +
#662870000000
0!
0'
#662880000000
1!
b100 %
1'
b100 +
#662890000000
0!
0'
#662900000000
1!
b101 %
1'
b101 +
#662910000000
0!
0'
#662920000000
1!
b110 %
1'
b110 +
#662930000000
0!
0'
#662940000000
1!
b111 %
1'
b111 +
#662950000000
0!
0'
#662960000000
1!
0$
b1000 %
1'
0*
b1000 +
#662970000000
0!
0'
#662980000000
1!
b1001 %
1'
b1001 +
#662990000000
0!
0'
#663000000000
1!
b0 %
1'
b0 +
#663010000000
0!
0'
#663020000000
1!
1$
b1 %
1'
1*
b1 +
#663030000000
0!
0'
#663040000000
1!
b10 %
1'
b10 +
#663050000000
0!
0'
#663060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#663070000000
0!
0'
#663080000000
1!
b100 %
1'
b100 +
#663090000000
0!
0'
#663100000000
1!
b101 %
1'
b101 +
#663110000000
0!
0'
#663120000000
1!
0$
b110 %
1'
0*
b110 +
#663130000000
0!
0'
#663140000000
1!
b111 %
1'
b111 +
#663150000000
0!
0'
#663160000000
1!
b1000 %
1'
b1000 +
#663170000000
0!
0'
#663180000000
1!
b1001 %
1'
b1001 +
#663190000000
0!
0'
#663200000000
1!
b0 %
1'
b0 +
#663210000000
0!
0'
#663220000000
1!
1$
b1 %
1'
1*
b1 +
#663230000000
0!
0'
#663240000000
1!
b10 %
1'
b10 +
#663250000000
0!
0'
#663260000000
1!
b11 %
1'
b11 +
#663270000000
1"
1(
#663280000000
0!
0"
b100 &
0'
0(
b100 ,
#663290000000
1!
b100 %
1'
b100 +
#663300000000
0!
0'
#663310000000
1!
b101 %
1'
b101 +
#663320000000
0!
0'
#663330000000
1!
b110 %
1'
b110 +
#663340000000
0!
0'
#663350000000
1!
b111 %
1'
b111 +
#663360000000
0!
0'
#663370000000
1!
0$
b1000 %
1'
0*
b1000 +
#663380000000
0!
0'
#663390000000
1!
b1001 %
1'
b1001 +
#663400000000
0!
0'
#663410000000
1!
b0 %
1'
b0 +
#663420000000
0!
0'
#663430000000
1!
1$
b1 %
1'
1*
b1 +
#663440000000
0!
0'
#663450000000
1!
b10 %
1'
b10 +
#663460000000
0!
0'
#663470000000
1!
b11 %
1'
b11 +
#663480000000
0!
0'
#663490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#663500000000
0!
0'
#663510000000
1!
b101 %
1'
b101 +
#663520000000
0!
0'
#663530000000
1!
0$
b110 %
1'
0*
b110 +
#663540000000
0!
0'
#663550000000
1!
b111 %
1'
b111 +
#663560000000
0!
0'
#663570000000
1!
b1000 %
1'
b1000 +
#663580000000
0!
0'
#663590000000
1!
b1001 %
1'
b1001 +
#663600000000
0!
0'
#663610000000
1!
b0 %
1'
b0 +
#663620000000
0!
0'
#663630000000
1!
1$
b1 %
1'
1*
b1 +
#663640000000
0!
0'
#663650000000
1!
b10 %
1'
b10 +
#663660000000
0!
0'
#663670000000
1!
b11 %
1'
b11 +
#663680000000
0!
0'
#663690000000
1!
b100 %
1'
b100 +
#663700000000
1"
1(
#663710000000
0!
0"
b100 &
0'
0(
b100 ,
#663720000000
1!
b101 %
1'
b101 +
#663730000000
0!
0'
#663740000000
1!
b110 %
1'
b110 +
#663750000000
0!
0'
#663760000000
1!
b111 %
1'
b111 +
#663770000000
0!
0'
#663780000000
1!
0$
b1000 %
1'
0*
b1000 +
#663790000000
0!
0'
#663800000000
1!
b1001 %
1'
b1001 +
#663810000000
0!
0'
#663820000000
1!
b0 %
1'
b0 +
#663830000000
0!
0'
#663840000000
1!
1$
b1 %
1'
1*
b1 +
#663850000000
0!
0'
#663860000000
1!
b10 %
1'
b10 +
#663870000000
0!
0'
#663880000000
1!
b11 %
1'
b11 +
#663890000000
0!
0'
#663900000000
1!
b100 %
1'
b100 +
#663910000000
0!
0'
#663920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#663930000000
0!
0'
#663940000000
1!
0$
b110 %
1'
0*
b110 +
#663950000000
0!
0'
#663960000000
1!
b111 %
1'
b111 +
#663970000000
0!
0'
#663980000000
1!
b1000 %
1'
b1000 +
#663990000000
0!
0'
#664000000000
1!
b1001 %
1'
b1001 +
#664010000000
0!
0'
#664020000000
1!
b0 %
1'
b0 +
#664030000000
0!
0'
#664040000000
1!
1$
b1 %
1'
1*
b1 +
#664050000000
0!
0'
#664060000000
1!
b10 %
1'
b10 +
#664070000000
0!
0'
#664080000000
1!
b11 %
1'
b11 +
#664090000000
0!
0'
#664100000000
1!
b100 %
1'
b100 +
#664110000000
0!
0'
#664120000000
1!
b101 %
1'
b101 +
#664130000000
1"
1(
#664140000000
0!
0"
b100 &
0'
0(
b100 ,
#664150000000
1!
b110 %
1'
b110 +
#664160000000
0!
0'
#664170000000
1!
b111 %
1'
b111 +
#664180000000
0!
0'
#664190000000
1!
0$
b1000 %
1'
0*
b1000 +
#664200000000
0!
0'
#664210000000
1!
b1001 %
1'
b1001 +
#664220000000
0!
0'
#664230000000
1!
b0 %
1'
b0 +
#664240000000
0!
0'
#664250000000
1!
1$
b1 %
1'
1*
b1 +
#664260000000
0!
0'
#664270000000
1!
b10 %
1'
b10 +
#664280000000
0!
0'
#664290000000
1!
b11 %
1'
b11 +
#664300000000
0!
0'
#664310000000
1!
b100 %
1'
b100 +
#664320000000
0!
0'
#664330000000
1!
b101 %
1'
b101 +
#664340000000
0!
0'
#664350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#664360000000
0!
0'
#664370000000
1!
b111 %
1'
b111 +
#664380000000
0!
0'
#664390000000
1!
b1000 %
1'
b1000 +
#664400000000
0!
0'
#664410000000
1!
b1001 %
1'
b1001 +
#664420000000
0!
0'
#664430000000
1!
b0 %
1'
b0 +
#664440000000
0!
0'
#664450000000
1!
1$
b1 %
1'
1*
b1 +
#664460000000
0!
0'
#664470000000
1!
b10 %
1'
b10 +
#664480000000
0!
0'
#664490000000
1!
b11 %
1'
b11 +
#664500000000
0!
0'
#664510000000
1!
b100 %
1'
b100 +
#664520000000
0!
0'
#664530000000
1!
b101 %
1'
b101 +
#664540000000
0!
0'
#664550000000
1!
0$
b110 %
1'
0*
b110 +
#664560000000
1"
1(
#664570000000
0!
0"
b100 &
0'
0(
b100 ,
#664580000000
1!
1$
b111 %
1'
1*
b111 +
#664590000000
0!
0'
#664600000000
1!
0$
b1000 %
1'
0*
b1000 +
#664610000000
0!
0'
#664620000000
1!
b1001 %
1'
b1001 +
#664630000000
0!
0'
#664640000000
1!
b0 %
1'
b0 +
#664650000000
0!
0'
#664660000000
1!
1$
b1 %
1'
1*
b1 +
#664670000000
0!
0'
#664680000000
1!
b10 %
1'
b10 +
#664690000000
0!
0'
#664700000000
1!
b11 %
1'
b11 +
#664710000000
0!
0'
#664720000000
1!
b100 %
1'
b100 +
#664730000000
0!
0'
#664740000000
1!
b101 %
1'
b101 +
#664750000000
0!
0'
#664760000000
1!
b110 %
1'
b110 +
#664770000000
0!
0'
#664780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#664790000000
0!
0'
#664800000000
1!
b1000 %
1'
b1000 +
#664810000000
0!
0'
#664820000000
1!
b1001 %
1'
b1001 +
#664830000000
0!
0'
#664840000000
1!
b0 %
1'
b0 +
#664850000000
0!
0'
#664860000000
1!
1$
b1 %
1'
1*
b1 +
#664870000000
0!
0'
#664880000000
1!
b10 %
1'
b10 +
#664890000000
0!
0'
#664900000000
1!
b11 %
1'
b11 +
#664910000000
0!
0'
#664920000000
1!
b100 %
1'
b100 +
#664930000000
0!
0'
#664940000000
1!
b101 %
1'
b101 +
#664950000000
0!
0'
#664960000000
1!
0$
b110 %
1'
0*
b110 +
#664970000000
0!
0'
#664980000000
1!
b111 %
1'
b111 +
#664990000000
1"
1(
#665000000000
0!
0"
b100 &
0'
0(
b100 ,
#665010000000
1!
b1000 %
1'
b1000 +
#665020000000
0!
0'
#665030000000
1!
b1001 %
1'
b1001 +
#665040000000
0!
0'
#665050000000
1!
b0 %
1'
b0 +
#665060000000
0!
0'
#665070000000
1!
1$
b1 %
1'
1*
b1 +
#665080000000
0!
0'
#665090000000
1!
b10 %
1'
b10 +
#665100000000
0!
0'
#665110000000
1!
b11 %
1'
b11 +
#665120000000
0!
0'
#665130000000
1!
b100 %
1'
b100 +
#665140000000
0!
0'
#665150000000
1!
b101 %
1'
b101 +
#665160000000
0!
0'
#665170000000
1!
b110 %
1'
b110 +
#665180000000
0!
0'
#665190000000
1!
b111 %
1'
b111 +
#665200000000
0!
0'
#665210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#665220000000
0!
0'
#665230000000
1!
b1001 %
1'
b1001 +
#665240000000
0!
0'
#665250000000
1!
b0 %
1'
b0 +
#665260000000
0!
0'
#665270000000
1!
1$
b1 %
1'
1*
b1 +
#665280000000
0!
0'
#665290000000
1!
b10 %
1'
b10 +
#665300000000
0!
0'
#665310000000
1!
b11 %
1'
b11 +
#665320000000
0!
0'
#665330000000
1!
b100 %
1'
b100 +
#665340000000
0!
0'
#665350000000
1!
b101 %
1'
b101 +
#665360000000
0!
0'
#665370000000
1!
0$
b110 %
1'
0*
b110 +
#665380000000
0!
0'
#665390000000
1!
b111 %
1'
b111 +
#665400000000
0!
0'
#665410000000
1!
b1000 %
1'
b1000 +
#665420000000
1"
1(
#665430000000
0!
0"
b100 &
0'
0(
b100 ,
#665440000000
1!
b1001 %
1'
b1001 +
#665450000000
0!
0'
#665460000000
1!
b0 %
1'
b0 +
#665470000000
0!
0'
#665480000000
1!
1$
b1 %
1'
1*
b1 +
#665490000000
0!
0'
#665500000000
1!
b10 %
1'
b10 +
#665510000000
0!
0'
#665520000000
1!
b11 %
1'
b11 +
#665530000000
0!
0'
#665540000000
1!
b100 %
1'
b100 +
#665550000000
0!
0'
#665560000000
1!
b101 %
1'
b101 +
#665570000000
0!
0'
#665580000000
1!
b110 %
1'
b110 +
#665590000000
0!
0'
#665600000000
1!
b111 %
1'
b111 +
#665610000000
0!
0'
#665620000000
1!
0$
b1000 %
1'
0*
b1000 +
#665630000000
0!
0'
#665640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#665650000000
0!
0'
#665660000000
1!
b0 %
1'
b0 +
#665670000000
0!
0'
#665680000000
1!
1$
b1 %
1'
1*
b1 +
#665690000000
0!
0'
#665700000000
1!
b10 %
1'
b10 +
#665710000000
0!
0'
#665720000000
1!
b11 %
1'
b11 +
#665730000000
0!
0'
#665740000000
1!
b100 %
1'
b100 +
#665750000000
0!
0'
#665760000000
1!
b101 %
1'
b101 +
#665770000000
0!
0'
#665780000000
1!
0$
b110 %
1'
0*
b110 +
#665790000000
0!
0'
#665800000000
1!
b111 %
1'
b111 +
#665810000000
0!
0'
#665820000000
1!
b1000 %
1'
b1000 +
#665830000000
0!
0'
#665840000000
1!
b1001 %
1'
b1001 +
#665850000000
1"
1(
#665860000000
0!
0"
b100 &
0'
0(
b100 ,
#665870000000
1!
b0 %
1'
b0 +
#665880000000
0!
0'
#665890000000
1!
1$
b1 %
1'
1*
b1 +
#665900000000
0!
0'
#665910000000
1!
b10 %
1'
b10 +
#665920000000
0!
0'
#665930000000
1!
b11 %
1'
b11 +
#665940000000
0!
0'
#665950000000
1!
b100 %
1'
b100 +
#665960000000
0!
0'
#665970000000
1!
b101 %
1'
b101 +
#665980000000
0!
0'
#665990000000
1!
b110 %
1'
b110 +
#666000000000
0!
0'
#666010000000
1!
b111 %
1'
b111 +
#666020000000
0!
0'
#666030000000
1!
0$
b1000 %
1'
0*
b1000 +
#666040000000
0!
0'
#666050000000
1!
b1001 %
1'
b1001 +
#666060000000
0!
0'
#666070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#666080000000
0!
0'
#666090000000
1!
1$
b1 %
1'
1*
b1 +
#666100000000
0!
0'
#666110000000
1!
b10 %
1'
b10 +
#666120000000
0!
0'
#666130000000
1!
b11 %
1'
b11 +
#666140000000
0!
0'
#666150000000
1!
b100 %
1'
b100 +
#666160000000
0!
0'
#666170000000
1!
b101 %
1'
b101 +
#666180000000
0!
0'
#666190000000
1!
0$
b110 %
1'
0*
b110 +
#666200000000
0!
0'
#666210000000
1!
b111 %
1'
b111 +
#666220000000
0!
0'
#666230000000
1!
b1000 %
1'
b1000 +
#666240000000
0!
0'
#666250000000
1!
b1001 %
1'
b1001 +
#666260000000
0!
0'
#666270000000
1!
b0 %
1'
b0 +
#666280000000
1"
1(
#666290000000
0!
0"
b100 &
0'
0(
b100 ,
#666300000000
1!
1$
b1 %
1'
1*
b1 +
#666310000000
0!
0'
#666320000000
1!
b10 %
1'
b10 +
#666330000000
0!
0'
#666340000000
1!
b11 %
1'
b11 +
#666350000000
0!
0'
#666360000000
1!
b100 %
1'
b100 +
#666370000000
0!
0'
#666380000000
1!
b101 %
1'
b101 +
#666390000000
0!
0'
#666400000000
1!
b110 %
1'
b110 +
#666410000000
0!
0'
#666420000000
1!
b111 %
1'
b111 +
#666430000000
0!
0'
#666440000000
1!
0$
b1000 %
1'
0*
b1000 +
#666450000000
0!
0'
#666460000000
1!
b1001 %
1'
b1001 +
#666470000000
0!
0'
#666480000000
1!
b0 %
1'
b0 +
#666490000000
0!
0'
#666500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#666510000000
0!
0'
#666520000000
1!
b10 %
1'
b10 +
#666530000000
0!
0'
#666540000000
1!
b11 %
1'
b11 +
#666550000000
0!
0'
#666560000000
1!
b100 %
1'
b100 +
#666570000000
0!
0'
#666580000000
1!
b101 %
1'
b101 +
#666590000000
0!
0'
#666600000000
1!
0$
b110 %
1'
0*
b110 +
#666610000000
0!
0'
#666620000000
1!
b111 %
1'
b111 +
#666630000000
0!
0'
#666640000000
1!
b1000 %
1'
b1000 +
#666650000000
0!
0'
#666660000000
1!
b1001 %
1'
b1001 +
#666670000000
0!
0'
#666680000000
1!
b0 %
1'
b0 +
#666690000000
0!
0'
#666700000000
1!
1$
b1 %
1'
1*
b1 +
#666710000000
1"
1(
#666720000000
0!
0"
b100 &
0'
0(
b100 ,
#666730000000
1!
b10 %
1'
b10 +
#666740000000
0!
0'
#666750000000
1!
b11 %
1'
b11 +
#666760000000
0!
0'
#666770000000
1!
b100 %
1'
b100 +
#666780000000
0!
0'
#666790000000
1!
b101 %
1'
b101 +
#666800000000
0!
0'
#666810000000
1!
b110 %
1'
b110 +
#666820000000
0!
0'
#666830000000
1!
b111 %
1'
b111 +
#666840000000
0!
0'
#666850000000
1!
0$
b1000 %
1'
0*
b1000 +
#666860000000
0!
0'
#666870000000
1!
b1001 %
1'
b1001 +
#666880000000
0!
0'
#666890000000
1!
b0 %
1'
b0 +
#666900000000
0!
0'
#666910000000
1!
1$
b1 %
1'
1*
b1 +
#666920000000
0!
0'
#666930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#666940000000
0!
0'
#666950000000
1!
b11 %
1'
b11 +
#666960000000
0!
0'
#666970000000
1!
b100 %
1'
b100 +
#666980000000
0!
0'
#666990000000
1!
b101 %
1'
b101 +
#667000000000
0!
0'
#667010000000
1!
0$
b110 %
1'
0*
b110 +
#667020000000
0!
0'
#667030000000
1!
b111 %
1'
b111 +
#667040000000
0!
0'
#667050000000
1!
b1000 %
1'
b1000 +
#667060000000
0!
0'
#667070000000
1!
b1001 %
1'
b1001 +
#667080000000
0!
0'
#667090000000
1!
b0 %
1'
b0 +
#667100000000
0!
0'
#667110000000
1!
1$
b1 %
1'
1*
b1 +
#667120000000
0!
0'
#667130000000
1!
b10 %
1'
b10 +
#667140000000
1"
1(
#667150000000
0!
0"
b100 &
0'
0(
b100 ,
#667160000000
1!
b11 %
1'
b11 +
#667170000000
0!
0'
#667180000000
1!
b100 %
1'
b100 +
#667190000000
0!
0'
#667200000000
1!
b101 %
1'
b101 +
#667210000000
0!
0'
#667220000000
1!
b110 %
1'
b110 +
#667230000000
0!
0'
#667240000000
1!
b111 %
1'
b111 +
#667250000000
0!
0'
#667260000000
1!
0$
b1000 %
1'
0*
b1000 +
#667270000000
0!
0'
#667280000000
1!
b1001 %
1'
b1001 +
#667290000000
0!
0'
#667300000000
1!
b0 %
1'
b0 +
#667310000000
0!
0'
#667320000000
1!
1$
b1 %
1'
1*
b1 +
#667330000000
0!
0'
#667340000000
1!
b10 %
1'
b10 +
#667350000000
0!
0'
#667360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#667370000000
0!
0'
#667380000000
1!
b100 %
1'
b100 +
#667390000000
0!
0'
#667400000000
1!
b101 %
1'
b101 +
#667410000000
0!
0'
#667420000000
1!
0$
b110 %
1'
0*
b110 +
#667430000000
0!
0'
#667440000000
1!
b111 %
1'
b111 +
#667450000000
0!
0'
#667460000000
1!
b1000 %
1'
b1000 +
#667470000000
0!
0'
#667480000000
1!
b1001 %
1'
b1001 +
#667490000000
0!
0'
#667500000000
1!
b0 %
1'
b0 +
#667510000000
0!
0'
#667520000000
1!
1$
b1 %
1'
1*
b1 +
#667530000000
0!
0'
#667540000000
1!
b10 %
1'
b10 +
#667550000000
0!
0'
#667560000000
1!
b11 %
1'
b11 +
#667570000000
1"
1(
#667580000000
0!
0"
b100 &
0'
0(
b100 ,
#667590000000
1!
b100 %
1'
b100 +
#667600000000
0!
0'
#667610000000
1!
b101 %
1'
b101 +
#667620000000
0!
0'
#667630000000
1!
b110 %
1'
b110 +
#667640000000
0!
0'
#667650000000
1!
b111 %
1'
b111 +
#667660000000
0!
0'
#667670000000
1!
0$
b1000 %
1'
0*
b1000 +
#667680000000
0!
0'
#667690000000
1!
b1001 %
1'
b1001 +
#667700000000
0!
0'
#667710000000
1!
b0 %
1'
b0 +
#667720000000
0!
0'
#667730000000
1!
1$
b1 %
1'
1*
b1 +
#667740000000
0!
0'
#667750000000
1!
b10 %
1'
b10 +
#667760000000
0!
0'
#667770000000
1!
b11 %
1'
b11 +
#667780000000
0!
0'
#667790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#667800000000
0!
0'
#667810000000
1!
b101 %
1'
b101 +
#667820000000
0!
0'
#667830000000
1!
0$
b110 %
1'
0*
b110 +
#667840000000
0!
0'
#667850000000
1!
b111 %
1'
b111 +
#667860000000
0!
0'
#667870000000
1!
b1000 %
1'
b1000 +
#667880000000
0!
0'
#667890000000
1!
b1001 %
1'
b1001 +
#667900000000
0!
0'
#667910000000
1!
b0 %
1'
b0 +
#667920000000
0!
0'
#667930000000
1!
1$
b1 %
1'
1*
b1 +
#667940000000
0!
0'
#667950000000
1!
b10 %
1'
b10 +
#667960000000
0!
0'
#667970000000
1!
b11 %
1'
b11 +
#667980000000
0!
0'
#667990000000
1!
b100 %
1'
b100 +
#668000000000
1"
1(
#668010000000
0!
0"
b100 &
0'
0(
b100 ,
#668020000000
1!
b101 %
1'
b101 +
#668030000000
0!
0'
#668040000000
1!
b110 %
1'
b110 +
#668050000000
0!
0'
#668060000000
1!
b111 %
1'
b111 +
#668070000000
0!
0'
#668080000000
1!
0$
b1000 %
1'
0*
b1000 +
#668090000000
0!
0'
#668100000000
1!
b1001 %
1'
b1001 +
#668110000000
0!
0'
#668120000000
1!
b0 %
1'
b0 +
#668130000000
0!
0'
#668140000000
1!
1$
b1 %
1'
1*
b1 +
#668150000000
0!
0'
#668160000000
1!
b10 %
1'
b10 +
#668170000000
0!
0'
#668180000000
1!
b11 %
1'
b11 +
#668190000000
0!
0'
#668200000000
1!
b100 %
1'
b100 +
#668210000000
0!
0'
#668220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#668230000000
0!
0'
#668240000000
1!
0$
b110 %
1'
0*
b110 +
#668250000000
0!
0'
#668260000000
1!
b111 %
1'
b111 +
#668270000000
0!
0'
#668280000000
1!
b1000 %
1'
b1000 +
#668290000000
0!
0'
#668300000000
1!
b1001 %
1'
b1001 +
#668310000000
0!
0'
#668320000000
1!
b0 %
1'
b0 +
#668330000000
0!
0'
#668340000000
1!
1$
b1 %
1'
1*
b1 +
#668350000000
0!
0'
#668360000000
1!
b10 %
1'
b10 +
#668370000000
0!
0'
#668380000000
1!
b11 %
1'
b11 +
#668390000000
0!
0'
#668400000000
1!
b100 %
1'
b100 +
#668410000000
0!
0'
#668420000000
1!
b101 %
1'
b101 +
#668430000000
1"
1(
#668440000000
0!
0"
b100 &
0'
0(
b100 ,
#668450000000
1!
b110 %
1'
b110 +
#668460000000
0!
0'
#668470000000
1!
b111 %
1'
b111 +
#668480000000
0!
0'
#668490000000
1!
0$
b1000 %
1'
0*
b1000 +
#668500000000
0!
0'
#668510000000
1!
b1001 %
1'
b1001 +
#668520000000
0!
0'
#668530000000
1!
b0 %
1'
b0 +
#668540000000
0!
0'
#668550000000
1!
1$
b1 %
1'
1*
b1 +
#668560000000
0!
0'
#668570000000
1!
b10 %
1'
b10 +
#668580000000
0!
0'
#668590000000
1!
b11 %
1'
b11 +
#668600000000
0!
0'
#668610000000
1!
b100 %
1'
b100 +
#668620000000
0!
0'
#668630000000
1!
b101 %
1'
b101 +
#668640000000
0!
0'
#668650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#668660000000
0!
0'
#668670000000
1!
b111 %
1'
b111 +
#668680000000
0!
0'
#668690000000
1!
b1000 %
1'
b1000 +
#668700000000
0!
0'
#668710000000
1!
b1001 %
1'
b1001 +
#668720000000
0!
0'
#668730000000
1!
b0 %
1'
b0 +
#668740000000
0!
0'
#668750000000
1!
1$
b1 %
1'
1*
b1 +
#668760000000
0!
0'
#668770000000
1!
b10 %
1'
b10 +
#668780000000
0!
0'
#668790000000
1!
b11 %
1'
b11 +
#668800000000
0!
0'
#668810000000
1!
b100 %
1'
b100 +
#668820000000
0!
0'
#668830000000
1!
b101 %
1'
b101 +
#668840000000
0!
0'
#668850000000
1!
0$
b110 %
1'
0*
b110 +
#668860000000
1"
1(
#668870000000
0!
0"
b100 &
0'
0(
b100 ,
#668880000000
1!
1$
b111 %
1'
1*
b111 +
#668890000000
0!
0'
#668900000000
1!
0$
b1000 %
1'
0*
b1000 +
#668910000000
0!
0'
#668920000000
1!
b1001 %
1'
b1001 +
#668930000000
0!
0'
#668940000000
1!
b0 %
1'
b0 +
#668950000000
0!
0'
#668960000000
1!
1$
b1 %
1'
1*
b1 +
#668970000000
0!
0'
#668980000000
1!
b10 %
1'
b10 +
#668990000000
0!
0'
#669000000000
1!
b11 %
1'
b11 +
#669010000000
0!
0'
#669020000000
1!
b100 %
1'
b100 +
#669030000000
0!
0'
#669040000000
1!
b101 %
1'
b101 +
#669050000000
0!
0'
#669060000000
1!
b110 %
1'
b110 +
#669070000000
0!
0'
#669080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#669090000000
0!
0'
#669100000000
1!
b1000 %
1'
b1000 +
#669110000000
0!
0'
#669120000000
1!
b1001 %
1'
b1001 +
#669130000000
0!
0'
#669140000000
1!
b0 %
1'
b0 +
#669150000000
0!
0'
#669160000000
1!
1$
b1 %
1'
1*
b1 +
#669170000000
0!
0'
#669180000000
1!
b10 %
1'
b10 +
#669190000000
0!
0'
#669200000000
1!
b11 %
1'
b11 +
#669210000000
0!
0'
#669220000000
1!
b100 %
1'
b100 +
#669230000000
0!
0'
#669240000000
1!
b101 %
1'
b101 +
#669250000000
0!
0'
#669260000000
1!
0$
b110 %
1'
0*
b110 +
#669270000000
0!
0'
#669280000000
1!
b111 %
1'
b111 +
#669290000000
1"
1(
#669300000000
0!
0"
b100 &
0'
0(
b100 ,
#669310000000
1!
b1000 %
1'
b1000 +
#669320000000
0!
0'
#669330000000
1!
b1001 %
1'
b1001 +
#669340000000
0!
0'
#669350000000
1!
b0 %
1'
b0 +
#669360000000
0!
0'
#669370000000
1!
1$
b1 %
1'
1*
b1 +
#669380000000
0!
0'
#669390000000
1!
b10 %
1'
b10 +
#669400000000
0!
0'
#669410000000
1!
b11 %
1'
b11 +
#669420000000
0!
0'
#669430000000
1!
b100 %
1'
b100 +
#669440000000
0!
0'
#669450000000
1!
b101 %
1'
b101 +
#669460000000
0!
0'
#669470000000
1!
b110 %
1'
b110 +
#669480000000
0!
0'
#669490000000
1!
b111 %
1'
b111 +
#669500000000
0!
0'
#669510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#669520000000
0!
0'
#669530000000
1!
b1001 %
1'
b1001 +
#669540000000
0!
0'
#669550000000
1!
b0 %
1'
b0 +
#669560000000
0!
0'
#669570000000
1!
1$
b1 %
1'
1*
b1 +
#669580000000
0!
0'
#669590000000
1!
b10 %
1'
b10 +
#669600000000
0!
0'
#669610000000
1!
b11 %
1'
b11 +
#669620000000
0!
0'
#669630000000
1!
b100 %
1'
b100 +
#669640000000
0!
0'
#669650000000
1!
b101 %
1'
b101 +
#669660000000
0!
0'
#669670000000
1!
0$
b110 %
1'
0*
b110 +
#669680000000
0!
0'
#669690000000
1!
b111 %
1'
b111 +
#669700000000
0!
0'
#669710000000
1!
b1000 %
1'
b1000 +
#669720000000
1"
1(
#669730000000
0!
0"
b100 &
0'
0(
b100 ,
#669740000000
1!
b1001 %
1'
b1001 +
#669750000000
0!
0'
#669760000000
1!
b0 %
1'
b0 +
#669770000000
0!
0'
#669780000000
1!
1$
b1 %
1'
1*
b1 +
#669790000000
0!
0'
#669800000000
1!
b10 %
1'
b10 +
#669810000000
0!
0'
#669820000000
1!
b11 %
1'
b11 +
#669830000000
0!
0'
#669840000000
1!
b100 %
1'
b100 +
#669850000000
0!
0'
#669860000000
1!
b101 %
1'
b101 +
#669870000000
0!
0'
#669880000000
1!
b110 %
1'
b110 +
#669890000000
0!
0'
#669900000000
1!
b111 %
1'
b111 +
#669910000000
0!
0'
#669920000000
1!
0$
b1000 %
1'
0*
b1000 +
#669930000000
0!
0'
#669940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#669950000000
0!
0'
#669960000000
1!
b0 %
1'
b0 +
#669970000000
0!
0'
#669980000000
1!
1$
b1 %
1'
1*
b1 +
#669990000000
0!
0'
#670000000000
1!
b10 %
1'
b10 +
#670010000000
0!
0'
#670020000000
1!
b11 %
1'
b11 +
#670030000000
0!
0'
#670040000000
1!
b100 %
1'
b100 +
#670050000000
0!
0'
#670060000000
1!
b101 %
1'
b101 +
#670070000000
0!
0'
#670080000000
1!
0$
b110 %
1'
0*
b110 +
#670090000000
0!
0'
#670100000000
1!
b111 %
1'
b111 +
#670110000000
0!
0'
#670120000000
1!
b1000 %
1'
b1000 +
#670130000000
0!
0'
#670140000000
1!
b1001 %
1'
b1001 +
#670150000000
1"
1(
#670160000000
0!
0"
b100 &
0'
0(
b100 ,
#670170000000
1!
b0 %
1'
b0 +
#670180000000
0!
0'
#670190000000
1!
1$
b1 %
1'
1*
b1 +
#670200000000
0!
0'
#670210000000
1!
b10 %
1'
b10 +
#670220000000
0!
0'
#670230000000
1!
b11 %
1'
b11 +
#670240000000
0!
0'
#670250000000
1!
b100 %
1'
b100 +
#670260000000
0!
0'
#670270000000
1!
b101 %
1'
b101 +
#670280000000
0!
0'
#670290000000
1!
b110 %
1'
b110 +
#670300000000
0!
0'
#670310000000
1!
b111 %
1'
b111 +
#670320000000
0!
0'
#670330000000
1!
0$
b1000 %
1'
0*
b1000 +
#670340000000
0!
0'
#670350000000
1!
b1001 %
1'
b1001 +
#670360000000
0!
0'
#670370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#670380000000
0!
0'
#670390000000
1!
1$
b1 %
1'
1*
b1 +
#670400000000
0!
0'
#670410000000
1!
b10 %
1'
b10 +
#670420000000
0!
0'
#670430000000
1!
b11 %
1'
b11 +
#670440000000
0!
0'
#670450000000
1!
b100 %
1'
b100 +
#670460000000
0!
0'
#670470000000
1!
b101 %
1'
b101 +
#670480000000
0!
0'
#670490000000
1!
0$
b110 %
1'
0*
b110 +
#670500000000
0!
0'
#670510000000
1!
b111 %
1'
b111 +
#670520000000
0!
0'
#670530000000
1!
b1000 %
1'
b1000 +
#670540000000
0!
0'
#670550000000
1!
b1001 %
1'
b1001 +
#670560000000
0!
0'
#670570000000
1!
b0 %
1'
b0 +
#670580000000
1"
1(
#670590000000
0!
0"
b100 &
0'
0(
b100 ,
#670600000000
1!
1$
b1 %
1'
1*
b1 +
#670610000000
0!
0'
#670620000000
1!
b10 %
1'
b10 +
#670630000000
0!
0'
#670640000000
1!
b11 %
1'
b11 +
#670650000000
0!
0'
#670660000000
1!
b100 %
1'
b100 +
#670670000000
0!
0'
#670680000000
1!
b101 %
1'
b101 +
#670690000000
0!
0'
#670700000000
1!
b110 %
1'
b110 +
#670710000000
0!
0'
#670720000000
1!
b111 %
1'
b111 +
#670730000000
0!
0'
#670740000000
1!
0$
b1000 %
1'
0*
b1000 +
#670750000000
0!
0'
#670760000000
1!
b1001 %
1'
b1001 +
#670770000000
0!
0'
#670780000000
1!
b0 %
1'
b0 +
#670790000000
0!
0'
#670800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#670810000000
0!
0'
#670820000000
1!
b10 %
1'
b10 +
#670830000000
0!
0'
#670840000000
1!
b11 %
1'
b11 +
#670850000000
0!
0'
#670860000000
1!
b100 %
1'
b100 +
#670870000000
0!
0'
#670880000000
1!
b101 %
1'
b101 +
#670890000000
0!
0'
#670900000000
1!
0$
b110 %
1'
0*
b110 +
#670910000000
0!
0'
#670920000000
1!
b111 %
1'
b111 +
#670930000000
0!
0'
#670940000000
1!
b1000 %
1'
b1000 +
#670950000000
0!
0'
#670960000000
1!
b1001 %
1'
b1001 +
#670970000000
0!
0'
#670980000000
1!
b0 %
1'
b0 +
#670990000000
0!
0'
#671000000000
1!
1$
b1 %
1'
1*
b1 +
#671010000000
1"
1(
#671020000000
0!
0"
b100 &
0'
0(
b100 ,
#671030000000
1!
b10 %
1'
b10 +
#671040000000
0!
0'
#671050000000
1!
b11 %
1'
b11 +
#671060000000
0!
0'
#671070000000
1!
b100 %
1'
b100 +
#671080000000
0!
0'
#671090000000
1!
b101 %
1'
b101 +
#671100000000
0!
0'
#671110000000
1!
b110 %
1'
b110 +
#671120000000
0!
0'
#671130000000
1!
b111 %
1'
b111 +
#671140000000
0!
0'
#671150000000
1!
0$
b1000 %
1'
0*
b1000 +
#671160000000
0!
0'
#671170000000
1!
b1001 %
1'
b1001 +
#671180000000
0!
0'
#671190000000
1!
b0 %
1'
b0 +
#671200000000
0!
0'
#671210000000
1!
1$
b1 %
1'
1*
b1 +
#671220000000
0!
0'
#671230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#671240000000
0!
0'
#671250000000
1!
b11 %
1'
b11 +
#671260000000
0!
0'
#671270000000
1!
b100 %
1'
b100 +
#671280000000
0!
0'
#671290000000
1!
b101 %
1'
b101 +
#671300000000
0!
0'
#671310000000
1!
0$
b110 %
1'
0*
b110 +
#671320000000
0!
0'
#671330000000
1!
b111 %
1'
b111 +
#671340000000
0!
0'
#671350000000
1!
b1000 %
1'
b1000 +
#671360000000
0!
0'
#671370000000
1!
b1001 %
1'
b1001 +
#671380000000
0!
0'
#671390000000
1!
b0 %
1'
b0 +
#671400000000
0!
0'
#671410000000
1!
1$
b1 %
1'
1*
b1 +
#671420000000
0!
0'
#671430000000
1!
b10 %
1'
b10 +
#671440000000
1"
1(
#671450000000
0!
0"
b100 &
0'
0(
b100 ,
#671460000000
1!
b11 %
1'
b11 +
#671470000000
0!
0'
#671480000000
1!
b100 %
1'
b100 +
#671490000000
0!
0'
#671500000000
1!
b101 %
1'
b101 +
#671510000000
0!
0'
#671520000000
1!
b110 %
1'
b110 +
#671530000000
0!
0'
#671540000000
1!
b111 %
1'
b111 +
#671550000000
0!
0'
#671560000000
1!
0$
b1000 %
1'
0*
b1000 +
#671570000000
0!
0'
#671580000000
1!
b1001 %
1'
b1001 +
#671590000000
0!
0'
#671600000000
1!
b0 %
1'
b0 +
#671610000000
0!
0'
#671620000000
1!
1$
b1 %
1'
1*
b1 +
#671630000000
0!
0'
#671640000000
1!
b10 %
1'
b10 +
#671650000000
0!
0'
#671660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#671670000000
0!
0'
#671680000000
1!
b100 %
1'
b100 +
#671690000000
0!
0'
#671700000000
1!
b101 %
1'
b101 +
#671710000000
0!
0'
#671720000000
1!
0$
b110 %
1'
0*
b110 +
#671730000000
0!
0'
#671740000000
1!
b111 %
1'
b111 +
#671750000000
0!
0'
#671760000000
1!
b1000 %
1'
b1000 +
#671770000000
0!
0'
#671780000000
1!
b1001 %
1'
b1001 +
#671790000000
0!
0'
#671800000000
1!
b0 %
1'
b0 +
#671810000000
0!
0'
#671820000000
1!
1$
b1 %
1'
1*
b1 +
#671830000000
0!
0'
#671840000000
1!
b10 %
1'
b10 +
#671850000000
0!
0'
#671860000000
1!
b11 %
1'
b11 +
#671870000000
1"
1(
#671880000000
0!
0"
b100 &
0'
0(
b100 ,
#671890000000
1!
b100 %
1'
b100 +
#671900000000
0!
0'
#671910000000
1!
b101 %
1'
b101 +
#671920000000
0!
0'
#671930000000
1!
b110 %
1'
b110 +
#671940000000
0!
0'
#671950000000
1!
b111 %
1'
b111 +
#671960000000
0!
0'
#671970000000
1!
0$
b1000 %
1'
0*
b1000 +
#671980000000
0!
0'
#671990000000
1!
b1001 %
1'
b1001 +
#672000000000
0!
0'
#672010000000
1!
b0 %
1'
b0 +
#672020000000
0!
0'
#672030000000
1!
1$
b1 %
1'
1*
b1 +
#672040000000
0!
0'
#672050000000
1!
b10 %
1'
b10 +
#672060000000
0!
0'
#672070000000
1!
b11 %
1'
b11 +
#672080000000
0!
0'
#672090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#672100000000
0!
0'
#672110000000
1!
b101 %
1'
b101 +
#672120000000
0!
0'
#672130000000
1!
0$
b110 %
1'
0*
b110 +
#672140000000
0!
0'
#672150000000
1!
b111 %
1'
b111 +
#672160000000
0!
0'
#672170000000
1!
b1000 %
1'
b1000 +
#672180000000
0!
0'
#672190000000
1!
b1001 %
1'
b1001 +
#672200000000
0!
0'
#672210000000
1!
b0 %
1'
b0 +
#672220000000
0!
0'
#672230000000
1!
1$
b1 %
1'
1*
b1 +
#672240000000
0!
0'
#672250000000
1!
b10 %
1'
b10 +
#672260000000
0!
0'
#672270000000
1!
b11 %
1'
b11 +
#672280000000
0!
0'
#672290000000
1!
b100 %
1'
b100 +
#672300000000
1"
1(
#672310000000
0!
0"
b100 &
0'
0(
b100 ,
#672320000000
1!
b101 %
1'
b101 +
#672330000000
0!
0'
#672340000000
1!
b110 %
1'
b110 +
#672350000000
0!
0'
#672360000000
1!
b111 %
1'
b111 +
#672370000000
0!
0'
#672380000000
1!
0$
b1000 %
1'
0*
b1000 +
#672390000000
0!
0'
#672400000000
1!
b1001 %
1'
b1001 +
#672410000000
0!
0'
#672420000000
1!
b0 %
1'
b0 +
#672430000000
0!
0'
#672440000000
1!
1$
b1 %
1'
1*
b1 +
#672450000000
0!
0'
#672460000000
1!
b10 %
1'
b10 +
#672470000000
0!
0'
#672480000000
1!
b11 %
1'
b11 +
#672490000000
0!
0'
#672500000000
1!
b100 %
1'
b100 +
#672510000000
0!
0'
#672520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#672530000000
0!
0'
#672540000000
1!
0$
b110 %
1'
0*
b110 +
#672550000000
0!
0'
#672560000000
1!
b111 %
1'
b111 +
#672570000000
0!
0'
#672580000000
1!
b1000 %
1'
b1000 +
#672590000000
0!
0'
#672600000000
1!
b1001 %
1'
b1001 +
#672610000000
0!
0'
#672620000000
1!
b0 %
1'
b0 +
#672630000000
0!
0'
#672640000000
1!
1$
b1 %
1'
1*
b1 +
#672650000000
0!
0'
#672660000000
1!
b10 %
1'
b10 +
#672670000000
0!
0'
#672680000000
1!
b11 %
1'
b11 +
#672690000000
0!
0'
#672700000000
1!
b100 %
1'
b100 +
#672710000000
0!
0'
#672720000000
1!
b101 %
1'
b101 +
#672730000000
1"
1(
#672740000000
0!
0"
b100 &
0'
0(
b100 ,
#672750000000
1!
b110 %
1'
b110 +
#672760000000
0!
0'
#672770000000
1!
b111 %
1'
b111 +
#672780000000
0!
0'
#672790000000
1!
0$
b1000 %
1'
0*
b1000 +
#672800000000
0!
0'
#672810000000
1!
b1001 %
1'
b1001 +
#672820000000
0!
0'
#672830000000
1!
b0 %
1'
b0 +
#672840000000
0!
0'
#672850000000
1!
1$
b1 %
1'
1*
b1 +
#672860000000
0!
0'
#672870000000
1!
b10 %
1'
b10 +
#672880000000
0!
0'
#672890000000
1!
b11 %
1'
b11 +
#672900000000
0!
0'
#672910000000
1!
b100 %
1'
b100 +
#672920000000
0!
0'
#672930000000
1!
b101 %
1'
b101 +
#672940000000
0!
0'
#672950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#672960000000
0!
0'
#672970000000
1!
b111 %
1'
b111 +
#672980000000
0!
0'
#672990000000
1!
b1000 %
1'
b1000 +
#673000000000
0!
0'
#673010000000
1!
b1001 %
1'
b1001 +
#673020000000
0!
0'
#673030000000
1!
b0 %
1'
b0 +
#673040000000
0!
0'
#673050000000
1!
1$
b1 %
1'
1*
b1 +
#673060000000
0!
0'
#673070000000
1!
b10 %
1'
b10 +
#673080000000
0!
0'
#673090000000
1!
b11 %
1'
b11 +
#673100000000
0!
0'
#673110000000
1!
b100 %
1'
b100 +
#673120000000
0!
0'
#673130000000
1!
b101 %
1'
b101 +
#673140000000
0!
0'
#673150000000
1!
0$
b110 %
1'
0*
b110 +
#673160000000
1"
1(
#673170000000
0!
0"
b100 &
0'
0(
b100 ,
#673180000000
1!
1$
b111 %
1'
1*
b111 +
#673190000000
0!
0'
#673200000000
1!
0$
b1000 %
1'
0*
b1000 +
#673210000000
0!
0'
#673220000000
1!
b1001 %
1'
b1001 +
#673230000000
0!
0'
#673240000000
1!
b0 %
1'
b0 +
#673250000000
0!
0'
#673260000000
1!
1$
b1 %
1'
1*
b1 +
#673270000000
0!
0'
#673280000000
1!
b10 %
1'
b10 +
#673290000000
0!
0'
#673300000000
1!
b11 %
1'
b11 +
#673310000000
0!
0'
#673320000000
1!
b100 %
1'
b100 +
#673330000000
0!
0'
#673340000000
1!
b101 %
1'
b101 +
#673350000000
0!
0'
#673360000000
1!
b110 %
1'
b110 +
#673370000000
0!
0'
#673380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#673390000000
0!
0'
#673400000000
1!
b1000 %
1'
b1000 +
#673410000000
0!
0'
#673420000000
1!
b1001 %
1'
b1001 +
#673430000000
0!
0'
#673440000000
1!
b0 %
1'
b0 +
#673450000000
0!
0'
#673460000000
1!
1$
b1 %
1'
1*
b1 +
#673470000000
0!
0'
#673480000000
1!
b10 %
1'
b10 +
#673490000000
0!
0'
#673500000000
1!
b11 %
1'
b11 +
#673510000000
0!
0'
#673520000000
1!
b100 %
1'
b100 +
#673530000000
0!
0'
#673540000000
1!
b101 %
1'
b101 +
#673550000000
0!
0'
#673560000000
1!
0$
b110 %
1'
0*
b110 +
#673570000000
0!
0'
#673580000000
1!
b111 %
1'
b111 +
#673590000000
1"
1(
#673600000000
0!
0"
b100 &
0'
0(
b100 ,
#673610000000
1!
b1000 %
1'
b1000 +
#673620000000
0!
0'
#673630000000
1!
b1001 %
1'
b1001 +
#673640000000
0!
0'
#673650000000
1!
b0 %
1'
b0 +
#673660000000
0!
0'
#673670000000
1!
1$
b1 %
1'
1*
b1 +
#673680000000
0!
0'
#673690000000
1!
b10 %
1'
b10 +
#673700000000
0!
0'
#673710000000
1!
b11 %
1'
b11 +
#673720000000
0!
0'
#673730000000
1!
b100 %
1'
b100 +
#673740000000
0!
0'
#673750000000
1!
b101 %
1'
b101 +
#673760000000
0!
0'
#673770000000
1!
b110 %
1'
b110 +
#673780000000
0!
0'
#673790000000
1!
b111 %
1'
b111 +
#673800000000
0!
0'
#673810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#673820000000
0!
0'
#673830000000
1!
b1001 %
1'
b1001 +
#673840000000
0!
0'
#673850000000
1!
b0 %
1'
b0 +
#673860000000
0!
0'
#673870000000
1!
1$
b1 %
1'
1*
b1 +
#673880000000
0!
0'
#673890000000
1!
b10 %
1'
b10 +
#673900000000
0!
0'
#673910000000
1!
b11 %
1'
b11 +
#673920000000
0!
0'
#673930000000
1!
b100 %
1'
b100 +
#673940000000
0!
0'
#673950000000
1!
b101 %
1'
b101 +
#673960000000
0!
0'
#673970000000
1!
0$
b110 %
1'
0*
b110 +
#673980000000
0!
0'
#673990000000
1!
b111 %
1'
b111 +
#674000000000
0!
0'
#674010000000
1!
b1000 %
1'
b1000 +
#674020000000
1"
1(
#674030000000
0!
0"
b100 &
0'
0(
b100 ,
#674040000000
1!
b1001 %
1'
b1001 +
#674050000000
0!
0'
#674060000000
1!
b0 %
1'
b0 +
#674070000000
0!
0'
#674080000000
1!
1$
b1 %
1'
1*
b1 +
#674090000000
0!
0'
#674100000000
1!
b10 %
1'
b10 +
#674110000000
0!
0'
#674120000000
1!
b11 %
1'
b11 +
#674130000000
0!
0'
#674140000000
1!
b100 %
1'
b100 +
#674150000000
0!
0'
#674160000000
1!
b101 %
1'
b101 +
#674170000000
0!
0'
#674180000000
1!
b110 %
1'
b110 +
#674190000000
0!
0'
#674200000000
1!
b111 %
1'
b111 +
#674210000000
0!
0'
#674220000000
1!
0$
b1000 %
1'
0*
b1000 +
#674230000000
0!
0'
#674240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#674250000000
0!
0'
#674260000000
1!
b0 %
1'
b0 +
#674270000000
0!
0'
#674280000000
1!
1$
b1 %
1'
1*
b1 +
#674290000000
0!
0'
#674300000000
1!
b10 %
1'
b10 +
#674310000000
0!
0'
#674320000000
1!
b11 %
1'
b11 +
#674330000000
0!
0'
#674340000000
1!
b100 %
1'
b100 +
#674350000000
0!
0'
#674360000000
1!
b101 %
1'
b101 +
#674370000000
0!
0'
#674380000000
1!
0$
b110 %
1'
0*
b110 +
#674390000000
0!
0'
#674400000000
1!
b111 %
1'
b111 +
#674410000000
0!
0'
#674420000000
1!
b1000 %
1'
b1000 +
#674430000000
0!
0'
#674440000000
1!
b1001 %
1'
b1001 +
#674450000000
1"
1(
#674460000000
0!
0"
b100 &
0'
0(
b100 ,
#674470000000
1!
b0 %
1'
b0 +
#674480000000
0!
0'
#674490000000
1!
1$
b1 %
1'
1*
b1 +
#674500000000
0!
0'
#674510000000
1!
b10 %
1'
b10 +
#674520000000
0!
0'
#674530000000
1!
b11 %
1'
b11 +
#674540000000
0!
0'
#674550000000
1!
b100 %
1'
b100 +
#674560000000
0!
0'
#674570000000
1!
b101 %
1'
b101 +
#674580000000
0!
0'
#674590000000
1!
b110 %
1'
b110 +
#674600000000
0!
0'
#674610000000
1!
b111 %
1'
b111 +
#674620000000
0!
0'
#674630000000
1!
0$
b1000 %
1'
0*
b1000 +
#674640000000
0!
0'
#674650000000
1!
b1001 %
1'
b1001 +
#674660000000
0!
0'
#674670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#674680000000
0!
0'
#674690000000
1!
1$
b1 %
1'
1*
b1 +
#674700000000
0!
0'
#674710000000
1!
b10 %
1'
b10 +
#674720000000
0!
0'
#674730000000
1!
b11 %
1'
b11 +
#674740000000
0!
0'
#674750000000
1!
b100 %
1'
b100 +
#674760000000
0!
0'
#674770000000
1!
b101 %
1'
b101 +
#674780000000
0!
0'
#674790000000
1!
0$
b110 %
1'
0*
b110 +
#674800000000
0!
0'
#674810000000
1!
b111 %
1'
b111 +
#674820000000
0!
0'
#674830000000
1!
b1000 %
1'
b1000 +
#674840000000
0!
0'
#674850000000
1!
b1001 %
1'
b1001 +
#674860000000
0!
0'
#674870000000
1!
b0 %
1'
b0 +
#674880000000
1"
1(
#674890000000
0!
0"
b100 &
0'
0(
b100 ,
#674900000000
1!
1$
b1 %
1'
1*
b1 +
#674910000000
0!
0'
#674920000000
1!
b10 %
1'
b10 +
#674930000000
0!
0'
#674940000000
1!
b11 %
1'
b11 +
#674950000000
0!
0'
#674960000000
1!
b100 %
1'
b100 +
#674970000000
0!
0'
#674980000000
1!
b101 %
1'
b101 +
#674990000000
0!
0'
#675000000000
1!
b110 %
1'
b110 +
#675010000000
0!
0'
#675020000000
1!
b111 %
1'
b111 +
#675030000000
0!
0'
#675040000000
1!
0$
b1000 %
1'
0*
b1000 +
#675050000000
0!
0'
#675060000000
1!
b1001 %
1'
b1001 +
#675070000000
0!
0'
#675080000000
1!
b0 %
1'
b0 +
#675090000000
0!
0'
#675100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#675110000000
0!
0'
#675120000000
1!
b10 %
1'
b10 +
#675130000000
0!
0'
#675140000000
1!
b11 %
1'
b11 +
#675150000000
0!
0'
#675160000000
1!
b100 %
1'
b100 +
#675170000000
0!
0'
#675180000000
1!
b101 %
1'
b101 +
#675190000000
0!
0'
#675200000000
1!
0$
b110 %
1'
0*
b110 +
#675210000000
0!
0'
#675220000000
1!
b111 %
1'
b111 +
#675230000000
0!
0'
#675240000000
1!
b1000 %
1'
b1000 +
#675250000000
0!
0'
#675260000000
1!
b1001 %
1'
b1001 +
#675270000000
0!
0'
#675280000000
1!
b0 %
1'
b0 +
#675290000000
0!
0'
#675300000000
1!
1$
b1 %
1'
1*
b1 +
#675310000000
1"
1(
#675320000000
0!
0"
b100 &
0'
0(
b100 ,
#675330000000
1!
b10 %
1'
b10 +
#675340000000
0!
0'
#675350000000
1!
b11 %
1'
b11 +
#675360000000
0!
0'
#675370000000
1!
b100 %
1'
b100 +
#675380000000
0!
0'
#675390000000
1!
b101 %
1'
b101 +
#675400000000
0!
0'
#675410000000
1!
b110 %
1'
b110 +
#675420000000
0!
0'
#675430000000
1!
b111 %
1'
b111 +
#675440000000
0!
0'
#675450000000
1!
0$
b1000 %
1'
0*
b1000 +
#675460000000
0!
0'
#675470000000
1!
b1001 %
1'
b1001 +
#675480000000
0!
0'
#675490000000
1!
b0 %
1'
b0 +
#675500000000
0!
0'
#675510000000
1!
1$
b1 %
1'
1*
b1 +
#675520000000
0!
0'
#675530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#675540000000
0!
0'
#675550000000
1!
b11 %
1'
b11 +
#675560000000
0!
0'
#675570000000
1!
b100 %
1'
b100 +
#675580000000
0!
0'
#675590000000
1!
b101 %
1'
b101 +
#675600000000
0!
0'
#675610000000
1!
0$
b110 %
1'
0*
b110 +
#675620000000
0!
0'
#675630000000
1!
b111 %
1'
b111 +
#675640000000
0!
0'
#675650000000
1!
b1000 %
1'
b1000 +
#675660000000
0!
0'
#675670000000
1!
b1001 %
1'
b1001 +
#675680000000
0!
0'
#675690000000
1!
b0 %
1'
b0 +
#675700000000
0!
0'
#675710000000
1!
1$
b1 %
1'
1*
b1 +
#675720000000
0!
0'
#675730000000
1!
b10 %
1'
b10 +
#675740000000
1"
1(
#675750000000
0!
0"
b100 &
0'
0(
b100 ,
#675760000000
1!
b11 %
1'
b11 +
#675770000000
0!
0'
#675780000000
1!
b100 %
1'
b100 +
#675790000000
0!
0'
#675800000000
1!
b101 %
1'
b101 +
#675810000000
0!
0'
#675820000000
1!
b110 %
1'
b110 +
#675830000000
0!
0'
#675840000000
1!
b111 %
1'
b111 +
#675850000000
0!
0'
#675860000000
1!
0$
b1000 %
1'
0*
b1000 +
#675870000000
0!
0'
#675880000000
1!
b1001 %
1'
b1001 +
#675890000000
0!
0'
#675900000000
1!
b0 %
1'
b0 +
#675910000000
0!
0'
#675920000000
1!
1$
b1 %
1'
1*
b1 +
#675930000000
0!
0'
#675940000000
1!
b10 %
1'
b10 +
#675950000000
0!
0'
#675960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#675970000000
0!
0'
#675980000000
1!
b100 %
1'
b100 +
#675990000000
0!
0'
#676000000000
1!
b101 %
1'
b101 +
#676010000000
0!
0'
#676020000000
1!
0$
b110 %
1'
0*
b110 +
#676030000000
0!
0'
#676040000000
1!
b111 %
1'
b111 +
#676050000000
0!
0'
#676060000000
1!
b1000 %
1'
b1000 +
#676070000000
0!
0'
#676080000000
1!
b1001 %
1'
b1001 +
#676090000000
0!
0'
#676100000000
1!
b0 %
1'
b0 +
#676110000000
0!
0'
#676120000000
1!
1$
b1 %
1'
1*
b1 +
#676130000000
0!
0'
#676140000000
1!
b10 %
1'
b10 +
#676150000000
0!
0'
#676160000000
1!
b11 %
1'
b11 +
#676170000000
1"
1(
#676180000000
0!
0"
b100 &
0'
0(
b100 ,
#676190000000
1!
b100 %
1'
b100 +
#676200000000
0!
0'
#676210000000
1!
b101 %
1'
b101 +
#676220000000
0!
0'
#676230000000
1!
b110 %
1'
b110 +
#676240000000
0!
0'
#676250000000
1!
b111 %
1'
b111 +
#676260000000
0!
0'
#676270000000
1!
0$
b1000 %
1'
0*
b1000 +
#676280000000
0!
0'
#676290000000
1!
b1001 %
1'
b1001 +
#676300000000
0!
0'
#676310000000
1!
b0 %
1'
b0 +
#676320000000
0!
0'
#676330000000
1!
1$
b1 %
1'
1*
b1 +
#676340000000
0!
0'
#676350000000
1!
b10 %
1'
b10 +
#676360000000
0!
0'
#676370000000
1!
b11 %
1'
b11 +
#676380000000
0!
0'
#676390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#676400000000
0!
0'
#676410000000
1!
b101 %
1'
b101 +
#676420000000
0!
0'
#676430000000
1!
0$
b110 %
1'
0*
b110 +
#676440000000
0!
0'
#676450000000
1!
b111 %
1'
b111 +
#676460000000
0!
0'
#676470000000
1!
b1000 %
1'
b1000 +
#676480000000
0!
0'
#676490000000
1!
b1001 %
1'
b1001 +
#676500000000
0!
0'
#676510000000
1!
b0 %
1'
b0 +
#676520000000
0!
0'
#676530000000
1!
1$
b1 %
1'
1*
b1 +
#676540000000
0!
0'
#676550000000
1!
b10 %
1'
b10 +
#676560000000
0!
0'
#676570000000
1!
b11 %
1'
b11 +
#676580000000
0!
0'
#676590000000
1!
b100 %
1'
b100 +
#676600000000
1"
1(
#676610000000
0!
0"
b100 &
0'
0(
b100 ,
#676620000000
1!
b101 %
1'
b101 +
#676630000000
0!
0'
#676640000000
1!
b110 %
1'
b110 +
#676650000000
0!
0'
#676660000000
1!
b111 %
1'
b111 +
#676670000000
0!
0'
#676680000000
1!
0$
b1000 %
1'
0*
b1000 +
#676690000000
0!
0'
#676700000000
1!
b1001 %
1'
b1001 +
#676710000000
0!
0'
#676720000000
1!
b0 %
1'
b0 +
#676730000000
0!
0'
#676740000000
1!
1$
b1 %
1'
1*
b1 +
#676750000000
0!
0'
#676760000000
1!
b10 %
1'
b10 +
#676770000000
0!
0'
#676780000000
1!
b11 %
1'
b11 +
#676790000000
0!
0'
#676800000000
1!
b100 %
1'
b100 +
#676810000000
0!
0'
#676820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#676830000000
0!
0'
#676840000000
1!
0$
b110 %
1'
0*
b110 +
#676850000000
0!
0'
#676860000000
1!
b111 %
1'
b111 +
#676870000000
0!
0'
#676880000000
1!
b1000 %
1'
b1000 +
#676890000000
0!
0'
#676900000000
1!
b1001 %
1'
b1001 +
#676910000000
0!
0'
#676920000000
1!
b0 %
1'
b0 +
#676930000000
0!
0'
#676940000000
1!
1$
b1 %
1'
1*
b1 +
#676950000000
0!
0'
#676960000000
1!
b10 %
1'
b10 +
#676970000000
0!
0'
#676980000000
1!
b11 %
1'
b11 +
#676990000000
0!
0'
#677000000000
1!
b100 %
1'
b100 +
#677010000000
0!
0'
#677020000000
1!
b101 %
1'
b101 +
#677030000000
1"
1(
#677040000000
0!
0"
b100 &
0'
0(
b100 ,
#677050000000
1!
b110 %
1'
b110 +
#677060000000
0!
0'
#677070000000
1!
b111 %
1'
b111 +
#677080000000
0!
0'
#677090000000
1!
0$
b1000 %
1'
0*
b1000 +
#677100000000
0!
0'
#677110000000
1!
b1001 %
1'
b1001 +
#677120000000
0!
0'
#677130000000
1!
b0 %
1'
b0 +
#677140000000
0!
0'
#677150000000
1!
1$
b1 %
1'
1*
b1 +
#677160000000
0!
0'
#677170000000
1!
b10 %
1'
b10 +
#677180000000
0!
0'
#677190000000
1!
b11 %
1'
b11 +
#677200000000
0!
0'
#677210000000
1!
b100 %
1'
b100 +
#677220000000
0!
0'
#677230000000
1!
b101 %
1'
b101 +
#677240000000
0!
0'
#677250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#677260000000
0!
0'
#677270000000
1!
b111 %
1'
b111 +
#677280000000
0!
0'
#677290000000
1!
b1000 %
1'
b1000 +
#677300000000
0!
0'
#677310000000
1!
b1001 %
1'
b1001 +
#677320000000
0!
0'
#677330000000
1!
b0 %
1'
b0 +
#677340000000
0!
0'
#677350000000
1!
1$
b1 %
1'
1*
b1 +
#677360000000
0!
0'
#677370000000
1!
b10 %
1'
b10 +
#677380000000
0!
0'
#677390000000
1!
b11 %
1'
b11 +
#677400000000
0!
0'
#677410000000
1!
b100 %
1'
b100 +
#677420000000
0!
0'
#677430000000
1!
b101 %
1'
b101 +
#677440000000
0!
0'
#677450000000
1!
0$
b110 %
1'
0*
b110 +
#677460000000
1"
1(
#677470000000
0!
0"
b100 &
0'
0(
b100 ,
#677480000000
1!
1$
b111 %
1'
1*
b111 +
#677490000000
0!
0'
#677500000000
1!
0$
b1000 %
1'
0*
b1000 +
#677510000000
0!
0'
#677520000000
1!
b1001 %
1'
b1001 +
#677530000000
0!
0'
#677540000000
1!
b0 %
1'
b0 +
#677550000000
0!
0'
#677560000000
1!
1$
b1 %
1'
1*
b1 +
#677570000000
0!
0'
#677580000000
1!
b10 %
1'
b10 +
#677590000000
0!
0'
#677600000000
1!
b11 %
1'
b11 +
#677610000000
0!
0'
#677620000000
1!
b100 %
1'
b100 +
#677630000000
0!
0'
#677640000000
1!
b101 %
1'
b101 +
#677650000000
0!
0'
#677660000000
1!
b110 %
1'
b110 +
#677670000000
0!
0'
#677680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#677690000000
0!
0'
#677700000000
1!
b1000 %
1'
b1000 +
#677710000000
0!
0'
#677720000000
1!
b1001 %
1'
b1001 +
#677730000000
0!
0'
#677740000000
1!
b0 %
1'
b0 +
#677750000000
0!
0'
#677760000000
1!
1$
b1 %
1'
1*
b1 +
#677770000000
0!
0'
#677780000000
1!
b10 %
1'
b10 +
#677790000000
0!
0'
#677800000000
1!
b11 %
1'
b11 +
#677810000000
0!
0'
#677820000000
1!
b100 %
1'
b100 +
#677830000000
0!
0'
#677840000000
1!
b101 %
1'
b101 +
#677850000000
0!
0'
#677860000000
1!
0$
b110 %
1'
0*
b110 +
#677870000000
0!
0'
#677880000000
1!
b111 %
1'
b111 +
#677890000000
1"
1(
#677900000000
0!
0"
b100 &
0'
0(
b100 ,
#677910000000
1!
b1000 %
1'
b1000 +
#677920000000
0!
0'
#677930000000
1!
b1001 %
1'
b1001 +
#677940000000
0!
0'
#677950000000
1!
b0 %
1'
b0 +
#677960000000
0!
0'
#677970000000
1!
1$
b1 %
1'
1*
b1 +
#677980000000
0!
0'
#677990000000
1!
b10 %
1'
b10 +
#678000000000
0!
0'
#678010000000
1!
b11 %
1'
b11 +
#678020000000
0!
0'
#678030000000
1!
b100 %
1'
b100 +
#678040000000
0!
0'
#678050000000
1!
b101 %
1'
b101 +
#678060000000
0!
0'
#678070000000
1!
b110 %
1'
b110 +
#678080000000
0!
0'
#678090000000
1!
b111 %
1'
b111 +
#678100000000
0!
0'
#678110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#678120000000
0!
0'
#678130000000
1!
b1001 %
1'
b1001 +
#678140000000
0!
0'
#678150000000
1!
b0 %
1'
b0 +
#678160000000
0!
0'
#678170000000
1!
1$
b1 %
1'
1*
b1 +
#678180000000
0!
0'
#678190000000
1!
b10 %
1'
b10 +
#678200000000
0!
0'
#678210000000
1!
b11 %
1'
b11 +
#678220000000
0!
0'
#678230000000
1!
b100 %
1'
b100 +
#678240000000
0!
0'
#678250000000
1!
b101 %
1'
b101 +
#678260000000
0!
0'
#678270000000
1!
0$
b110 %
1'
0*
b110 +
#678280000000
0!
0'
#678290000000
1!
b111 %
1'
b111 +
#678300000000
0!
0'
#678310000000
1!
b1000 %
1'
b1000 +
#678320000000
1"
1(
#678330000000
0!
0"
b100 &
0'
0(
b100 ,
#678340000000
1!
b1001 %
1'
b1001 +
#678350000000
0!
0'
#678360000000
1!
b0 %
1'
b0 +
#678370000000
0!
0'
#678380000000
1!
1$
b1 %
1'
1*
b1 +
#678390000000
0!
0'
#678400000000
1!
b10 %
1'
b10 +
#678410000000
0!
0'
#678420000000
1!
b11 %
1'
b11 +
#678430000000
0!
0'
#678440000000
1!
b100 %
1'
b100 +
#678450000000
0!
0'
#678460000000
1!
b101 %
1'
b101 +
#678470000000
0!
0'
#678480000000
1!
b110 %
1'
b110 +
#678490000000
0!
0'
#678500000000
1!
b111 %
1'
b111 +
#678510000000
0!
0'
#678520000000
1!
0$
b1000 %
1'
0*
b1000 +
#678530000000
0!
0'
#678540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#678550000000
0!
0'
#678560000000
1!
b0 %
1'
b0 +
#678570000000
0!
0'
#678580000000
1!
1$
b1 %
1'
1*
b1 +
#678590000000
0!
0'
#678600000000
1!
b10 %
1'
b10 +
#678610000000
0!
0'
#678620000000
1!
b11 %
1'
b11 +
#678630000000
0!
0'
#678640000000
1!
b100 %
1'
b100 +
#678650000000
0!
0'
#678660000000
1!
b101 %
1'
b101 +
#678670000000
0!
0'
#678680000000
1!
0$
b110 %
1'
0*
b110 +
#678690000000
0!
0'
#678700000000
1!
b111 %
1'
b111 +
#678710000000
0!
0'
#678720000000
1!
b1000 %
1'
b1000 +
#678730000000
0!
0'
#678740000000
1!
b1001 %
1'
b1001 +
#678750000000
1"
1(
#678760000000
0!
0"
b100 &
0'
0(
b100 ,
#678770000000
1!
b0 %
1'
b0 +
#678780000000
0!
0'
#678790000000
1!
1$
b1 %
1'
1*
b1 +
#678800000000
0!
0'
#678810000000
1!
b10 %
1'
b10 +
#678820000000
0!
0'
#678830000000
1!
b11 %
1'
b11 +
#678840000000
0!
0'
#678850000000
1!
b100 %
1'
b100 +
#678860000000
0!
0'
#678870000000
1!
b101 %
1'
b101 +
#678880000000
0!
0'
#678890000000
1!
b110 %
1'
b110 +
#678900000000
0!
0'
#678910000000
1!
b111 %
1'
b111 +
#678920000000
0!
0'
#678930000000
1!
0$
b1000 %
1'
0*
b1000 +
#678940000000
0!
0'
#678950000000
1!
b1001 %
1'
b1001 +
#678960000000
0!
0'
#678970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#678980000000
0!
0'
#678990000000
1!
1$
b1 %
1'
1*
b1 +
#679000000000
0!
0'
#679010000000
1!
b10 %
1'
b10 +
#679020000000
0!
0'
#679030000000
1!
b11 %
1'
b11 +
#679040000000
0!
0'
#679050000000
1!
b100 %
1'
b100 +
#679060000000
0!
0'
#679070000000
1!
b101 %
1'
b101 +
#679080000000
0!
0'
#679090000000
1!
0$
b110 %
1'
0*
b110 +
#679100000000
0!
0'
#679110000000
1!
b111 %
1'
b111 +
#679120000000
0!
0'
#679130000000
1!
b1000 %
1'
b1000 +
#679140000000
0!
0'
#679150000000
1!
b1001 %
1'
b1001 +
#679160000000
0!
0'
#679170000000
1!
b0 %
1'
b0 +
#679180000000
1"
1(
#679190000000
0!
0"
b100 &
0'
0(
b100 ,
#679200000000
1!
1$
b1 %
1'
1*
b1 +
#679210000000
0!
0'
#679220000000
1!
b10 %
1'
b10 +
#679230000000
0!
0'
#679240000000
1!
b11 %
1'
b11 +
#679250000000
0!
0'
#679260000000
1!
b100 %
1'
b100 +
#679270000000
0!
0'
#679280000000
1!
b101 %
1'
b101 +
#679290000000
0!
0'
#679300000000
1!
b110 %
1'
b110 +
#679310000000
0!
0'
#679320000000
1!
b111 %
1'
b111 +
#679330000000
0!
0'
#679340000000
1!
0$
b1000 %
1'
0*
b1000 +
#679350000000
0!
0'
#679360000000
1!
b1001 %
1'
b1001 +
#679370000000
0!
0'
#679380000000
1!
b0 %
1'
b0 +
#679390000000
0!
0'
#679400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#679410000000
0!
0'
#679420000000
1!
b10 %
1'
b10 +
#679430000000
0!
0'
#679440000000
1!
b11 %
1'
b11 +
#679450000000
0!
0'
#679460000000
1!
b100 %
1'
b100 +
#679470000000
0!
0'
#679480000000
1!
b101 %
1'
b101 +
#679490000000
0!
0'
#679500000000
1!
0$
b110 %
1'
0*
b110 +
#679510000000
0!
0'
#679520000000
1!
b111 %
1'
b111 +
#679530000000
0!
0'
#679540000000
1!
b1000 %
1'
b1000 +
#679550000000
0!
0'
#679560000000
1!
b1001 %
1'
b1001 +
#679570000000
0!
0'
#679580000000
1!
b0 %
1'
b0 +
#679590000000
0!
0'
#679600000000
1!
1$
b1 %
1'
1*
b1 +
#679610000000
1"
1(
#679620000000
0!
0"
b100 &
0'
0(
b100 ,
#679630000000
1!
b10 %
1'
b10 +
#679640000000
0!
0'
#679650000000
1!
b11 %
1'
b11 +
#679660000000
0!
0'
#679670000000
1!
b100 %
1'
b100 +
#679680000000
0!
0'
#679690000000
1!
b101 %
1'
b101 +
#679700000000
0!
0'
#679710000000
1!
b110 %
1'
b110 +
#679720000000
0!
0'
#679730000000
1!
b111 %
1'
b111 +
#679740000000
0!
0'
#679750000000
1!
0$
b1000 %
1'
0*
b1000 +
#679760000000
0!
0'
#679770000000
1!
b1001 %
1'
b1001 +
#679780000000
0!
0'
#679790000000
1!
b0 %
1'
b0 +
#679800000000
0!
0'
#679810000000
1!
1$
b1 %
1'
1*
b1 +
#679820000000
0!
0'
#679830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#679840000000
0!
0'
#679850000000
1!
b11 %
1'
b11 +
#679860000000
0!
0'
#679870000000
1!
b100 %
1'
b100 +
#679880000000
0!
0'
#679890000000
1!
b101 %
1'
b101 +
#679900000000
0!
0'
#679910000000
1!
0$
b110 %
1'
0*
b110 +
#679920000000
0!
0'
#679930000000
1!
b111 %
1'
b111 +
#679940000000
0!
0'
#679950000000
1!
b1000 %
1'
b1000 +
#679960000000
0!
0'
#679970000000
1!
b1001 %
1'
b1001 +
#679980000000
0!
0'
#679990000000
1!
b0 %
1'
b0 +
#680000000000
0!
0'
#680010000000
1!
1$
b1 %
1'
1*
b1 +
#680020000000
0!
0'
#680030000000
1!
b10 %
1'
b10 +
#680040000000
1"
1(
#680050000000
0!
0"
b100 &
0'
0(
b100 ,
#680060000000
1!
b11 %
1'
b11 +
#680070000000
0!
0'
#680080000000
1!
b100 %
1'
b100 +
#680090000000
0!
0'
#680100000000
1!
b101 %
1'
b101 +
#680110000000
0!
0'
#680120000000
1!
b110 %
1'
b110 +
#680130000000
0!
0'
#680140000000
1!
b111 %
1'
b111 +
#680150000000
0!
0'
#680160000000
1!
0$
b1000 %
1'
0*
b1000 +
#680170000000
0!
0'
#680180000000
1!
b1001 %
1'
b1001 +
#680190000000
0!
0'
#680200000000
1!
b0 %
1'
b0 +
#680210000000
0!
0'
#680220000000
1!
1$
b1 %
1'
1*
b1 +
#680230000000
0!
0'
#680240000000
1!
b10 %
1'
b10 +
#680250000000
0!
0'
#680260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#680270000000
0!
0'
#680280000000
1!
b100 %
1'
b100 +
#680290000000
0!
0'
#680300000000
1!
b101 %
1'
b101 +
#680310000000
0!
0'
#680320000000
1!
0$
b110 %
1'
0*
b110 +
#680330000000
0!
0'
#680340000000
1!
b111 %
1'
b111 +
#680350000000
0!
0'
#680360000000
1!
b1000 %
1'
b1000 +
#680370000000
0!
0'
#680380000000
1!
b1001 %
1'
b1001 +
#680390000000
0!
0'
#680400000000
1!
b0 %
1'
b0 +
#680410000000
0!
0'
#680420000000
1!
1$
b1 %
1'
1*
b1 +
#680430000000
0!
0'
#680440000000
1!
b10 %
1'
b10 +
#680450000000
0!
0'
#680460000000
1!
b11 %
1'
b11 +
#680470000000
1"
1(
#680480000000
0!
0"
b100 &
0'
0(
b100 ,
#680490000000
1!
b100 %
1'
b100 +
#680500000000
0!
0'
#680510000000
1!
b101 %
1'
b101 +
#680520000000
0!
0'
#680530000000
1!
b110 %
1'
b110 +
#680540000000
0!
0'
#680550000000
1!
b111 %
1'
b111 +
#680560000000
0!
0'
#680570000000
1!
0$
b1000 %
1'
0*
b1000 +
#680580000000
0!
0'
#680590000000
1!
b1001 %
1'
b1001 +
#680600000000
0!
0'
#680610000000
1!
b0 %
1'
b0 +
#680620000000
0!
0'
#680630000000
1!
1$
b1 %
1'
1*
b1 +
#680640000000
0!
0'
#680650000000
1!
b10 %
1'
b10 +
#680660000000
0!
0'
#680670000000
1!
b11 %
1'
b11 +
#680680000000
0!
0'
#680690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#680700000000
0!
0'
#680710000000
1!
b101 %
1'
b101 +
#680720000000
0!
0'
#680730000000
1!
0$
b110 %
1'
0*
b110 +
#680740000000
0!
0'
#680750000000
1!
b111 %
1'
b111 +
#680760000000
0!
0'
#680770000000
1!
b1000 %
1'
b1000 +
#680780000000
0!
0'
#680790000000
1!
b1001 %
1'
b1001 +
#680800000000
0!
0'
#680810000000
1!
b0 %
1'
b0 +
#680820000000
0!
0'
#680830000000
1!
1$
b1 %
1'
1*
b1 +
#680840000000
0!
0'
#680850000000
1!
b10 %
1'
b10 +
#680860000000
0!
0'
#680870000000
1!
b11 %
1'
b11 +
#680880000000
0!
0'
#680890000000
1!
b100 %
1'
b100 +
#680900000000
1"
1(
#680910000000
0!
0"
b100 &
0'
0(
b100 ,
#680920000000
1!
b101 %
1'
b101 +
#680930000000
0!
0'
#680940000000
1!
b110 %
1'
b110 +
#680950000000
0!
0'
#680960000000
1!
b111 %
1'
b111 +
#680970000000
0!
0'
#680980000000
1!
0$
b1000 %
1'
0*
b1000 +
#680990000000
0!
0'
#681000000000
1!
b1001 %
1'
b1001 +
#681010000000
0!
0'
#681020000000
1!
b0 %
1'
b0 +
#681030000000
0!
0'
#681040000000
1!
1$
b1 %
1'
1*
b1 +
#681050000000
0!
0'
#681060000000
1!
b10 %
1'
b10 +
#681070000000
0!
0'
#681080000000
1!
b11 %
1'
b11 +
#681090000000
0!
0'
#681100000000
1!
b100 %
1'
b100 +
#681110000000
0!
0'
#681120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#681130000000
0!
0'
#681140000000
1!
0$
b110 %
1'
0*
b110 +
#681150000000
0!
0'
#681160000000
1!
b111 %
1'
b111 +
#681170000000
0!
0'
#681180000000
1!
b1000 %
1'
b1000 +
#681190000000
0!
0'
#681200000000
1!
b1001 %
1'
b1001 +
#681210000000
0!
0'
#681220000000
1!
b0 %
1'
b0 +
#681230000000
0!
0'
#681240000000
1!
1$
b1 %
1'
1*
b1 +
#681250000000
0!
0'
#681260000000
1!
b10 %
1'
b10 +
#681270000000
0!
0'
#681280000000
1!
b11 %
1'
b11 +
#681290000000
0!
0'
#681300000000
1!
b100 %
1'
b100 +
#681310000000
0!
0'
#681320000000
1!
b101 %
1'
b101 +
#681330000000
1"
1(
#681340000000
0!
0"
b100 &
0'
0(
b100 ,
#681350000000
1!
b110 %
1'
b110 +
#681360000000
0!
0'
#681370000000
1!
b111 %
1'
b111 +
#681380000000
0!
0'
#681390000000
1!
0$
b1000 %
1'
0*
b1000 +
#681400000000
0!
0'
#681410000000
1!
b1001 %
1'
b1001 +
#681420000000
0!
0'
#681430000000
1!
b0 %
1'
b0 +
#681440000000
0!
0'
#681450000000
1!
1$
b1 %
1'
1*
b1 +
#681460000000
0!
0'
#681470000000
1!
b10 %
1'
b10 +
#681480000000
0!
0'
#681490000000
1!
b11 %
1'
b11 +
#681500000000
0!
0'
#681510000000
1!
b100 %
1'
b100 +
#681520000000
0!
0'
#681530000000
1!
b101 %
1'
b101 +
#681540000000
0!
0'
#681550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#681560000000
0!
0'
#681570000000
1!
b111 %
1'
b111 +
#681580000000
0!
0'
#681590000000
1!
b1000 %
1'
b1000 +
#681600000000
0!
0'
#681610000000
1!
b1001 %
1'
b1001 +
#681620000000
0!
0'
#681630000000
1!
b0 %
1'
b0 +
#681640000000
0!
0'
#681650000000
1!
1$
b1 %
1'
1*
b1 +
#681660000000
0!
0'
#681670000000
1!
b10 %
1'
b10 +
#681680000000
0!
0'
#681690000000
1!
b11 %
1'
b11 +
#681700000000
0!
0'
#681710000000
1!
b100 %
1'
b100 +
#681720000000
0!
0'
#681730000000
1!
b101 %
1'
b101 +
#681740000000
0!
0'
#681750000000
1!
0$
b110 %
1'
0*
b110 +
#681760000000
1"
1(
#681770000000
0!
0"
b100 &
0'
0(
b100 ,
#681780000000
1!
1$
b111 %
1'
1*
b111 +
#681790000000
0!
0'
#681800000000
1!
0$
b1000 %
1'
0*
b1000 +
#681810000000
0!
0'
#681820000000
1!
b1001 %
1'
b1001 +
#681830000000
0!
0'
#681840000000
1!
b0 %
1'
b0 +
#681850000000
0!
0'
#681860000000
1!
1$
b1 %
1'
1*
b1 +
#681870000000
0!
0'
#681880000000
1!
b10 %
1'
b10 +
#681890000000
0!
0'
#681900000000
1!
b11 %
1'
b11 +
#681910000000
0!
0'
#681920000000
1!
b100 %
1'
b100 +
#681930000000
0!
0'
#681940000000
1!
b101 %
1'
b101 +
#681950000000
0!
0'
#681960000000
1!
b110 %
1'
b110 +
#681970000000
0!
0'
#681980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#681990000000
0!
0'
#682000000000
1!
b1000 %
1'
b1000 +
#682010000000
0!
0'
#682020000000
1!
b1001 %
1'
b1001 +
#682030000000
0!
0'
#682040000000
1!
b0 %
1'
b0 +
#682050000000
0!
0'
#682060000000
1!
1$
b1 %
1'
1*
b1 +
#682070000000
0!
0'
#682080000000
1!
b10 %
1'
b10 +
#682090000000
0!
0'
#682100000000
1!
b11 %
1'
b11 +
#682110000000
0!
0'
#682120000000
1!
b100 %
1'
b100 +
#682130000000
0!
0'
#682140000000
1!
b101 %
1'
b101 +
#682150000000
0!
0'
#682160000000
1!
0$
b110 %
1'
0*
b110 +
#682170000000
0!
0'
#682180000000
1!
b111 %
1'
b111 +
#682190000000
1"
1(
#682200000000
0!
0"
b100 &
0'
0(
b100 ,
#682210000000
1!
b1000 %
1'
b1000 +
#682220000000
0!
0'
#682230000000
1!
b1001 %
1'
b1001 +
#682240000000
0!
0'
#682250000000
1!
b0 %
1'
b0 +
#682260000000
0!
0'
#682270000000
1!
1$
b1 %
1'
1*
b1 +
#682280000000
0!
0'
#682290000000
1!
b10 %
1'
b10 +
#682300000000
0!
0'
#682310000000
1!
b11 %
1'
b11 +
#682320000000
0!
0'
#682330000000
1!
b100 %
1'
b100 +
#682340000000
0!
0'
#682350000000
1!
b101 %
1'
b101 +
#682360000000
0!
0'
#682370000000
1!
b110 %
1'
b110 +
#682380000000
0!
0'
#682390000000
1!
b111 %
1'
b111 +
#682400000000
0!
0'
#682410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#682420000000
0!
0'
#682430000000
1!
b1001 %
1'
b1001 +
#682440000000
0!
0'
#682450000000
1!
b0 %
1'
b0 +
#682460000000
0!
0'
#682470000000
1!
1$
b1 %
1'
1*
b1 +
#682480000000
0!
0'
#682490000000
1!
b10 %
1'
b10 +
#682500000000
0!
0'
#682510000000
1!
b11 %
1'
b11 +
#682520000000
0!
0'
#682530000000
1!
b100 %
1'
b100 +
#682540000000
0!
0'
#682550000000
1!
b101 %
1'
b101 +
#682560000000
0!
0'
#682570000000
1!
0$
b110 %
1'
0*
b110 +
#682580000000
0!
0'
#682590000000
1!
b111 %
1'
b111 +
#682600000000
0!
0'
#682610000000
1!
b1000 %
1'
b1000 +
#682620000000
1"
1(
#682630000000
0!
0"
b100 &
0'
0(
b100 ,
#682640000000
1!
b1001 %
1'
b1001 +
#682650000000
0!
0'
#682660000000
1!
b0 %
1'
b0 +
#682670000000
0!
0'
#682680000000
1!
1$
b1 %
1'
1*
b1 +
#682690000000
0!
0'
#682700000000
1!
b10 %
1'
b10 +
#682710000000
0!
0'
#682720000000
1!
b11 %
1'
b11 +
#682730000000
0!
0'
#682740000000
1!
b100 %
1'
b100 +
#682750000000
0!
0'
#682760000000
1!
b101 %
1'
b101 +
#682770000000
0!
0'
#682780000000
1!
b110 %
1'
b110 +
#682790000000
0!
0'
#682800000000
1!
b111 %
1'
b111 +
#682810000000
0!
0'
#682820000000
1!
0$
b1000 %
1'
0*
b1000 +
#682830000000
0!
0'
#682840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#682850000000
0!
0'
#682860000000
1!
b0 %
1'
b0 +
#682870000000
0!
0'
#682880000000
1!
1$
b1 %
1'
1*
b1 +
#682890000000
0!
0'
#682900000000
1!
b10 %
1'
b10 +
#682910000000
0!
0'
#682920000000
1!
b11 %
1'
b11 +
#682930000000
0!
0'
#682940000000
1!
b100 %
1'
b100 +
#682950000000
0!
0'
#682960000000
1!
b101 %
1'
b101 +
#682970000000
0!
0'
#682980000000
1!
0$
b110 %
1'
0*
b110 +
#682990000000
0!
0'
#683000000000
1!
b111 %
1'
b111 +
#683010000000
0!
0'
#683020000000
1!
b1000 %
1'
b1000 +
#683030000000
0!
0'
#683040000000
1!
b1001 %
1'
b1001 +
#683050000000
1"
1(
#683060000000
0!
0"
b100 &
0'
0(
b100 ,
#683070000000
1!
b0 %
1'
b0 +
#683080000000
0!
0'
#683090000000
1!
1$
b1 %
1'
1*
b1 +
#683100000000
0!
0'
#683110000000
1!
b10 %
1'
b10 +
#683120000000
0!
0'
#683130000000
1!
b11 %
1'
b11 +
#683140000000
0!
0'
#683150000000
1!
b100 %
1'
b100 +
#683160000000
0!
0'
#683170000000
1!
b101 %
1'
b101 +
#683180000000
0!
0'
#683190000000
1!
b110 %
1'
b110 +
#683200000000
0!
0'
#683210000000
1!
b111 %
1'
b111 +
#683220000000
0!
0'
#683230000000
1!
0$
b1000 %
1'
0*
b1000 +
#683240000000
0!
0'
#683250000000
1!
b1001 %
1'
b1001 +
#683260000000
0!
0'
#683270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#683280000000
0!
0'
#683290000000
1!
1$
b1 %
1'
1*
b1 +
#683300000000
0!
0'
#683310000000
1!
b10 %
1'
b10 +
#683320000000
0!
0'
#683330000000
1!
b11 %
1'
b11 +
#683340000000
0!
0'
#683350000000
1!
b100 %
1'
b100 +
#683360000000
0!
0'
#683370000000
1!
b101 %
1'
b101 +
#683380000000
0!
0'
#683390000000
1!
0$
b110 %
1'
0*
b110 +
#683400000000
0!
0'
#683410000000
1!
b111 %
1'
b111 +
#683420000000
0!
0'
#683430000000
1!
b1000 %
1'
b1000 +
#683440000000
0!
0'
#683450000000
1!
b1001 %
1'
b1001 +
#683460000000
0!
0'
#683470000000
1!
b0 %
1'
b0 +
#683480000000
1"
1(
#683490000000
0!
0"
b100 &
0'
0(
b100 ,
#683500000000
1!
1$
b1 %
1'
1*
b1 +
#683510000000
0!
0'
#683520000000
1!
b10 %
1'
b10 +
#683530000000
0!
0'
#683540000000
1!
b11 %
1'
b11 +
#683550000000
0!
0'
#683560000000
1!
b100 %
1'
b100 +
#683570000000
0!
0'
#683580000000
1!
b101 %
1'
b101 +
#683590000000
0!
0'
#683600000000
1!
b110 %
1'
b110 +
#683610000000
0!
0'
#683620000000
1!
b111 %
1'
b111 +
#683630000000
0!
0'
#683640000000
1!
0$
b1000 %
1'
0*
b1000 +
#683650000000
0!
0'
#683660000000
1!
b1001 %
1'
b1001 +
#683670000000
0!
0'
#683680000000
1!
b0 %
1'
b0 +
#683690000000
0!
0'
#683700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#683710000000
0!
0'
#683720000000
1!
b10 %
1'
b10 +
#683730000000
0!
0'
#683740000000
1!
b11 %
1'
b11 +
#683750000000
0!
0'
#683760000000
1!
b100 %
1'
b100 +
#683770000000
0!
0'
#683780000000
1!
b101 %
1'
b101 +
#683790000000
0!
0'
#683800000000
1!
0$
b110 %
1'
0*
b110 +
#683810000000
0!
0'
#683820000000
1!
b111 %
1'
b111 +
#683830000000
0!
0'
#683840000000
1!
b1000 %
1'
b1000 +
#683850000000
0!
0'
#683860000000
1!
b1001 %
1'
b1001 +
#683870000000
0!
0'
#683880000000
1!
b0 %
1'
b0 +
#683890000000
0!
0'
#683900000000
1!
1$
b1 %
1'
1*
b1 +
#683910000000
1"
1(
#683920000000
0!
0"
b100 &
0'
0(
b100 ,
#683930000000
1!
b10 %
1'
b10 +
#683940000000
0!
0'
#683950000000
1!
b11 %
1'
b11 +
#683960000000
0!
0'
#683970000000
1!
b100 %
1'
b100 +
#683980000000
0!
0'
#683990000000
1!
b101 %
1'
b101 +
#684000000000
0!
0'
#684010000000
1!
b110 %
1'
b110 +
#684020000000
0!
0'
#684030000000
1!
b111 %
1'
b111 +
#684040000000
0!
0'
#684050000000
1!
0$
b1000 %
1'
0*
b1000 +
#684060000000
0!
0'
#684070000000
1!
b1001 %
1'
b1001 +
#684080000000
0!
0'
#684090000000
1!
b0 %
1'
b0 +
#684100000000
0!
0'
#684110000000
1!
1$
b1 %
1'
1*
b1 +
#684120000000
0!
0'
#684130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#684140000000
0!
0'
#684150000000
1!
b11 %
1'
b11 +
#684160000000
0!
0'
#684170000000
1!
b100 %
1'
b100 +
#684180000000
0!
0'
#684190000000
1!
b101 %
1'
b101 +
#684200000000
0!
0'
#684210000000
1!
0$
b110 %
1'
0*
b110 +
#684220000000
0!
0'
#684230000000
1!
b111 %
1'
b111 +
#684240000000
0!
0'
#684250000000
1!
b1000 %
1'
b1000 +
#684260000000
0!
0'
#684270000000
1!
b1001 %
1'
b1001 +
#684280000000
0!
0'
#684290000000
1!
b0 %
1'
b0 +
#684300000000
0!
0'
#684310000000
1!
1$
b1 %
1'
1*
b1 +
#684320000000
0!
0'
#684330000000
1!
b10 %
1'
b10 +
#684340000000
1"
1(
#684350000000
0!
0"
b100 &
0'
0(
b100 ,
#684360000000
1!
b11 %
1'
b11 +
#684370000000
0!
0'
#684380000000
1!
b100 %
1'
b100 +
#684390000000
0!
0'
#684400000000
1!
b101 %
1'
b101 +
#684410000000
0!
0'
#684420000000
1!
b110 %
1'
b110 +
#684430000000
0!
0'
#684440000000
1!
b111 %
1'
b111 +
#684450000000
0!
0'
#684460000000
1!
0$
b1000 %
1'
0*
b1000 +
#684470000000
0!
0'
#684480000000
1!
b1001 %
1'
b1001 +
#684490000000
0!
0'
#684500000000
1!
b0 %
1'
b0 +
#684510000000
0!
0'
#684520000000
1!
1$
b1 %
1'
1*
b1 +
#684530000000
0!
0'
#684540000000
1!
b10 %
1'
b10 +
#684550000000
0!
0'
#684560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#684570000000
0!
0'
#684580000000
1!
b100 %
1'
b100 +
#684590000000
0!
0'
#684600000000
1!
b101 %
1'
b101 +
#684610000000
0!
0'
#684620000000
1!
0$
b110 %
1'
0*
b110 +
#684630000000
0!
0'
#684640000000
1!
b111 %
1'
b111 +
#684650000000
0!
0'
#684660000000
1!
b1000 %
1'
b1000 +
#684670000000
0!
0'
#684680000000
1!
b1001 %
1'
b1001 +
#684690000000
0!
0'
#684700000000
1!
b0 %
1'
b0 +
#684710000000
0!
0'
#684720000000
1!
1$
b1 %
1'
1*
b1 +
#684730000000
0!
0'
#684740000000
1!
b10 %
1'
b10 +
#684750000000
0!
0'
#684760000000
1!
b11 %
1'
b11 +
#684770000000
1"
1(
#684780000000
0!
0"
b100 &
0'
0(
b100 ,
#684790000000
1!
b100 %
1'
b100 +
#684800000000
0!
0'
#684810000000
1!
b101 %
1'
b101 +
#684820000000
0!
0'
#684830000000
1!
b110 %
1'
b110 +
#684840000000
0!
0'
#684850000000
1!
b111 %
1'
b111 +
#684860000000
0!
0'
#684870000000
1!
0$
b1000 %
1'
0*
b1000 +
#684880000000
0!
0'
#684890000000
1!
b1001 %
1'
b1001 +
#684900000000
0!
0'
#684910000000
1!
b0 %
1'
b0 +
#684920000000
0!
0'
#684930000000
1!
1$
b1 %
1'
1*
b1 +
#684940000000
0!
0'
#684950000000
1!
b10 %
1'
b10 +
#684960000000
0!
0'
#684970000000
1!
b11 %
1'
b11 +
#684980000000
0!
0'
#684990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#685000000000
0!
0'
#685010000000
1!
b101 %
1'
b101 +
#685020000000
0!
0'
#685030000000
1!
0$
b110 %
1'
0*
b110 +
#685040000000
0!
0'
#685050000000
1!
b111 %
1'
b111 +
#685060000000
0!
0'
#685070000000
1!
b1000 %
1'
b1000 +
#685080000000
0!
0'
#685090000000
1!
b1001 %
1'
b1001 +
#685100000000
0!
0'
#685110000000
1!
b0 %
1'
b0 +
#685120000000
0!
0'
#685130000000
1!
1$
b1 %
1'
1*
b1 +
#685140000000
0!
0'
#685150000000
1!
b10 %
1'
b10 +
#685160000000
0!
0'
#685170000000
1!
b11 %
1'
b11 +
#685180000000
0!
0'
#685190000000
1!
b100 %
1'
b100 +
#685200000000
1"
1(
#685210000000
0!
0"
b100 &
0'
0(
b100 ,
#685220000000
1!
b101 %
1'
b101 +
#685230000000
0!
0'
#685240000000
1!
b110 %
1'
b110 +
#685250000000
0!
0'
#685260000000
1!
b111 %
1'
b111 +
#685270000000
0!
0'
#685280000000
1!
0$
b1000 %
1'
0*
b1000 +
#685290000000
0!
0'
#685300000000
1!
b1001 %
1'
b1001 +
#685310000000
0!
0'
#685320000000
1!
b0 %
1'
b0 +
#685330000000
0!
0'
#685340000000
1!
1$
b1 %
1'
1*
b1 +
#685350000000
0!
0'
#685360000000
1!
b10 %
1'
b10 +
#685370000000
0!
0'
#685380000000
1!
b11 %
1'
b11 +
#685390000000
0!
0'
#685400000000
1!
b100 %
1'
b100 +
#685410000000
0!
0'
#685420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#685430000000
0!
0'
#685440000000
1!
0$
b110 %
1'
0*
b110 +
#685450000000
0!
0'
#685460000000
1!
b111 %
1'
b111 +
#685470000000
0!
0'
#685480000000
1!
b1000 %
1'
b1000 +
#685490000000
0!
0'
#685500000000
1!
b1001 %
1'
b1001 +
#685510000000
0!
0'
#685520000000
1!
b0 %
1'
b0 +
#685530000000
0!
0'
#685540000000
1!
1$
b1 %
1'
1*
b1 +
#685550000000
0!
0'
#685560000000
1!
b10 %
1'
b10 +
#685570000000
0!
0'
#685580000000
1!
b11 %
1'
b11 +
#685590000000
0!
0'
#685600000000
1!
b100 %
1'
b100 +
#685610000000
0!
0'
#685620000000
1!
b101 %
1'
b101 +
#685630000000
1"
1(
#685640000000
0!
0"
b100 &
0'
0(
b100 ,
#685650000000
1!
b110 %
1'
b110 +
#685660000000
0!
0'
#685670000000
1!
b111 %
1'
b111 +
#685680000000
0!
0'
#685690000000
1!
0$
b1000 %
1'
0*
b1000 +
#685700000000
0!
0'
#685710000000
1!
b1001 %
1'
b1001 +
#685720000000
0!
0'
#685730000000
1!
b0 %
1'
b0 +
#685740000000
0!
0'
#685750000000
1!
1$
b1 %
1'
1*
b1 +
#685760000000
0!
0'
#685770000000
1!
b10 %
1'
b10 +
#685780000000
0!
0'
#685790000000
1!
b11 %
1'
b11 +
#685800000000
0!
0'
#685810000000
1!
b100 %
1'
b100 +
#685820000000
0!
0'
#685830000000
1!
b101 %
1'
b101 +
#685840000000
0!
0'
#685850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#685860000000
0!
0'
#685870000000
1!
b111 %
1'
b111 +
#685880000000
0!
0'
#685890000000
1!
b1000 %
1'
b1000 +
#685900000000
0!
0'
#685910000000
1!
b1001 %
1'
b1001 +
#685920000000
0!
0'
#685930000000
1!
b0 %
1'
b0 +
#685940000000
0!
0'
#685950000000
1!
1$
b1 %
1'
1*
b1 +
#685960000000
0!
0'
#685970000000
1!
b10 %
1'
b10 +
#685980000000
0!
0'
#685990000000
1!
b11 %
1'
b11 +
#686000000000
0!
0'
#686010000000
1!
b100 %
1'
b100 +
#686020000000
0!
0'
#686030000000
1!
b101 %
1'
b101 +
#686040000000
0!
0'
#686050000000
1!
0$
b110 %
1'
0*
b110 +
#686060000000
1"
1(
#686070000000
0!
0"
b100 &
0'
0(
b100 ,
#686080000000
1!
1$
b111 %
1'
1*
b111 +
#686090000000
0!
0'
#686100000000
1!
0$
b1000 %
1'
0*
b1000 +
#686110000000
0!
0'
#686120000000
1!
b1001 %
1'
b1001 +
#686130000000
0!
0'
#686140000000
1!
b0 %
1'
b0 +
#686150000000
0!
0'
#686160000000
1!
1$
b1 %
1'
1*
b1 +
#686170000000
0!
0'
#686180000000
1!
b10 %
1'
b10 +
#686190000000
0!
0'
#686200000000
1!
b11 %
1'
b11 +
#686210000000
0!
0'
#686220000000
1!
b100 %
1'
b100 +
#686230000000
0!
0'
#686240000000
1!
b101 %
1'
b101 +
#686250000000
0!
0'
#686260000000
1!
b110 %
1'
b110 +
#686270000000
0!
0'
#686280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#686290000000
0!
0'
#686300000000
1!
b1000 %
1'
b1000 +
#686310000000
0!
0'
#686320000000
1!
b1001 %
1'
b1001 +
#686330000000
0!
0'
#686340000000
1!
b0 %
1'
b0 +
#686350000000
0!
0'
#686360000000
1!
1$
b1 %
1'
1*
b1 +
#686370000000
0!
0'
#686380000000
1!
b10 %
1'
b10 +
#686390000000
0!
0'
#686400000000
1!
b11 %
1'
b11 +
#686410000000
0!
0'
#686420000000
1!
b100 %
1'
b100 +
#686430000000
0!
0'
#686440000000
1!
b101 %
1'
b101 +
#686450000000
0!
0'
#686460000000
1!
0$
b110 %
1'
0*
b110 +
#686470000000
0!
0'
#686480000000
1!
b111 %
1'
b111 +
#686490000000
1"
1(
#686500000000
0!
0"
b100 &
0'
0(
b100 ,
#686510000000
1!
b1000 %
1'
b1000 +
#686520000000
0!
0'
#686530000000
1!
b1001 %
1'
b1001 +
#686540000000
0!
0'
#686550000000
1!
b0 %
1'
b0 +
#686560000000
0!
0'
#686570000000
1!
1$
b1 %
1'
1*
b1 +
#686580000000
0!
0'
#686590000000
1!
b10 %
1'
b10 +
#686600000000
0!
0'
#686610000000
1!
b11 %
1'
b11 +
#686620000000
0!
0'
#686630000000
1!
b100 %
1'
b100 +
#686640000000
0!
0'
#686650000000
1!
b101 %
1'
b101 +
#686660000000
0!
0'
#686670000000
1!
b110 %
1'
b110 +
#686680000000
0!
0'
#686690000000
1!
b111 %
1'
b111 +
#686700000000
0!
0'
#686710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#686720000000
0!
0'
#686730000000
1!
b1001 %
1'
b1001 +
#686740000000
0!
0'
#686750000000
1!
b0 %
1'
b0 +
#686760000000
0!
0'
#686770000000
1!
1$
b1 %
1'
1*
b1 +
#686780000000
0!
0'
#686790000000
1!
b10 %
1'
b10 +
#686800000000
0!
0'
#686810000000
1!
b11 %
1'
b11 +
#686820000000
0!
0'
#686830000000
1!
b100 %
1'
b100 +
#686840000000
0!
0'
#686850000000
1!
b101 %
1'
b101 +
#686860000000
0!
0'
#686870000000
1!
0$
b110 %
1'
0*
b110 +
#686880000000
0!
0'
#686890000000
1!
b111 %
1'
b111 +
#686900000000
0!
0'
#686910000000
1!
b1000 %
1'
b1000 +
#686920000000
1"
1(
#686930000000
0!
0"
b100 &
0'
0(
b100 ,
#686940000000
1!
b1001 %
1'
b1001 +
#686950000000
0!
0'
#686960000000
1!
b0 %
1'
b0 +
#686970000000
0!
0'
#686980000000
1!
1$
b1 %
1'
1*
b1 +
#686990000000
0!
0'
#687000000000
1!
b10 %
1'
b10 +
#687010000000
0!
0'
#687020000000
1!
b11 %
1'
b11 +
#687030000000
0!
0'
#687040000000
1!
b100 %
1'
b100 +
#687050000000
0!
0'
#687060000000
1!
b101 %
1'
b101 +
#687070000000
0!
0'
#687080000000
1!
b110 %
1'
b110 +
#687090000000
0!
0'
#687100000000
1!
b111 %
1'
b111 +
#687110000000
0!
0'
#687120000000
1!
0$
b1000 %
1'
0*
b1000 +
#687130000000
0!
0'
#687140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#687150000000
0!
0'
#687160000000
1!
b0 %
1'
b0 +
#687170000000
0!
0'
#687180000000
1!
1$
b1 %
1'
1*
b1 +
#687190000000
0!
0'
#687200000000
1!
b10 %
1'
b10 +
#687210000000
0!
0'
#687220000000
1!
b11 %
1'
b11 +
#687230000000
0!
0'
#687240000000
1!
b100 %
1'
b100 +
#687250000000
0!
0'
#687260000000
1!
b101 %
1'
b101 +
#687270000000
0!
0'
#687280000000
1!
0$
b110 %
1'
0*
b110 +
#687290000000
0!
0'
#687300000000
1!
b111 %
1'
b111 +
#687310000000
0!
0'
#687320000000
1!
b1000 %
1'
b1000 +
#687330000000
0!
0'
#687340000000
1!
b1001 %
1'
b1001 +
#687350000000
1"
1(
#687360000000
0!
0"
b100 &
0'
0(
b100 ,
#687370000000
1!
b0 %
1'
b0 +
#687380000000
0!
0'
#687390000000
1!
1$
b1 %
1'
1*
b1 +
#687400000000
0!
0'
#687410000000
1!
b10 %
1'
b10 +
#687420000000
0!
0'
#687430000000
1!
b11 %
1'
b11 +
#687440000000
0!
0'
#687450000000
1!
b100 %
1'
b100 +
#687460000000
0!
0'
#687470000000
1!
b101 %
1'
b101 +
#687480000000
0!
0'
#687490000000
1!
b110 %
1'
b110 +
#687500000000
0!
0'
#687510000000
1!
b111 %
1'
b111 +
#687520000000
0!
0'
#687530000000
1!
0$
b1000 %
1'
0*
b1000 +
#687540000000
0!
0'
#687550000000
1!
b1001 %
1'
b1001 +
#687560000000
0!
0'
#687570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#687580000000
0!
0'
#687590000000
1!
1$
b1 %
1'
1*
b1 +
#687600000000
0!
0'
#687610000000
1!
b10 %
1'
b10 +
#687620000000
0!
0'
#687630000000
1!
b11 %
1'
b11 +
#687640000000
0!
0'
#687650000000
1!
b100 %
1'
b100 +
#687660000000
0!
0'
#687670000000
1!
b101 %
1'
b101 +
#687680000000
0!
0'
#687690000000
1!
0$
b110 %
1'
0*
b110 +
#687700000000
0!
0'
#687710000000
1!
b111 %
1'
b111 +
#687720000000
0!
0'
#687730000000
1!
b1000 %
1'
b1000 +
#687740000000
0!
0'
#687750000000
1!
b1001 %
1'
b1001 +
#687760000000
0!
0'
#687770000000
1!
b0 %
1'
b0 +
#687780000000
1"
1(
#687790000000
0!
0"
b100 &
0'
0(
b100 ,
#687800000000
1!
1$
b1 %
1'
1*
b1 +
#687810000000
0!
0'
#687820000000
1!
b10 %
1'
b10 +
#687830000000
0!
0'
#687840000000
1!
b11 %
1'
b11 +
#687850000000
0!
0'
#687860000000
1!
b100 %
1'
b100 +
#687870000000
0!
0'
#687880000000
1!
b101 %
1'
b101 +
#687890000000
0!
0'
#687900000000
1!
b110 %
1'
b110 +
#687910000000
0!
0'
#687920000000
1!
b111 %
1'
b111 +
#687930000000
0!
0'
#687940000000
1!
0$
b1000 %
1'
0*
b1000 +
#687950000000
0!
0'
#687960000000
1!
b1001 %
1'
b1001 +
#687970000000
0!
0'
#687980000000
1!
b0 %
1'
b0 +
#687990000000
0!
0'
#688000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#688010000000
0!
0'
#688020000000
1!
b10 %
1'
b10 +
#688030000000
0!
0'
#688040000000
1!
b11 %
1'
b11 +
#688050000000
0!
0'
#688060000000
1!
b100 %
1'
b100 +
#688070000000
0!
0'
#688080000000
1!
b101 %
1'
b101 +
#688090000000
0!
0'
#688100000000
1!
0$
b110 %
1'
0*
b110 +
#688110000000
0!
0'
#688120000000
1!
b111 %
1'
b111 +
#688130000000
0!
0'
#688140000000
1!
b1000 %
1'
b1000 +
#688150000000
0!
0'
#688160000000
1!
b1001 %
1'
b1001 +
#688170000000
0!
0'
#688180000000
1!
b0 %
1'
b0 +
#688190000000
0!
0'
#688200000000
1!
1$
b1 %
1'
1*
b1 +
#688210000000
1"
1(
#688220000000
0!
0"
b100 &
0'
0(
b100 ,
#688230000000
1!
b10 %
1'
b10 +
#688240000000
0!
0'
#688250000000
1!
b11 %
1'
b11 +
#688260000000
0!
0'
#688270000000
1!
b100 %
1'
b100 +
#688280000000
0!
0'
#688290000000
1!
b101 %
1'
b101 +
#688300000000
0!
0'
#688310000000
1!
b110 %
1'
b110 +
#688320000000
0!
0'
#688330000000
1!
b111 %
1'
b111 +
#688340000000
0!
0'
#688350000000
1!
0$
b1000 %
1'
0*
b1000 +
#688360000000
0!
0'
#688370000000
1!
b1001 %
1'
b1001 +
#688380000000
0!
0'
#688390000000
1!
b0 %
1'
b0 +
#688400000000
0!
0'
#688410000000
1!
1$
b1 %
1'
1*
b1 +
#688420000000
0!
0'
#688430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#688440000000
0!
0'
#688450000000
1!
b11 %
1'
b11 +
#688460000000
0!
0'
#688470000000
1!
b100 %
1'
b100 +
#688480000000
0!
0'
#688490000000
1!
b101 %
1'
b101 +
#688500000000
0!
0'
#688510000000
1!
0$
b110 %
1'
0*
b110 +
#688520000000
0!
0'
#688530000000
1!
b111 %
1'
b111 +
#688540000000
0!
0'
#688550000000
1!
b1000 %
1'
b1000 +
#688560000000
0!
0'
#688570000000
1!
b1001 %
1'
b1001 +
#688580000000
0!
0'
#688590000000
1!
b0 %
1'
b0 +
#688600000000
0!
0'
#688610000000
1!
1$
b1 %
1'
1*
b1 +
#688620000000
0!
0'
#688630000000
1!
b10 %
1'
b10 +
#688640000000
1"
1(
#688650000000
0!
0"
b100 &
0'
0(
b100 ,
#688660000000
1!
b11 %
1'
b11 +
#688670000000
0!
0'
#688680000000
1!
b100 %
1'
b100 +
#688690000000
0!
0'
#688700000000
1!
b101 %
1'
b101 +
#688710000000
0!
0'
#688720000000
1!
b110 %
1'
b110 +
#688730000000
0!
0'
#688740000000
1!
b111 %
1'
b111 +
#688750000000
0!
0'
#688760000000
1!
0$
b1000 %
1'
0*
b1000 +
#688770000000
0!
0'
#688780000000
1!
b1001 %
1'
b1001 +
#688790000000
0!
0'
#688800000000
1!
b0 %
1'
b0 +
#688810000000
0!
0'
#688820000000
1!
1$
b1 %
1'
1*
b1 +
#688830000000
0!
0'
#688840000000
1!
b10 %
1'
b10 +
#688850000000
0!
0'
#688860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#688870000000
0!
0'
#688880000000
1!
b100 %
1'
b100 +
#688890000000
0!
0'
#688900000000
1!
b101 %
1'
b101 +
#688910000000
0!
0'
#688920000000
1!
0$
b110 %
1'
0*
b110 +
#688930000000
0!
0'
#688940000000
1!
b111 %
1'
b111 +
#688950000000
0!
0'
#688960000000
1!
b1000 %
1'
b1000 +
#688970000000
0!
0'
#688980000000
1!
b1001 %
1'
b1001 +
#688990000000
0!
0'
#689000000000
1!
b0 %
1'
b0 +
#689010000000
0!
0'
#689020000000
1!
1$
b1 %
1'
1*
b1 +
#689030000000
0!
0'
#689040000000
1!
b10 %
1'
b10 +
#689050000000
0!
0'
#689060000000
1!
b11 %
1'
b11 +
#689070000000
1"
1(
#689080000000
0!
0"
b100 &
0'
0(
b100 ,
#689090000000
1!
b100 %
1'
b100 +
#689100000000
0!
0'
#689110000000
1!
b101 %
1'
b101 +
#689120000000
0!
0'
#689130000000
1!
b110 %
1'
b110 +
#689140000000
0!
0'
#689150000000
1!
b111 %
1'
b111 +
#689160000000
0!
0'
#689170000000
1!
0$
b1000 %
1'
0*
b1000 +
#689180000000
0!
0'
#689190000000
1!
b1001 %
1'
b1001 +
#689200000000
0!
0'
#689210000000
1!
b0 %
1'
b0 +
#689220000000
0!
0'
#689230000000
1!
1$
b1 %
1'
1*
b1 +
#689240000000
0!
0'
#689250000000
1!
b10 %
1'
b10 +
#689260000000
0!
0'
#689270000000
1!
b11 %
1'
b11 +
#689280000000
0!
0'
#689290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#689300000000
0!
0'
#689310000000
1!
b101 %
1'
b101 +
#689320000000
0!
0'
#689330000000
1!
0$
b110 %
1'
0*
b110 +
#689340000000
0!
0'
#689350000000
1!
b111 %
1'
b111 +
#689360000000
0!
0'
#689370000000
1!
b1000 %
1'
b1000 +
#689380000000
0!
0'
#689390000000
1!
b1001 %
1'
b1001 +
#689400000000
0!
0'
#689410000000
1!
b0 %
1'
b0 +
#689420000000
0!
0'
#689430000000
1!
1$
b1 %
1'
1*
b1 +
#689440000000
0!
0'
#689450000000
1!
b10 %
1'
b10 +
#689460000000
0!
0'
#689470000000
1!
b11 %
1'
b11 +
#689480000000
0!
0'
#689490000000
1!
b100 %
1'
b100 +
#689500000000
1"
1(
#689510000000
0!
0"
b100 &
0'
0(
b100 ,
#689520000000
1!
b101 %
1'
b101 +
#689530000000
0!
0'
#689540000000
1!
b110 %
1'
b110 +
#689550000000
0!
0'
#689560000000
1!
b111 %
1'
b111 +
#689570000000
0!
0'
#689580000000
1!
0$
b1000 %
1'
0*
b1000 +
#689590000000
0!
0'
#689600000000
1!
b1001 %
1'
b1001 +
#689610000000
0!
0'
#689620000000
1!
b0 %
1'
b0 +
#689630000000
0!
0'
#689640000000
1!
1$
b1 %
1'
1*
b1 +
#689650000000
0!
0'
#689660000000
1!
b10 %
1'
b10 +
#689670000000
0!
0'
#689680000000
1!
b11 %
1'
b11 +
#689690000000
0!
0'
#689700000000
1!
b100 %
1'
b100 +
#689710000000
0!
0'
#689720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#689730000000
0!
0'
#689740000000
1!
0$
b110 %
1'
0*
b110 +
#689750000000
0!
0'
#689760000000
1!
b111 %
1'
b111 +
#689770000000
0!
0'
#689780000000
1!
b1000 %
1'
b1000 +
#689790000000
0!
0'
#689800000000
1!
b1001 %
1'
b1001 +
#689810000000
0!
0'
#689820000000
1!
b0 %
1'
b0 +
#689830000000
0!
0'
#689840000000
1!
1$
b1 %
1'
1*
b1 +
#689850000000
0!
0'
#689860000000
1!
b10 %
1'
b10 +
#689870000000
0!
0'
#689880000000
1!
b11 %
1'
b11 +
#689890000000
0!
0'
#689900000000
1!
b100 %
1'
b100 +
#689910000000
0!
0'
#689920000000
1!
b101 %
1'
b101 +
#689930000000
1"
1(
#689940000000
0!
0"
b100 &
0'
0(
b100 ,
#689950000000
1!
b110 %
1'
b110 +
#689960000000
0!
0'
#689970000000
1!
b111 %
1'
b111 +
#689980000000
0!
0'
#689990000000
1!
0$
b1000 %
1'
0*
b1000 +
#690000000000
0!
0'
#690010000000
1!
b1001 %
1'
b1001 +
#690020000000
0!
0'
#690030000000
1!
b0 %
1'
b0 +
#690040000000
0!
0'
#690050000000
1!
1$
b1 %
1'
1*
b1 +
#690060000000
0!
0'
#690070000000
1!
b10 %
1'
b10 +
#690080000000
0!
0'
#690090000000
1!
b11 %
1'
b11 +
#690100000000
0!
0'
#690110000000
1!
b100 %
1'
b100 +
#690120000000
0!
0'
#690130000000
1!
b101 %
1'
b101 +
#690140000000
0!
0'
#690150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#690160000000
0!
0'
#690170000000
1!
b111 %
1'
b111 +
#690180000000
0!
0'
#690190000000
1!
b1000 %
1'
b1000 +
#690200000000
0!
0'
#690210000000
1!
b1001 %
1'
b1001 +
#690220000000
0!
0'
#690230000000
1!
b0 %
1'
b0 +
#690240000000
0!
0'
#690250000000
1!
1$
b1 %
1'
1*
b1 +
#690260000000
0!
0'
#690270000000
1!
b10 %
1'
b10 +
#690280000000
0!
0'
#690290000000
1!
b11 %
1'
b11 +
#690300000000
0!
0'
#690310000000
1!
b100 %
1'
b100 +
#690320000000
0!
0'
#690330000000
1!
b101 %
1'
b101 +
#690340000000
0!
0'
#690350000000
1!
0$
b110 %
1'
0*
b110 +
#690360000000
1"
1(
#690370000000
0!
0"
b100 &
0'
0(
b100 ,
#690380000000
1!
1$
b111 %
1'
1*
b111 +
#690390000000
0!
0'
#690400000000
1!
0$
b1000 %
1'
0*
b1000 +
#690410000000
0!
0'
#690420000000
1!
b1001 %
1'
b1001 +
#690430000000
0!
0'
#690440000000
1!
b0 %
1'
b0 +
#690450000000
0!
0'
#690460000000
1!
1$
b1 %
1'
1*
b1 +
#690470000000
0!
0'
#690480000000
1!
b10 %
1'
b10 +
#690490000000
0!
0'
#690500000000
1!
b11 %
1'
b11 +
#690510000000
0!
0'
#690520000000
1!
b100 %
1'
b100 +
#690530000000
0!
0'
#690540000000
1!
b101 %
1'
b101 +
#690550000000
0!
0'
#690560000000
1!
b110 %
1'
b110 +
#690570000000
0!
0'
#690580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#690590000000
0!
0'
#690600000000
1!
b1000 %
1'
b1000 +
#690610000000
0!
0'
#690620000000
1!
b1001 %
1'
b1001 +
#690630000000
0!
0'
#690640000000
1!
b0 %
1'
b0 +
#690650000000
0!
0'
#690660000000
1!
1$
b1 %
1'
1*
b1 +
#690670000000
0!
0'
#690680000000
1!
b10 %
1'
b10 +
#690690000000
0!
0'
#690700000000
1!
b11 %
1'
b11 +
#690710000000
0!
0'
#690720000000
1!
b100 %
1'
b100 +
#690730000000
0!
0'
#690740000000
1!
b101 %
1'
b101 +
#690750000000
0!
0'
#690760000000
1!
0$
b110 %
1'
0*
b110 +
#690770000000
0!
0'
#690780000000
1!
b111 %
1'
b111 +
#690790000000
1"
1(
#690800000000
0!
0"
b100 &
0'
0(
b100 ,
#690810000000
1!
b1000 %
1'
b1000 +
#690820000000
0!
0'
#690830000000
1!
b1001 %
1'
b1001 +
#690840000000
0!
0'
#690850000000
1!
b0 %
1'
b0 +
#690860000000
0!
0'
#690870000000
1!
1$
b1 %
1'
1*
b1 +
#690880000000
0!
0'
#690890000000
1!
b10 %
1'
b10 +
#690900000000
0!
0'
#690910000000
1!
b11 %
1'
b11 +
#690920000000
0!
0'
#690930000000
1!
b100 %
1'
b100 +
#690940000000
0!
0'
#690950000000
1!
b101 %
1'
b101 +
#690960000000
0!
0'
#690970000000
1!
b110 %
1'
b110 +
#690980000000
0!
0'
#690990000000
1!
b111 %
1'
b111 +
#691000000000
0!
0'
#691010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#691020000000
0!
0'
#691030000000
1!
b1001 %
1'
b1001 +
#691040000000
0!
0'
#691050000000
1!
b0 %
1'
b0 +
#691060000000
0!
0'
#691070000000
1!
1$
b1 %
1'
1*
b1 +
#691080000000
0!
0'
#691090000000
1!
b10 %
1'
b10 +
#691100000000
0!
0'
#691110000000
1!
b11 %
1'
b11 +
#691120000000
0!
0'
#691130000000
1!
b100 %
1'
b100 +
#691140000000
0!
0'
#691150000000
1!
b101 %
1'
b101 +
#691160000000
0!
0'
#691170000000
1!
0$
b110 %
1'
0*
b110 +
#691180000000
0!
0'
#691190000000
1!
b111 %
1'
b111 +
#691200000000
0!
0'
#691210000000
1!
b1000 %
1'
b1000 +
#691220000000
1"
1(
#691230000000
0!
0"
b100 &
0'
0(
b100 ,
#691240000000
1!
b1001 %
1'
b1001 +
#691250000000
0!
0'
#691260000000
1!
b0 %
1'
b0 +
#691270000000
0!
0'
#691280000000
1!
1$
b1 %
1'
1*
b1 +
#691290000000
0!
0'
#691300000000
1!
b10 %
1'
b10 +
#691310000000
0!
0'
#691320000000
1!
b11 %
1'
b11 +
#691330000000
0!
0'
#691340000000
1!
b100 %
1'
b100 +
#691350000000
0!
0'
#691360000000
1!
b101 %
1'
b101 +
#691370000000
0!
0'
#691380000000
1!
b110 %
1'
b110 +
#691390000000
0!
0'
#691400000000
1!
b111 %
1'
b111 +
#691410000000
0!
0'
#691420000000
1!
0$
b1000 %
1'
0*
b1000 +
#691430000000
0!
0'
#691440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#691450000000
0!
0'
#691460000000
1!
b0 %
1'
b0 +
#691470000000
0!
0'
#691480000000
1!
1$
b1 %
1'
1*
b1 +
#691490000000
0!
0'
#691500000000
1!
b10 %
1'
b10 +
#691510000000
0!
0'
#691520000000
1!
b11 %
1'
b11 +
#691530000000
0!
0'
#691540000000
1!
b100 %
1'
b100 +
#691550000000
0!
0'
#691560000000
1!
b101 %
1'
b101 +
#691570000000
0!
0'
#691580000000
1!
0$
b110 %
1'
0*
b110 +
#691590000000
0!
0'
#691600000000
1!
b111 %
1'
b111 +
#691610000000
0!
0'
#691620000000
1!
b1000 %
1'
b1000 +
#691630000000
0!
0'
#691640000000
1!
b1001 %
1'
b1001 +
#691650000000
1"
1(
#691660000000
0!
0"
b100 &
0'
0(
b100 ,
#691670000000
1!
b0 %
1'
b0 +
#691680000000
0!
0'
#691690000000
1!
1$
b1 %
1'
1*
b1 +
#691700000000
0!
0'
#691710000000
1!
b10 %
1'
b10 +
#691720000000
0!
0'
#691730000000
1!
b11 %
1'
b11 +
#691740000000
0!
0'
#691750000000
1!
b100 %
1'
b100 +
#691760000000
0!
0'
#691770000000
1!
b101 %
1'
b101 +
#691780000000
0!
0'
#691790000000
1!
b110 %
1'
b110 +
#691800000000
0!
0'
#691810000000
1!
b111 %
1'
b111 +
#691820000000
0!
0'
#691830000000
1!
0$
b1000 %
1'
0*
b1000 +
#691840000000
0!
0'
#691850000000
1!
b1001 %
1'
b1001 +
#691860000000
0!
0'
#691870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#691880000000
0!
0'
#691890000000
1!
1$
b1 %
1'
1*
b1 +
#691900000000
0!
0'
#691910000000
1!
b10 %
1'
b10 +
#691920000000
0!
0'
#691930000000
1!
b11 %
1'
b11 +
#691940000000
0!
0'
#691950000000
1!
b100 %
1'
b100 +
#691960000000
0!
0'
#691970000000
1!
b101 %
1'
b101 +
#691980000000
0!
0'
#691990000000
1!
0$
b110 %
1'
0*
b110 +
#692000000000
0!
0'
#692010000000
1!
b111 %
1'
b111 +
#692020000000
0!
0'
#692030000000
1!
b1000 %
1'
b1000 +
#692040000000
0!
0'
#692050000000
1!
b1001 %
1'
b1001 +
#692060000000
0!
0'
#692070000000
1!
b0 %
1'
b0 +
#692080000000
1"
1(
#692090000000
0!
0"
b100 &
0'
0(
b100 ,
#692100000000
1!
1$
b1 %
1'
1*
b1 +
#692110000000
0!
0'
#692120000000
1!
b10 %
1'
b10 +
#692130000000
0!
0'
#692140000000
1!
b11 %
1'
b11 +
#692150000000
0!
0'
#692160000000
1!
b100 %
1'
b100 +
#692170000000
0!
0'
#692180000000
1!
b101 %
1'
b101 +
#692190000000
0!
0'
#692200000000
1!
b110 %
1'
b110 +
#692210000000
0!
0'
#692220000000
1!
b111 %
1'
b111 +
#692230000000
0!
0'
#692240000000
1!
0$
b1000 %
1'
0*
b1000 +
#692250000000
0!
0'
#692260000000
1!
b1001 %
1'
b1001 +
#692270000000
0!
0'
#692280000000
1!
b0 %
1'
b0 +
#692290000000
0!
0'
#692300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#692310000000
0!
0'
#692320000000
1!
b10 %
1'
b10 +
#692330000000
0!
0'
#692340000000
1!
b11 %
1'
b11 +
#692350000000
0!
0'
#692360000000
1!
b100 %
1'
b100 +
#692370000000
0!
0'
#692380000000
1!
b101 %
1'
b101 +
#692390000000
0!
0'
#692400000000
1!
0$
b110 %
1'
0*
b110 +
#692410000000
0!
0'
#692420000000
1!
b111 %
1'
b111 +
#692430000000
0!
0'
#692440000000
1!
b1000 %
1'
b1000 +
#692450000000
0!
0'
#692460000000
1!
b1001 %
1'
b1001 +
#692470000000
0!
0'
#692480000000
1!
b0 %
1'
b0 +
#692490000000
0!
0'
#692500000000
1!
1$
b1 %
1'
1*
b1 +
#692510000000
1"
1(
#692520000000
0!
0"
b100 &
0'
0(
b100 ,
#692530000000
1!
b10 %
1'
b10 +
#692540000000
0!
0'
#692550000000
1!
b11 %
1'
b11 +
#692560000000
0!
0'
#692570000000
1!
b100 %
1'
b100 +
#692580000000
0!
0'
#692590000000
1!
b101 %
1'
b101 +
#692600000000
0!
0'
#692610000000
1!
b110 %
1'
b110 +
#692620000000
0!
0'
#692630000000
1!
b111 %
1'
b111 +
#692640000000
0!
0'
#692650000000
1!
0$
b1000 %
1'
0*
b1000 +
#692660000000
0!
0'
#692670000000
1!
b1001 %
1'
b1001 +
#692680000000
0!
0'
#692690000000
1!
b0 %
1'
b0 +
#692700000000
0!
0'
#692710000000
1!
1$
b1 %
1'
1*
b1 +
#692720000000
0!
0'
#692730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#692740000000
0!
0'
#692750000000
1!
b11 %
1'
b11 +
#692760000000
0!
0'
#692770000000
1!
b100 %
1'
b100 +
#692780000000
0!
0'
#692790000000
1!
b101 %
1'
b101 +
#692800000000
0!
0'
#692810000000
1!
0$
b110 %
1'
0*
b110 +
#692820000000
0!
0'
#692830000000
1!
b111 %
1'
b111 +
#692840000000
0!
0'
#692850000000
1!
b1000 %
1'
b1000 +
#692860000000
0!
0'
#692870000000
1!
b1001 %
1'
b1001 +
#692880000000
0!
0'
#692890000000
1!
b0 %
1'
b0 +
#692900000000
0!
0'
#692910000000
1!
1$
b1 %
1'
1*
b1 +
#692920000000
0!
0'
#692930000000
1!
b10 %
1'
b10 +
#692940000000
1"
1(
#692950000000
0!
0"
b100 &
0'
0(
b100 ,
#692960000000
1!
b11 %
1'
b11 +
#692970000000
0!
0'
#692980000000
1!
b100 %
1'
b100 +
#692990000000
0!
0'
#693000000000
1!
b101 %
1'
b101 +
#693010000000
0!
0'
#693020000000
1!
b110 %
1'
b110 +
#693030000000
0!
0'
#693040000000
1!
b111 %
1'
b111 +
#693050000000
0!
0'
#693060000000
1!
0$
b1000 %
1'
0*
b1000 +
#693070000000
0!
0'
#693080000000
1!
b1001 %
1'
b1001 +
#693090000000
0!
0'
#693100000000
1!
b0 %
1'
b0 +
#693110000000
0!
0'
#693120000000
1!
1$
b1 %
1'
1*
b1 +
#693130000000
0!
0'
#693140000000
1!
b10 %
1'
b10 +
#693150000000
0!
0'
#693160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#693170000000
0!
0'
#693180000000
1!
b100 %
1'
b100 +
#693190000000
0!
0'
#693200000000
1!
b101 %
1'
b101 +
#693210000000
0!
0'
#693220000000
1!
0$
b110 %
1'
0*
b110 +
#693230000000
0!
0'
#693240000000
1!
b111 %
1'
b111 +
#693250000000
0!
0'
#693260000000
1!
b1000 %
1'
b1000 +
#693270000000
0!
0'
#693280000000
1!
b1001 %
1'
b1001 +
#693290000000
0!
0'
#693300000000
1!
b0 %
1'
b0 +
#693310000000
0!
0'
#693320000000
1!
1$
b1 %
1'
1*
b1 +
#693330000000
0!
0'
#693340000000
1!
b10 %
1'
b10 +
#693350000000
0!
0'
#693360000000
1!
b11 %
1'
b11 +
#693370000000
1"
1(
#693380000000
0!
0"
b100 &
0'
0(
b100 ,
#693390000000
1!
b100 %
1'
b100 +
#693400000000
0!
0'
#693410000000
1!
b101 %
1'
b101 +
#693420000000
0!
0'
#693430000000
1!
b110 %
1'
b110 +
#693440000000
0!
0'
#693450000000
1!
b111 %
1'
b111 +
#693460000000
0!
0'
#693470000000
1!
0$
b1000 %
1'
0*
b1000 +
#693480000000
0!
0'
#693490000000
1!
b1001 %
1'
b1001 +
#693500000000
0!
0'
#693510000000
1!
b0 %
1'
b0 +
#693520000000
0!
0'
#693530000000
1!
1$
b1 %
1'
1*
b1 +
#693540000000
0!
0'
#693550000000
1!
b10 %
1'
b10 +
#693560000000
0!
0'
#693570000000
1!
b11 %
1'
b11 +
#693580000000
0!
0'
#693590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#693600000000
0!
0'
#693610000000
1!
b101 %
1'
b101 +
#693620000000
0!
0'
#693630000000
1!
0$
b110 %
1'
0*
b110 +
#693640000000
0!
0'
#693650000000
1!
b111 %
1'
b111 +
#693660000000
0!
0'
#693670000000
1!
b1000 %
1'
b1000 +
#693680000000
0!
0'
#693690000000
1!
b1001 %
1'
b1001 +
#693700000000
0!
0'
#693710000000
1!
b0 %
1'
b0 +
#693720000000
0!
0'
#693730000000
1!
1$
b1 %
1'
1*
b1 +
#693740000000
0!
0'
#693750000000
1!
b10 %
1'
b10 +
#693760000000
0!
0'
#693770000000
1!
b11 %
1'
b11 +
#693780000000
0!
0'
#693790000000
1!
b100 %
1'
b100 +
#693800000000
1"
1(
#693810000000
0!
0"
b100 &
0'
0(
b100 ,
#693820000000
1!
b101 %
1'
b101 +
#693830000000
0!
0'
#693840000000
1!
b110 %
1'
b110 +
#693850000000
0!
0'
#693860000000
1!
b111 %
1'
b111 +
#693870000000
0!
0'
#693880000000
1!
0$
b1000 %
1'
0*
b1000 +
#693890000000
0!
0'
#693900000000
1!
b1001 %
1'
b1001 +
#693910000000
0!
0'
#693920000000
1!
b0 %
1'
b0 +
#693930000000
0!
0'
#693940000000
1!
1$
b1 %
1'
1*
b1 +
#693950000000
0!
0'
#693960000000
1!
b10 %
1'
b10 +
#693970000000
0!
0'
#693980000000
1!
b11 %
1'
b11 +
#693990000000
0!
0'
#694000000000
1!
b100 %
1'
b100 +
#694010000000
0!
0'
#694020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#694030000000
0!
0'
#694040000000
1!
0$
b110 %
1'
0*
b110 +
#694050000000
0!
0'
#694060000000
1!
b111 %
1'
b111 +
#694070000000
0!
0'
#694080000000
1!
b1000 %
1'
b1000 +
#694090000000
0!
0'
#694100000000
1!
b1001 %
1'
b1001 +
#694110000000
0!
0'
#694120000000
1!
b0 %
1'
b0 +
#694130000000
0!
0'
#694140000000
1!
1$
b1 %
1'
1*
b1 +
#694150000000
0!
0'
#694160000000
1!
b10 %
1'
b10 +
#694170000000
0!
0'
#694180000000
1!
b11 %
1'
b11 +
#694190000000
0!
0'
#694200000000
1!
b100 %
1'
b100 +
#694210000000
0!
0'
#694220000000
1!
b101 %
1'
b101 +
#694230000000
1"
1(
#694240000000
0!
0"
b100 &
0'
0(
b100 ,
#694250000000
1!
b110 %
1'
b110 +
#694260000000
0!
0'
#694270000000
1!
b111 %
1'
b111 +
#694280000000
0!
0'
#694290000000
1!
0$
b1000 %
1'
0*
b1000 +
#694300000000
0!
0'
#694310000000
1!
b1001 %
1'
b1001 +
#694320000000
0!
0'
#694330000000
1!
b0 %
1'
b0 +
#694340000000
0!
0'
#694350000000
1!
1$
b1 %
1'
1*
b1 +
#694360000000
0!
0'
#694370000000
1!
b10 %
1'
b10 +
#694380000000
0!
0'
#694390000000
1!
b11 %
1'
b11 +
#694400000000
0!
0'
#694410000000
1!
b100 %
1'
b100 +
#694420000000
0!
0'
#694430000000
1!
b101 %
1'
b101 +
#694440000000
0!
0'
#694450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#694460000000
0!
0'
#694470000000
1!
b111 %
1'
b111 +
#694480000000
0!
0'
#694490000000
1!
b1000 %
1'
b1000 +
#694500000000
0!
0'
#694510000000
1!
b1001 %
1'
b1001 +
#694520000000
0!
0'
#694530000000
1!
b0 %
1'
b0 +
#694540000000
0!
0'
#694550000000
1!
1$
b1 %
1'
1*
b1 +
#694560000000
0!
0'
#694570000000
1!
b10 %
1'
b10 +
#694580000000
0!
0'
#694590000000
1!
b11 %
1'
b11 +
#694600000000
0!
0'
#694610000000
1!
b100 %
1'
b100 +
#694620000000
0!
0'
#694630000000
1!
b101 %
1'
b101 +
#694640000000
0!
0'
#694650000000
1!
0$
b110 %
1'
0*
b110 +
#694660000000
1"
1(
#694670000000
0!
0"
b100 &
0'
0(
b100 ,
#694680000000
1!
1$
b111 %
1'
1*
b111 +
#694690000000
0!
0'
#694700000000
1!
0$
b1000 %
1'
0*
b1000 +
#694710000000
0!
0'
#694720000000
1!
b1001 %
1'
b1001 +
#694730000000
0!
0'
#694740000000
1!
b0 %
1'
b0 +
#694750000000
0!
0'
#694760000000
1!
1$
b1 %
1'
1*
b1 +
#694770000000
0!
0'
#694780000000
1!
b10 %
1'
b10 +
#694790000000
0!
0'
#694800000000
1!
b11 %
1'
b11 +
#694810000000
0!
0'
#694820000000
1!
b100 %
1'
b100 +
#694830000000
0!
0'
#694840000000
1!
b101 %
1'
b101 +
#694850000000
0!
0'
#694860000000
1!
b110 %
1'
b110 +
#694870000000
0!
0'
#694880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#694890000000
0!
0'
#694900000000
1!
b1000 %
1'
b1000 +
#694910000000
0!
0'
#694920000000
1!
b1001 %
1'
b1001 +
#694930000000
0!
0'
#694940000000
1!
b0 %
1'
b0 +
#694950000000
0!
0'
#694960000000
1!
1$
b1 %
1'
1*
b1 +
#694970000000
0!
0'
#694980000000
1!
b10 %
1'
b10 +
#694990000000
0!
0'
#695000000000
1!
b11 %
1'
b11 +
#695010000000
0!
0'
#695020000000
1!
b100 %
1'
b100 +
#695030000000
0!
0'
#695040000000
1!
b101 %
1'
b101 +
#695050000000
0!
0'
#695060000000
1!
0$
b110 %
1'
0*
b110 +
#695070000000
0!
0'
#695080000000
1!
b111 %
1'
b111 +
#695090000000
1"
1(
#695100000000
0!
0"
b100 &
0'
0(
b100 ,
#695110000000
1!
b1000 %
1'
b1000 +
#695120000000
0!
0'
#695130000000
1!
b1001 %
1'
b1001 +
#695140000000
0!
0'
#695150000000
1!
b0 %
1'
b0 +
#695160000000
0!
0'
#695170000000
1!
1$
b1 %
1'
1*
b1 +
#695180000000
0!
0'
#695190000000
1!
b10 %
1'
b10 +
#695200000000
0!
0'
#695210000000
1!
b11 %
1'
b11 +
#695220000000
0!
0'
#695230000000
1!
b100 %
1'
b100 +
#695240000000
0!
0'
#695250000000
1!
b101 %
1'
b101 +
#695260000000
0!
0'
#695270000000
1!
b110 %
1'
b110 +
#695280000000
0!
0'
#695290000000
1!
b111 %
1'
b111 +
#695300000000
0!
0'
#695310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#695320000000
0!
0'
#695330000000
1!
b1001 %
1'
b1001 +
#695340000000
0!
0'
#695350000000
1!
b0 %
1'
b0 +
#695360000000
0!
0'
#695370000000
1!
1$
b1 %
1'
1*
b1 +
#695380000000
0!
0'
#695390000000
1!
b10 %
1'
b10 +
#695400000000
0!
0'
#695410000000
1!
b11 %
1'
b11 +
#695420000000
0!
0'
#695430000000
1!
b100 %
1'
b100 +
#695440000000
0!
0'
#695450000000
1!
b101 %
1'
b101 +
#695460000000
0!
0'
#695470000000
1!
0$
b110 %
1'
0*
b110 +
#695480000000
0!
0'
#695490000000
1!
b111 %
1'
b111 +
#695500000000
0!
0'
#695510000000
1!
b1000 %
1'
b1000 +
#695520000000
1"
1(
#695530000000
0!
0"
b100 &
0'
0(
b100 ,
#695540000000
1!
b1001 %
1'
b1001 +
#695550000000
0!
0'
#695560000000
1!
b0 %
1'
b0 +
#695570000000
0!
0'
#695580000000
1!
1$
b1 %
1'
1*
b1 +
#695590000000
0!
0'
#695600000000
1!
b10 %
1'
b10 +
#695610000000
0!
0'
#695620000000
1!
b11 %
1'
b11 +
#695630000000
0!
0'
#695640000000
1!
b100 %
1'
b100 +
#695650000000
0!
0'
#695660000000
1!
b101 %
1'
b101 +
#695670000000
0!
0'
#695680000000
1!
b110 %
1'
b110 +
#695690000000
0!
0'
#695700000000
1!
b111 %
1'
b111 +
#695710000000
0!
0'
#695720000000
1!
0$
b1000 %
1'
0*
b1000 +
#695730000000
0!
0'
#695740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#695750000000
0!
0'
#695760000000
1!
b0 %
1'
b0 +
#695770000000
0!
0'
#695780000000
1!
1$
b1 %
1'
1*
b1 +
#695790000000
0!
0'
#695800000000
1!
b10 %
1'
b10 +
#695810000000
0!
0'
#695820000000
1!
b11 %
1'
b11 +
#695830000000
0!
0'
#695840000000
1!
b100 %
1'
b100 +
#695850000000
0!
0'
#695860000000
1!
b101 %
1'
b101 +
#695870000000
0!
0'
#695880000000
1!
0$
b110 %
1'
0*
b110 +
#695890000000
0!
0'
#695900000000
1!
b111 %
1'
b111 +
#695910000000
0!
0'
#695920000000
1!
b1000 %
1'
b1000 +
#695930000000
0!
0'
#695940000000
1!
b1001 %
1'
b1001 +
#695950000000
1"
1(
#695960000000
0!
0"
b100 &
0'
0(
b100 ,
#695970000000
1!
b0 %
1'
b0 +
#695980000000
0!
0'
#695990000000
1!
1$
b1 %
1'
1*
b1 +
#696000000000
0!
0'
#696010000000
1!
b10 %
1'
b10 +
#696020000000
0!
0'
#696030000000
1!
b11 %
1'
b11 +
#696040000000
0!
0'
#696050000000
1!
b100 %
1'
b100 +
#696060000000
0!
0'
#696070000000
1!
b101 %
1'
b101 +
#696080000000
0!
0'
#696090000000
1!
b110 %
1'
b110 +
#696100000000
0!
0'
#696110000000
1!
b111 %
1'
b111 +
#696120000000
0!
0'
#696130000000
1!
0$
b1000 %
1'
0*
b1000 +
#696140000000
0!
0'
#696150000000
1!
b1001 %
1'
b1001 +
#696160000000
0!
0'
#696170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#696180000000
0!
0'
#696190000000
1!
1$
b1 %
1'
1*
b1 +
#696200000000
0!
0'
#696210000000
1!
b10 %
1'
b10 +
#696220000000
0!
0'
#696230000000
1!
b11 %
1'
b11 +
#696240000000
0!
0'
#696250000000
1!
b100 %
1'
b100 +
#696260000000
0!
0'
#696270000000
1!
b101 %
1'
b101 +
#696280000000
0!
0'
#696290000000
1!
0$
b110 %
1'
0*
b110 +
#696300000000
0!
0'
#696310000000
1!
b111 %
1'
b111 +
#696320000000
0!
0'
#696330000000
1!
b1000 %
1'
b1000 +
#696340000000
0!
0'
#696350000000
1!
b1001 %
1'
b1001 +
#696360000000
0!
0'
#696370000000
1!
b0 %
1'
b0 +
#696380000000
1"
1(
#696390000000
0!
0"
b100 &
0'
0(
b100 ,
#696400000000
1!
1$
b1 %
1'
1*
b1 +
#696410000000
0!
0'
#696420000000
1!
b10 %
1'
b10 +
#696430000000
0!
0'
#696440000000
1!
b11 %
1'
b11 +
#696450000000
0!
0'
#696460000000
1!
b100 %
1'
b100 +
#696470000000
0!
0'
#696480000000
1!
b101 %
1'
b101 +
#696490000000
0!
0'
#696500000000
1!
b110 %
1'
b110 +
#696510000000
0!
0'
#696520000000
1!
b111 %
1'
b111 +
#696530000000
0!
0'
#696540000000
1!
0$
b1000 %
1'
0*
b1000 +
#696550000000
0!
0'
#696560000000
1!
b1001 %
1'
b1001 +
#696570000000
0!
0'
#696580000000
1!
b0 %
1'
b0 +
#696590000000
0!
0'
#696600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#696610000000
0!
0'
#696620000000
1!
b10 %
1'
b10 +
#696630000000
0!
0'
#696640000000
1!
b11 %
1'
b11 +
#696650000000
0!
0'
#696660000000
1!
b100 %
1'
b100 +
#696670000000
0!
0'
#696680000000
1!
b101 %
1'
b101 +
#696690000000
0!
0'
#696700000000
1!
0$
b110 %
1'
0*
b110 +
#696710000000
0!
0'
#696720000000
1!
b111 %
1'
b111 +
#696730000000
0!
0'
#696740000000
1!
b1000 %
1'
b1000 +
#696750000000
0!
0'
#696760000000
1!
b1001 %
1'
b1001 +
#696770000000
0!
0'
#696780000000
1!
b0 %
1'
b0 +
#696790000000
0!
0'
#696800000000
1!
1$
b1 %
1'
1*
b1 +
#696810000000
1"
1(
#696820000000
0!
0"
b100 &
0'
0(
b100 ,
#696830000000
1!
b10 %
1'
b10 +
#696840000000
0!
0'
#696850000000
1!
b11 %
1'
b11 +
#696860000000
0!
0'
#696870000000
1!
b100 %
1'
b100 +
#696880000000
0!
0'
#696890000000
1!
b101 %
1'
b101 +
#696900000000
0!
0'
#696910000000
1!
b110 %
1'
b110 +
#696920000000
0!
0'
#696930000000
1!
b111 %
1'
b111 +
#696940000000
0!
0'
#696950000000
1!
0$
b1000 %
1'
0*
b1000 +
#696960000000
0!
0'
#696970000000
1!
b1001 %
1'
b1001 +
#696980000000
0!
0'
#696990000000
1!
b0 %
1'
b0 +
#697000000000
0!
0'
#697010000000
1!
1$
b1 %
1'
1*
b1 +
#697020000000
0!
0'
#697030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#697040000000
0!
0'
#697050000000
1!
b11 %
1'
b11 +
#697060000000
0!
0'
#697070000000
1!
b100 %
1'
b100 +
#697080000000
0!
0'
#697090000000
1!
b101 %
1'
b101 +
#697100000000
0!
0'
#697110000000
1!
0$
b110 %
1'
0*
b110 +
#697120000000
0!
0'
#697130000000
1!
b111 %
1'
b111 +
#697140000000
0!
0'
#697150000000
1!
b1000 %
1'
b1000 +
#697160000000
0!
0'
#697170000000
1!
b1001 %
1'
b1001 +
#697180000000
0!
0'
#697190000000
1!
b0 %
1'
b0 +
#697200000000
0!
0'
#697210000000
1!
1$
b1 %
1'
1*
b1 +
#697220000000
0!
0'
#697230000000
1!
b10 %
1'
b10 +
#697240000000
1"
1(
#697250000000
0!
0"
b100 &
0'
0(
b100 ,
#697260000000
1!
b11 %
1'
b11 +
#697270000000
0!
0'
#697280000000
1!
b100 %
1'
b100 +
#697290000000
0!
0'
#697300000000
1!
b101 %
1'
b101 +
#697310000000
0!
0'
#697320000000
1!
b110 %
1'
b110 +
#697330000000
0!
0'
#697340000000
1!
b111 %
1'
b111 +
#697350000000
0!
0'
#697360000000
1!
0$
b1000 %
1'
0*
b1000 +
#697370000000
0!
0'
#697380000000
1!
b1001 %
1'
b1001 +
#697390000000
0!
0'
#697400000000
1!
b0 %
1'
b0 +
#697410000000
0!
0'
#697420000000
1!
1$
b1 %
1'
1*
b1 +
#697430000000
0!
0'
#697440000000
1!
b10 %
1'
b10 +
#697450000000
0!
0'
#697460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#697470000000
0!
0'
#697480000000
1!
b100 %
1'
b100 +
#697490000000
0!
0'
#697500000000
1!
b101 %
1'
b101 +
#697510000000
0!
0'
#697520000000
1!
0$
b110 %
1'
0*
b110 +
#697530000000
0!
0'
#697540000000
1!
b111 %
1'
b111 +
#697550000000
0!
0'
#697560000000
1!
b1000 %
1'
b1000 +
#697570000000
0!
0'
#697580000000
1!
b1001 %
1'
b1001 +
#697590000000
0!
0'
#697600000000
1!
b0 %
1'
b0 +
#697610000000
0!
0'
#697620000000
1!
1$
b1 %
1'
1*
b1 +
#697630000000
0!
0'
#697640000000
1!
b10 %
1'
b10 +
#697650000000
0!
0'
#697660000000
1!
b11 %
1'
b11 +
#697670000000
1"
1(
#697680000000
0!
0"
b100 &
0'
0(
b100 ,
#697690000000
1!
b100 %
1'
b100 +
#697700000000
0!
0'
#697710000000
1!
b101 %
1'
b101 +
#697720000000
0!
0'
#697730000000
1!
b110 %
1'
b110 +
#697740000000
0!
0'
#697750000000
1!
b111 %
1'
b111 +
#697760000000
0!
0'
#697770000000
1!
0$
b1000 %
1'
0*
b1000 +
#697780000000
0!
0'
#697790000000
1!
b1001 %
1'
b1001 +
#697800000000
0!
0'
#697810000000
1!
b0 %
1'
b0 +
#697820000000
0!
0'
#697830000000
1!
1$
b1 %
1'
1*
b1 +
#697840000000
0!
0'
#697850000000
1!
b10 %
1'
b10 +
#697860000000
0!
0'
#697870000000
1!
b11 %
1'
b11 +
#697880000000
0!
0'
#697890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#697900000000
0!
0'
#697910000000
1!
b101 %
1'
b101 +
#697920000000
0!
0'
#697930000000
1!
0$
b110 %
1'
0*
b110 +
#697940000000
0!
0'
#697950000000
1!
b111 %
1'
b111 +
#697960000000
0!
0'
#697970000000
1!
b1000 %
1'
b1000 +
#697980000000
0!
0'
#697990000000
1!
b1001 %
1'
b1001 +
#698000000000
0!
0'
#698010000000
1!
b0 %
1'
b0 +
#698020000000
0!
0'
#698030000000
1!
1$
b1 %
1'
1*
b1 +
#698040000000
0!
0'
#698050000000
1!
b10 %
1'
b10 +
#698060000000
0!
0'
#698070000000
1!
b11 %
1'
b11 +
#698080000000
0!
0'
#698090000000
1!
b100 %
1'
b100 +
#698100000000
1"
1(
#698110000000
0!
0"
b100 &
0'
0(
b100 ,
#698120000000
1!
b101 %
1'
b101 +
#698130000000
0!
0'
#698140000000
1!
b110 %
1'
b110 +
#698150000000
0!
0'
#698160000000
1!
b111 %
1'
b111 +
#698170000000
0!
0'
#698180000000
1!
0$
b1000 %
1'
0*
b1000 +
#698190000000
0!
0'
#698200000000
1!
b1001 %
1'
b1001 +
#698210000000
0!
0'
#698220000000
1!
b0 %
1'
b0 +
#698230000000
0!
0'
#698240000000
1!
1$
b1 %
1'
1*
b1 +
#698250000000
0!
0'
#698260000000
1!
b10 %
1'
b10 +
#698270000000
0!
0'
#698280000000
1!
b11 %
1'
b11 +
#698290000000
0!
0'
#698300000000
1!
b100 %
1'
b100 +
#698310000000
0!
0'
#698320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#698330000000
0!
0'
#698340000000
1!
0$
b110 %
1'
0*
b110 +
#698350000000
0!
0'
#698360000000
1!
b111 %
1'
b111 +
#698370000000
0!
0'
#698380000000
1!
b1000 %
1'
b1000 +
#698390000000
0!
0'
#698400000000
1!
b1001 %
1'
b1001 +
#698410000000
0!
0'
#698420000000
1!
b0 %
1'
b0 +
#698430000000
0!
0'
#698440000000
1!
1$
b1 %
1'
1*
b1 +
#698450000000
0!
0'
#698460000000
1!
b10 %
1'
b10 +
#698470000000
0!
0'
#698480000000
1!
b11 %
1'
b11 +
#698490000000
0!
0'
#698500000000
1!
b100 %
1'
b100 +
#698510000000
0!
0'
#698520000000
1!
b101 %
1'
b101 +
#698530000000
1"
1(
#698540000000
0!
0"
b100 &
0'
0(
b100 ,
#698550000000
1!
b110 %
1'
b110 +
#698560000000
0!
0'
#698570000000
1!
b111 %
1'
b111 +
#698580000000
0!
0'
#698590000000
1!
0$
b1000 %
1'
0*
b1000 +
#698600000000
0!
0'
#698610000000
1!
b1001 %
1'
b1001 +
#698620000000
0!
0'
#698630000000
1!
b0 %
1'
b0 +
#698640000000
0!
0'
#698650000000
1!
1$
b1 %
1'
1*
b1 +
#698660000000
0!
0'
#698670000000
1!
b10 %
1'
b10 +
#698680000000
0!
0'
#698690000000
1!
b11 %
1'
b11 +
#698700000000
0!
0'
#698710000000
1!
b100 %
1'
b100 +
#698720000000
0!
0'
#698730000000
1!
b101 %
1'
b101 +
#698740000000
0!
0'
#698750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#698760000000
0!
0'
#698770000000
1!
b111 %
1'
b111 +
#698780000000
0!
0'
#698790000000
1!
b1000 %
1'
b1000 +
#698800000000
0!
0'
#698810000000
1!
b1001 %
1'
b1001 +
#698820000000
0!
0'
#698830000000
1!
b0 %
1'
b0 +
#698840000000
0!
0'
#698850000000
1!
1$
b1 %
1'
1*
b1 +
#698860000000
0!
0'
#698870000000
1!
b10 %
1'
b10 +
#698880000000
0!
0'
#698890000000
1!
b11 %
1'
b11 +
#698900000000
0!
0'
#698910000000
1!
b100 %
1'
b100 +
#698920000000
0!
0'
#698930000000
1!
b101 %
1'
b101 +
#698940000000
0!
0'
#698950000000
1!
0$
b110 %
1'
0*
b110 +
#698960000000
1"
1(
#698970000000
0!
0"
b100 &
0'
0(
b100 ,
#698980000000
1!
1$
b111 %
1'
1*
b111 +
#698990000000
0!
0'
#699000000000
1!
0$
b1000 %
1'
0*
b1000 +
#699010000000
0!
0'
#699020000000
1!
b1001 %
1'
b1001 +
#699030000000
0!
0'
#699040000000
1!
b0 %
1'
b0 +
#699050000000
0!
0'
#699060000000
1!
1$
b1 %
1'
1*
b1 +
#699070000000
0!
0'
#699080000000
1!
b10 %
1'
b10 +
#699090000000
0!
0'
#699100000000
1!
b11 %
1'
b11 +
#699110000000
0!
0'
#699120000000
1!
b100 %
1'
b100 +
#699130000000
0!
0'
#699140000000
1!
b101 %
1'
b101 +
#699150000000
0!
0'
#699160000000
1!
b110 %
1'
b110 +
#699170000000
0!
0'
#699180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#699190000000
0!
0'
#699200000000
1!
b1000 %
1'
b1000 +
#699210000000
0!
0'
#699220000000
1!
b1001 %
1'
b1001 +
#699230000000
0!
0'
#699240000000
1!
b0 %
1'
b0 +
#699250000000
0!
0'
#699260000000
1!
1$
b1 %
1'
1*
b1 +
#699270000000
0!
0'
#699280000000
1!
b10 %
1'
b10 +
#699290000000
0!
0'
#699300000000
1!
b11 %
1'
b11 +
#699310000000
0!
0'
#699320000000
1!
b100 %
1'
b100 +
#699330000000
0!
0'
#699340000000
1!
b101 %
1'
b101 +
#699350000000
0!
0'
#699360000000
1!
0$
b110 %
1'
0*
b110 +
#699370000000
0!
0'
#699380000000
1!
b111 %
1'
b111 +
#699390000000
1"
1(
#699400000000
0!
0"
b100 &
0'
0(
b100 ,
#699410000000
1!
b1000 %
1'
b1000 +
#699420000000
0!
0'
#699430000000
1!
b1001 %
1'
b1001 +
#699440000000
0!
0'
#699450000000
1!
b0 %
1'
b0 +
#699460000000
0!
0'
#699470000000
1!
1$
b1 %
1'
1*
b1 +
#699480000000
0!
0'
#699490000000
1!
b10 %
1'
b10 +
#699500000000
0!
0'
#699510000000
1!
b11 %
1'
b11 +
#699520000000
0!
0'
#699530000000
1!
b100 %
1'
b100 +
#699540000000
0!
0'
#699550000000
1!
b101 %
1'
b101 +
#699560000000
0!
0'
#699570000000
1!
b110 %
1'
b110 +
#699580000000
0!
0'
#699590000000
1!
b111 %
1'
b111 +
#699600000000
0!
0'
#699610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#699620000000
0!
0'
#699630000000
1!
b1001 %
1'
b1001 +
#699640000000
0!
0'
#699650000000
1!
b0 %
1'
b0 +
#699660000000
0!
0'
#699670000000
1!
1$
b1 %
1'
1*
b1 +
#699680000000
0!
0'
#699690000000
1!
b10 %
1'
b10 +
#699700000000
0!
0'
#699710000000
1!
b11 %
1'
b11 +
#699720000000
0!
0'
#699730000000
1!
b100 %
1'
b100 +
#699740000000
0!
0'
#699750000000
1!
b101 %
1'
b101 +
#699760000000
0!
0'
#699770000000
1!
0$
b110 %
1'
0*
b110 +
#699780000000
0!
0'
#699790000000
1!
b111 %
1'
b111 +
#699800000000
0!
0'
#699810000000
1!
b1000 %
1'
b1000 +
#699820000000
1"
1(
#699830000000
0!
0"
b100 &
0'
0(
b100 ,
#699840000000
1!
b1001 %
1'
b1001 +
#699850000000
0!
0'
#699860000000
1!
b0 %
1'
b0 +
#699870000000
0!
0'
#699880000000
1!
1$
b1 %
1'
1*
b1 +
#699890000000
0!
0'
#699900000000
1!
b10 %
1'
b10 +
#699910000000
0!
0'
#699920000000
1!
b11 %
1'
b11 +
#699930000000
0!
0'
#699940000000
1!
b100 %
1'
b100 +
#699950000000
0!
0'
#699960000000
1!
b101 %
1'
b101 +
#699970000000
0!
0'
#699980000000
1!
b110 %
1'
b110 +
#699990000000
0!
0'
#700000000000
1!
b111 %
1'
b111 +
#700010000000
0!
0'
#700020000000
1!
0$
b1000 %
1'
0*
b1000 +
#700030000000
0!
0'
#700040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#700050000000
0!
0'
#700060000000
1!
b0 %
1'
b0 +
#700070000000
0!
0'
#700080000000
1!
1$
b1 %
1'
1*
b1 +
#700090000000
0!
0'
#700100000000
1!
b10 %
1'
b10 +
#700110000000
0!
0'
#700120000000
1!
b11 %
1'
b11 +
#700130000000
0!
0'
#700140000000
1!
b100 %
1'
b100 +
#700150000000
0!
0'
#700160000000
1!
b101 %
1'
b101 +
#700170000000
0!
0'
#700180000000
1!
0$
b110 %
1'
0*
b110 +
#700190000000
0!
0'
#700200000000
1!
b111 %
1'
b111 +
#700210000000
0!
0'
#700220000000
1!
b1000 %
1'
b1000 +
#700230000000
0!
0'
#700240000000
1!
b1001 %
1'
b1001 +
#700250000000
1"
1(
#700260000000
0!
0"
b100 &
0'
0(
b100 ,
#700270000000
1!
b0 %
1'
b0 +
#700280000000
0!
0'
#700290000000
1!
1$
b1 %
1'
1*
b1 +
#700300000000
0!
0'
#700310000000
1!
b10 %
1'
b10 +
#700320000000
0!
0'
#700330000000
1!
b11 %
1'
b11 +
#700340000000
0!
0'
#700350000000
1!
b100 %
1'
b100 +
#700360000000
0!
0'
#700370000000
1!
b101 %
1'
b101 +
#700380000000
0!
0'
#700390000000
1!
b110 %
1'
b110 +
#700400000000
0!
0'
#700410000000
1!
b111 %
1'
b111 +
#700420000000
0!
0'
#700430000000
1!
0$
b1000 %
1'
0*
b1000 +
#700440000000
0!
0'
#700450000000
1!
b1001 %
1'
b1001 +
#700460000000
0!
0'
#700470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#700480000000
0!
0'
#700490000000
1!
1$
b1 %
1'
1*
b1 +
#700500000000
0!
0'
#700510000000
1!
b10 %
1'
b10 +
#700520000000
0!
0'
#700530000000
1!
b11 %
1'
b11 +
#700540000000
0!
0'
#700550000000
1!
b100 %
1'
b100 +
#700560000000
0!
0'
#700570000000
1!
b101 %
1'
b101 +
#700580000000
0!
0'
#700590000000
1!
0$
b110 %
1'
0*
b110 +
#700600000000
0!
0'
#700610000000
1!
b111 %
1'
b111 +
#700620000000
0!
0'
#700630000000
1!
b1000 %
1'
b1000 +
#700640000000
0!
0'
#700650000000
1!
b1001 %
1'
b1001 +
#700660000000
0!
0'
#700670000000
1!
b0 %
1'
b0 +
#700680000000
1"
1(
#700690000000
0!
0"
b100 &
0'
0(
b100 ,
#700700000000
1!
1$
b1 %
1'
1*
b1 +
#700710000000
0!
0'
#700720000000
1!
b10 %
1'
b10 +
#700730000000
0!
0'
#700740000000
1!
b11 %
1'
b11 +
#700750000000
0!
0'
#700760000000
1!
b100 %
1'
b100 +
#700770000000
0!
0'
#700780000000
1!
b101 %
1'
b101 +
#700790000000
0!
0'
#700800000000
1!
b110 %
1'
b110 +
#700810000000
0!
0'
#700820000000
1!
b111 %
1'
b111 +
#700830000000
0!
0'
#700840000000
1!
0$
b1000 %
1'
0*
b1000 +
#700850000000
0!
0'
#700860000000
1!
b1001 %
1'
b1001 +
#700870000000
0!
0'
#700880000000
1!
b0 %
1'
b0 +
#700890000000
0!
0'
#700900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#700910000000
0!
0'
#700920000000
1!
b10 %
1'
b10 +
#700930000000
0!
0'
#700940000000
1!
b11 %
1'
b11 +
#700950000000
0!
0'
#700960000000
1!
b100 %
1'
b100 +
#700970000000
0!
0'
#700980000000
1!
b101 %
1'
b101 +
#700990000000
0!
0'
#701000000000
1!
0$
b110 %
1'
0*
b110 +
#701010000000
0!
0'
#701020000000
1!
b111 %
1'
b111 +
#701030000000
0!
0'
#701040000000
1!
b1000 %
1'
b1000 +
#701050000000
0!
0'
#701060000000
1!
b1001 %
1'
b1001 +
#701070000000
0!
0'
#701080000000
1!
b0 %
1'
b0 +
#701090000000
0!
0'
#701100000000
1!
1$
b1 %
1'
1*
b1 +
#701110000000
1"
1(
#701120000000
0!
0"
b100 &
0'
0(
b100 ,
#701130000000
1!
b10 %
1'
b10 +
#701140000000
0!
0'
#701150000000
1!
b11 %
1'
b11 +
#701160000000
0!
0'
#701170000000
1!
b100 %
1'
b100 +
#701180000000
0!
0'
#701190000000
1!
b101 %
1'
b101 +
#701200000000
0!
0'
#701210000000
1!
b110 %
1'
b110 +
#701220000000
0!
0'
#701230000000
1!
b111 %
1'
b111 +
#701240000000
0!
0'
#701250000000
1!
0$
b1000 %
1'
0*
b1000 +
#701260000000
0!
0'
#701270000000
1!
b1001 %
1'
b1001 +
#701280000000
0!
0'
#701290000000
1!
b0 %
1'
b0 +
#701300000000
0!
0'
#701310000000
1!
1$
b1 %
1'
1*
b1 +
#701320000000
0!
0'
#701330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#701340000000
0!
0'
#701350000000
1!
b11 %
1'
b11 +
#701360000000
0!
0'
#701370000000
1!
b100 %
1'
b100 +
#701380000000
0!
0'
#701390000000
1!
b101 %
1'
b101 +
#701400000000
0!
0'
#701410000000
1!
0$
b110 %
1'
0*
b110 +
#701420000000
0!
0'
#701430000000
1!
b111 %
1'
b111 +
#701440000000
0!
0'
#701450000000
1!
b1000 %
1'
b1000 +
#701460000000
0!
0'
#701470000000
1!
b1001 %
1'
b1001 +
#701480000000
0!
0'
#701490000000
1!
b0 %
1'
b0 +
#701500000000
0!
0'
#701510000000
1!
1$
b1 %
1'
1*
b1 +
#701520000000
0!
0'
#701530000000
1!
b10 %
1'
b10 +
#701540000000
1"
1(
#701550000000
0!
0"
b100 &
0'
0(
b100 ,
#701560000000
1!
b11 %
1'
b11 +
#701570000000
0!
0'
#701580000000
1!
b100 %
1'
b100 +
#701590000000
0!
0'
#701600000000
1!
b101 %
1'
b101 +
#701610000000
0!
0'
#701620000000
1!
b110 %
1'
b110 +
#701630000000
0!
0'
#701640000000
1!
b111 %
1'
b111 +
#701650000000
0!
0'
#701660000000
1!
0$
b1000 %
1'
0*
b1000 +
#701670000000
0!
0'
#701680000000
1!
b1001 %
1'
b1001 +
#701690000000
0!
0'
#701700000000
1!
b0 %
1'
b0 +
#701710000000
0!
0'
#701720000000
1!
1$
b1 %
1'
1*
b1 +
#701730000000
0!
0'
#701740000000
1!
b10 %
1'
b10 +
#701750000000
0!
0'
#701760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#701770000000
0!
0'
#701780000000
1!
b100 %
1'
b100 +
#701790000000
0!
0'
#701800000000
1!
b101 %
1'
b101 +
#701810000000
0!
0'
#701820000000
1!
0$
b110 %
1'
0*
b110 +
#701830000000
0!
0'
#701840000000
1!
b111 %
1'
b111 +
#701850000000
0!
0'
#701860000000
1!
b1000 %
1'
b1000 +
#701870000000
0!
0'
#701880000000
1!
b1001 %
1'
b1001 +
#701890000000
0!
0'
#701900000000
1!
b0 %
1'
b0 +
#701910000000
0!
0'
#701920000000
1!
1$
b1 %
1'
1*
b1 +
#701930000000
0!
0'
#701940000000
1!
b10 %
1'
b10 +
#701950000000
0!
0'
#701960000000
1!
b11 %
1'
b11 +
#701970000000
1"
1(
#701980000000
0!
0"
b100 &
0'
0(
b100 ,
#701990000000
1!
b100 %
1'
b100 +
#702000000000
0!
0'
#702010000000
1!
b101 %
1'
b101 +
#702020000000
0!
0'
#702030000000
1!
b110 %
1'
b110 +
#702040000000
0!
0'
#702050000000
1!
b111 %
1'
b111 +
#702060000000
0!
0'
#702070000000
1!
0$
b1000 %
1'
0*
b1000 +
#702080000000
0!
0'
#702090000000
1!
b1001 %
1'
b1001 +
#702100000000
0!
0'
#702110000000
1!
b0 %
1'
b0 +
#702120000000
0!
0'
#702130000000
1!
1$
b1 %
1'
1*
b1 +
#702140000000
0!
0'
#702150000000
1!
b10 %
1'
b10 +
#702160000000
0!
0'
#702170000000
1!
b11 %
1'
b11 +
#702180000000
0!
0'
#702190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#702200000000
0!
0'
#702210000000
1!
b101 %
1'
b101 +
#702220000000
0!
0'
#702230000000
1!
0$
b110 %
1'
0*
b110 +
#702240000000
0!
0'
#702250000000
1!
b111 %
1'
b111 +
#702260000000
0!
0'
#702270000000
1!
b1000 %
1'
b1000 +
#702280000000
0!
0'
#702290000000
1!
b1001 %
1'
b1001 +
#702300000000
0!
0'
#702310000000
1!
b0 %
1'
b0 +
#702320000000
0!
0'
#702330000000
1!
1$
b1 %
1'
1*
b1 +
#702340000000
0!
0'
#702350000000
1!
b10 %
1'
b10 +
#702360000000
0!
0'
#702370000000
1!
b11 %
1'
b11 +
#702380000000
0!
0'
#702390000000
1!
b100 %
1'
b100 +
#702400000000
1"
1(
#702410000000
0!
0"
b100 &
0'
0(
b100 ,
#702420000000
1!
b101 %
1'
b101 +
#702430000000
0!
0'
#702440000000
1!
b110 %
1'
b110 +
#702450000000
0!
0'
#702460000000
1!
b111 %
1'
b111 +
#702470000000
0!
0'
#702480000000
1!
0$
b1000 %
1'
0*
b1000 +
#702490000000
0!
0'
#702500000000
1!
b1001 %
1'
b1001 +
#702510000000
0!
0'
#702520000000
1!
b0 %
1'
b0 +
#702530000000
0!
0'
#702540000000
1!
1$
b1 %
1'
1*
b1 +
#702550000000
0!
0'
#702560000000
1!
b10 %
1'
b10 +
#702570000000
0!
0'
#702580000000
1!
b11 %
1'
b11 +
#702590000000
0!
0'
#702600000000
1!
b100 %
1'
b100 +
#702610000000
0!
0'
#702620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#702630000000
0!
0'
#702640000000
1!
0$
b110 %
1'
0*
b110 +
#702650000000
0!
0'
#702660000000
1!
b111 %
1'
b111 +
#702670000000
0!
0'
#702680000000
1!
b1000 %
1'
b1000 +
#702690000000
0!
0'
#702700000000
1!
b1001 %
1'
b1001 +
#702710000000
0!
0'
#702720000000
1!
b0 %
1'
b0 +
#702730000000
0!
0'
#702740000000
1!
1$
b1 %
1'
1*
b1 +
#702750000000
0!
0'
#702760000000
1!
b10 %
1'
b10 +
#702770000000
0!
0'
#702780000000
1!
b11 %
1'
b11 +
#702790000000
0!
0'
#702800000000
1!
b100 %
1'
b100 +
#702810000000
0!
0'
#702820000000
1!
b101 %
1'
b101 +
#702830000000
1"
1(
#702840000000
0!
0"
b100 &
0'
0(
b100 ,
#702850000000
1!
b110 %
1'
b110 +
#702860000000
0!
0'
#702870000000
1!
b111 %
1'
b111 +
#702880000000
0!
0'
#702890000000
1!
0$
b1000 %
1'
0*
b1000 +
#702900000000
0!
0'
#702910000000
1!
b1001 %
1'
b1001 +
#702920000000
0!
0'
#702930000000
1!
b0 %
1'
b0 +
#702940000000
0!
0'
#702950000000
1!
1$
b1 %
1'
1*
b1 +
#702960000000
0!
0'
#702970000000
1!
b10 %
1'
b10 +
#702980000000
0!
0'
#702990000000
1!
b11 %
1'
b11 +
#703000000000
0!
0'
#703010000000
1!
b100 %
1'
b100 +
#703020000000
0!
0'
#703030000000
1!
b101 %
1'
b101 +
#703040000000
0!
0'
#703050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#703060000000
0!
0'
#703070000000
1!
b111 %
1'
b111 +
#703080000000
0!
0'
#703090000000
1!
b1000 %
1'
b1000 +
#703100000000
0!
0'
#703110000000
1!
b1001 %
1'
b1001 +
#703120000000
0!
0'
#703130000000
1!
b0 %
1'
b0 +
#703140000000
0!
0'
#703150000000
1!
1$
b1 %
1'
1*
b1 +
#703160000000
0!
0'
#703170000000
1!
b10 %
1'
b10 +
#703180000000
0!
0'
#703190000000
1!
b11 %
1'
b11 +
#703200000000
0!
0'
#703210000000
1!
b100 %
1'
b100 +
#703220000000
0!
0'
#703230000000
1!
b101 %
1'
b101 +
#703240000000
0!
0'
#703250000000
1!
0$
b110 %
1'
0*
b110 +
#703260000000
1"
1(
#703270000000
0!
0"
b100 &
0'
0(
b100 ,
#703280000000
1!
1$
b111 %
1'
1*
b111 +
#703290000000
0!
0'
#703300000000
1!
0$
b1000 %
1'
0*
b1000 +
#703310000000
0!
0'
#703320000000
1!
b1001 %
1'
b1001 +
#703330000000
0!
0'
#703340000000
1!
b0 %
1'
b0 +
#703350000000
0!
0'
#703360000000
1!
1$
b1 %
1'
1*
b1 +
#703370000000
0!
0'
#703380000000
1!
b10 %
1'
b10 +
#703390000000
0!
0'
#703400000000
1!
b11 %
1'
b11 +
#703410000000
0!
0'
#703420000000
1!
b100 %
1'
b100 +
#703430000000
0!
0'
#703440000000
1!
b101 %
1'
b101 +
#703450000000
0!
0'
#703460000000
1!
b110 %
1'
b110 +
#703470000000
0!
0'
#703480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#703490000000
0!
0'
#703500000000
1!
b1000 %
1'
b1000 +
#703510000000
0!
0'
#703520000000
1!
b1001 %
1'
b1001 +
#703530000000
0!
0'
#703540000000
1!
b0 %
1'
b0 +
#703550000000
0!
0'
#703560000000
1!
1$
b1 %
1'
1*
b1 +
#703570000000
0!
0'
#703580000000
1!
b10 %
1'
b10 +
#703590000000
0!
0'
#703600000000
1!
b11 %
1'
b11 +
#703610000000
0!
0'
#703620000000
1!
b100 %
1'
b100 +
#703630000000
0!
0'
#703640000000
1!
b101 %
1'
b101 +
#703650000000
0!
0'
#703660000000
1!
0$
b110 %
1'
0*
b110 +
#703670000000
0!
0'
#703680000000
1!
b111 %
1'
b111 +
#703690000000
1"
1(
#703700000000
0!
0"
b100 &
0'
0(
b100 ,
#703710000000
1!
b1000 %
1'
b1000 +
#703720000000
0!
0'
#703730000000
1!
b1001 %
1'
b1001 +
#703740000000
0!
0'
#703750000000
1!
b0 %
1'
b0 +
#703760000000
0!
0'
#703770000000
1!
1$
b1 %
1'
1*
b1 +
#703780000000
0!
0'
#703790000000
1!
b10 %
1'
b10 +
#703800000000
0!
0'
#703810000000
1!
b11 %
1'
b11 +
#703820000000
0!
0'
#703830000000
1!
b100 %
1'
b100 +
#703840000000
0!
0'
#703850000000
1!
b101 %
1'
b101 +
#703860000000
0!
0'
#703870000000
1!
b110 %
1'
b110 +
#703880000000
0!
0'
#703890000000
1!
b111 %
1'
b111 +
#703900000000
0!
0'
#703910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#703920000000
0!
0'
#703930000000
1!
b1001 %
1'
b1001 +
#703940000000
0!
0'
#703950000000
1!
b0 %
1'
b0 +
#703960000000
0!
0'
#703970000000
1!
1$
b1 %
1'
1*
b1 +
#703980000000
0!
0'
#703990000000
1!
b10 %
1'
b10 +
#704000000000
0!
0'
#704010000000
1!
b11 %
1'
b11 +
#704020000000
0!
0'
#704030000000
1!
b100 %
1'
b100 +
#704040000000
0!
0'
#704050000000
1!
b101 %
1'
b101 +
#704060000000
0!
0'
#704070000000
1!
0$
b110 %
1'
0*
b110 +
#704080000000
0!
0'
#704090000000
1!
b111 %
1'
b111 +
#704100000000
0!
0'
#704110000000
1!
b1000 %
1'
b1000 +
#704120000000
1"
1(
#704130000000
0!
0"
b100 &
0'
0(
b100 ,
#704140000000
1!
b1001 %
1'
b1001 +
#704150000000
0!
0'
#704160000000
1!
b0 %
1'
b0 +
#704170000000
0!
0'
#704180000000
1!
1$
b1 %
1'
1*
b1 +
#704190000000
0!
0'
#704200000000
1!
b10 %
1'
b10 +
#704210000000
0!
0'
#704220000000
1!
b11 %
1'
b11 +
#704230000000
0!
0'
#704240000000
1!
b100 %
1'
b100 +
#704250000000
0!
0'
#704260000000
1!
b101 %
1'
b101 +
#704270000000
0!
0'
#704280000000
1!
b110 %
1'
b110 +
#704290000000
0!
0'
#704300000000
1!
b111 %
1'
b111 +
#704310000000
0!
0'
#704320000000
1!
0$
b1000 %
1'
0*
b1000 +
#704330000000
0!
0'
#704340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#704350000000
0!
0'
#704360000000
1!
b0 %
1'
b0 +
#704370000000
0!
0'
#704380000000
1!
1$
b1 %
1'
1*
b1 +
#704390000000
0!
0'
#704400000000
1!
b10 %
1'
b10 +
#704410000000
0!
0'
#704420000000
1!
b11 %
1'
b11 +
#704430000000
0!
0'
#704440000000
1!
b100 %
1'
b100 +
#704450000000
0!
0'
#704460000000
1!
b101 %
1'
b101 +
#704470000000
0!
0'
#704480000000
1!
0$
b110 %
1'
0*
b110 +
#704490000000
0!
0'
#704500000000
1!
b111 %
1'
b111 +
#704510000000
0!
0'
#704520000000
1!
b1000 %
1'
b1000 +
#704530000000
0!
0'
#704540000000
1!
b1001 %
1'
b1001 +
#704550000000
1"
1(
#704560000000
0!
0"
b100 &
0'
0(
b100 ,
#704570000000
1!
b0 %
1'
b0 +
#704580000000
0!
0'
#704590000000
1!
1$
b1 %
1'
1*
b1 +
#704600000000
0!
0'
#704610000000
1!
b10 %
1'
b10 +
#704620000000
0!
0'
#704630000000
1!
b11 %
1'
b11 +
#704640000000
0!
0'
#704650000000
1!
b100 %
1'
b100 +
#704660000000
0!
0'
#704670000000
1!
b101 %
1'
b101 +
#704680000000
0!
0'
#704690000000
1!
b110 %
1'
b110 +
#704700000000
0!
0'
#704710000000
1!
b111 %
1'
b111 +
#704720000000
0!
0'
#704730000000
1!
0$
b1000 %
1'
0*
b1000 +
#704740000000
0!
0'
#704750000000
1!
b1001 %
1'
b1001 +
#704760000000
0!
0'
#704770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#704780000000
0!
0'
#704790000000
1!
1$
b1 %
1'
1*
b1 +
#704800000000
0!
0'
#704810000000
1!
b10 %
1'
b10 +
#704820000000
0!
0'
#704830000000
1!
b11 %
1'
b11 +
#704840000000
0!
0'
#704850000000
1!
b100 %
1'
b100 +
#704860000000
0!
0'
#704870000000
1!
b101 %
1'
b101 +
#704880000000
0!
0'
#704890000000
1!
0$
b110 %
1'
0*
b110 +
#704900000000
0!
0'
#704910000000
1!
b111 %
1'
b111 +
#704920000000
0!
0'
#704930000000
1!
b1000 %
1'
b1000 +
#704940000000
0!
0'
#704950000000
1!
b1001 %
1'
b1001 +
#704960000000
0!
0'
#704970000000
1!
b0 %
1'
b0 +
#704980000000
1"
1(
#704990000000
0!
0"
b100 &
0'
0(
b100 ,
#705000000000
1!
1$
b1 %
1'
1*
b1 +
#705010000000
0!
0'
#705020000000
1!
b10 %
1'
b10 +
#705030000000
0!
0'
#705040000000
1!
b11 %
1'
b11 +
#705050000000
0!
0'
#705060000000
1!
b100 %
1'
b100 +
#705070000000
0!
0'
#705080000000
1!
b101 %
1'
b101 +
#705090000000
0!
0'
#705100000000
1!
b110 %
1'
b110 +
#705110000000
0!
0'
#705120000000
1!
b111 %
1'
b111 +
#705130000000
0!
0'
#705140000000
1!
0$
b1000 %
1'
0*
b1000 +
#705150000000
0!
0'
#705160000000
1!
b1001 %
1'
b1001 +
#705170000000
0!
0'
#705180000000
1!
b0 %
1'
b0 +
#705190000000
0!
0'
#705200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#705210000000
0!
0'
#705220000000
1!
b10 %
1'
b10 +
#705230000000
0!
0'
#705240000000
1!
b11 %
1'
b11 +
#705250000000
0!
0'
#705260000000
1!
b100 %
1'
b100 +
#705270000000
0!
0'
#705280000000
1!
b101 %
1'
b101 +
#705290000000
0!
0'
#705300000000
1!
0$
b110 %
1'
0*
b110 +
#705310000000
0!
0'
#705320000000
1!
b111 %
1'
b111 +
#705330000000
0!
0'
#705340000000
1!
b1000 %
1'
b1000 +
#705350000000
0!
0'
#705360000000
1!
b1001 %
1'
b1001 +
#705370000000
0!
0'
#705380000000
1!
b0 %
1'
b0 +
#705390000000
0!
0'
#705400000000
1!
1$
b1 %
1'
1*
b1 +
#705410000000
1"
1(
#705420000000
0!
0"
b100 &
0'
0(
b100 ,
#705430000000
1!
b10 %
1'
b10 +
#705440000000
0!
0'
#705450000000
1!
b11 %
1'
b11 +
#705460000000
0!
0'
#705470000000
1!
b100 %
1'
b100 +
#705480000000
0!
0'
#705490000000
1!
b101 %
1'
b101 +
#705500000000
0!
0'
#705510000000
1!
b110 %
1'
b110 +
#705520000000
0!
0'
#705530000000
1!
b111 %
1'
b111 +
#705540000000
0!
0'
#705550000000
1!
0$
b1000 %
1'
0*
b1000 +
#705560000000
0!
0'
#705570000000
1!
b1001 %
1'
b1001 +
#705580000000
0!
0'
#705590000000
1!
b0 %
1'
b0 +
#705600000000
0!
0'
#705610000000
1!
1$
b1 %
1'
1*
b1 +
#705620000000
0!
0'
#705630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#705640000000
0!
0'
#705650000000
1!
b11 %
1'
b11 +
#705660000000
0!
0'
#705670000000
1!
b100 %
1'
b100 +
#705680000000
0!
0'
#705690000000
1!
b101 %
1'
b101 +
#705700000000
0!
0'
#705710000000
1!
0$
b110 %
1'
0*
b110 +
#705720000000
0!
0'
#705730000000
1!
b111 %
1'
b111 +
#705740000000
0!
0'
#705750000000
1!
b1000 %
1'
b1000 +
#705760000000
0!
0'
#705770000000
1!
b1001 %
1'
b1001 +
#705780000000
0!
0'
#705790000000
1!
b0 %
1'
b0 +
#705800000000
0!
0'
#705810000000
1!
1$
b1 %
1'
1*
b1 +
#705820000000
0!
0'
#705830000000
1!
b10 %
1'
b10 +
#705840000000
1"
1(
#705850000000
0!
0"
b100 &
0'
0(
b100 ,
#705860000000
1!
b11 %
1'
b11 +
#705870000000
0!
0'
#705880000000
1!
b100 %
1'
b100 +
#705890000000
0!
0'
#705900000000
1!
b101 %
1'
b101 +
#705910000000
0!
0'
#705920000000
1!
b110 %
1'
b110 +
#705930000000
0!
0'
#705940000000
1!
b111 %
1'
b111 +
#705950000000
0!
0'
#705960000000
1!
0$
b1000 %
1'
0*
b1000 +
#705970000000
0!
0'
#705980000000
1!
b1001 %
1'
b1001 +
#705990000000
0!
0'
#706000000000
1!
b0 %
1'
b0 +
#706010000000
0!
0'
#706020000000
1!
1$
b1 %
1'
1*
b1 +
#706030000000
0!
0'
#706040000000
1!
b10 %
1'
b10 +
#706050000000
0!
0'
#706060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#706070000000
0!
0'
#706080000000
1!
b100 %
1'
b100 +
#706090000000
0!
0'
#706100000000
1!
b101 %
1'
b101 +
#706110000000
0!
0'
#706120000000
1!
0$
b110 %
1'
0*
b110 +
#706130000000
0!
0'
#706140000000
1!
b111 %
1'
b111 +
#706150000000
0!
0'
#706160000000
1!
b1000 %
1'
b1000 +
#706170000000
0!
0'
#706180000000
1!
b1001 %
1'
b1001 +
#706190000000
0!
0'
#706200000000
1!
b0 %
1'
b0 +
#706210000000
0!
0'
#706220000000
1!
1$
b1 %
1'
1*
b1 +
#706230000000
0!
0'
#706240000000
1!
b10 %
1'
b10 +
#706250000000
0!
0'
#706260000000
1!
b11 %
1'
b11 +
#706270000000
1"
1(
#706280000000
0!
0"
b100 &
0'
0(
b100 ,
#706290000000
1!
b100 %
1'
b100 +
#706300000000
0!
0'
#706310000000
1!
b101 %
1'
b101 +
#706320000000
0!
0'
#706330000000
1!
b110 %
1'
b110 +
#706340000000
0!
0'
#706350000000
1!
b111 %
1'
b111 +
#706360000000
0!
0'
#706370000000
1!
0$
b1000 %
1'
0*
b1000 +
#706380000000
0!
0'
#706390000000
1!
b1001 %
1'
b1001 +
#706400000000
0!
0'
#706410000000
1!
b0 %
1'
b0 +
#706420000000
0!
0'
#706430000000
1!
1$
b1 %
1'
1*
b1 +
#706440000000
0!
0'
#706450000000
1!
b10 %
1'
b10 +
#706460000000
0!
0'
#706470000000
1!
b11 %
1'
b11 +
#706480000000
0!
0'
#706490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#706500000000
0!
0'
#706510000000
1!
b101 %
1'
b101 +
#706520000000
0!
0'
#706530000000
1!
0$
b110 %
1'
0*
b110 +
#706540000000
0!
0'
#706550000000
1!
b111 %
1'
b111 +
#706560000000
0!
0'
#706570000000
1!
b1000 %
1'
b1000 +
#706580000000
0!
0'
#706590000000
1!
b1001 %
1'
b1001 +
#706600000000
0!
0'
#706610000000
1!
b0 %
1'
b0 +
#706620000000
0!
0'
#706630000000
1!
1$
b1 %
1'
1*
b1 +
#706640000000
0!
0'
#706650000000
1!
b10 %
1'
b10 +
#706660000000
0!
0'
#706670000000
1!
b11 %
1'
b11 +
#706680000000
0!
0'
#706690000000
1!
b100 %
1'
b100 +
#706700000000
1"
1(
#706710000000
0!
0"
b100 &
0'
0(
b100 ,
#706720000000
1!
b101 %
1'
b101 +
#706730000000
0!
0'
#706740000000
1!
b110 %
1'
b110 +
#706750000000
0!
0'
#706760000000
1!
b111 %
1'
b111 +
#706770000000
0!
0'
#706780000000
1!
0$
b1000 %
1'
0*
b1000 +
#706790000000
0!
0'
#706800000000
1!
b1001 %
1'
b1001 +
#706810000000
0!
0'
#706820000000
1!
b0 %
1'
b0 +
#706830000000
0!
0'
#706840000000
1!
1$
b1 %
1'
1*
b1 +
#706850000000
0!
0'
#706860000000
1!
b10 %
1'
b10 +
#706870000000
0!
0'
#706880000000
1!
b11 %
1'
b11 +
#706890000000
0!
0'
#706900000000
1!
b100 %
1'
b100 +
#706910000000
0!
0'
#706920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#706930000000
0!
0'
#706940000000
1!
0$
b110 %
1'
0*
b110 +
#706950000000
0!
0'
#706960000000
1!
b111 %
1'
b111 +
#706970000000
0!
0'
#706980000000
1!
b1000 %
1'
b1000 +
#706990000000
0!
0'
#707000000000
1!
b1001 %
1'
b1001 +
#707010000000
0!
0'
#707020000000
1!
b0 %
1'
b0 +
#707030000000
0!
0'
#707040000000
1!
1$
b1 %
1'
1*
b1 +
#707050000000
0!
0'
#707060000000
1!
b10 %
1'
b10 +
#707070000000
0!
0'
#707080000000
1!
b11 %
1'
b11 +
#707090000000
0!
0'
#707100000000
1!
b100 %
1'
b100 +
#707110000000
0!
0'
#707120000000
1!
b101 %
1'
b101 +
#707130000000
1"
1(
#707140000000
0!
0"
b100 &
0'
0(
b100 ,
#707150000000
1!
b110 %
1'
b110 +
#707160000000
0!
0'
#707170000000
1!
b111 %
1'
b111 +
#707180000000
0!
0'
#707190000000
1!
0$
b1000 %
1'
0*
b1000 +
#707200000000
0!
0'
#707210000000
1!
b1001 %
1'
b1001 +
#707220000000
0!
0'
#707230000000
1!
b0 %
1'
b0 +
#707240000000
0!
0'
#707250000000
1!
1$
b1 %
1'
1*
b1 +
#707260000000
0!
0'
#707270000000
1!
b10 %
1'
b10 +
#707280000000
0!
0'
#707290000000
1!
b11 %
1'
b11 +
#707300000000
0!
0'
#707310000000
1!
b100 %
1'
b100 +
#707320000000
0!
0'
#707330000000
1!
b101 %
1'
b101 +
#707340000000
0!
0'
#707350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#707360000000
0!
0'
#707370000000
1!
b111 %
1'
b111 +
#707380000000
0!
0'
#707390000000
1!
b1000 %
1'
b1000 +
#707400000000
0!
0'
#707410000000
1!
b1001 %
1'
b1001 +
#707420000000
0!
0'
#707430000000
1!
b0 %
1'
b0 +
#707440000000
0!
0'
#707450000000
1!
1$
b1 %
1'
1*
b1 +
#707460000000
0!
0'
#707470000000
1!
b10 %
1'
b10 +
#707480000000
0!
0'
#707490000000
1!
b11 %
1'
b11 +
#707500000000
0!
0'
#707510000000
1!
b100 %
1'
b100 +
#707520000000
0!
0'
#707530000000
1!
b101 %
1'
b101 +
#707540000000
0!
0'
#707550000000
1!
0$
b110 %
1'
0*
b110 +
#707560000000
1"
1(
#707570000000
0!
0"
b100 &
0'
0(
b100 ,
#707580000000
1!
1$
b111 %
1'
1*
b111 +
#707590000000
0!
0'
#707600000000
1!
0$
b1000 %
1'
0*
b1000 +
#707610000000
0!
0'
#707620000000
1!
b1001 %
1'
b1001 +
#707630000000
0!
0'
#707640000000
1!
b0 %
1'
b0 +
#707650000000
0!
0'
#707660000000
1!
1$
b1 %
1'
1*
b1 +
#707670000000
0!
0'
#707680000000
1!
b10 %
1'
b10 +
#707690000000
0!
0'
#707700000000
1!
b11 %
1'
b11 +
#707710000000
0!
0'
#707720000000
1!
b100 %
1'
b100 +
#707730000000
0!
0'
#707740000000
1!
b101 %
1'
b101 +
#707750000000
0!
0'
#707760000000
1!
b110 %
1'
b110 +
#707770000000
0!
0'
#707780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#707790000000
0!
0'
#707800000000
1!
b1000 %
1'
b1000 +
#707810000000
0!
0'
#707820000000
1!
b1001 %
1'
b1001 +
#707830000000
0!
0'
#707840000000
1!
b0 %
1'
b0 +
#707850000000
0!
0'
#707860000000
1!
1$
b1 %
1'
1*
b1 +
#707870000000
0!
0'
#707880000000
1!
b10 %
1'
b10 +
#707890000000
0!
0'
#707900000000
1!
b11 %
1'
b11 +
#707910000000
0!
0'
#707920000000
1!
b100 %
1'
b100 +
#707930000000
0!
0'
#707940000000
1!
b101 %
1'
b101 +
#707950000000
0!
0'
#707960000000
1!
0$
b110 %
1'
0*
b110 +
#707970000000
0!
0'
#707980000000
1!
b111 %
1'
b111 +
#707990000000
1"
1(
#708000000000
0!
0"
b100 &
0'
0(
b100 ,
#708010000000
1!
b1000 %
1'
b1000 +
#708020000000
0!
0'
#708030000000
1!
b1001 %
1'
b1001 +
#708040000000
0!
0'
#708050000000
1!
b0 %
1'
b0 +
#708060000000
0!
0'
#708070000000
1!
1$
b1 %
1'
1*
b1 +
#708080000000
0!
0'
#708090000000
1!
b10 %
1'
b10 +
#708100000000
0!
0'
#708110000000
1!
b11 %
1'
b11 +
#708120000000
0!
0'
#708130000000
1!
b100 %
1'
b100 +
#708140000000
0!
0'
#708150000000
1!
b101 %
1'
b101 +
#708160000000
0!
0'
#708170000000
1!
b110 %
1'
b110 +
#708180000000
0!
0'
#708190000000
1!
b111 %
1'
b111 +
#708200000000
0!
0'
#708210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#708220000000
0!
0'
#708230000000
1!
b1001 %
1'
b1001 +
#708240000000
0!
0'
#708250000000
1!
b0 %
1'
b0 +
#708260000000
0!
0'
#708270000000
1!
1$
b1 %
1'
1*
b1 +
#708280000000
0!
0'
#708290000000
1!
b10 %
1'
b10 +
#708300000000
0!
0'
#708310000000
1!
b11 %
1'
b11 +
#708320000000
0!
0'
#708330000000
1!
b100 %
1'
b100 +
#708340000000
0!
0'
#708350000000
1!
b101 %
1'
b101 +
#708360000000
0!
0'
#708370000000
1!
0$
b110 %
1'
0*
b110 +
#708380000000
0!
0'
#708390000000
1!
b111 %
1'
b111 +
#708400000000
0!
0'
#708410000000
1!
b1000 %
1'
b1000 +
#708420000000
1"
1(
#708430000000
0!
0"
b100 &
0'
0(
b100 ,
#708440000000
1!
b1001 %
1'
b1001 +
#708450000000
0!
0'
#708460000000
1!
b0 %
1'
b0 +
#708470000000
0!
0'
#708480000000
1!
1$
b1 %
1'
1*
b1 +
#708490000000
0!
0'
#708500000000
1!
b10 %
1'
b10 +
#708510000000
0!
0'
#708520000000
1!
b11 %
1'
b11 +
#708530000000
0!
0'
#708540000000
1!
b100 %
1'
b100 +
#708550000000
0!
0'
#708560000000
1!
b101 %
1'
b101 +
#708570000000
0!
0'
#708580000000
1!
b110 %
1'
b110 +
#708590000000
0!
0'
#708600000000
1!
b111 %
1'
b111 +
#708610000000
0!
0'
#708620000000
1!
0$
b1000 %
1'
0*
b1000 +
#708630000000
0!
0'
#708640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#708650000000
0!
0'
#708660000000
1!
b0 %
1'
b0 +
#708670000000
0!
0'
#708680000000
1!
1$
b1 %
1'
1*
b1 +
#708690000000
0!
0'
#708700000000
1!
b10 %
1'
b10 +
#708710000000
0!
0'
#708720000000
1!
b11 %
1'
b11 +
#708730000000
0!
0'
#708740000000
1!
b100 %
1'
b100 +
#708750000000
0!
0'
#708760000000
1!
b101 %
1'
b101 +
#708770000000
0!
0'
#708780000000
1!
0$
b110 %
1'
0*
b110 +
#708790000000
0!
0'
#708800000000
1!
b111 %
1'
b111 +
#708810000000
0!
0'
#708820000000
1!
b1000 %
1'
b1000 +
#708830000000
0!
0'
#708840000000
1!
b1001 %
1'
b1001 +
#708850000000
1"
1(
#708860000000
0!
0"
b100 &
0'
0(
b100 ,
#708870000000
1!
b0 %
1'
b0 +
#708880000000
0!
0'
#708890000000
1!
1$
b1 %
1'
1*
b1 +
#708900000000
0!
0'
#708910000000
1!
b10 %
1'
b10 +
#708920000000
0!
0'
#708930000000
1!
b11 %
1'
b11 +
#708940000000
0!
0'
#708950000000
1!
b100 %
1'
b100 +
#708960000000
0!
0'
#708970000000
1!
b101 %
1'
b101 +
#708980000000
0!
0'
#708990000000
1!
b110 %
1'
b110 +
#709000000000
0!
0'
#709010000000
1!
b111 %
1'
b111 +
#709020000000
0!
0'
#709030000000
1!
0$
b1000 %
1'
0*
b1000 +
#709040000000
0!
0'
#709050000000
1!
b1001 %
1'
b1001 +
#709060000000
0!
0'
#709070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#709080000000
0!
0'
#709090000000
1!
1$
b1 %
1'
1*
b1 +
#709100000000
0!
0'
#709110000000
1!
b10 %
1'
b10 +
#709120000000
0!
0'
#709130000000
1!
b11 %
1'
b11 +
#709140000000
0!
0'
#709150000000
1!
b100 %
1'
b100 +
#709160000000
0!
0'
#709170000000
1!
b101 %
1'
b101 +
#709180000000
0!
0'
#709190000000
1!
0$
b110 %
1'
0*
b110 +
#709200000000
0!
0'
#709210000000
1!
b111 %
1'
b111 +
#709220000000
0!
0'
#709230000000
1!
b1000 %
1'
b1000 +
#709240000000
0!
0'
#709250000000
1!
b1001 %
1'
b1001 +
#709260000000
0!
0'
#709270000000
1!
b0 %
1'
b0 +
#709280000000
1"
1(
#709290000000
0!
0"
b100 &
0'
0(
b100 ,
#709300000000
1!
1$
b1 %
1'
1*
b1 +
#709310000000
0!
0'
#709320000000
1!
b10 %
1'
b10 +
#709330000000
0!
0'
#709340000000
1!
b11 %
1'
b11 +
#709350000000
0!
0'
#709360000000
1!
b100 %
1'
b100 +
#709370000000
0!
0'
#709380000000
1!
b101 %
1'
b101 +
#709390000000
0!
0'
#709400000000
1!
b110 %
1'
b110 +
#709410000000
0!
0'
#709420000000
1!
b111 %
1'
b111 +
#709430000000
0!
0'
#709440000000
1!
0$
b1000 %
1'
0*
b1000 +
#709450000000
0!
0'
#709460000000
1!
b1001 %
1'
b1001 +
#709470000000
0!
0'
#709480000000
1!
b0 %
1'
b0 +
#709490000000
0!
0'
#709500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#709510000000
0!
0'
#709520000000
1!
b10 %
1'
b10 +
#709530000000
0!
0'
#709540000000
1!
b11 %
1'
b11 +
#709550000000
0!
0'
#709560000000
1!
b100 %
1'
b100 +
#709570000000
0!
0'
#709580000000
1!
b101 %
1'
b101 +
#709590000000
0!
0'
#709600000000
1!
0$
b110 %
1'
0*
b110 +
#709610000000
0!
0'
#709620000000
1!
b111 %
1'
b111 +
#709630000000
0!
0'
#709640000000
1!
b1000 %
1'
b1000 +
#709650000000
0!
0'
#709660000000
1!
b1001 %
1'
b1001 +
#709670000000
0!
0'
#709680000000
1!
b0 %
1'
b0 +
#709690000000
0!
0'
#709700000000
1!
1$
b1 %
1'
1*
b1 +
#709710000000
1"
1(
#709720000000
0!
0"
b100 &
0'
0(
b100 ,
#709730000000
1!
b10 %
1'
b10 +
#709740000000
0!
0'
#709750000000
1!
b11 %
1'
b11 +
#709760000000
0!
0'
#709770000000
1!
b100 %
1'
b100 +
#709780000000
0!
0'
#709790000000
1!
b101 %
1'
b101 +
#709800000000
0!
0'
#709810000000
1!
b110 %
1'
b110 +
#709820000000
0!
0'
#709830000000
1!
b111 %
1'
b111 +
#709840000000
0!
0'
#709850000000
1!
0$
b1000 %
1'
0*
b1000 +
#709860000000
0!
0'
#709870000000
1!
b1001 %
1'
b1001 +
#709880000000
0!
0'
#709890000000
1!
b0 %
1'
b0 +
#709900000000
0!
0'
#709910000000
1!
1$
b1 %
1'
1*
b1 +
#709920000000
0!
0'
#709930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#709940000000
0!
0'
#709950000000
1!
b11 %
1'
b11 +
#709960000000
0!
0'
#709970000000
1!
b100 %
1'
b100 +
#709980000000
0!
0'
#709990000000
1!
b101 %
1'
b101 +
#710000000000
0!
0'
#710010000000
1!
0$
b110 %
1'
0*
b110 +
#710020000000
0!
0'
#710030000000
1!
b111 %
1'
b111 +
#710040000000
0!
0'
#710050000000
1!
b1000 %
1'
b1000 +
#710060000000
0!
0'
#710070000000
1!
b1001 %
1'
b1001 +
#710080000000
0!
0'
#710090000000
1!
b0 %
1'
b0 +
#710100000000
0!
0'
#710110000000
1!
1$
b1 %
1'
1*
b1 +
#710120000000
0!
0'
#710130000000
1!
b10 %
1'
b10 +
#710140000000
1"
1(
#710150000000
0!
0"
b100 &
0'
0(
b100 ,
#710160000000
1!
b11 %
1'
b11 +
#710170000000
0!
0'
#710180000000
1!
b100 %
1'
b100 +
#710190000000
0!
0'
#710200000000
1!
b101 %
1'
b101 +
#710210000000
0!
0'
#710220000000
1!
b110 %
1'
b110 +
#710230000000
0!
0'
#710240000000
1!
b111 %
1'
b111 +
#710250000000
0!
0'
#710260000000
1!
0$
b1000 %
1'
0*
b1000 +
#710270000000
0!
0'
#710280000000
1!
b1001 %
1'
b1001 +
#710290000000
0!
0'
#710300000000
1!
b0 %
1'
b0 +
#710310000000
0!
0'
#710320000000
1!
1$
b1 %
1'
1*
b1 +
#710330000000
0!
0'
#710340000000
1!
b10 %
1'
b10 +
#710350000000
0!
0'
#710360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#710370000000
0!
0'
#710380000000
1!
b100 %
1'
b100 +
#710390000000
0!
0'
#710400000000
1!
b101 %
1'
b101 +
#710410000000
0!
0'
#710420000000
1!
0$
b110 %
1'
0*
b110 +
#710430000000
0!
0'
#710440000000
1!
b111 %
1'
b111 +
#710450000000
0!
0'
#710460000000
1!
b1000 %
1'
b1000 +
#710470000000
0!
0'
#710480000000
1!
b1001 %
1'
b1001 +
#710490000000
0!
0'
#710500000000
1!
b0 %
1'
b0 +
#710510000000
0!
0'
#710520000000
1!
1$
b1 %
1'
1*
b1 +
#710530000000
0!
0'
#710540000000
1!
b10 %
1'
b10 +
#710550000000
0!
0'
#710560000000
1!
b11 %
1'
b11 +
#710570000000
1"
1(
#710580000000
0!
0"
b100 &
0'
0(
b100 ,
#710590000000
1!
b100 %
1'
b100 +
#710600000000
0!
0'
#710610000000
1!
b101 %
1'
b101 +
#710620000000
0!
0'
#710630000000
1!
b110 %
1'
b110 +
#710640000000
0!
0'
#710650000000
1!
b111 %
1'
b111 +
#710660000000
0!
0'
#710670000000
1!
0$
b1000 %
1'
0*
b1000 +
#710680000000
0!
0'
#710690000000
1!
b1001 %
1'
b1001 +
#710700000000
0!
0'
#710710000000
1!
b0 %
1'
b0 +
#710720000000
0!
0'
#710730000000
1!
1$
b1 %
1'
1*
b1 +
#710740000000
0!
0'
#710750000000
1!
b10 %
1'
b10 +
#710760000000
0!
0'
#710770000000
1!
b11 %
1'
b11 +
#710780000000
0!
0'
#710790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#710800000000
0!
0'
#710810000000
1!
b101 %
1'
b101 +
#710820000000
0!
0'
#710830000000
1!
0$
b110 %
1'
0*
b110 +
#710840000000
0!
0'
#710850000000
1!
b111 %
1'
b111 +
#710860000000
0!
0'
#710870000000
1!
b1000 %
1'
b1000 +
#710880000000
0!
0'
#710890000000
1!
b1001 %
1'
b1001 +
#710900000000
0!
0'
#710910000000
1!
b0 %
1'
b0 +
#710920000000
0!
0'
#710930000000
1!
1$
b1 %
1'
1*
b1 +
#710940000000
0!
0'
#710950000000
1!
b10 %
1'
b10 +
#710960000000
0!
0'
#710970000000
1!
b11 %
1'
b11 +
#710980000000
0!
0'
#710990000000
1!
b100 %
1'
b100 +
#711000000000
1"
1(
#711010000000
0!
0"
b100 &
0'
0(
b100 ,
#711020000000
1!
b101 %
1'
b101 +
#711030000000
0!
0'
#711040000000
1!
b110 %
1'
b110 +
#711050000000
0!
0'
#711060000000
1!
b111 %
1'
b111 +
#711070000000
0!
0'
#711080000000
1!
0$
b1000 %
1'
0*
b1000 +
#711090000000
0!
0'
#711100000000
1!
b1001 %
1'
b1001 +
#711110000000
0!
0'
#711120000000
1!
b0 %
1'
b0 +
#711130000000
0!
0'
#711140000000
1!
1$
b1 %
1'
1*
b1 +
#711150000000
0!
0'
#711160000000
1!
b10 %
1'
b10 +
#711170000000
0!
0'
#711180000000
1!
b11 %
1'
b11 +
#711190000000
0!
0'
#711200000000
1!
b100 %
1'
b100 +
#711210000000
0!
0'
#711220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#711230000000
0!
0'
#711240000000
1!
0$
b110 %
1'
0*
b110 +
#711250000000
0!
0'
#711260000000
1!
b111 %
1'
b111 +
#711270000000
0!
0'
#711280000000
1!
b1000 %
1'
b1000 +
#711290000000
0!
0'
#711300000000
1!
b1001 %
1'
b1001 +
#711310000000
0!
0'
#711320000000
1!
b0 %
1'
b0 +
#711330000000
0!
0'
#711340000000
1!
1$
b1 %
1'
1*
b1 +
#711350000000
0!
0'
#711360000000
1!
b10 %
1'
b10 +
#711370000000
0!
0'
#711380000000
1!
b11 %
1'
b11 +
#711390000000
0!
0'
#711400000000
1!
b100 %
1'
b100 +
#711410000000
0!
0'
#711420000000
1!
b101 %
1'
b101 +
#711430000000
1"
1(
#711440000000
0!
0"
b100 &
0'
0(
b100 ,
#711450000000
1!
b110 %
1'
b110 +
#711460000000
0!
0'
#711470000000
1!
b111 %
1'
b111 +
#711480000000
0!
0'
#711490000000
1!
0$
b1000 %
1'
0*
b1000 +
#711500000000
0!
0'
#711510000000
1!
b1001 %
1'
b1001 +
#711520000000
0!
0'
#711530000000
1!
b0 %
1'
b0 +
#711540000000
0!
0'
#711550000000
1!
1$
b1 %
1'
1*
b1 +
#711560000000
0!
0'
#711570000000
1!
b10 %
1'
b10 +
#711580000000
0!
0'
#711590000000
1!
b11 %
1'
b11 +
#711600000000
0!
0'
#711610000000
1!
b100 %
1'
b100 +
#711620000000
0!
0'
#711630000000
1!
b101 %
1'
b101 +
#711640000000
0!
0'
#711650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#711660000000
0!
0'
#711670000000
1!
b111 %
1'
b111 +
#711680000000
0!
0'
#711690000000
1!
b1000 %
1'
b1000 +
#711700000000
0!
0'
#711710000000
1!
b1001 %
1'
b1001 +
#711720000000
0!
0'
#711730000000
1!
b0 %
1'
b0 +
#711740000000
0!
0'
#711750000000
1!
1$
b1 %
1'
1*
b1 +
#711760000000
0!
0'
#711770000000
1!
b10 %
1'
b10 +
#711780000000
0!
0'
#711790000000
1!
b11 %
1'
b11 +
#711800000000
0!
0'
#711810000000
1!
b100 %
1'
b100 +
#711820000000
0!
0'
#711830000000
1!
b101 %
1'
b101 +
#711840000000
0!
0'
#711850000000
1!
0$
b110 %
1'
0*
b110 +
#711860000000
1"
1(
#711870000000
0!
0"
b100 &
0'
0(
b100 ,
#711880000000
1!
1$
b111 %
1'
1*
b111 +
#711890000000
0!
0'
#711900000000
1!
0$
b1000 %
1'
0*
b1000 +
#711910000000
0!
0'
#711920000000
1!
b1001 %
1'
b1001 +
#711930000000
0!
0'
#711940000000
1!
b0 %
1'
b0 +
#711950000000
0!
0'
#711960000000
1!
1$
b1 %
1'
1*
b1 +
#711970000000
0!
0'
#711980000000
1!
b10 %
1'
b10 +
#711990000000
0!
0'
#712000000000
1!
b11 %
1'
b11 +
#712010000000
0!
0'
#712020000000
1!
b100 %
1'
b100 +
#712030000000
0!
0'
#712040000000
1!
b101 %
1'
b101 +
#712050000000
0!
0'
#712060000000
1!
b110 %
1'
b110 +
#712070000000
0!
0'
#712080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#712090000000
0!
0'
#712100000000
1!
b1000 %
1'
b1000 +
#712110000000
0!
0'
#712120000000
1!
b1001 %
1'
b1001 +
#712130000000
0!
0'
#712140000000
1!
b0 %
1'
b0 +
#712150000000
0!
0'
#712160000000
1!
1$
b1 %
1'
1*
b1 +
#712170000000
0!
0'
#712180000000
1!
b10 %
1'
b10 +
#712190000000
0!
0'
#712200000000
1!
b11 %
1'
b11 +
#712210000000
0!
0'
#712220000000
1!
b100 %
1'
b100 +
#712230000000
0!
0'
#712240000000
1!
b101 %
1'
b101 +
#712250000000
0!
0'
#712260000000
1!
0$
b110 %
1'
0*
b110 +
#712270000000
0!
0'
#712280000000
1!
b111 %
1'
b111 +
#712290000000
1"
1(
#712300000000
0!
0"
b100 &
0'
0(
b100 ,
#712310000000
1!
b1000 %
1'
b1000 +
#712320000000
0!
0'
#712330000000
1!
b1001 %
1'
b1001 +
#712340000000
0!
0'
#712350000000
1!
b0 %
1'
b0 +
#712360000000
0!
0'
#712370000000
1!
1$
b1 %
1'
1*
b1 +
#712380000000
0!
0'
#712390000000
1!
b10 %
1'
b10 +
#712400000000
0!
0'
#712410000000
1!
b11 %
1'
b11 +
#712420000000
0!
0'
#712430000000
1!
b100 %
1'
b100 +
#712440000000
0!
0'
#712450000000
1!
b101 %
1'
b101 +
#712460000000
0!
0'
#712470000000
1!
b110 %
1'
b110 +
#712480000000
0!
0'
#712490000000
1!
b111 %
1'
b111 +
#712500000000
0!
0'
#712510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#712520000000
0!
0'
#712530000000
1!
b1001 %
1'
b1001 +
#712540000000
0!
0'
#712550000000
1!
b0 %
1'
b0 +
#712560000000
0!
0'
#712570000000
1!
1$
b1 %
1'
1*
b1 +
#712580000000
0!
0'
#712590000000
1!
b10 %
1'
b10 +
#712600000000
0!
0'
#712610000000
1!
b11 %
1'
b11 +
#712620000000
0!
0'
#712630000000
1!
b100 %
1'
b100 +
#712640000000
0!
0'
#712650000000
1!
b101 %
1'
b101 +
#712660000000
0!
0'
#712670000000
1!
0$
b110 %
1'
0*
b110 +
#712680000000
0!
0'
#712690000000
1!
b111 %
1'
b111 +
#712700000000
0!
0'
#712710000000
1!
b1000 %
1'
b1000 +
#712720000000
1"
1(
#712730000000
0!
0"
b100 &
0'
0(
b100 ,
#712740000000
1!
b1001 %
1'
b1001 +
#712750000000
0!
0'
#712760000000
1!
b0 %
1'
b0 +
#712770000000
0!
0'
#712780000000
1!
1$
b1 %
1'
1*
b1 +
#712790000000
0!
0'
#712800000000
1!
b10 %
1'
b10 +
#712810000000
0!
0'
#712820000000
1!
b11 %
1'
b11 +
#712830000000
0!
0'
#712840000000
1!
b100 %
1'
b100 +
#712850000000
0!
0'
#712860000000
1!
b101 %
1'
b101 +
#712870000000
0!
0'
#712880000000
1!
b110 %
1'
b110 +
#712890000000
0!
0'
#712900000000
1!
b111 %
1'
b111 +
#712910000000
0!
0'
#712920000000
1!
0$
b1000 %
1'
0*
b1000 +
#712930000000
0!
0'
#712940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#712950000000
0!
0'
#712960000000
1!
b0 %
1'
b0 +
#712970000000
0!
0'
#712980000000
1!
1$
b1 %
1'
1*
b1 +
#712990000000
0!
0'
#713000000000
1!
b10 %
1'
b10 +
#713010000000
0!
0'
#713020000000
1!
b11 %
1'
b11 +
#713030000000
0!
0'
#713040000000
1!
b100 %
1'
b100 +
#713050000000
0!
0'
#713060000000
1!
b101 %
1'
b101 +
#713070000000
0!
0'
#713080000000
1!
0$
b110 %
1'
0*
b110 +
#713090000000
0!
0'
#713100000000
1!
b111 %
1'
b111 +
#713110000000
0!
0'
#713120000000
1!
b1000 %
1'
b1000 +
#713130000000
0!
0'
#713140000000
1!
b1001 %
1'
b1001 +
#713150000000
1"
1(
#713160000000
0!
0"
b100 &
0'
0(
b100 ,
#713170000000
1!
b0 %
1'
b0 +
#713180000000
0!
0'
#713190000000
1!
1$
b1 %
1'
1*
b1 +
#713200000000
0!
0'
#713210000000
1!
b10 %
1'
b10 +
#713220000000
0!
0'
#713230000000
1!
b11 %
1'
b11 +
#713240000000
0!
0'
#713250000000
1!
b100 %
1'
b100 +
#713260000000
0!
0'
#713270000000
1!
b101 %
1'
b101 +
#713280000000
0!
0'
#713290000000
1!
b110 %
1'
b110 +
#713300000000
0!
0'
#713310000000
1!
b111 %
1'
b111 +
#713320000000
0!
0'
#713330000000
1!
0$
b1000 %
1'
0*
b1000 +
#713340000000
0!
0'
#713350000000
1!
b1001 %
1'
b1001 +
#713360000000
0!
0'
#713370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#713380000000
0!
0'
#713390000000
1!
1$
b1 %
1'
1*
b1 +
#713400000000
0!
0'
#713410000000
1!
b10 %
1'
b10 +
#713420000000
0!
0'
#713430000000
1!
b11 %
1'
b11 +
#713440000000
0!
0'
#713450000000
1!
b100 %
1'
b100 +
#713460000000
0!
0'
#713470000000
1!
b101 %
1'
b101 +
#713480000000
0!
0'
#713490000000
1!
0$
b110 %
1'
0*
b110 +
#713500000000
0!
0'
#713510000000
1!
b111 %
1'
b111 +
#713520000000
0!
0'
#713530000000
1!
b1000 %
1'
b1000 +
#713540000000
0!
0'
#713550000000
1!
b1001 %
1'
b1001 +
#713560000000
0!
0'
#713570000000
1!
b0 %
1'
b0 +
#713580000000
1"
1(
#713590000000
0!
0"
b100 &
0'
0(
b100 ,
#713600000000
1!
1$
b1 %
1'
1*
b1 +
#713610000000
0!
0'
#713620000000
1!
b10 %
1'
b10 +
#713630000000
0!
0'
#713640000000
1!
b11 %
1'
b11 +
#713650000000
0!
0'
#713660000000
1!
b100 %
1'
b100 +
#713670000000
0!
0'
#713680000000
1!
b101 %
1'
b101 +
#713690000000
0!
0'
#713700000000
1!
b110 %
1'
b110 +
#713710000000
0!
0'
#713720000000
1!
b111 %
1'
b111 +
#713730000000
0!
0'
#713740000000
1!
0$
b1000 %
1'
0*
b1000 +
#713750000000
0!
0'
#713760000000
1!
b1001 %
1'
b1001 +
#713770000000
0!
0'
#713780000000
1!
b0 %
1'
b0 +
#713790000000
0!
0'
#713800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#713810000000
0!
0'
#713820000000
1!
b10 %
1'
b10 +
#713830000000
0!
0'
#713840000000
1!
b11 %
1'
b11 +
#713850000000
0!
0'
#713860000000
1!
b100 %
1'
b100 +
#713870000000
0!
0'
#713880000000
1!
b101 %
1'
b101 +
#713890000000
0!
0'
#713900000000
1!
0$
b110 %
1'
0*
b110 +
#713910000000
0!
0'
#713920000000
1!
b111 %
1'
b111 +
#713930000000
0!
0'
#713940000000
1!
b1000 %
1'
b1000 +
#713950000000
0!
0'
#713960000000
1!
b1001 %
1'
b1001 +
#713970000000
0!
0'
#713980000000
1!
b0 %
1'
b0 +
#713990000000
0!
0'
#714000000000
1!
1$
b1 %
1'
1*
b1 +
#714010000000
1"
1(
#714020000000
0!
0"
b100 &
0'
0(
b100 ,
#714030000000
1!
b10 %
1'
b10 +
#714040000000
0!
0'
#714050000000
1!
b11 %
1'
b11 +
#714060000000
0!
0'
#714070000000
1!
b100 %
1'
b100 +
#714080000000
0!
0'
#714090000000
1!
b101 %
1'
b101 +
#714100000000
0!
0'
#714110000000
1!
b110 %
1'
b110 +
#714120000000
0!
0'
#714130000000
1!
b111 %
1'
b111 +
#714140000000
0!
0'
#714150000000
1!
0$
b1000 %
1'
0*
b1000 +
#714160000000
0!
0'
#714170000000
1!
b1001 %
1'
b1001 +
#714180000000
0!
0'
#714190000000
1!
b0 %
1'
b0 +
#714200000000
0!
0'
#714210000000
1!
1$
b1 %
1'
1*
b1 +
#714220000000
0!
0'
#714230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#714240000000
0!
0'
#714250000000
1!
b11 %
1'
b11 +
#714260000000
0!
0'
#714270000000
1!
b100 %
1'
b100 +
#714280000000
0!
0'
#714290000000
1!
b101 %
1'
b101 +
#714300000000
0!
0'
#714310000000
1!
0$
b110 %
1'
0*
b110 +
#714320000000
0!
0'
#714330000000
1!
b111 %
1'
b111 +
#714340000000
0!
0'
#714350000000
1!
b1000 %
1'
b1000 +
#714360000000
0!
0'
#714370000000
1!
b1001 %
1'
b1001 +
#714380000000
0!
0'
#714390000000
1!
b0 %
1'
b0 +
#714400000000
0!
0'
#714410000000
1!
1$
b1 %
1'
1*
b1 +
#714420000000
0!
0'
#714430000000
1!
b10 %
1'
b10 +
#714440000000
1"
1(
#714450000000
0!
0"
b100 &
0'
0(
b100 ,
#714460000000
1!
b11 %
1'
b11 +
#714470000000
0!
0'
#714480000000
1!
b100 %
1'
b100 +
#714490000000
0!
0'
#714500000000
1!
b101 %
1'
b101 +
#714510000000
0!
0'
#714520000000
1!
b110 %
1'
b110 +
#714530000000
0!
0'
#714540000000
1!
b111 %
1'
b111 +
#714550000000
0!
0'
#714560000000
1!
0$
b1000 %
1'
0*
b1000 +
#714570000000
0!
0'
#714580000000
1!
b1001 %
1'
b1001 +
#714590000000
0!
0'
#714600000000
1!
b0 %
1'
b0 +
#714610000000
0!
0'
#714620000000
1!
1$
b1 %
1'
1*
b1 +
#714630000000
0!
0'
#714640000000
1!
b10 %
1'
b10 +
#714650000000
0!
0'
#714660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#714670000000
0!
0'
#714680000000
1!
b100 %
1'
b100 +
#714690000000
0!
0'
#714700000000
1!
b101 %
1'
b101 +
#714710000000
0!
0'
#714720000000
1!
0$
b110 %
1'
0*
b110 +
#714730000000
0!
0'
#714740000000
1!
b111 %
1'
b111 +
#714750000000
0!
0'
#714760000000
1!
b1000 %
1'
b1000 +
#714770000000
0!
0'
#714780000000
1!
b1001 %
1'
b1001 +
#714790000000
0!
0'
#714800000000
1!
b0 %
1'
b0 +
#714810000000
0!
0'
#714820000000
1!
1$
b1 %
1'
1*
b1 +
#714830000000
0!
0'
#714840000000
1!
b10 %
1'
b10 +
#714850000000
0!
0'
#714860000000
1!
b11 %
1'
b11 +
#714870000000
1"
1(
#714880000000
0!
0"
b100 &
0'
0(
b100 ,
#714890000000
1!
b100 %
1'
b100 +
#714900000000
0!
0'
#714910000000
1!
b101 %
1'
b101 +
#714920000000
0!
0'
#714930000000
1!
b110 %
1'
b110 +
#714940000000
0!
0'
#714950000000
1!
b111 %
1'
b111 +
#714960000000
0!
0'
#714970000000
1!
0$
b1000 %
1'
0*
b1000 +
#714980000000
0!
0'
#714990000000
1!
b1001 %
1'
b1001 +
#715000000000
0!
0'
#715010000000
1!
b0 %
1'
b0 +
#715020000000
0!
0'
#715030000000
1!
1$
b1 %
1'
1*
b1 +
#715040000000
0!
0'
#715050000000
1!
b10 %
1'
b10 +
#715060000000
0!
0'
#715070000000
1!
b11 %
1'
b11 +
#715080000000
0!
0'
#715090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#715100000000
0!
0'
#715110000000
1!
b101 %
1'
b101 +
#715120000000
0!
0'
#715130000000
1!
0$
b110 %
1'
0*
b110 +
#715140000000
0!
0'
#715150000000
1!
b111 %
1'
b111 +
#715160000000
0!
0'
#715170000000
1!
b1000 %
1'
b1000 +
#715180000000
0!
0'
#715190000000
1!
b1001 %
1'
b1001 +
#715200000000
0!
0'
#715210000000
1!
b0 %
1'
b0 +
#715220000000
0!
0'
#715230000000
1!
1$
b1 %
1'
1*
b1 +
#715240000000
0!
0'
#715250000000
1!
b10 %
1'
b10 +
#715260000000
0!
0'
#715270000000
1!
b11 %
1'
b11 +
#715280000000
0!
0'
#715290000000
1!
b100 %
1'
b100 +
#715300000000
1"
1(
#715310000000
0!
0"
b100 &
0'
0(
b100 ,
#715320000000
1!
b101 %
1'
b101 +
#715330000000
0!
0'
#715340000000
1!
b110 %
1'
b110 +
#715350000000
0!
0'
#715360000000
1!
b111 %
1'
b111 +
#715370000000
0!
0'
#715380000000
1!
0$
b1000 %
1'
0*
b1000 +
#715390000000
0!
0'
#715400000000
1!
b1001 %
1'
b1001 +
#715410000000
0!
0'
#715420000000
1!
b0 %
1'
b0 +
#715430000000
0!
0'
#715440000000
1!
1$
b1 %
1'
1*
b1 +
#715450000000
0!
0'
#715460000000
1!
b10 %
1'
b10 +
#715470000000
0!
0'
#715480000000
1!
b11 %
1'
b11 +
#715490000000
0!
0'
#715500000000
1!
b100 %
1'
b100 +
#715510000000
0!
0'
#715520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#715530000000
0!
0'
#715540000000
1!
0$
b110 %
1'
0*
b110 +
#715550000000
0!
0'
#715560000000
1!
b111 %
1'
b111 +
#715570000000
0!
0'
#715580000000
1!
b1000 %
1'
b1000 +
#715590000000
0!
0'
#715600000000
1!
b1001 %
1'
b1001 +
#715610000000
0!
0'
#715620000000
1!
b0 %
1'
b0 +
#715630000000
0!
0'
#715640000000
1!
1$
b1 %
1'
1*
b1 +
#715650000000
0!
0'
#715660000000
1!
b10 %
1'
b10 +
#715670000000
0!
0'
#715680000000
1!
b11 %
1'
b11 +
#715690000000
0!
0'
#715700000000
1!
b100 %
1'
b100 +
#715710000000
0!
0'
#715720000000
1!
b101 %
1'
b101 +
#715730000000
1"
1(
#715740000000
0!
0"
b100 &
0'
0(
b100 ,
#715750000000
1!
b110 %
1'
b110 +
#715760000000
0!
0'
#715770000000
1!
b111 %
1'
b111 +
#715780000000
0!
0'
#715790000000
1!
0$
b1000 %
1'
0*
b1000 +
#715800000000
0!
0'
#715810000000
1!
b1001 %
1'
b1001 +
#715820000000
0!
0'
#715830000000
1!
b0 %
1'
b0 +
#715840000000
0!
0'
#715850000000
1!
1$
b1 %
1'
1*
b1 +
#715860000000
0!
0'
#715870000000
1!
b10 %
1'
b10 +
#715880000000
0!
0'
#715890000000
1!
b11 %
1'
b11 +
#715900000000
0!
0'
#715910000000
1!
b100 %
1'
b100 +
#715920000000
0!
0'
#715930000000
1!
b101 %
1'
b101 +
#715940000000
0!
0'
#715950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#715960000000
0!
0'
#715970000000
1!
b111 %
1'
b111 +
#715980000000
0!
0'
#715990000000
1!
b1000 %
1'
b1000 +
#716000000000
0!
0'
#716010000000
1!
b1001 %
1'
b1001 +
#716020000000
0!
0'
#716030000000
1!
b0 %
1'
b0 +
#716040000000
0!
0'
#716050000000
1!
1$
b1 %
1'
1*
b1 +
#716060000000
0!
0'
#716070000000
1!
b10 %
1'
b10 +
#716080000000
0!
0'
#716090000000
1!
b11 %
1'
b11 +
#716100000000
0!
0'
#716110000000
1!
b100 %
1'
b100 +
#716120000000
0!
0'
#716130000000
1!
b101 %
1'
b101 +
#716140000000
0!
0'
#716150000000
1!
0$
b110 %
1'
0*
b110 +
#716160000000
1"
1(
#716170000000
0!
0"
b100 &
0'
0(
b100 ,
#716180000000
1!
1$
b111 %
1'
1*
b111 +
#716190000000
0!
0'
#716200000000
1!
0$
b1000 %
1'
0*
b1000 +
#716210000000
0!
0'
#716220000000
1!
b1001 %
1'
b1001 +
#716230000000
0!
0'
#716240000000
1!
b0 %
1'
b0 +
#716250000000
0!
0'
#716260000000
1!
1$
b1 %
1'
1*
b1 +
#716270000000
0!
0'
#716280000000
1!
b10 %
1'
b10 +
#716290000000
0!
0'
#716300000000
1!
b11 %
1'
b11 +
#716310000000
0!
0'
#716320000000
1!
b100 %
1'
b100 +
#716330000000
0!
0'
#716340000000
1!
b101 %
1'
b101 +
#716350000000
0!
0'
#716360000000
1!
b110 %
1'
b110 +
#716370000000
0!
0'
#716380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#716390000000
0!
0'
#716400000000
1!
b1000 %
1'
b1000 +
#716410000000
0!
0'
#716420000000
1!
b1001 %
1'
b1001 +
#716430000000
0!
0'
#716440000000
1!
b0 %
1'
b0 +
#716450000000
0!
0'
#716460000000
1!
1$
b1 %
1'
1*
b1 +
#716470000000
0!
0'
#716480000000
1!
b10 %
1'
b10 +
#716490000000
0!
0'
#716500000000
1!
b11 %
1'
b11 +
#716510000000
0!
0'
#716520000000
1!
b100 %
1'
b100 +
#716530000000
0!
0'
#716540000000
1!
b101 %
1'
b101 +
#716550000000
0!
0'
#716560000000
1!
0$
b110 %
1'
0*
b110 +
#716570000000
0!
0'
#716580000000
1!
b111 %
1'
b111 +
#716590000000
1"
1(
#716600000000
0!
0"
b100 &
0'
0(
b100 ,
#716610000000
1!
b1000 %
1'
b1000 +
#716620000000
0!
0'
#716630000000
1!
b1001 %
1'
b1001 +
#716640000000
0!
0'
#716650000000
1!
b0 %
1'
b0 +
#716660000000
0!
0'
#716670000000
1!
1$
b1 %
1'
1*
b1 +
#716680000000
0!
0'
#716690000000
1!
b10 %
1'
b10 +
#716700000000
0!
0'
#716710000000
1!
b11 %
1'
b11 +
#716720000000
0!
0'
#716730000000
1!
b100 %
1'
b100 +
#716740000000
0!
0'
#716750000000
1!
b101 %
1'
b101 +
#716760000000
0!
0'
#716770000000
1!
b110 %
1'
b110 +
#716780000000
0!
0'
#716790000000
1!
b111 %
1'
b111 +
#716800000000
0!
0'
#716810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#716820000000
0!
0'
#716830000000
1!
b1001 %
1'
b1001 +
#716840000000
0!
0'
#716850000000
1!
b0 %
1'
b0 +
#716860000000
0!
0'
#716870000000
1!
1$
b1 %
1'
1*
b1 +
#716880000000
0!
0'
#716890000000
1!
b10 %
1'
b10 +
#716900000000
0!
0'
#716910000000
1!
b11 %
1'
b11 +
#716920000000
0!
0'
#716930000000
1!
b100 %
1'
b100 +
#716940000000
0!
0'
#716950000000
1!
b101 %
1'
b101 +
#716960000000
0!
0'
#716970000000
1!
0$
b110 %
1'
0*
b110 +
#716980000000
0!
0'
#716990000000
1!
b111 %
1'
b111 +
#717000000000
0!
0'
#717010000000
1!
b1000 %
1'
b1000 +
#717020000000
1"
1(
#717030000000
0!
0"
b100 &
0'
0(
b100 ,
#717040000000
1!
b1001 %
1'
b1001 +
#717050000000
0!
0'
#717060000000
1!
b0 %
1'
b0 +
#717070000000
0!
0'
#717080000000
1!
1$
b1 %
1'
1*
b1 +
#717090000000
0!
0'
#717100000000
1!
b10 %
1'
b10 +
#717110000000
0!
0'
#717120000000
1!
b11 %
1'
b11 +
#717130000000
0!
0'
#717140000000
1!
b100 %
1'
b100 +
#717150000000
0!
0'
#717160000000
1!
b101 %
1'
b101 +
#717170000000
0!
0'
#717180000000
1!
b110 %
1'
b110 +
#717190000000
0!
0'
#717200000000
1!
b111 %
1'
b111 +
#717210000000
0!
0'
#717220000000
1!
0$
b1000 %
1'
0*
b1000 +
#717230000000
0!
0'
#717240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#717250000000
0!
0'
#717260000000
1!
b0 %
1'
b0 +
#717270000000
0!
0'
#717280000000
1!
1$
b1 %
1'
1*
b1 +
#717290000000
0!
0'
#717300000000
1!
b10 %
1'
b10 +
#717310000000
0!
0'
#717320000000
1!
b11 %
1'
b11 +
#717330000000
0!
0'
#717340000000
1!
b100 %
1'
b100 +
#717350000000
0!
0'
#717360000000
1!
b101 %
1'
b101 +
#717370000000
0!
0'
#717380000000
1!
0$
b110 %
1'
0*
b110 +
#717390000000
0!
0'
#717400000000
1!
b111 %
1'
b111 +
#717410000000
0!
0'
#717420000000
1!
b1000 %
1'
b1000 +
#717430000000
0!
0'
#717440000000
1!
b1001 %
1'
b1001 +
#717450000000
1"
1(
#717460000000
0!
0"
b100 &
0'
0(
b100 ,
#717470000000
1!
b0 %
1'
b0 +
#717480000000
0!
0'
#717490000000
1!
1$
b1 %
1'
1*
b1 +
#717500000000
0!
0'
#717510000000
1!
b10 %
1'
b10 +
#717520000000
0!
0'
#717530000000
1!
b11 %
1'
b11 +
#717540000000
0!
0'
#717550000000
1!
b100 %
1'
b100 +
#717560000000
0!
0'
#717570000000
1!
b101 %
1'
b101 +
#717580000000
0!
0'
#717590000000
1!
b110 %
1'
b110 +
#717600000000
0!
0'
#717610000000
1!
b111 %
1'
b111 +
#717620000000
0!
0'
#717630000000
1!
0$
b1000 %
1'
0*
b1000 +
#717640000000
0!
0'
#717650000000
1!
b1001 %
1'
b1001 +
#717660000000
0!
0'
#717670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#717680000000
0!
0'
#717690000000
1!
1$
b1 %
1'
1*
b1 +
#717700000000
0!
0'
#717710000000
1!
b10 %
1'
b10 +
#717720000000
0!
0'
#717730000000
1!
b11 %
1'
b11 +
#717740000000
0!
0'
#717750000000
1!
b100 %
1'
b100 +
#717760000000
0!
0'
#717770000000
1!
b101 %
1'
b101 +
#717780000000
0!
0'
#717790000000
1!
0$
b110 %
1'
0*
b110 +
#717800000000
0!
0'
#717810000000
1!
b111 %
1'
b111 +
#717820000000
0!
0'
#717830000000
1!
b1000 %
1'
b1000 +
#717840000000
0!
0'
#717850000000
1!
b1001 %
1'
b1001 +
#717860000000
0!
0'
#717870000000
1!
b0 %
1'
b0 +
#717880000000
1"
1(
#717890000000
0!
0"
b100 &
0'
0(
b100 ,
#717900000000
1!
1$
b1 %
1'
1*
b1 +
#717910000000
0!
0'
#717920000000
1!
b10 %
1'
b10 +
#717930000000
0!
0'
#717940000000
1!
b11 %
1'
b11 +
#717950000000
0!
0'
#717960000000
1!
b100 %
1'
b100 +
#717970000000
0!
0'
#717980000000
1!
b101 %
1'
b101 +
#717990000000
0!
0'
#718000000000
1!
b110 %
1'
b110 +
#718010000000
0!
0'
#718020000000
1!
b111 %
1'
b111 +
#718030000000
0!
0'
#718040000000
1!
0$
b1000 %
1'
0*
b1000 +
#718050000000
0!
0'
#718060000000
1!
b1001 %
1'
b1001 +
#718070000000
0!
0'
#718080000000
1!
b0 %
1'
b0 +
#718090000000
0!
0'
#718100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#718110000000
0!
0'
#718120000000
1!
b10 %
1'
b10 +
#718130000000
0!
0'
#718140000000
1!
b11 %
1'
b11 +
#718150000000
0!
0'
#718160000000
1!
b100 %
1'
b100 +
#718170000000
0!
0'
#718180000000
1!
b101 %
1'
b101 +
#718190000000
0!
0'
#718200000000
1!
0$
b110 %
1'
0*
b110 +
#718210000000
0!
0'
#718220000000
1!
b111 %
1'
b111 +
#718230000000
0!
0'
#718240000000
1!
b1000 %
1'
b1000 +
#718250000000
0!
0'
#718260000000
1!
b1001 %
1'
b1001 +
#718270000000
0!
0'
#718280000000
1!
b0 %
1'
b0 +
#718290000000
0!
0'
#718300000000
1!
1$
b1 %
1'
1*
b1 +
#718310000000
1"
1(
#718320000000
0!
0"
b100 &
0'
0(
b100 ,
#718330000000
1!
b10 %
1'
b10 +
#718340000000
0!
0'
#718350000000
1!
b11 %
1'
b11 +
#718360000000
0!
0'
#718370000000
1!
b100 %
1'
b100 +
#718380000000
0!
0'
#718390000000
1!
b101 %
1'
b101 +
#718400000000
0!
0'
#718410000000
1!
b110 %
1'
b110 +
#718420000000
0!
0'
#718430000000
1!
b111 %
1'
b111 +
#718440000000
0!
0'
#718450000000
1!
0$
b1000 %
1'
0*
b1000 +
#718460000000
0!
0'
#718470000000
1!
b1001 %
1'
b1001 +
#718480000000
0!
0'
#718490000000
1!
b0 %
1'
b0 +
#718500000000
0!
0'
#718510000000
1!
1$
b1 %
1'
1*
b1 +
#718520000000
0!
0'
#718530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#718540000000
0!
0'
#718550000000
1!
b11 %
1'
b11 +
#718560000000
0!
0'
#718570000000
1!
b100 %
1'
b100 +
#718580000000
0!
0'
#718590000000
1!
b101 %
1'
b101 +
#718600000000
0!
0'
#718610000000
1!
0$
b110 %
1'
0*
b110 +
#718620000000
0!
0'
#718630000000
1!
b111 %
1'
b111 +
#718640000000
0!
0'
#718650000000
1!
b1000 %
1'
b1000 +
#718660000000
0!
0'
#718670000000
1!
b1001 %
1'
b1001 +
#718680000000
0!
0'
#718690000000
1!
b0 %
1'
b0 +
#718700000000
0!
0'
#718710000000
1!
1$
b1 %
1'
1*
b1 +
#718720000000
0!
0'
#718730000000
1!
b10 %
1'
b10 +
#718740000000
1"
1(
#718750000000
0!
0"
b100 &
0'
0(
b100 ,
#718760000000
1!
b11 %
1'
b11 +
#718770000000
0!
0'
#718780000000
1!
b100 %
1'
b100 +
#718790000000
0!
0'
#718800000000
1!
b101 %
1'
b101 +
#718810000000
0!
0'
#718820000000
1!
b110 %
1'
b110 +
#718830000000
0!
0'
#718840000000
1!
b111 %
1'
b111 +
#718850000000
0!
0'
#718860000000
1!
0$
b1000 %
1'
0*
b1000 +
#718870000000
0!
0'
#718880000000
1!
b1001 %
1'
b1001 +
#718890000000
0!
0'
#718900000000
1!
b0 %
1'
b0 +
#718910000000
0!
0'
#718920000000
1!
1$
b1 %
1'
1*
b1 +
#718930000000
0!
0'
#718940000000
1!
b10 %
1'
b10 +
#718950000000
0!
0'
#718960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#718970000000
0!
0'
#718980000000
1!
b100 %
1'
b100 +
#718990000000
0!
0'
#719000000000
1!
b101 %
1'
b101 +
#719010000000
0!
0'
#719020000000
1!
0$
b110 %
1'
0*
b110 +
#719030000000
0!
0'
#719040000000
1!
b111 %
1'
b111 +
#719050000000
0!
0'
#719060000000
1!
b1000 %
1'
b1000 +
#719070000000
0!
0'
#719080000000
1!
b1001 %
1'
b1001 +
#719090000000
0!
0'
#719100000000
1!
b0 %
1'
b0 +
#719110000000
0!
0'
#719120000000
1!
1$
b1 %
1'
1*
b1 +
#719130000000
0!
0'
#719140000000
1!
b10 %
1'
b10 +
#719150000000
0!
0'
#719160000000
1!
b11 %
1'
b11 +
#719170000000
1"
1(
#719180000000
0!
0"
b100 &
0'
0(
b100 ,
#719190000000
1!
b100 %
1'
b100 +
#719200000000
0!
0'
#719210000000
1!
b101 %
1'
b101 +
#719220000000
0!
0'
#719230000000
1!
b110 %
1'
b110 +
#719240000000
0!
0'
#719250000000
1!
b111 %
1'
b111 +
#719260000000
0!
0'
#719270000000
1!
0$
b1000 %
1'
0*
b1000 +
#719280000000
0!
0'
#719290000000
1!
b1001 %
1'
b1001 +
#719300000000
0!
0'
#719310000000
1!
b0 %
1'
b0 +
#719320000000
0!
0'
#719330000000
1!
1$
b1 %
1'
1*
b1 +
#719340000000
0!
0'
#719350000000
1!
b10 %
1'
b10 +
#719360000000
0!
0'
#719370000000
1!
b11 %
1'
b11 +
#719380000000
0!
0'
#719390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#719400000000
0!
0'
#719410000000
1!
b101 %
1'
b101 +
#719420000000
0!
0'
#719430000000
1!
0$
b110 %
1'
0*
b110 +
#719440000000
0!
0'
#719450000000
1!
b111 %
1'
b111 +
#719460000000
0!
0'
#719470000000
1!
b1000 %
1'
b1000 +
#719480000000
0!
0'
#719490000000
1!
b1001 %
1'
b1001 +
#719500000000
0!
0'
#719510000000
1!
b0 %
1'
b0 +
#719520000000
0!
0'
#719530000000
1!
1$
b1 %
1'
1*
b1 +
#719540000000
0!
0'
#719550000000
1!
b10 %
1'
b10 +
#719560000000
0!
0'
#719570000000
1!
b11 %
1'
b11 +
#719580000000
0!
0'
#719590000000
1!
b100 %
1'
b100 +
#719600000000
1"
1(
#719610000000
0!
0"
b100 &
0'
0(
b100 ,
#719620000000
1!
b101 %
1'
b101 +
#719630000000
0!
0'
#719640000000
1!
b110 %
1'
b110 +
#719650000000
0!
0'
#719660000000
1!
b111 %
1'
b111 +
#719670000000
0!
0'
#719680000000
1!
0$
b1000 %
1'
0*
b1000 +
#719690000000
0!
0'
#719700000000
1!
b1001 %
1'
b1001 +
#719710000000
0!
0'
#719720000000
1!
b0 %
1'
b0 +
#719730000000
0!
0'
#719740000000
1!
1$
b1 %
1'
1*
b1 +
#719750000000
0!
0'
#719760000000
1!
b10 %
1'
b10 +
#719770000000
0!
0'
#719780000000
1!
b11 %
1'
b11 +
#719790000000
0!
0'
#719800000000
1!
b100 %
1'
b100 +
#719810000000
0!
0'
#719820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#719830000000
0!
0'
#719840000000
1!
0$
b110 %
1'
0*
b110 +
#719850000000
0!
0'
#719860000000
1!
b111 %
1'
b111 +
#719870000000
0!
0'
#719880000000
1!
b1000 %
1'
b1000 +
#719890000000
0!
0'
#719900000000
1!
b1001 %
1'
b1001 +
#719910000000
0!
0'
#719920000000
1!
b0 %
1'
b0 +
#719930000000
0!
0'
#719940000000
1!
1$
b1 %
1'
1*
b1 +
#719950000000
0!
0'
#719960000000
1!
b10 %
1'
b10 +
#719970000000
0!
0'
#719980000000
1!
b11 %
1'
b11 +
#719990000000
0!
0'
#720000000000
1!
b100 %
1'
b100 +
#720010000000
0!
0'
#720020000000
1!
b101 %
1'
b101 +
#720030000000
1"
1(
#720040000000
0!
0"
b100 &
0'
0(
b100 ,
#720050000000
1!
b110 %
1'
b110 +
#720060000000
0!
0'
#720070000000
1!
b111 %
1'
b111 +
#720080000000
0!
0'
#720090000000
1!
0$
b1000 %
1'
0*
b1000 +
#720100000000
0!
0'
#720110000000
1!
b1001 %
1'
b1001 +
#720120000000
0!
0'
#720130000000
1!
b0 %
1'
b0 +
#720140000000
0!
0'
#720150000000
1!
1$
b1 %
1'
1*
b1 +
#720160000000
0!
0'
#720170000000
1!
b10 %
1'
b10 +
#720180000000
0!
0'
#720190000000
1!
b11 %
1'
b11 +
#720200000000
0!
0'
#720210000000
1!
b100 %
1'
b100 +
#720220000000
0!
0'
#720230000000
1!
b101 %
1'
b101 +
#720240000000
0!
0'
#720250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#720260000000
0!
0'
#720270000000
1!
b111 %
1'
b111 +
#720280000000
0!
0'
#720290000000
1!
b1000 %
1'
b1000 +
#720300000000
0!
0'
#720310000000
1!
b1001 %
1'
b1001 +
#720320000000
0!
0'
#720330000000
1!
b0 %
1'
b0 +
#720340000000
0!
0'
#720350000000
1!
1$
b1 %
1'
1*
b1 +
#720360000000
0!
0'
#720370000000
1!
b10 %
1'
b10 +
#720380000000
0!
0'
#720390000000
1!
b11 %
1'
b11 +
#720400000000
0!
0'
#720410000000
1!
b100 %
1'
b100 +
#720420000000
0!
0'
#720430000000
1!
b101 %
1'
b101 +
#720440000000
0!
0'
#720450000000
1!
0$
b110 %
1'
0*
b110 +
#720460000000
1"
1(
#720470000000
0!
0"
b100 &
0'
0(
b100 ,
#720480000000
1!
1$
b111 %
1'
1*
b111 +
#720490000000
0!
0'
#720500000000
1!
0$
b1000 %
1'
0*
b1000 +
#720510000000
0!
0'
#720520000000
1!
b1001 %
1'
b1001 +
#720530000000
0!
0'
#720540000000
1!
b0 %
1'
b0 +
#720550000000
0!
0'
#720560000000
1!
1$
b1 %
1'
1*
b1 +
#720570000000
0!
0'
#720580000000
1!
b10 %
1'
b10 +
#720590000000
0!
0'
#720600000000
1!
b11 %
1'
b11 +
#720610000000
0!
0'
#720620000000
1!
b100 %
1'
b100 +
#720630000000
0!
0'
#720640000000
1!
b101 %
1'
b101 +
#720650000000
0!
0'
#720660000000
1!
b110 %
1'
b110 +
#720670000000
0!
0'
#720680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#720690000000
0!
0'
#720700000000
1!
b1000 %
1'
b1000 +
#720710000000
0!
0'
#720720000000
1!
b1001 %
1'
b1001 +
#720730000000
0!
0'
#720740000000
1!
b0 %
1'
b0 +
#720750000000
0!
0'
#720760000000
1!
1$
b1 %
1'
1*
b1 +
#720770000000
0!
0'
#720780000000
1!
b10 %
1'
b10 +
#720790000000
0!
0'
#720800000000
1!
b11 %
1'
b11 +
#720810000000
0!
0'
#720820000000
1!
b100 %
1'
b100 +
#720830000000
0!
0'
#720840000000
1!
b101 %
1'
b101 +
#720850000000
0!
0'
#720860000000
1!
0$
b110 %
1'
0*
b110 +
#720870000000
0!
0'
#720880000000
1!
b111 %
1'
b111 +
#720890000000
1"
1(
#720900000000
0!
0"
b100 &
0'
0(
b100 ,
#720910000000
1!
b1000 %
1'
b1000 +
#720920000000
0!
0'
#720930000000
1!
b1001 %
1'
b1001 +
#720940000000
0!
0'
#720950000000
1!
b0 %
1'
b0 +
#720960000000
0!
0'
#720970000000
1!
1$
b1 %
1'
1*
b1 +
#720980000000
0!
0'
#720990000000
1!
b10 %
1'
b10 +
#721000000000
0!
0'
#721010000000
1!
b11 %
1'
b11 +
#721020000000
0!
0'
#721030000000
1!
b100 %
1'
b100 +
#721040000000
0!
0'
#721050000000
1!
b101 %
1'
b101 +
#721060000000
0!
0'
#721070000000
1!
b110 %
1'
b110 +
#721080000000
0!
0'
#721090000000
1!
b111 %
1'
b111 +
#721100000000
0!
0'
#721110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#721120000000
0!
0'
#721130000000
1!
b1001 %
1'
b1001 +
#721140000000
0!
0'
#721150000000
1!
b0 %
1'
b0 +
#721160000000
0!
0'
#721170000000
1!
1$
b1 %
1'
1*
b1 +
#721180000000
0!
0'
#721190000000
1!
b10 %
1'
b10 +
#721200000000
0!
0'
#721210000000
1!
b11 %
1'
b11 +
#721220000000
0!
0'
#721230000000
1!
b100 %
1'
b100 +
#721240000000
0!
0'
#721250000000
1!
b101 %
1'
b101 +
#721260000000
0!
0'
#721270000000
1!
0$
b110 %
1'
0*
b110 +
#721280000000
0!
0'
#721290000000
1!
b111 %
1'
b111 +
#721300000000
0!
0'
#721310000000
1!
b1000 %
1'
b1000 +
#721320000000
1"
1(
#721330000000
0!
0"
b100 &
0'
0(
b100 ,
#721340000000
1!
b1001 %
1'
b1001 +
#721350000000
0!
0'
#721360000000
1!
b0 %
1'
b0 +
#721370000000
0!
0'
#721380000000
1!
1$
b1 %
1'
1*
b1 +
#721390000000
0!
0'
#721400000000
1!
b10 %
1'
b10 +
#721410000000
0!
0'
#721420000000
1!
b11 %
1'
b11 +
#721430000000
0!
0'
#721440000000
1!
b100 %
1'
b100 +
#721450000000
0!
0'
#721460000000
1!
b101 %
1'
b101 +
#721470000000
0!
0'
#721480000000
1!
b110 %
1'
b110 +
#721490000000
0!
0'
#721500000000
1!
b111 %
1'
b111 +
#721510000000
0!
0'
#721520000000
1!
0$
b1000 %
1'
0*
b1000 +
#721530000000
0!
0'
#721540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#721550000000
0!
0'
#721560000000
1!
b0 %
1'
b0 +
#721570000000
0!
0'
#721580000000
1!
1$
b1 %
1'
1*
b1 +
#721590000000
0!
0'
#721600000000
1!
b10 %
1'
b10 +
#721610000000
0!
0'
#721620000000
1!
b11 %
1'
b11 +
#721630000000
0!
0'
#721640000000
1!
b100 %
1'
b100 +
#721650000000
0!
0'
#721660000000
1!
b101 %
1'
b101 +
#721670000000
0!
0'
#721680000000
1!
0$
b110 %
1'
0*
b110 +
#721690000000
0!
0'
#721700000000
1!
b111 %
1'
b111 +
#721710000000
0!
0'
#721720000000
1!
b1000 %
1'
b1000 +
#721730000000
0!
0'
#721740000000
1!
b1001 %
1'
b1001 +
#721750000000
1"
1(
#721760000000
0!
0"
b100 &
0'
0(
b100 ,
#721770000000
1!
b0 %
1'
b0 +
#721780000000
0!
0'
#721790000000
1!
1$
b1 %
1'
1*
b1 +
#721800000000
0!
0'
#721810000000
1!
b10 %
1'
b10 +
#721820000000
0!
0'
#721830000000
1!
b11 %
1'
b11 +
#721840000000
0!
0'
#721850000000
1!
b100 %
1'
b100 +
#721860000000
0!
0'
#721870000000
1!
b101 %
1'
b101 +
#721880000000
0!
0'
#721890000000
1!
b110 %
1'
b110 +
#721900000000
0!
0'
#721910000000
1!
b111 %
1'
b111 +
#721920000000
0!
0'
#721930000000
1!
0$
b1000 %
1'
0*
b1000 +
#721940000000
0!
0'
#721950000000
1!
b1001 %
1'
b1001 +
#721960000000
0!
0'
#721970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#721980000000
0!
0'
#721990000000
1!
1$
b1 %
1'
1*
b1 +
#722000000000
0!
0'
#722010000000
1!
b10 %
1'
b10 +
#722020000000
0!
0'
#722030000000
1!
b11 %
1'
b11 +
#722040000000
0!
0'
#722050000000
1!
b100 %
1'
b100 +
#722060000000
0!
0'
#722070000000
1!
b101 %
1'
b101 +
#722080000000
0!
0'
#722090000000
1!
0$
b110 %
1'
0*
b110 +
#722100000000
0!
0'
#722110000000
1!
b111 %
1'
b111 +
#722120000000
0!
0'
#722130000000
1!
b1000 %
1'
b1000 +
#722140000000
0!
0'
#722150000000
1!
b1001 %
1'
b1001 +
#722160000000
0!
0'
#722170000000
1!
b0 %
1'
b0 +
#722180000000
1"
1(
#722190000000
0!
0"
b100 &
0'
0(
b100 ,
#722200000000
1!
1$
b1 %
1'
1*
b1 +
#722210000000
0!
0'
#722220000000
1!
b10 %
1'
b10 +
#722230000000
0!
0'
#722240000000
1!
b11 %
1'
b11 +
#722250000000
0!
0'
#722260000000
1!
b100 %
1'
b100 +
#722270000000
0!
0'
#722280000000
1!
b101 %
1'
b101 +
#722290000000
0!
0'
#722300000000
1!
b110 %
1'
b110 +
#722310000000
0!
0'
#722320000000
1!
b111 %
1'
b111 +
#722330000000
0!
0'
#722340000000
1!
0$
b1000 %
1'
0*
b1000 +
#722350000000
0!
0'
#722360000000
1!
b1001 %
1'
b1001 +
#722370000000
0!
0'
#722380000000
1!
b0 %
1'
b0 +
#722390000000
0!
0'
#722400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#722410000000
0!
0'
#722420000000
1!
b10 %
1'
b10 +
#722430000000
0!
0'
#722440000000
1!
b11 %
1'
b11 +
#722450000000
0!
0'
#722460000000
1!
b100 %
1'
b100 +
#722470000000
0!
0'
#722480000000
1!
b101 %
1'
b101 +
#722490000000
0!
0'
#722500000000
1!
0$
b110 %
1'
0*
b110 +
#722510000000
0!
0'
#722520000000
1!
b111 %
1'
b111 +
#722530000000
0!
0'
#722540000000
1!
b1000 %
1'
b1000 +
#722550000000
0!
0'
#722560000000
1!
b1001 %
1'
b1001 +
#722570000000
0!
0'
#722580000000
1!
b0 %
1'
b0 +
#722590000000
0!
0'
#722600000000
1!
1$
b1 %
1'
1*
b1 +
#722610000000
1"
1(
#722620000000
0!
0"
b100 &
0'
0(
b100 ,
#722630000000
1!
b10 %
1'
b10 +
#722640000000
0!
0'
#722650000000
1!
b11 %
1'
b11 +
#722660000000
0!
0'
#722670000000
1!
b100 %
1'
b100 +
#722680000000
0!
0'
#722690000000
1!
b101 %
1'
b101 +
#722700000000
0!
0'
#722710000000
1!
b110 %
1'
b110 +
#722720000000
0!
0'
#722730000000
1!
b111 %
1'
b111 +
#722740000000
0!
0'
#722750000000
1!
0$
b1000 %
1'
0*
b1000 +
#722760000000
0!
0'
#722770000000
1!
b1001 %
1'
b1001 +
#722780000000
0!
0'
#722790000000
1!
b0 %
1'
b0 +
#722800000000
0!
0'
#722810000000
1!
1$
b1 %
1'
1*
b1 +
#722820000000
0!
0'
#722830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#722840000000
0!
0'
#722850000000
1!
b11 %
1'
b11 +
#722860000000
0!
0'
#722870000000
1!
b100 %
1'
b100 +
#722880000000
0!
0'
#722890000000
1!
b101 %
1'
b101 +
#722900000000
0!
0'
#722910000000
1!
0$
b110 %
1'
0*
b110 +
#722920000000
0!
0'
#722930000000
1!
b111 %
1'
b111 +
#722940000000
0!
0'
#722950000000
1!
b1000 %
1'
b1000 +
#722960000000
0!
0'
#722970000000
1!
b1001 %
1'
b1001 +
#722980000000
0!
0'
#722990000000
1!
b0 %
1'
b0 +
#723000000000
0!
0'
#723010000000
1!
1$
b1 %
1'
1*
b1 +
#723020000000
0!
0'
#723030000000
1!
b10 %
1'
b10 +
#723040000000
1"
1(
#723050000000
0!
0"
b100 &
0'
0(
b100 ,
#723060000000
1!
b11 %
1'
b11 +
#723070000000
0!
0'
#723080000000
1!
b100 %
1'
b100 +
#723090000000
0!
0'
#723100000000
1!
b101 %
1'
b101 +
#723110000000
0!
0'
#723120000000
1!
b110 %
1'
b110 +
#723130000000
0!
0'
#723140000000
1!
b111 %
1'
b111 +
#723150000000
0!
0'
#723160000000
1!
0$
b1000 %
1'
0*
b1000 +
#723170000000
0!
0'
#723180000000
1!
b1001 %
1'
b1001 +
#723190000000
0!
0'
#723200000000
1!
b0 %
1'
b0 +
#723210000000
0!
0'
#723220000000
1!
1$
b1 %
1'
1*
b1 +
#723230000000
0!
0'
#723240000000
1!
b10 %
1'
b10 +
#723250000000
0!
0'
#723260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#723270000000
0!
0'
#723280000000
1!
b100 %
1'
b100 +
#723290000000
0!
0'
#723300000000
1!
b101 %
1'
b101 +
#723310000000
0!
0'
#723320000000
1!
0$
b110 %
1'
0*
b110 +
#723330000000
0!
0'
#723340000000
1!
b111 %
1'
b111 +
#723350000000
0!
0'
#723360000000
1!
b1000 %
1'
b1000 +
#723370000000
0!
0'
#723380000000
1!
b1001 %
1'
b1001 +
#723390000000
0!
0'
#723400000000
1!
b0 %
1'
b0 +
#723410000000
0!
0'
#723420000000
1!
1$
b1 %
1'
1*
b1 +
#723430000000
0!
0'
#723440000000
1!
b10 %
1'
b10 +
#723450000000
0!
0'
#723460000000
1!
b11 %
1'
b11 +
#723470000000
1"
1(
#723480000000
0!
0"
b100 &
0'
0(
b100 ,
#723490000000
1!
b100 %
1'
b100 +
#723500000000
0!
0'
#723510000000
1!
b101 %
1'
b101 +
#723520000000
0!
0'
#723530000000
1!
b110 %
1'
b110 +
#723540000000
0!
0'
#723550000000
1!
b111 %
1'
b111 +
#723560000000
0!
0'
#723570000000
1!
0$
b1000 %
1'
0*
b1000 +
#723580000000
0!
0'
#723590000000
1!
b1001 %
1'
b1001 +
#723600000000
0!
0'
#723610000000
1!
b0 %
1'
b0 +
#723620000000
0!
0'
#723630000000
1!
1$
b1 %
1'
1*
b1 +
#723640000000
0!
0'
#723650000000
1!
b10 %
1'
b10 +
#723660000000
0!
0'
#723670000000
1!
b11 %
1'
b11 +
#723680000000
0!
0'
#723690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#723700000000
0!
0'
#723710000000
1!
b101 %
1'
b101 +
#723720000000
0!
0'
#723730000000
1!
0$
b110 %
1'
0*
b110 +
#723740000000
0!
0'
#723750000000
1!
b111 %
1'
b111 +
#723760000000
0!
0'
#723770000000
1!
b1000 %
1'
b1000 +
#723780000000
0!
0'
#723790000000
1!
b1001 %
1'
b1001 +
#723800000000
0!
0'
#723810000000
1!
b0 %
1'
b0 +
#723820000000
0!
0'
#723830000000
1!
1$
b1 %
1'
1*
b1 +
#723840000000
0!
0'
#723850000000
1!
b10 %
1'
b10 +
#723860000000
0!
0'
#723870000000
1!
b11 %
1'
b11 +
#723880000000
0!
0'
#723890000000
1!
b100 %
1'
b100 +
#723900000000
1"
1(
#723910000000
0!
0"
b100 &
0'
0(
b100 ,
#723920000000
1!
b101 %
1'
b101 +
#723930000000
0!
0'
#723940000000
1!
b110 %
1'
b110 +
#723950000000
0!
0'
#723960000000
1!
b111 %
1'
b111 +
#723970000000
0!
0'
#723980000000
1!
0$
b1000 %
1'
0*
b1000 +
#723990000000
0!
0'
#724000000000
1!
b1001 %
1'
b1001 +
#724010000000
0!
0'
#724020000000
1!
b0 %
1'
b0 +
#724030000000
0!
0'
#724040000000
1!
1$
b1 %
1'
1*
b1 +
#724050000000
0!
0'
#724060000000
1!
b10 %
1'
b10 +
#724070000000
0!
0'
#724080000000
1!
b11 %
1'
b11 +
#724090000000
0!
0'
#724100000000
1!
b100 %
1'
b100 +
#724110000000
0!
0'
#724120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#724130000000
0!
0'
#724140000000
1!
0$
b110 %
1'
0*
b110 +
#724150000000
0!
0'
#724160000000
1!
b111 %
1'
b111 +
#724170000000
0!
0'
#724180000000
1!
b1000 %
1'
b1000 +
#724190000000
0!
0'
#724200000000
1!
b1001 %
1'
b1001 +
#724210000000
0!
0'
#724220000000
1!
b0 %
1'
b0 +
#724230000000
0!
0'
#724240000000
1!
1$
b1 %
1'
1*
b1 +
#724250000000
0!
0'
#724260000000
1!
b10 %
1'
b10 +
#724270000000
0!
0'
#724280000000
1!
b11 %
1'
b11 +
#724290000000
0!
0'
#724300000000
1!
b100 %
1'
b100 +
#724310000000
0!
0'
#724320000000
1!
b101 %
1'
b101 +
#724330000000
1"
1(
#724340000000
0!
0"
b100 &
0'
0(
b100 ,
#724350000000
1!
b110 %
1'
b110 +
#724360000000
0!
0'
#724370000000
1!
b111 %
1'
b111 +
#724380000000
0!
0'
#724390000000
1!
0$
b1000 %
1'
0*
b1000 +
#724400000000
0!
0'
#724410000000
1!
b1001 %
1'
b1001 +
#724420000000
0!
0'
#724430000000
1!
b0 %
1'
b0 +
#724440000000
0!
0'
#724450000000
1!
1$
b1 %
1'
1*
b1 +
#724460000000
0!
0'
#724470000000
1!
b10 %
1'
b10 +
#724480000000
0!
0'
#724490000000
1!
b11 %
1'
b11 +
#724500000000
0!
0'
#724510000000
1!
b100 %
1'
b100 +
#724520000000
0!
0'
#724530000000
1!
b101 %
1'
b101 +
#724540000000
0!
0'
#724550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#724560000000
0!
0'
#724570000000
1!
b111 %
1'
b111 +
#724580000000
0!
0'
#724590000000
1!
b1000 %
1'
b1000 +
#724600000000
0!
0'
#724610000000
1!
b1001 %
1'
b1001 +
#724620000000
0!
0'
#724630000000
1!
b0 %
1'
b0 +
#724640000000
0!
0'
#724650000000
1!
1$
b1 %
1'
1*
b1 +
#724660000000
0!
0'
#724670000000
1!
b10 %
1'
b10 +
#724680000000
0!
0'
#724690000000
1!
b11 %
1'
b11 +
#724700000000
0!
0'
#724710000000
1!
b100 %
1'
b100 +
#724720000000
0!
0'
#724730000000
1!
b101 %
1'
b101 +
#724740000000
0!
0'
#724750000000
1!
0$
b110 %
1'
0*
b110 +
#724760000000
1"
1(
#724770000000
0!
0"
b100 &
0'
0(
b100 ,
#724780000000
1!
1$
b111 %
1'
1*
b111 +
#724790000000
0!
0'
#724800000000
1!
0$
b1000 %
1'
0*
b1000 +
#724810000000
0!
0'
#724820000000
1!
b1001 %
1'
b1001 +
#724830000000
0!
0'
#724840000000
1!
b0 %
1'
b0 +
#724850000000
0!
0'
#724860000000
1!
1$
b1 %
1'
1*
b1 +
#724870000000
0!
0'
#724880000000
1!
b10 %
1'
b10 +
#724890000000
0!
0'
#724900000000
1!
b11 %
1'
b11 +
#724910000000
0!
0'
#724920000000
1!
b100 %
1'
b100 +
#724930000000
0!
0'
#724940000000
1!
b101 %
1'
b101 +
#724950000000
0!
0'
#724960000000
1!
b110 %
1'
b110 +
#724970000000
0!
0'
#724980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#724990000000
0!
0'
#725000000000
1!
b1000 %
1'
b1000 +
#725010000000
0!
0'
#725020000000
1!
b1001 %
1'
b1001 +
#725030000000
0!
0'
#725040000000
1!
b0 %
1'
b0 +
#725050000000
0!
0'
#725060000000
1!
1$
b1 %
1'
1*
b1 +
#725070000000
0!
0'
#725080000000
1!
b10 %
1'
b10 +
#725090000000
0!
0'
#725100000000
1!
b11 %
1'
b11 +
#725110000000
0!
0'
#725120000000
1!
b100 %
1'
b100 +
#725130000000
0!
0'
#725140000000
1!
b101 %
1'
b101 +
#725150000000
0!
0'
#725160000000
1!
0$
b110 %
1'
0*
b110 +
#725170000000
0!
0'
#725180000000
1!
b111 %
1'
b111 +
#725190000000
1"
1(
#725200000000
0!
0"
b100 &
0'
0(
b100 ,
#725210000000
1!
b1000 %
1'
b1000 +
#725220000000
0!
0'
#725230000000
1!
b1001 %
1'
b1001 +
#725240000000
0!
0'
#725250000000
1!
b0 %
1'
b0 +
#725260000000
0!
0'
#725270000000
1!
1$
b1 %
1'
1*
b1 +
#725280000000
0!
0'
#725290000000
1!
b10 %
1'
b10 +
#725300000000
0!
0'
#725310000000
1!
b11 %
1'
b11 +
#725320000000
0!
0'
#725330000000
1!
b100 %
1'
b100 +
#725340000000
0!
0'
#725350000000
1!
b101 %
1'
b101 +
#725360000000
0!
0'
#725370000000
1!
b110 %
1'
b110 +
#725380000000
0!
0'
#725390000000
1!
b111 %
1'
b111 +
#725400000000
0!
0'
#725410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#725420000000
0!
0'
#725430000000
1!
b1001 %
1'
b1001 +
#725440000000
0!
0'
#725450000000
1!
b0 %
1'
b0 +
#725460000000
0!
0'
#725470000000
1!
1$
b1 %
1'
1*
b1 +
#725480000000
0!
0'
#725490000000
1!
b10 %
1'
b10 +
#725500000000
0!
0'
#725510000000
1!
b11 %
1'
b11 +
#725520000000
0!
0'
#725530000000
1!
b100 %
1'
b100 +
#725540000000
0!
0'
#725550000000
1!
b101 %
1'
b101 +
#725560000000
0!
0'
#725570000000
1!
0$
b110 %
1'
0*
b110 +
#725580000000
0!
0'
#725590000000
1!
b111 %
1'
b111 +
#725600000000
0!
0'
#725610000000
1!
b1000 %
1'
b1000 +
#725620000000
1"
1(
#725630000000
0!
0"
b100 &
0'
0(
b100 ,
#725640000000
1!
b1001 %
1'
b1001 +
#725650000000
0!
0'
#725660000000
1!
b0 %
1'
b0 +
#725670000000
0!
0'
#725680000000
1!
1$
b1 %
1'
1*
b1 +
#725690000000
0!
0'
#725700000000
1!
b10 %
1'
b10 +
#725710000000
0!
0'
#725720000000
1!
b11 %
1'
b11 +
#725730000000
0!
0'
#725740000000
1!
b100 %
1'
b100 +
#725750000000
0!
0'
#725760000000
1!
b101 %
1'
b101 +
#725770000000
0!
0'
#725780000000
1!
b110 %
1'
b110 +
#725790000000
0!
0'
#725800000000
1!
b111 %
1'
b111 +
#725810000000
0!
0'
#725820000000
1!
0$
b1000 %
1'
0*
b1000 +
#725830000000
0!
0'
#725840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#725850000000
0!
0'
#725860000000
1!
b0 %
1'
b0 +
#725870000000
0!
0'
#725880000000
1!
1$
b1 %
1'
1*
b1 +
#725890000000
0!
0'
#725900000000
1!
b10 %
1'
b10 +
#725910000000
0!
0'
#725920000000
1!
b11 %
1'
b11 +
#725930000000
0!
0'
#725940000000
1!
b100 %
1'
b100 +
#725950000000
0!
0'
#725960000000
1!
b101 %
1'
b101 +
#725970000000
0!
0'
#725980000000
1!
0$
b110 %
1'
0*
b110 +
#725990000000
0!
0'
#726000000000
1!
b111 %
1'
b111 +
#726010000000
0!
0'
#726020000000
1!
b1000 %
1'
b1000 +
#726030000000
0!
0'
#726040000000
1!
b1001 %
1'
b1001 +
#726050000000
1"
1(
#726060000000
0!
0"
b100 &
0'
0(
b100 ,
#726070000000
1!
b0 %
1'
b0 +
#726080000000
0!
0'
#726090000000
1!
1$
b1 %
1'
1*
b1 +
#726100000000
0!
0'
#726110000000
1!
b10 %
1'
b10 +
#726120000000
0!
0'
#726130000000
1!
b11 %
1'
b11 +
#726140000000
0!
0'
#726150000000
1!
b100 %
1'
b100 +
#726160000000
0!
0'
#726170000000
1!
b101 %
1'
b101 +
#726180000000
0!
0'
#726190000000
1!
b110 %
1'
b110 +
#726200000000
0!
0'
#726210000000
1!
b111 %
1'
b111 +
#726220000000
0!
0'
#726230000000
1!
0$
b1000 %
1'
0*
b1000 +
#726240000000
0!
0'
#726250000000
1!
b1001 %
1'
b1001 +
#726260000000
0!
0'
#726270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#726280000000
0!
0'
#726290000000
1!
1$
b1 %
1'
1*
b1 +
#726300000000
0!
0'
#726310000000
1!
b10 %
1'
b10 +
#726320000000
0!
0'
#726330000000
1!
b11 %
1'
b11 +
#726340000000
0!
0'
#726350000000
1!
b100 %
1'
b100 +
#726360000000
0!
0'
#726370000000
1!
b101 %
1'
b101 +
#726380000000
0!
0'
#726390000000
1!
0$
b110 %
1'
0*
b110 +
#726400000000
0!
0'
#726410000000
1!
b111 %
1'
b111 +
#726420000000
0!
0'
#726430000000
1!
b1000 %
1'
b1000 +
#726440000000
0!
0'
#726450000000
1!
b1001 %
1'
b1001 +
#726460000000
0!
0'
#726470000000
1!
b0 %
1'
b0 +
#726480000000
1"
1(
#726490000000
0!
0"
b100 &
0'
0(
b100 ,
#726500000000
1!
1$
b1 %
1'
1*
b1 +
#726510000000
0!
0'
#726520000000
1!
b10 %
1'
b10 +
#726530000000
0!
0'
#726540000000
1!
b11 %
1'
b11 +
#726550000000
0!
0'
#726560000000
1!
b100 %
1'
b100 +
#726570000000
0!
0'
#726580000000
1!
b101 %
1'
b101 +
#726590000000
0!
0'
#726600000000
1!
b110 %
1'
b110 +
#726610000000
0!
0'
#726620000000
1!
b111 %
1'
b111 +
#726630000000
0!
0'
#726640000000
1!
0$
b1000 %
1'
0*
b1000 +
#726650000000
0!
0'
#726660000000
1!
b1001 %
1'
b1001 +
#726670000000
0!
0'
#726680000000
1!
b0 %
1'
b0 +
#726690000000
0!
0'
#726700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#726710000000
0!
0'
#726720000000
1!
b10 %
1'
b10 +
#726730000000
0!
0'
#726740000000
1!
b11 %
1'
b11 +
#726750000000
0!
0'
#726760000000
1!
b100 %
1'
b100 +
#726770000000
0!
0'
#726780000000
1!
b101 %
1'
b101 +
#726790000000
0!
0'
#726800000000
1!
0$
b110 %
1'
0*
b110 +
#726810000000
0!
0'
#726820000000
1!
b111 %
1'
b111 +
#726830000000
0!
0'
#726840000000
1!
b1000 %
1'
b1000 +
#726850000000
0!
0'
#726860000000
1!
b1001 %
1'
b1001 +
#726870000000
0!
0'
#726880000000
1!
b0 %
1'
b0 +
#726890000000
0!
0'
#726900000000
1!
1$
b1 %
1'
1*
b1 +
#726910000000
1"
1(
#726920000000
0!
0"
b100 &
0'
0(
b100 ,
#726930000000
1!
b10 %
1'
b10 +
#726940000000
0!
0'
#726950000000
1!
b11 %
1'
b11 +
#726960000000
0!
0'
#726970000000
1!
b100 %
1'
b100 +
#726980000000
0!
0'
#726990000000
1!
b101 %
1'
b101 +
#727000000000
0!
0'
#727010000000
1!
b110 %
1'
b110 +
#727020000000
0!
0'
#727030000000
1!
b111 %
1'
b111 +
#727040000000
0!
0'
#727050000000
1!
0$
b1000 %
1'
0*
b1000 +
#727060000000
0!
0'
#727070000000
1!
b1001 %
1'
b1001 +
#727080000000
0!
0'
#727090000000
1!
b0 %
1'
b0 +
#727100000000
0!
0'
#727110000000
1!
1$
b1 %
1'
1*
b1 +
#727120000000
0!
0'
#727130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#727140000000
0!
0'
#727150000000
1!
b11 %
1'
b11 +
#727160000000
0!
0'
#727170000000
1!
b100 %
1'
b100 +
#727180000000
0!
0'
#727190000000
1!
b101 %
1'
b101 +
#727200000000
0!
0'
#727210000000
1!
0$
b110 %
1'
0*
b110 +
#727220000000
0!
0'
#727230000000
1!
b111 %
1'
b111 +
#727240000000
0!
0'
#727250000000
1!
b1000 %
1'
b1000 +
#727260000000
0!
0'
#727270000000
1!
b1001 %
1'
b1001 +
#727280000000
0!
0'
#727290000000
1!
b0 %
1'
b0 +
#727300000000
0!
0'
#727310000000
1!
1$
b1 %
1'
1*
b1 +
#727320000000
0!
0'
#727330000000
1!
b10 %
1'
b10 +
#727340000000
1"
1(
#727350000000
0!
0"
b100 &
0'
0(
b100 ,
#727360000000
1!
b11 %
1'
b11 +
#727370000000
0!
0'
#727380000000
1!
b100 %
1'
b100 +
#727390000000
0!
0'
#727400000000
1!
b101 %
1'
b101 +
#727410000000
0!
0'
#727420000000
1!
b110 %
1'
b110 +
#727430000000
0!
0'
#727440000000
1!
b111 %
1'
b111 +
#727450000000
0!
0'
#727460000000
1!
0$
b1000 %
1'
0*
b1000 +
#727470000000
0!
0'
#727480000000
1!
b1001 %
1'
b1001 +
#727490000000
0!
0'
#727500000000
1!
b0 %
1'
b0 +
#727510000000
0!
0'
#727520000000
1!
1$
b1 %
1'
1*
b1 +
#727530000000
0!
0'
#727540000000
1!
b10 %
1'
b10 +
#727550000000
0!
0'
#727560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#727570000000
0!
0'
#727580000000
1!
b100 %
1'
b100 +
#727590000000
0!
0'
#727600000000
1!
b101 %
1'
b101 +
#727610000000
0!
0'
#727620000000
1!
0$
b110 %
1'
0*
b110 +
#727630000000
0!
0'
#727640000000
1!
b111 %
1'
b111 +
#727650000000
0!
0'
#727660000000
1!
b1000 %
1'
b1000 +
#727670000000
0!
0'
#727680000000
1!
b1001 %
1'
b1001 +
#727690000000
0!
0'
#727700000000
1!
b0 %
1'
b0 +
#727710000000
0!
0'
#727720000000
1!
1$
b1 %
1'
1*
b1 +
#727730000000
0!
0'
#727740000000
1!
b10 %
1'
b10 +
#727750000000
0!
0'
#727760000000
1!
b11 %
1'
b11 +
#727770000000
1"
1(
#727780000000
0!
0"
b100 &
0'
0(
b100 ,
#727790000000
1!
b100 %
1'
b100 +
#727800000000
0!
0'
#727810000000
1!
b101 %
1'
b101 +
#727820000000
0!
0'
#727830000000
1!
b110 %
1'
b110 +
#727840000000
0!
0'
#727850000000
1!
b111 %
1'
b111 +
#727860000000
0!
0'
#727870000000
1!
0$
b1000 %
1'
0*
b1000 +
#727880000000
0!
0'
#727890000000
1!
b1001 %
1'
b1001 +
#727900000000
0!
0'
#727910000000
1!
b0 %
1'
b0 +
#727920000000
0!
0'
#727930000000
1!
1$
b1 %
1'
1*
b1 +
#727940000000
0!
0'
#727950000000
1!
b10 %
1'
b10 +
#727960000000
0!
0'
#727970000000
1!
b11 %
1'
b11 +
#727980000000
0!
0'
#727990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#728000000000
0!
0'
#728010000000
1!
b101 %
1'
b101 +
#728020000000
0!
0'
#728030000000
1!
0$
b110 %
1'
0*
b110 +
#728040000000
0!
0'
#728050000000
1!
b111 %
1'
b111 +
#728060000000
0!
0'
#728070000000
1!
b1000 %
1'
b1000 +
#728080000000
0!
0'
#728090000000
1!
b1001 %
1'
b1001 +
#728100000000
0!
0'
#728110000000
1!
b0 %
1'
b0 +
#728120000000
0!
0'
#728130000000
1!
1$
b1 %
1'
1*
b1 +
#728140000000
0!
0'
#728150000000
1!
b10 %
1'
b10 +
#728160000000
0!
0'
#728170000000
1!
b11 %
1'
b11 +
#728180000000
0!
0'
#728190000000
1!
b100 %
1'
b100 +
#728200000000
1"
1(
#728210000000
0!
0"
b100 &
0'
0(
b100 ,
#728220000000
1!
b101 %
1'
b101 +
#728230000000
0!
0'
#728240000000
1!
b110 %
1'
b110 +
#728250000000
0!
0'
#728260000000
1!
b111 %
1'
b111 +
#728270000000
0!
0'
#728280000000
1!
0$
b1000 %
1'
0*
b1000 +
#728290000000
0!
0'
#728300000000
1!
b1001 %
1'
b1001 +
#728310000000
0!
0'
#728320000000
1!
b0 %
1'
b0 +
#728330000000
0!
0'
#728340000000
1!
1$
b1 %
1'
1*
b1 +
#728350000000
0!
0'
#728360000000
1!
b10 %
1'
b10 +
#728370000000
0!
0'
#728380000000
1!
b11 %
1'
b11 +
#728390000000
0!
0'
#728400000000
1!
b100 %
1'
b100 +
#728410000000
0!
0'
#728420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#728430000000
0!
0'
#728440000000
1!
0$
b110 %
1'
0*
b110 +
#728450000000
0!
0'
#728460000000
1!
b111 %
1'
b111 +
#728470000000
0!
0'
#728480000000
1!
b1000 %
1'
b1000 +
#728490000000
0!
0'
#728500000000
1!
b1001 %
1'
b1001 +
#728510000000
0!
0'
#728520000000
1!
b0 %
1'
b0 +
#728530000000
0!
0'
#728540000000
1!
1$
b1 %
1'
1*
b1 +
#728550000000
0!
0'
#728560000000
1!
b10 %
1'
b10 +
#728570000000
0!
0'
#728580000000
1!
b11 %
1'
b11 +
#728590000000
0!
0'
#728600000000
1!
b100 %
1'
b100 +
#728610000000
0!
0'
#728620000000
1!
b101 %
1'
b101 +
#728630000000
1"
1(
#728640000000
0!
0"
b100 &
0'
0(
b100 ,
#728650000000
1!
b110 %
1'
b110 +
#728660000000
0!
0'
#728670000000
1!
b111 %
1'
b111 +
#728680000000
0!
0'
#728690000000
1!
0$
b1000 %
1'
0*
b1000 +
#728700000000
0!
0'
#728710000000
1!
b1001 %
1'
b1001 +
#728720000000
0!
0'
#728730000000
1!
b0 %
1'
b0 +
#728740000000
0!
0'
#728750000000
1!
1$
b1 %
1'
1*
b1 +
#728760000000
0!
0'
#728770000000
1!
b10 %
1'
b10 +
#728780000000
0!
0'
#728790000000
1!
b11 %
1'
b11 +
#728800000000
0!
0'
#728810000000
1!
b100 %
1'
b100 +
#728820000000
0!
0'
#728830000000
1!
b101 %
1'
b101 +
#728840000000
0!
0'
#728850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#728860000000
0!
0'
#728870000000
1!
b111 %
1'
b111 +
#728880000000
0!
0'
#728890000000
1!
b1000 %
1'
b1000 +
#728900000000
0!
0'
#728910000000
1!
b1001 %
1'
b1001 +
#728920000000
0!
0'
#728930000000
1!
b0 %
1'
b0 +
#728940000000
0!
0'
#728950000000
1!
1$
b1 %
1'
1*
b1 +
#728960000000
0!
0'
#728970000000
1!
b10 %
1'
b10 +
#728980000000
0!
0'
#728990000000
1!
b11 %
1'
b11 +
#729000000000
0!
0'
#729010000000
1!
b100 %
1'
b100 +
#729020000000
0!
0'
#729030000000
1!
b101 %
1'
b101 +
#729040000000
0!
0'
#729050000000
1!
0$
b110 %
1'
0*
b110 +
#729060000000
1"
1(
#729070000000
0!
0"
b100 &
0'
0(
b100 ,
#729080000000
1!
1$
b111 %
1'
1*
b111 +
#729090000000
0!
0'
#729100000000
1!
0$
b1000 %
1'
0*
b1000 +
#729110000000
0!
0'
#729120000000
1!
b1001 %
1'
b1001 +
#729130000000
0!
0'
#729140000000
1!
b0 %
1'
b0 +
#729150000000
0!
0'
#729160000000
1!
1$
b1 %
1'
1*
b1 +
#729170000000
0!
0'
#729180000000
1!
b10 %
1'
b10 +
#729190000000
0!
0'
#729200000000
1!
b11 %
1'
b11 +
#729210000000
0!
0'
#729220000000
1!
b100 %
1'
b100 +
#729230000000
0!
0'
#729240000000
1!
b101 %
1'
b101 +
#729250000000
0!
0'
#729260000000
1!
b110 %
1'
b110 +
#729270000000
0!
0'
#729280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#729290000000
0!
0'
#729300000000
1!
b1000 %
1'
b1000 +
#729310000000
0!
0'
#729320000000
1!
b1001 %
1'
b1001 +
#729330000000
0!
0'
#729340000000
1!
b0 %
1'
b0 +
#729350000000
0!
0'
#729360000000
1!
1$
b1 %
1'
1*
b1 +
#729370000000
0!
0'
#729380000000
1!
b10 %
1'
b10 +
#729390000000
0!
0'
#729400000000
1!
b11 %
1'
b11 +
#729410000000
0!
0'
#729420000000
1!
b100 %
1'
b100 +
#729430000000
0!
0'
#729440000000
1!
b101 %
1'
b101 +
#729450000000
0!
0'
#729460000000
1!
0$
b110 %
1'
0*
b110 +
#729470000000
0!
0'
#729480000000
1!
b111 %
1'
b111 +
#729490000000
1"
1(
#729500000000
0!
0"
b100 &
0'
0(
b100 ,
#729510000000
1!
b1000 %
1'
b1000 +
#729520000000
0!
0'
#729530000000
1!
b1001 %
1'
b1001 +
#729540000000
0!
0'
#729550000000
1!
b0 %
1'
b0 +
#729560000000
0!
0'
#729570000000
1!
1$
b1 %
1'
1*
b1 +
#729580000000
0!
0'
#729590000000
1!
b10 %
1'
b10 +
#729600000000
0!
0'
#729610000000
1!
b11 %
1'
b11 +
#729620000000
0!
0'
#729630000000
1!
b100 %
1'
b100 +
#729640000000
0!
0'
#729650000000
1!
b101 %
1'
b101 +
#729660000000
0!
0'
#729670000000
1!
b110 %
1'
b110 +
#729680000000
0!
0'
#729690000000
1!
b111 %
1'
b111 +
#729700000000
0!
0'
#729710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#729720000000
0!
0'
#729730000000
1!
b1001 %
1'
b1001 +
#729740000000
0!
0'
#729750000000
1!
b0 %
1'
b0 +
#729760000000
0!
0'
#729770000000
1!
1$
b1 %
1'
1*
b1 +
#729780000000
0!
0'
#729790000000
1!
b10 %
1'
b10 +
#729800000000
0!
0'
#729810000000
1!
b11 %
1'
b11 +
#729820000000
0!
0'
#729830000000
1!
b100 %
1'
b100 +
#729840000000
0!
0'
#729850000000
1!
b101 %
1'
b101 +
#729860000000
0!
0'
#729870000000
1!
0$
b110 %
1'
0*
b110 +
#729880000000
0!
0'
#729890000000
1!
b111 %
1'
b111 +
#729900000000
0!
0'
#729910000000
1!
b1000 %
1'
b1000 +
#729920000000
1"
1(
#729930000000
0!
0"
b100 &
0'
0(
b100 ,
#729940000000
1!
b1001 %
1'
b1001 +
#729950000000
0!
0'
#729960000000
1!
b0 %
1'
b0 +
#729970000000
0!
0'
#729980000000
1!
1$
b1 %
1'
1*
b1 +
#729990000000
0!
0'
#730000000000
1!
b10 %
1'
b10 +
#730010000000
0!
0'
#730020000000
1!
b11 %
1'
b11 +
#730030000000
0!
0'
#730040000000
1!
b100 %
1'
b100 +
#730050000000
0!
0'
#730060000000
1!
b101 %
1'
b101 +
#730070000000
0!
0'
#730080000000
1!
b110 %
1'
b110 +
#730090000000
0!
0'
#730100000000
1!
b111 %
1'
b111 +
#730110000000
0!
0'
#730120000000
1!
0$
b1000 %
1'
0*
b1000 +
#730130000000
0!
0'
#730140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#730150000000
0!
0'
#730160000000
1!
b0 %
1'
b0 +
#730170000000
0!
0'
#730180000000
1!
1$
b1 %
1'
1*
b1 +
#730190000000
0!
0'
#730200000000
1!
b10 %
1'
b10 +
#730210000000
0!
0'
#730220000000
1!
b11 %
1'
b11 +
#730230000000
0!
0'
#730240000000
1!
b100 %
1'
b100 +
#730250000000
0!
0'
#730260000000
1!
b101 %
1'
b101 +
#730270000000
0!
0'
#730280000000
1!
0$
b110 %
1'
0*
b110 +
#730290000000
0!
0'
#730300000000
1!
b111 %
1'
b111 +
#730310000000
0!
0'
#730320000000
1!
b1000 %
1'
b1000 +
#730330000000
0!
0'
#730340000000
1!
b1001 %
1'
b1001 +
#730350000000
1"
1(
#730360000000
0!
0"
b100 &
0'
0(
b100 ,
#730370000000
1!
b0 %
1'
b0 +
#730380000000
0!
0'
#730390000000
1!
1$
b1 %
1'
1*
b1 +
#730400000000
0!
0'
#730410000000
1!
b10 %
1'
b10 +
#730420000000
0!
0'
#730430000000
1!
b11 %
1'
b11 +
#730440000000
0!
0'
#730450000000
1!
b100 %
1'
b100 +
#730460000000
0!
0'
#730470000000
1!
b101 %
1'
b101 +
#730480000000
0!
0'
#730490000000
1!
b110 %
1'
b110 +
#730500000000
0!
0'
#730510000000
1!
b111 %
1'
b111 +
#730520000000
0!
0'
#730530000000
1!
0$
b1000 %
1'
0*
b1000 +
#730540000000
0!
0'
#730550000000
1!
b1001 %
1'
b1001 +
#730560000000
0!
0'
#730570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#730580000000
0!
0'
#730590000000
1!
1$
b1 %
1'
1*
b1 +
#730600000000
0!
0'
#730610000000
1!
b10 %
1'
b10 +
#730620000000
0!
0'
#730630000000
1!
b11 %
1'
b11 +
#730640000000
0!
0'
#730650000000
1!
b100 %
1'
b100 +
#730660000000
0!
0'
#730670000000
1!
b101 %
1'
b101 +
#730680000000
0!
0'
#730690000000
1!
0$
b110 %
1'
0*
b110 +
#730700000000
0!
0'
#730710000000
1!
b111 %
1'
b111 +
#730720000000
0!
0'
#730730000000
1!
b1000 %
1'
b1000 +
#730740000000
0!
0'
#730750000000
1!
b1001 %
1'
b1001 +
#730760000000
0!
0'
#730770000000
1!
b0 %
1'
b0 +
#730780000000
1"
1(
#730790000000
0!
0"
b100 &
0'
0(
b100 ,
#730800000000
1!
1$
b1 %
1'
1*
b1 +
#730810000000
0!
0'
#730820000000
1!
b10 %
1'
b10 +
#730830000000
0!
0'
#730840000000
1!
b11 %
1'
b11 +
#730850000000
0!
0'
#730860000000
1!
b100 %
1'
b100 +
#730870000000
0!
0'
#730880000000
1!
b101 %
1'
b101 +
#730890000000
0!
0'
#730900000000
1!
b110 %
1'
b110 +
#730910000000
0!
0'
#730920000000
1!
b111 %
1'
b111 +
#730930000000
0!
0'
#730940000000
1!
0$
b1000 %
1'
0*
b1000 +
#730950000000
0!
0'
#730960000000
1!
b1001 %
1'
b1001 +
#730970000000
0!
0'
#730980000000
1!
b0 %
1'
b0 +
#730990000000
0!
0'
#731000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#731010000000
0!
0'
#731020000000
1!
b10 %
1'
b10 +
#731030000000
0!
0'
#731040000000
1!
b11 %
1'
b11 +
#731050000000
0!
0'
#731060000000
1!
b100 %
1'
b100 +
#731070000000
0!
0'
#731080000000
1!
b101 %
1'
b101 +
#731090000000
0!
0'
#731100000000
1!
0$
b110 %
1'
0*
b110 +
#731110000000
0!
0'
#731120000000
1!
b111 %
1'
b111 +
#731130000000
0!
0'
#731140000000
1!
b1000 %
1'
b1000 +
#731150000000
0!
0'
#731160000000
1!
b1001 %
1'
b1001 +
#731170000000
0!
0'
#731180000000
1!
b0 %
1'
b0 +
#731190000000
0!
0'
#731200000000
1!
1$
b1 %
1'
1*
b1 +
#731210000000
1"
1(
#731220000000
0!
0"
b100 &
0'
0(
b100 ,
#731230000000
1!
b10 %
1'
b10 +
#731240000000
0!
0'
#731250000000
1!
b11 %
1'
b11 +
#731260000000
0!
0'
#731270000000
1!
b100 %
1'
b100 +
#731280000000
0!
0'
#731290000000
1!
b101 %
1'
b101 +
#731300000000
0!
0'
#731310000000
1!
b110 %
1'
b110 +
#731320000000
0!
0'
#731330000000
1!
b111 %
1'
b111 +
#731340000000
0!
0'
#731350000000
1!
0$
b1000 %
1'
0*
b1000 +
#731360000000
0!
0'
#731370000000
1!
b1001 %
1'
b1001 +
#731380000000
0!
0'
#731390000000
1!
b0 %
1'
b0 +
#731400000000
0!
0'
#731410000000
1!
1$
b1 %
1'
1*
b1 +
#731420000000
0!
0'
#731430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#731440000000
0!
0'
#731450000000
1!
b11 %
1'
b11 +
#731460000000
0!
0'
#731470000000
1!
b100 %
1'
b100 +
#731480000000
0!
0'
#731490000000
1!
b101 %
1'
b101 +
#731500000000
0!
0'
#731510000000
1!
0$
b110 %
1'
0*
b110 +
#731520000000
0!
0'
#731530000000
1!
b111 %
1'
b111 +
#731540000000
0!
0'
#731550000000
1!
b1000 %
1'
b1000 +
#731560000000
0!
0'
#731570000000
1!
b1001 %
1'
b1001 +
#731580000000
0!
0'
#731590000000
1!
b0 %
1'
b0 +
#731600000000
0!
0'
#731610000000
1!
1$
b1 %
1'
1*
b1 +
#731620000000
0!
0'
#731630000000
1!
b10 %
1'
b10 +
#731640000000
1"
1(
#731650000000
0!
0"
b100 &
0'
0(
b100 ,
#731660000000
1!
b11 %
1'
b11 +
#731670000000
0!
0'
#731680000000
1!
b100 %
1'
b100 +
#731690000000
0!
0'
#731700000000
1!
b101 %
1'
b101 +
#731710000000
0!
0'
#731720000000
1!
b110 %
1'
b110 +
#731730000000
0!
0'
#731740000000
1!
b111 %
1'
b111 +
#731750000000
0!
0'
#731760000000
1!
0$
b1000 %
1'
0*
b1000 +
#731770000000
0!
0'
#731780000000
1!
b1001 %
1'
b1001 +
#731790000000
0!
0'
#731800000000
1!
b0 %
1'
b0 +
#731810000000
0!
0'
#731820000000
1!
1$
b1 %
1'
1*
b1 +
#731830000000
0!
0'
#731840000000
1!
b10 %
1'
b10 +
#731850000000
0!
0'
#731860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#731870000000
0!
0'
#731880000000
1!
b100 %
1'
b100 +
#731890000000
0!
0'
#731900000000
1!
b101 %
1'
b101 +
#731910000000
0!
0'
#731920000000
1!
0$
b110 %
1'
0*
b110 +
#731930000000
0!
0'
#731940000000
1!
b111 %
1'
b111 +
#731950000000
0!
0'
#731960000000
1!
b1000 %
1'
b1000 +
#731970000000
0!
0'
#731980000000
1!
b1001 %
1'
b1001 +
#731990000000
0!
0'
#732000000000
1!
b0 %
1'
b0 +
#732010000000
0!
0'
#732020000000
1!
1$
b1 %
1'
1*
b1 +
#732030000000
0!
0'
#732040000000
1!
b10 %
1'
b10 +
#732050000000
0!
0'
#732060000000
1!
b11 %
1'
b11 +
#732070000000
1"
1(
#732080000000
0!
0"
b100 &
0'
0(
b100 ,
#732090000000
1!
b100 %
1'
b100 +
#732100000000
0!
0'
#732110000000
1!
b101 %
1'
b101 +
#732120000000
0!
0'
#732130000000
1!
b110 %
1'
b110 +
#732140000000
0!
0'
#732150000000
1!
b111 %
1'
b111 +
#732160000000
0!
0'
#732170000000
1!
0$
b1000 %
1'
0*
b1000 +
#732180000000
0!
0'
#732190000000
1!
b1001 %
1'
b1001 +
#732200000000
0!
0'
#732210000000
1!
b0 %
1'
b0 +
#732220000000
0!
0'
#732230000000
1!
1$
b1 %
1'
1*
b1 +
#732240000000
0!
0'
#732250000000
1!
b10 %
1'
b10 +
#732260000000
0!
0'
#732270000000
1!
b11 %
1'
b11 +
#732280000000
0!
0'
#732290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#732300000000
0!
0'
#732310000000
1!
b101 %
1'
b101 +
#732320000000
0!
0'
#732330000000
1!
0$
b110 %
1'
0*
b110 +
#732340000000
0!
0'
#732350000000
1!
b111 %
1'
b111 +
#732360000000
0!
0'
#732370000000
1!
b1000 %
1'
b1000 +
#732380000000
0!
0'
#732390000000
1!
b1001 %
1'
b1001 +
#732400000000
0!
0'
#732410000000
1!
b0 %
1'
b0 +
#732420000000
0!
0'
#732430000000
1!
1$
b1 %
1'
1*
b1 +
#732440000000
0!
0'
#732450000000
1!
b10 %
1'
b10 +
#732460000000
0!
0'
#732470000000
1!
b11 %
1'
b11 +
#732480000000
0!
0'
#732490000000
1!
b100 %
1'
b100 +
#732500000000
1"
1(
#732510000000
0!
0"
b100 &
0'
0(
b100 ,
#732520000000
1!
b101 %
1'
b101 +
#732530000000
0!
0'
#732540000000
1!
b110 %
1'
b110 +
#732550000000
0!
0'
#732560000000
1!
b111 %
1'
b111 +
#732570000000
0!
0'
#732580000000
1!
0$
b1000 %
1'
0*
b1000 +
#732590000000
0!
0'
#732600000000
1!
b1001 %
1'
b1001 +
#732610000000
0!
0'
#732620000000
1!
b0 %
1'
b0 +
#732630000000
0!
0'
#732640000000
1!
1$
b1 %
1'
1*
b1 +
#732650000000
0!
0'
#732660000000
1!
b10 %
1'
b10 +
#732670000000
0!
0'
#732680000000
1!
b11 %
1'
b11 +
#732690000000
0!
0'
#732700000000
1!
b100 %
1'
b100 +
#732710000000
0!
0'
#732720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#732730000000
0!
0'
#732740000000
1!
0$
b110 %
1'
0*
b110 +
#732750000000
0!
0'
#732760000000
1!
b111 %
1'
b111 +
#732770000000
0!
0'
#732780000000
1!
b1000 %
1'
b1000 +
#732790000000
0!
0'
#732800000000
1!
b1001 %
1'
b1001 +
#732810000000
0!
0'
#732820000000
1!
b0 %
1'
b0 +
#732830000000
0!
0'
#732840000000
1!
1$
b1 %
1'
1*
b1 +
#732850000000
0!
0'
#732860000000
1!
b10 %
1'
b10 +
#732870000000
0!
0'
#732880000000
1!
b11 %
1'
b11 +
#732890000000
0!
0'
#732900000000
1!
b100 %
1'
b100 +
#732910000000
0!
0'
#732920000000
1!
b101 %
1'
b101 +
#732930000000
1"
1(
#732940000000
0!
0"
b100 &
0'
0(
b100 ,
#732950000000
1!
b110 %
1'
b110 +
#732960000000
0!
0'
#732970000000
1!
b111 %
1'
b111 +
#732980000000
0!
0'
#732990000000
1!
0$
b1000 %
1'
0*
b1000 +
#733000000000
0!
0'
#733010000000
1!
b1001 %
1'
b1001 +
#733020000000
0!
0'
#733030000000
1!
b0 %
1'
b0 +
#733040000000
0!
0'
#733050000000
1!
1$
b1 %
1'
1*
b1 +
#733060000000
0!
0'
#733070000000
1!
b10 %
1'
b10 +
#733080000000
0!
0'
#733090000000
1!
b11 %
1'
b11 +
#733100000000
0!
0'
#733110000000
1!
b100 %
1'
b100 +
#733120000000
0!
0'
#733130000000
1!
b101 %
1'
b101 +
#733140000000
0!
0'
#733150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#733160000000
0!
0'
#733170000000
1!
b111 %
1'
b111 +
#733180000000
0!
0'
#733190000000
1!
b1000 %
1'
b1000 +
#733200000000
0!
0'
#733210000000
1!
b1001 %
1'
b1001 +
#733220000000
0!
0'
#733230000000
1!
b0 %
1'
b0 +
#733240000000
0!
0'
#733250000000
1!
1$
b1 %
1'
1*
b1 +
#733260000000
0!
0'
#733270000000
1!
b10 %
1'
b10 +
#733280000000
0!
0'
#733290000000
1!
b11 %
1'
b11 +
#733300000000
0!
0'
#733310000000
1!
b100 %
1'
b100 +
#733320000000
0!
0'
#733330000000
1!
b101 %
1'
b101 +
#733340000000
0!
0'
#733350000000
1!
0$
b110 %
1'
0*
b110 +
#733360000000
1"
1(
#733370000000
0!
0"
b100 &
0'
0(
b100 ,
#733380000000
1!
1$
b111 %
1'
1*
b111 +
#733390000000
0!
0'
#733400000000
1!
0$
b1000 %
1'
0*
b1000 +
#733410000000
0!
0'
#733420000000
1!
b1001 %
1'
b1001 +
#733430000000
0!
0'
#733440000000
1!
b0 %
1'
b0 +
#733450000000
0!
0'
#733460000000
1!
1$
b1 %
1'
1*
b1 +
#733470000000
0!
0'
#733480000000
1!
b10 %
1'
b10 +
#733490000000
0!
0'
#733500000000
1!
b11 %
1'
b11 +
#733510000000
0!
0'
#733520000000
1!
b100 %
1'
b100 +
#733530000000
0!
0'
#733540000000
1!
b101 %
1'
b101 +
#733550000000
0!
0'
#733560000000
1!
b110 %
1'
b110 +
#733570000000
0!
0'
#733580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#733590000000
0!
0'
#733600000000
1!
b1000 %
1'
b1000 +
#733610000000
0!
0'
#733620000000
1!
b1001 %
1'
b1001 +
#733630000000
0!
0'
#733640000000
1!
b0 %
1'
b0 +
#733650000000
0!
0'
#733660000000
1!
1$
b1 %
1'
1*
b1 +
#733670000000
0!
0'
#733680000000
1!
b10 %
1'
b10 +
#733690000000
0!
0'
#733700000000
1!
b11 %
1'
b11 +
#733710000000
0!
0'
#733720000000
1!
b100 %
1'
b100 +
#733730000000
0!
0'
#733740000000
1!
b101 %
1'
b101 +
#733750000000
0!
0'
#733760000000
1!
0$
b110 %
1'
0*
b110 +
#733770000000
0!
0'
#733780000000
1!
b111 %
1'
b111 +
#733790000000
1"
1(
#733800000000
0!
0"
b100 &
0'
0(
b100 ,
#733810000000
1!
b1000 %
1'
b1000 +
#733820000000
0!
0'
#733830000000
1!
b1001 %
1'
b1001 +
#733840000000
0!
0'
#733850000000
1!
b0 %
1'
b0 +
#733860000000
0!
0'
#733870000000
1!
1$
b1 %
1'
1*
b1 +
#733880000000
0!
0'
#733890000000
1!
b10 %
1'
b10 +
#733900000000
0!
0'
#733910000000
1!
b11 %
1'
b11 +
#733920000000
0!
0'
#733930000000
1!
b100 %
1'
b100 +
#733940000000
0!
0'
#733950000000
1!
b101 %
1'
b101 +
#733960000000
0!
0'
#733970000000
1!
b110 %
1'
b110 +
#733980000000
0!
0'
#733990000000
1!
b111 %
1'
b111 +
#734000000000
0!
0'
#734010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#734020000000
0!
0'
#734030000000
1!
b1001 %
1'
b1001 +
#734040000000
0!
0'
#734050000000
1!
b0 %
1'
b0 +
#734060000000
0!
0'
#734070000000
1!
1$
b1 %
1'
1*
b1 +
#734080000000
0!
0'
#734090000000
1!
b10 %
1'
b10 +
#734100000000
0!
0'
#734110000000
1!
b11 %
1'
b11 +
#734120000000
0!
0'
#734130000000
1!
b100 %
1'
b100 +
#734140000000
0!
0'
#734150000000
1!
b101 %
1'
b101 +
#734160000000
0!
0'
#734170000000
1!
0$
b110 %
1'
0*
b110 +
#734180000000
0!
0'
#734190000000
1!
b111 %
1'
b111 +
#734200000000
0!
0'
#734210000000
1!
b1000 %
1'
b1000 +
#734220000000
1"
1(
#734230000000
0!
0"
b100 &
0'
0(
b100 ,
#734240000000
1!
b1001 %
1'
b1001 +
#734250000000
0!
0'
#734260000000
1!
b0 %
1'
b0 +
#734270000000
0!
0'
#734280000000
1!
1$
b1 %
1'
1*
b1 +
#734290000000
0!
0'
#734300000000
1!
b10 %
1'
b10 +
#734310000000
0!
0'
#734320000000
1!
b11 %
1'
b11 +
#734330000000
0!
0'
#734340000000
1!
b100 %
1'
b100 +
#734350000000
0!
0'
#734360000000
1!
b101 %
1'
b101 +
#734370000000
0!
0'
#734380000000
1!
b110 %
1'
b110 +
#734390000000
0!
0'
#734400000000
1!
b111 %
1'
b111 +
#734410000000
0!
0'
#734420000000
1!
0$
b1000 %
1'
0*
b1000 +
#734430000000
0!
0'
#734440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#734450000000
0!
0'
#734460000000
1!
b0 %
1'
b0 +
#734470000000
0!
0'
#734480000000
1!
1$
b1 %
1'
1*
b1 +
#734490000000
0!
0'
#734500000000
1!
b10 %
1'
b10 +
#734510000000
0!
0'
#734520000000
1!
b11 %
1'
b11 +
#734530000000
0!
0'
#734540000000
1!
b100 %
1'
b100 +
#734550000000
0!
0'
#734560000000
1!
b101 %
1'
b101 +
#734570000000
0!
0'
#734580000000
1!
0$
b110 %
1'
0*
b110 +
#734590000000
0!
0'
#734600000000
1!
b111 %
1'
b111 +
#734610000000
0!
0'
#734620000000
1!
b1000 %
1'
b1000 +
#734630000000
0!
0'
#734640000000
1!
b1001 %
1'
b1001 +
#734650000000
1"
1(
#734660000000
0!
0"
b100 &
0'
0(
b100 ,
#734670000000
1!
b0 %
1'
b0 +
#734680000000
0!
0'
#734690000000
1!
1$
b1 %
1'
1*
b1 +
#734700000000
0!
0'
#734710000000
1!
b10 %
1'
b10 +
#734720000000
0!
0'
#734730000000
1!
b11 %
1'
b11 +
#734740000000
0!
0'
#734750000000
1!
b100 %
1'
b100 +
#734760000000
0!
0'
#734770000000
1!
b101 %
1'
b101 +
#734780000000
0!
0'
#734790000000
1!
b110 %
1'
b110 +
#734800000000
0!
0'
#734810000000
1!
b111 %
1'
b111 +
#734820000000
0!
0'
#734830000000
1!
0$
b1000 %
1'
0*
b1000 +
#734840000000
0!
0'
#734850000000
1!
b1001 %
1'
b1001 +
#734860000000
0!
0'
#734870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#734880000000
0!
0'
#734890000000
1!
1$
b1 %
1'
1*
b1 +
#734900000000
0!
0'
#734910000000
1!
b10 %
1'
b10 +
#734920000000
0!
0'
#734930000000
1!
b11 %
1'
b11 +
#734940000000
0!
0'
#734950000000
1!
b100 %
1'
b100 +
#734960000000
0!
0'
#734970000000
1!
b101 %
1'
b101 +
#734980000000
0!
0'
#734990000000
1!
0$
b110 %
1'
0*
b110 +
#735000000000
0!
0'
#735010000000
1!
b111 %
1'
b111 +
#735020000000
0!
0'
#735030000000
1!
b1000 %
1'
b1000 +
#735040000000
0!
0'
#735050000000
1!
b1001 %
1'
b1001 +
#735060000000
0!
0'
#735070000000
1!
b0 %
1'
b0 +
#735080000000
1"
1(
#735090000000
0!
0"
b100 &
0'
0(
b100 ,
#735100000000
1!
1$
b1 %
1'
1*
b1 +
#735110000000
0!
0'
#735120000000
1!
b10 %
1'
b10 +
#735130000000
0!
0'
#735140000000
1!
b11 %
1'
b11 +
#735150000000
0!
0'
#735160000000
1!
b100 %
1'
b100 +
#735170000000
0!
0'
#735180000000
1!
b101 %
1'
b101 +
#735190000000
0!
0'
#735200000000
1!
b110 %
1'
b110 +
#735210000000
0!
0'
#735220000000
1!
b111 %
1'
b111 +
#735230000000
0!
0'
#735240000000
1!
0$
b1000 %
1'
0*
b1000 +
#735250000000
0!
0'
#735260000000
1!
b1001 %
1'
b1001 +
#735270000000
0!
0'
#735280000000
1!
b0 %
1'
b0 +
#735290000000
0!
0'
#735300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#735310000000
0!
0'
#735320000000
1!
b10 %
1'
b10 +
#735330000000
0!
0'
#735340000000
1!
b11 %
1'
b11 +
#735350000000
0!
0'
#735360000000
1!
b100 %
1'
b100 +
#735370000000
0!
0'
#735380000000
1!
b101 %
1'
b101 +
#735390000000
0!
0'
#735400000000
1!
0$
b110 %
1'
0*
b110 +
#735410000000
0!
0'
#735420000000
1!
b111 %
1'
b111 +
#735430000000
0!
0'
#735440000000
1!
b1000 %
1'
b1000 +
#735450000000
0!
0'
#735460000000
1!
b1001 %
1'
b1001 +
#735470000000
0!
0'
#735480000000
1!
b0 %
1'
b0 +
#735490000000
0!
0'
#735500000000
1!
1$
b1 %
1'
1*
b1 +
#735510000000
1"
1(
#735520000000
0!
0"
b100 &
0'
0(
b100 ,
#735530000000
1!
b10 %
1'
b10 +
#735540000000
0!
0'
#735550000000
1!
b11 %
1'
b11 +
#735560000000
0!
0'
#735570000000
1!
b100 %
1'
b100 +
#735580000000
0!
0'
#735590000000
1!
b101 %
1'
b101 +
#735600000000
0!
0'
#735610000000
1!
b110 %
1'
b110 +
#735620000000
0!
0'
#735630000000
1!
b111 %
1'
b111 +
#735640000000
0!
0'
#735650000000
1!
0$
b1000 %
1'
0*
b1000 +
#735660000000
0!
0'
#735670000000
1!
b1001 %
1'
b1001 +
#735680000000
0!
0'
#735690000000
1!
b0 %
1'
b0 +
#735700000000
0!
0'
#735710000000
1!
1$
b1 %
1'
1*
b1 +
#735720000000
0!
0'
#735730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#735740000000
0!
0'
#735750000000
1!
b11 %
1'
b11 +
#735760000000
0!
0'
#735770000000
1!
b100 %
1'
b100 +
#735780000000
0!
0'
#735790000000
1!
b101 %
1'
b101 +
#735800000000
0!
0'
#735810000000
1!
0$
b110 %
1'
0*
b110 +
#735820000000
0!
0'
#735830000000
1!
b111 %
1'
b111 +
#735840000000
0!
0'
#735850000000
1!
b1000 %
1'
b1000 +
#735860000000
0!
0'
#735870000000
1!
b1001 %
1'
b1001 +
#735880000000
0!
0'
#735890000000
1!
b0 %
1'
b0 +
#735900000000
0!
0'
#735910000000
1!
1$
b1 %
1'
1*
b1 +
#735920000000
0!
0'
#735930000000
1!
b10 %
1'
b10 +
#735940000000
1"
1(
#735950000000
0!
0"
b100 &
0'
0(
b100 ,
#735960000000
1!
b11 %
1'
b11 +
#735970000000
0!
0'
#735980000000
1!
b100 %
1'
b100 +
#735990000000
0!
0'
#736000000000
1!
b101 %
1'
b101 +
#736010000000
0!
0'
#736020000000
1!
b110 %
1'
b110 +
#736030000000
0!
0'
#736040000000
1!
b111 %
1'
b111 +
#736050000000
0!
0'
#736060000000
1!
0$
b1000 %
1'
0*
b1000 +
#736070000000
0!
0'
#736080000000
1!
b1001 %
1'
b1001 +
#736090000000
0!
0'
#736100000000
1!
b0 %
1'
b0 +
#736110000000
0!
0'
#736120000000
1!
1$
b1 %
1'
1*
b1 +
#736130000000
0!
0'
#736140000000
1!
b10 %
1'
b10 +
#736150000000
0!
0'
#736160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#736170000000
0!
0'
#736180000000
1!
b100 %
1'
b100 +
#736190000000
0!
0'
#736200000000
1!
b101 %
1'
b101 +
#736210000000
0!
0'
#736220000000
1!
0$
b110 %
1'
0*
b110 +
#736230000000
0!
0'
#736240000000
1!
b111 %
1'
b111 +
#736250000000
0!
0'
#736260000000
1!
b1000 %
1'
b1000 +
#736270000000
0!
0'
#736280000000
1!
b1001 %
1'
b1001 +
#736290000000
0!
0'
#736300000000
1!
b0 %
1'
b0 +
#736310000000
0!
0'
#736320000000
1!
1$
b1 %
1'
1*
b1 +
#736330000000
0!
0'
#736340000000
1!
b10 %
1'
b10 +
#736350000000
0!
0'
#736360000000
1!
b11 %
1'
b11 +
#736370000000
1"
1(
#736380000000
0!
0"
b100 &
0'
0(
b100 ,
#736390000000
1!
b100 %
1'
b100 +
#736400000000
0!
0'
#736410000000
1!
b101 %
1'
b101 +
#736420000000
0!
0'
#736430000000
1!
b110 %
1'
b110 +
#736440000000
0!
0'
#736450000000
1!
b111 %
1'
b111 +
#736460000000
0!
0'
#736470000000
1!
0$
b1000 %
1'
0*
b1000 +
#736480000000
0!
0'
#736490000000
1!
b1001 %
1'
b1001 +
#736500000000
0!
0'
#736510000000
1!
b0 %
1'
b0 +
#736520000000
0!
0'
#736530000000
1!
1$
b1 %
1'
1*
b1 +
#736540000000
0!
0'
#736550000000
1!
b10 %
1'
b10 +
#736560000000
0!
0'
#736570000000
1!
b11 %
1'
b11 +
#736580000000
0!
0'
#736590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#736600000000
0!
0'
#736610000000
1!
b101 %
1'
b101 +
#736620000000
0!
0'
#736630000000
1!
0$
b110 %
1'
0*
b110 +
#736640000000
0!
0'
#736650000000
1!
b111 %
1'
b111 +
#736660000000
0!
0'
#736670000000
1!
b1000 %
1'
b1000 +
#736680000000
0!
0'
#736690000000
1!
b1001 %
1'
b1001 +
#736700000000
0!
0'
#736710000000
1!
b0 %
1'
b0 +
#736720000000
0!
0'
#736730000000
1!
1$
b1 %
1'
1*
b1 +
#736740000000
0!
0'
#736750000000
1!
b10 %
1'
b10 +
#736760000000
0!
0'
#736770000000
1!
b11 %
1'
b11 +
#736780000000
0!
0'
#736790000000
1!
b100 %
1'
b100 +
#736800000000
1"
1(
#736810000000
0!
0"
b100 &
0'
0(
b100 ,
#736820000000
1!
b101 %
1'
b101 +
#736830000000
0!
0'
#736840000000
1!
b110 %
1'
b110 +
#736850000000
0!
0'
#736860000000
1!
b111 %
1'
b111 +
#736870000000
0!
0'
#736880000000
1!
0$
b1000 %
1'
0*
b1000 +
#736890000000
0!
0'
#736900000000
1!
b1001 %
1'
b1001 +
#736910000000
0!
0'
#736920000000
1!
b0 %
1'
b0 +
#736930000000
0!
0'
#736940000000
1!
1$
b1 %
1'
1*
b1 +
#736950000000
0!
0'
#736960000000
1!
b10 %
1'
b10 +
#736970000000
0!
0'
#736980000000
1!
b11 %
1'
b11 +
#736990000000
0!
0'
#737000000000
1!
b100 %
1'
b100 +
#737010000000
0!
0'
#737020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#737030000000
0!
0'
#737040000000
1!
0$
b110 %
1'
0*
b110 +
#737050000000
0!
0'
#737060000000
1!
b111 %
1'
b111 +
#737070000000
0!
0'
#737080000000
1!
b1000 %
1'
b1000 +
#737090000000
0!
0'
#737100000000
1!
b1001 %
1'
b1001 +
#737110000000
0!
0'
#737120000000
1!
b0 %
1'
b0 +
#737130000000
0!
0'
#737140000000
1!
1$
b1 %
1'
1*
b1 +
#737150000000
0!
0'
#737160000000
1!
b10 %
1'
b10 +
#737170000000
0!
0'
#737180000000
1!
b11 %
1'
b11 +
#737190000000
0!
0'
#737200000000
1!
b100 %
1'
b100 +
#737210000000
0!
0'
#737220000000
1!
b101 %
1'
b101 +
#737230000000
1"
1(
#737240000000
0!
0"
b100 &
0'
0(
b100 ,
#737250000000
1!
b110 %
1'
b110 +
#737260000000
0!
0'
#737270000000
1!
b111 %
1'
b111 +
#737280000000
0!
0'
#737290000000
1!
0$
b1000 %
1'
0*
b1000 +
#737300000000
0!
0'
#737310000000
1!
b1001 %
1'
b1001 +
#737320000000
0!
0'
#737330000000
1!
b0 %
1'
b0 +
#737340000000
0!
0'
#737350000000
1!
1$
b1 %
1'
1*
b1 +
#737360000000
0!
0'
#737370000000
1!
b10 %
1'
b10 +
#737380000000
0!
0'
#737390000000
1!
b11 %
1'
b11 +
#737400000000
0!
0'
#737410000000
1!
b100 %
1'
b100 +
#737420000000
0!
0'
#737430000000
1!
b101 %
1'
b101 +
#737440000000
0!
0'
#737450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#737460000000
0!
0'
#737470000000
1!
b111 %
1'
b111 +
#737480000000
0!
0'
#737490000000
1!
b1000 %
1'
b1000 +
#737500000000
0!
0'
#737510000000
1!
b1001 %
1'
b1001 +
#737520000000
0!
0'
#737530000000
1!
b0 %
1'
b0 +
#737540000000
0!
0'
#737550000000
1!
1$
b1 %
1'
1*
b1 +
#737560000000
0!
0'
#737570000000
1!
b10 %
1'
b10 +
#737580000000
0!
0'
#737590000000
1!
b11 %
1'
b11 +
#737600000000
0!
0'
#737610000000
1!
b100 %
1'
b100 +
#737620000000
0!
0'
#737630000000
1!
b101 %
1'
b101 +
#737640000000
0!
0'
#737650000000
1!
0$
b110 %
1'
0*
b110 +
#737660000000
1"
1(
#737670000000
0!
0"
b100 &
0'
0(
b100 ,
#737680000000
1!
1$
b111 %
1'
1*
b111 +
#737690000000
0!
0'
#737700000000
1!
0$
b1000 %
1'
0*
b1000 +
#737710000000
0!
0'
#737720000000
1!
b1001 %
1'
b1001 +
#737730000000
0!
0'
#737740000000
1!
b0 %
1'
b0 +
#737750000000
0!
0'
#737760000000
1!
1$
b1 %
1'
1*
b1 +
#737770000000
0!
0'
#737780000000
1!
b10 %
1'
b10 +
#737790000000
0!
0'
#737800000000
1!
b11 %
1'
b11 +
#737810000000
0!
0'
#737820000000
1!
b100 %
1'
b100 +
#737830000000
0!
0'
#737840000000
1!
b101 %
1'
b101 +
#737850000000
0!
0'
#737860000000
1!
b110 %
1'
b110 +
#737870000000
0!
0'
#737880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#737890000000
0!
0'
#737900000000
1!
b1000 %
1'
b1000 +
#737910000000
0!
0'
#737920000000
1!
b1001 %
1'
b1001 +
#737930000000
0!
0'
#737940000000
1!
b0 %
1'
b0 +
#737950000000
0!
0'
#737960000000
1!
1$
b1 %
1'
1*
b1 +
#737970000000
0!
0'
#737980000000
1!
b10 %
1'
b10 +
#737990000000
0!
0'
#738000000000
1!
b11 %
1'
b11 +
#738010000000
0!
0'
#738020000000
1!
b100 %
1'
b100 +
#738030000000
0!
0'
#738040000000
1!
b101 %
1'
b101 +
#738050000000
0!
0'
#738060000000
1!
0$
b110 %
1'
0*
b110 +
#738070000000
0!
0'
#738080000000
1!
b111 %
1'
b111 +
#738090000000
1"
1(
#738100000000
0!
0"
b100 &
0'
0(
b100 ,
#738110000000
1!
b1000 %
1'
b1000 +
#738120000000
0!
0'
#738130000000
1!
b1001 %
1'
b1001 +
#738140000000
0!
0'
#738150000000
1!
b0 %
1'
b0 +
#738160000000
0!
0'
#738170000000
1!
1$
b1 %
1'
1*
b1 +
#738180000000
0!
0'
#738190000000
1!
b10 %
1'
b10 +
#738200000000
0!
0'
#738210000000
1!
b11 %
1'
b11 +
#738220000000
0!
0'
#738230000000
1!
b100 %
1'
b100 +
#738240000000
0!
0'
#738250000000
1!
b101 %
1'
b101 +
#738260000000
0!
0'
#738270000000
1!
b110 %
1'
b110 +
#738280000000
0!
0'
#738290000000
1!
b111 %
1'
b111 +
#738300000000
0!
0'
#738310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#738320000000
0!
0'
#738330000000
1!
b1001 %
1'
b1001 +
#738340000000
0!
0'
#738350000000
1!
b0 %
1'
b0 +
#738360000000
0!
0'
#738370000000
1!
1$
b1 %
1'
1*
b1 +
#738380000000
0!
0'
#738390000000
1!
b10 %
1'
b10 +
#738400000000
0!
0'
#738410000000
1!
b11 %
1'
b11 +
#738420000000
0!
0'
#738430000000
1!
b100 %
1'
b100 +
#738440000000
0!
0'
#738450000000
1!
b101 %
1'
b101 +
#738460000000
0!
0'
#738470000000
1!
0$
b110 %
1'
0*
b110 +
#738480000000
0!
0'
#738490000000
1!
b111 %
1'
b111 +
#738500000000
0!
0'
#738510000000
1!
b1000 %
1'
b1000 +
#738520000000
1"
1(
#738530000000
0!
0"
b100 &
0'
0(
b100 ,
#738540000000
1!
b1001 %
1'
b1001 +
#738550000000
0!
0'
#738560000000
1!
b0 %
1'
b0 +
#738570000000
0!
0'
#738580000000
1!
1$
b1 %
1'
1*
b1 +
#738590000000
0!
0'
#738600000000
1!
b10 %
1'
b10 +
#738610000000
0!
0'
#738620000000
1!
b11 %
1'
b11 +
#738630000000
0!
0'
#738640000000
1!
b100 %
1'
b100 +
#738650000000
0!
0'
#738660000000
1!
b101 %
1'
b101 +
#738670000000
0!
0'
#738680000000
1!
b110 %
1'
b110 +
#738690000000
0!
0'
#738700000000
1!
b111 %
1'
b111 +
#738710000000
0!
0'
#738720000000
1!
0$
b1000 %
1'
0*
b1000 +
#738730000000
0!
0'
#738740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#738750000000
0!
0'
#738760000000
1!
b0 %
1'
b0 +
#738770000000
0!
0'
#738780000000
1!
1$
b1 %
1'
1*
b1 +
#738790000000
0!
0'
#738800000000
1!
b10 %
1'
b10 +
#738810000000
0!
0'
#738820000000
1!
b11 %
1'
b11 +
#738830000000
0!
0'
#738840000000
1!
b100 %
1'
b100 +
#738850000000
0!
0'
#738860000000
1!
b101 %
1'
b101 +
#738870000000
0!
0'
#738880000000
1!
0$
b110 %
1'
0*
b110 +
#738890000000
0!
0'
#738900000000
1!
b111 %
1'
b111 +
#738910000000
0!
0'
#738920000000
1!
b1000 %
1'
b1000 +
#738930000000
0!
0'
#738940000000
1!
b1001 %
1'
b1001 +
#738950000000
1"
1(
#738960000000
0!
0"
b100 &
0'
0(
b100 ,
#738970000000
1!
b0 %
1'
b0 +
#738980000000
0!
0'
#738990000000
1!
1$
b1 %
1'
1*
b1 +
#739000000000
0!
0'
#739010000000
1!
b10 %
1'
b10 +
#739020000000
0!
0'
#739030000000
1!
b11 %
1'
b11 +
#739040000000
0!
0'
#739050000000
1!
b100 %
1'
b100 +
#739060000000
0!
0'
#739070000000
1!
b101 %
1'
b101 +
#739080000000
0!
0'
#739090000000
1!
b110 %
1'
b110 +
#739100000000
0!
0'
#739110000000
1!
b111 %
1'
b111 +
#739120000000
0!
0'
#739130000000
1!
0$
b1000 %
1'
0*
b1000 +
#739140000000
0!
0'
#739150000000
1!
b1001 %
1'
b1001 +
#739160000000
0!
0'
#739170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#739180000000
0!
0'
#739190000000
1!
1$
b1 %
1'
1*
b1 +
#739200000000
0!
0'
#739210000000
1!
b10 %
1'
b10 +
#739220000000
0!
0'
#739230000000
1!
b11 %
1'
b11 +
#739240000000
0!
0'
#739250000000
1!
b100 %
1'
b100 +
#739260000000
0!
0'
#739270000000
1!
b101 %
1'
b101 +
#739280000000
0!
0'
#739290000000
1!
0$
b110 %
1'
0*
b110 +
#739300000000
0!
0'
#739310000000
1!
b111 %
1'
b111 +
#739320000000
0!
0'
#739330000000
1!
b1000 %
1'
b1000 +
#739340000000
0!
0'
#739350000000
1!
b1001 %
1'
b1001 +
#739360000000
0!
0'
#739370000000
1!
b0 %
1'
b0 +
#739380000000
1"
1(
#739390000000
0!
0"
b100 &
0'
0(
b100 ,
#739400000000
1!
1$
b1 %
1'
1*
b1 +
#739410000000
0!
0'
#739420000000
1!
b10 %
1'
b10 +
#739430000000
0!
0'
#739440000000
1!
b11 %
1'
b11 +
#739450000000
0!
0'
#739460000000
1!
b100 %
1'
b100 +
#739470000000
0!
0'
#739480000000
1!
b101 %
1'
b101 +
#739490000000
0!
0'
#739500000000
1!
b110 %
1'
b110 +
#739510000000
0!
0'
#739520000000
1!
b111 %
1'
b111 +
#739530000000
0!
0'
#739540000000
1!
0$
b1000 %
1'
0*
b1000 +
#739550000000
0!
0'
#739560000000
1!
b1001 %
1'
b1001 +
#739570000000
0!
0'
#739580000000
1!
b0 %
1'
b0 +
#739590000000
0!
0'
#739600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#739610000000
0!
0'
#739620000000
1!
b10 %
1'
b10 +
#739630000000
0!
0'
#739640000000
1!
b11 %
1'
b11 +
#739650000000
0!
0'
#739660000000
1!
b100 %
1'
b100 +
#739670000000
0!
0'
#739680000000
1!
b101 %
1'
b101 +
#739690000000
0!
0'
#739700000000
1!
0$
b110 %
1'
0*
b110 +
#739710000000
0!
0'
#739720000000
1!
b111 %
1'
b111 +
#739730000000
0!
0'
#739740000000
1!
b1000 %
1'
b1000 +
#739750000000
0!
0'
#739760000000
1!
b1001 %
1'
b1001 +
#739770000000
0!
0'
#739780000000
1!
b0 %
1'
b0 +
#739790000000
0!
0'
#739800000000
1!
1$
b1 %
1'
1*
b1 +
#739810000000
1"
1(
#739820000000
0!
0"
b100 &
0'
0(
b100 ,
#739830000000
1!
b10 %
1'
b10 +
#739840000000
0!
0'
#739850000000
1!
b11 %
1'
b11 +
#739860000000
0!
0'
#739870000000
1!
b100 %
1'
b100 +
#739880000000
0!
0'
#739890000000
1!
b101 %
1'
b101 +
#739900000000
0!
0'
#739910000000
1!
b110 %
1'
b110 +
#739920000000
0!
0'
#739930000000
1!
b111 %
1'
b111 +
#739940000000
0!
0'
#739950000000
1!
0$
b1000 %
1'
0*
b1000 +
#739960000000
0!
0'
#739970000000
1!
b1001 %
1'
b1001 +
#739980000000
0!
0'
#739990000000
1!
b0 %
1'
b0 +
#740000000000
0!
0'
#740010000000
1!
1$
b1 %
1'
1*
b1 +
#740020000000
0!
0'
#740030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#740040000000
0!
0'
#740050000000
1!
b11 %
1'
b11 +
#740060000000
0!
0'
#740070000000
1!
b100 %
1'
b100 +
#740080000000
0!
0'
#740090000000
1!
b101 %
1'
b101 +
#740100000000
0!
0'
#740110000000
1!
0$
b110 %
1'
0*
b110 +
#740120000000
0!
0'
#740130000000
1!
b111 %
1'
b111 +
#740140000000
0!
0'
#740150000000
1!
b1000 %
1'
b1000 +
#740160000000
0!
0'
#740170000000
1!
b1001 %
1'
b1001 +
#740180000000
0!
0'
#740190000000
1!
b0 %
1'
b0 +
#740200000000
0!
0'
#740210000000
1!
1$
b1 %
1'
1*
b1 +
#740220000000
0!
0'
#740230000000
1!
b10 %
1'
b10 +
#740240000000
1"
1(
#740250000000
0!
0"
b100 &
0'
0(
b100 ,
#740260000000
1!
b11 %
1'
b11 +
#740270000000
0!
0'
#740280000000
1!
b100 %
1'
b100 +
#740290000000
0!
0'
#740300000000
1!
b101 %
1'
b101 +
#740310000000
0!
0'
#740320000000
1!
b110 %
1'
b110 +
#740330000000
0!
0'
#740340000000
1!
b111 %
1'
b111 +
#740350000000
0!
0'
#740360000000
1!
0$
b1000 %
1'
0*
b1000 +
#740370000000
0!
0'
#740380000000
1!
b1001 %
1'
b1001 +
#740390000000
0!
0'
#740400000000
1!
b0 %
1'
b0 +
#740410000000
0!
0'
#740420000000
1!
1$
b1 %
1'
1*
b1 +
#740430000000
0!
0'
#740440000000
1!
b10 %
1'
b10 +
#740450000000
0!
0'
#740460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#740470000000
0!
0'
#740480000000
1!
b100 %
1'
b100 +
#740490000000
0!
0'
#740500000000
1!
b101 %
1'
b101 +
#740510000000
0!
0'
#740520000000
1!
0$
b110 %
1'
0*
b110 +
#740530000000
0!
0'
#740540000000
1!
b111 %
1'
b111 +
#740550000000
0!
0'
#740560000000
1!
b1000 %
1'
b1000 +
#740570000000
0!
0'
#740580000000
1!
b1001 %
1'
b1001 +
#740590000000
0!
0'
#740600000000
1!
b0 %
1'
b0 +
#740610000000
0!
0'
#740620000000
1!
1$
b1 %
1'
1*
b1 +
#740630000000
0!
0'
#740640000000
1!
b10 %
1'
b10 +
#740650000000
0!
0'
#740660000000
1!
b11 %
1'
b11 +
#740670000000
1"
1(
#740680000000
0!
0"
b100 &
0'
0(
b100 ,
#740690000000
1!
b100 %
1'
b100 +
#740700000000
0!
0'
#740710000000
1!
b101 %
1'
b101 +
#740720000000
0!
0'
#740730000000
1!
b110 %
1'
b110 +
#740740000000
0!
0'
#740750000000
1!
b111 %
1'
b111 +
#740760000000
0!
0'
#740770000000
1!
0$
b1000 %
1'
0*
b1000 +
#740780000000
0!
0'
#740790000000
1!
b1001 %
1'
b1001 +
#740800000000
0!
0'
#740810000000
1!
b0 %
1'
b0 +
#740820000000
0!
0'
#740830000000
1!
1$
b1 %
1'
1*
b1 +
#740840000000
0!
0'
#740850000000
1!
b10 %
1'
b10 +
#740860000000
0!
0'
#740870000000
1!
b11 %
1'
b11 +
#740880000000
0!
0'
#740890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#740900000000
0!
0'
#740910000000
1!
b101 %
1'
b101 +
#740920000000
0!
0'
#740930000000
1!
0$
b110 %
1'
0*
b110 +
#740940000000
0!
0'
#740950000000
1!
b111 %
1'
b111 +
#740960000000
0!
0'
#740970000000
1!
b1000 %
1'
b1000 +
#740980000000
0!
0'
#740990000000
1!
b1001 %
1'
b1001 +
#741000000000
0!
0'
#741010000000
1!
b0 %
1'
b0 +
#741020000000
0!
0'
#741030000000
1!
1$
b1 %
1'
1*
b1 +
#741040000000
0!
0'
#741050000000
1!
b10 %
1'
b10 +
#741060000000
0!
0'
#741070000000
1!
b11 %
1'
b11 +
#741080000000
0!
0'
#741090000000
1!
b100 %
1'
b100 +
#741100000000
1"
1(
#741110000000
0!
0"
b100 &
0'
0(
b100 ,
#741120000000
1!
b101 %
1'
b101 +
#741130000000
0!
0'
#741140000000
1!
b110 %
1'
b110 +
#741150000000
0!
0'
#741160000000
1!
b111 %
1'
b111 +
#741170000000
0!
0'
#741180000000
1!
0$
b1000 %
1'
0*
b1000 +
#741190000000
0!
0'
#741200000000
1!
b1001 %
1'
b1001 +
#741210000000
0!
0'
#741220000000
1!
b0 %
1'
b0 +
#741230000000
0!
0'
#741240000000
1!
1$
b1 %
1'
1*
b1 +
#741250000000
0!
0'
#741260000000
1!
b10 %
1'
b10 +
#741270000000
0!
0'
#741280000000
1!
b11 %
1'
b11 +
#741290000000
0!
0'
#741300000000
1!
b100 %
1'
b100 +
#741310000000
0!
0'
#741320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#741330000000
0!
0'
#741340000000
1!
0$
b110 %
1'
0*
b110 +
#741350000000
0!
0'
#741360000000
1!
b111 %
1'
b111 +
#741370000000
0!
0'
#741380000000
1!
b1000 %
1'
b1000 +
#741390000000
0!
0'
#741400000000
1!
b1001 %
1'
b1001 +
#741410000000
0!
0'
#741420000000
1!
b0 %
1'
b0 +
#741430000000
0!
0'
#741440000000
1!
1$
b1 %
1'
1*
b1 +
#741450000000
0!
0'
#741460000000
1!
b10 %
1'
b10 +
#741470000000
0!
0'
#741480000000
1!
b11 %
1'
b11 +
#741490000000
0!
0'
#741500000000
1!
b100 %
1'
b100 +
#741510000000
0!
0'
#741520000000
1!
b101 %
1'
b101 +
#741530000000
1"
1(
#741540000000
0!
0"
b100 &
0'
0(
b100 ,
#741550000000
1!
b110 %
1'
b110 +
#741560000000
0!
0'
#741570000000
1!
b111 %
1'
b111 +
#741580000000
0!
0'
#741590000000
1!
0$
b1000 %
1'
0*
b1000 +
#741600000000
0!
0'
#741610000000
1!
b1001 %
1'
b1001 +
#741620000000
0!
0'
#741630000000
1!
b0 %
1'
b0 +
#741640000000
0!
0'
#741650000000
1!
1$
b1 %
1'
1*
b1 +
#741660000000
0!
0'
#741670000000
1!
b10 %
1'
b10 +
#741680000000
0!
0'
#741690000000
1!
b11 %
1'
b11 +
#741700000000
0!
0'
#741710000000
1!
b100 %
1'
b100 +
#741720000000
0!
0'
#741730000000
1!
b101 %
1'
b101 +
#741740000000
0!
0'
#741750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#741760000000
0!
0'
#741770000000
1!
b111 %
1'
b111 +
#741780000000
0!
0'
#741790000000
1!
b1000 %
1'
b1000 +
#741800000000
0!
0'
#741810000000
1!
b1001 %
1'
b1001 +
#741820000000
0!
0'
#741830000000
1!
b0 %
1'
b0 +
#741840000000
0!
0'
#741850000000
1!
1$
b1 %
1'
1*
b1 +
#741860000000
0!
0'
#741870000000
1!
b10 %
1'
b10 +
#741880000000
0!
0'
#741890000000
1!
b11 %
1'
b11 +
#741900000000
0!
0'
#741910000000
1!
b100 %
1'
b100 +
#741920000000
0!
0'
#741930000000
1!
b101 %
1'
b101 +
#741940000000
0!
0'
#741950000000
1!
0$
b110 %
1'
0*
b110 +
#741960000000
1"
1(
#741970000000
0!
0"
b100 &
0'
0(
b100 ,
#741980000000
1!
1$
b111 %
1'
1*
b111 +
#741990000000
0!
0'
#742000000000
1!
0$
b1000 %
1'
0*
b1000 +
#742010000000
0!
0'
#742020000000
1!
b1001 %
1'
b1001 +
#742030000000
0!
0'
#742040000000
1!
b0 %
1'
b0 +
#742050000000
0!
0'
#742060000000
1!
1$
b1 %
1'
1*
b1 +
#742070000000
0!
0'
#742080000000
1!
b10 %
1'
b10 +
#742090000000
0!
0'
#742100000000
1!
b11 %
1'
b11 +
#742110000000
0!
0'
#742120000000
1!
b100 %
1'
b100 +
#742130000000
0!
0'
#742140000000
1!
b101 %
1'
b101 +
#742150000000
0!
0'
#742160000000
1!
b110 %
1'
b110 +
#742170000000
0!
0'
#742180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#742190000000
0!
0'
#742200000000
1!
b1000 %
1'
b1000 +
#742210000000
0!
0'
#742220000000
1!
b1001 %
1'
b1001 +
#742230000000
0!
0'
#742240000000
1!
b0 %
1'
b0 +
#742250000000
0!
0'
#742260000000
1!
1$
b1 %
1'
1*
b1 +
#742270000000
0!
0'
#742280000000
1!
b10 %
1'
b10 +
#742290000000
0!
0'
#742300000000
1!
b11 %
1'
b11 +
#742310000000
0!
0'
#742320000000
1!
b100 %
1'
b100 +
#742330000000
0!
0'
#742340000000
1!
b101 %
1'
b101 +
#742350000000
0!
0'
#742360000000
1!
0$
b110 %
1'
0*
b110 +
#742370000000
0!
0'
#742380000000
1!
b111 %
1'
b111 +
#742390000000
1"
1(
#742400000000
0!
0"
b100 &
0'
0(
b100 ,
#742410000000
1!
b1000 %
1'
b1000 +
#742420000000
0!
0'
#742430000000
1!
b1001 %
1'
b1001 +
#742440000000
0!
0'
#742450000000
1!
b0 %
1'
b0 +
#742460000000
0!
0'
#742470000000
1!
1$
b1 %
1'
1*
b1 +
#742480000000
0!
0'
#742490000000
1!
b10 %
1'
b10 +
#742500000000
0!
0'
#742510000000
1!
b11 %
1'
b11 +
#742520000000
0!
0'
#742530000000
1!
b100 %
1'
b100 +
#742540000000
0!
0'
#742550000000
1!
b101 %
1'
b101 +
#742560000000
0!
0'
#742570000000
1!
b110 %
1'
b110 +
#742580000000
0!
0'
#742590000000
1!
b111 %
1'
b111 +
#742600000000
0!
0'
#742610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#742620000000
0!
0'
#742630000000
1!
b1001 %
1'
b1001 +
#742640000000
0!
0'
#742650000000
1!
b0 %
1'
b0 +
#742660000000
0!
0'
#742670000000
1!
1$
b1 %
1'
1*
b1 +
#742680000000
0!
0'
#742690000000
1!
b10 %
1'
b10 +
#742700000000
0!
0'
#742710000000
1!
b11 %
1'
b11 +
#742720000000
0!
0'
#742730000000
1!
b100 %
1'
b100 +
#742740000000
0!
0'
#742750000000
1!
b101 %
1'
b101 +
#742760000000
0!
0'
#742770000000
1!
0$
b110 %
1'
0*
b110 +
#742780000000
0!
0'
#742790000000
1!
b111 %
1'
b111 +
#742800000000
0!
0'
#742810000000
1!
b1000 %
1'
b1000 +
#742820000000
1"
1(
#742830000000
0!
0"
b100 &
0'
0(
b100 ,
#742840000000
1!
b1001 %
1'
b1001 +
#742850000000
0!
0'
#742860000000
1!
b0 %
1'
b0 +
#742870000000
0!
0'
#742880000000
1!
1$
b1 %
1'
1*
b1 +
#742890000000
0!
0'
#742900000000
1!
b10 %
1'
b10 +
#742910000000
0!
0'
#742920000000
1!
b11 %
1'
b11 +
#742930000000
0!
0'
#742940000000
1!
b100 %
1'
b100 +
#742950000000
0!
0'
#742960000000
1!
b101 %
1'
b101 +
#742970000000
0!
0'
#742980000000
1!
b110 %
1'
b110 +
#742990000000
0!
0'
#743000000000
1!
b111 %
1'
b111 +
#743010000000
0!
0'
#743020000000
1!
0$
b1000 %
1'
0*
b1000 +
#743030000000
0!
0'
#743040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#743050000000
0!
0'
#743060000000
1!
b0 %
1'
b0 +
#743070000000
0!
0'
#743080000000
1!
1$
b1 %
1'
1*
b1 +
#743090000000
0!
0'
#743100000000
1!
b10 %
1'
b10 +
#743110000000
0!
0'
#743120000000
1!
b11 %
1'
b11 +
#743130000000
0!
0'
#743140000000
1!
b100 %
1'
b100 +
#743150000000
0!
0'
#743160000000
1!
b101 %
1'
b101 +
#743170000000
0!
0'
#743180000000
1!
0$
b110 %
1'
0*
b110 +
#743190000000
0!
0'
#743200000000
1!
b111 %
1'
b111 +
#743210000000
0!
0'
#743220000000
1!
b1000 %
1'
b1000 +
#743230000000
0!
0'
#743240000000
1!
b1001 %
1'
b1001 +
#743250000000
1"
1(
#743260000000
0!
0"
b100 &
0'
0(
b100 ,
#743270000000
1!
b0 %
1'
b0 +
#743280000000
0!
0'
#743290000000
1!
1$
b1 %
1'
1*
b1 +
#743300000000
0!
0'
#743310000000
1!
b10 %
1'
b10 +
#743320000000
0!
0'
#743330000000
1!
b11 %
1'
b11 +
#743340000000
0!
0'
#743350000000
1!
b100 %
1'
b100 +
#743360000000
0!
0'
#743370000000
1!
b101 %
1'
b101 +
#743380000000
0!
0'
#743390000000
1!
b110 %
1'
b110 +
#743400000000
0!
0'
#743410000000
1!
b111 %
1'
b111 +
#743420000000
0!
0'
#743430000000
1!
0$
b1000 %
1'
0*
b1000 +
#743440000000
0!
0'
#743450000000
1!
b1001 %
1'
b1001 +
#743460000000
0!
0'
#743470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#743480000000
0!
0'
#743490000000
1!
1$
b1 %
1'
1*
b1 +
#743500000000
0!
0'
#743510000000
1!
b10 %
1'
b10 +
#743520000000
0!
0'
#743530000000
1!
b11 %
1'
b11 +
#743540000000
0!
0'
#743550000000
1!
b100 %
1'
b100 +
#743560000000
0!
0'
#743570000000
1!
b101 %
1'
b101 +
#743580000000
0!
0'
#743590000000
1!
0$
b110 %
1'
0*
b110 +
#743600000000
0!
0'
#743610000000
1!
b111 %
1'
b111 +
#743620000000
0!
0'
#743630000000
1!
b1000 %
1'
b1000 +
#743640000000
0!
0'
#743650000000
1!
b1001 %
1'
b1001 +
#743660000000
0!
0'
#743670000000
1!
b0 %
1'
b0 +
#743680000000
1"
1(
#743690000000
0!
0"
b100 &
0'
0(
b100 ,
#743700000000
1!
1$
b1 %
1'
1*
b1 +
#743710000000
0!
0'
#743720000000
1!
b10 %
1'
b10 +
#743730000000
0!
0'
#743740000000
1!
b11 %
1'
b11 +
#743750000000
0!
0'
#743760000000
1!
b100 %
1'
b100 +
#743770000000
0!
0'
#743780000000
1!
b101 %
1'
b101 +
#743790000000
0!
0'
#743800000000
1!
b110 %
1'
b110 +
#743810000000
0!
0'
#743820000000
1!
b111 %
1'
b111 +
#743830000000
0!
0'
#743840000000
1!
0$
b1000 %
1'
0*
b1000 +
#743850000000
0!
0'
#743860000000
1!
b1001 %
1'
b1001 +
#743870000000
0!
0'
#743880000000
1!
b0 %
1'
b0 +
#743890000000
0!
0'
#743900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#743910000000
0!
0'
#743920000000
1!
b10 %
1'
b10 +
#743930000000
0!
0'
#743940000000
1!
b11 %
1'
b11 +
#743950000000
0!
0'
#743960000000
1!
b100 %
1'
b100 +
#743970000000
0!
0'
#743980000000
1!
b101 %
1'
b101 +
#743990000000
0!
0'
#744000000000
1!
0$
b110 %
1'
0*
b110 +
#744010000000
0!
0'
#744020000000
1!
b111 %
1'
b111 +
#744030000000
0!
0'
#744040000000
1!
b1000 %
1'
b1000 +
#744050000000
0!
0'
#744060000000
1!
b1001 %
1'
b1001 +
#744070000000
0!
0'
#744080000000
1!
b0 %
1'
b0 +
#744090000000
0!
0'
#744100000000
1!
1$
b1 %
1'
1*
b1 +
#744110000000
1"
1(
#744120000000
0!
0"
b100 &
0'
0(
b100 ,
#744130000000
1!
b10 %
1'
b10 +
#744140000000
0!
0'
#744150000000
1!
b11 %
1'
b11 +
#744160000000
0!
0'
#744170000000
1!
b100 %
1'
b100 +
#744180000000
0!
0'
#744190000000
1!
b101 %
1'
b101 +
#744200000000
0!
0'
#744210000000
1!
b110 %
1'
b110 +
#744220000000
0!
0'
#744230000000
1!
b111 %
1'
b111 +
#744240000000
0!
0'
#744250000000
1!
0$
b1000 %
1'
0*
b1000 +
#744260000000
0!
0'
#744270000000
1!
b1001 %
1'
b1001 +
#744280000000
0!
0'
#744290000000
1!
b0 %
1'
b0 +
#744300000000
0!
0'
#744310000000
1!
1$
b1 %
1'
1*
b1 +
#744320000000
0!
0'
#744330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#744340000000
0!
0'
#744350000000
1!
b11 %
1'
b11 +
#744360000000
0!
0'
#744370000000
1!
b100 %
1'
b100 +
#744380000000
0!
0'
#744390000000
1!
b101 %
1'
b101 +
#744400000000
0!
0'
#744410000000
1!
0$
b110 %
1'
0*
b110 +
#744420000000
0!
0'
#744430000000
1!
b111 %
1'
b111 +
#744440000000
0!
0'
#744450000000
1!
b1000 %
1'
b1000 +
#744460000000
0!
0'
#744470000000
1!
b1001 %
1'
b1001 +
#744480000000
0!
0'
#744490000000
1!
b0 %
1'
b0 +
#744500000000
0!
0'
#744510000000
1!
1$
b1 %
1'
1*
b1 +
#744520000000
0!
0'
#744530000000
1!
b10 %
1'
b10 +
#744540000000
1"
1(
#744550000000
0!
0"
b100 &
0'
0(
b100 ,
#744560000000
1!
b11 %
1'
b11 +
#744570000000
0!
0'
#744580000000
1!
b100 %
1'
b100 +
#744590000000
0!
0'
#744600000000
1!
b101 %
1'
b101 +
#744610000000
0!
0'
#744620000000
1!
b110 %
1'
b110 +
#744630000000
0!
0'
#744640000000
1!
b111 %
1'
b111 +
#744650000000
0!
0'
#744660000000
1!
0$
b1000 %
1'
0*
b1000 +
#744670000000
0!
0'
#744680000000
1!
b1001 %
1'
b1001 +
#744690000000
0!
0'
#744700000000
1!
b0 %
1'
b0 +
#744710000000
0!
0'
#744720000000
1!
1$
b1 %
1'
1*
b1 +
#744730000000
0!
0'
#744740000000
1!
b10 %
1'
b10 +
#744750000000
0!
0'
#744760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#744770000000
0!
0'
#744780000000
1!
b100 %
1'
b100 +
#744790000000
0!
0'
#744800000000
1!
b101 %
1'
b101 +
#744810000000
0!
0'
#744820000000
1!
0$
b110 %
1'
0*
b110 +
#744830000000
0!
0'
#744840000000
1!
b111 %
1'
b111 +
#744850000000
0!
0'
#744860000000
1!
b1000 %
1'
b1000 +
#744870000000
0!
0'
#744880000000
1!
b1001 %
1'
b1001 +
#744890000000
0!
0'
#744900000000
1!
b0 %
1'
b0 +
#744910000000
0!
0'
#744920000000
1!
1$
b1 %
1'
1*
b1 +
#744930000000
0!
0'
#744940000000
1!
b10 %
1'
b10 +
#744950000000
0!
0'
#744960000000
1!
b11 %
1'
b11 +
#744970000000
1"
1(
#744980000000
0!
0"
b100 &
0'
0(
b100 ,
#744990000000
1!
b100 %
1'
b100 +
#745000000000
0!
0'
#745010000000
1!
b101 %
1'
b101 +
#745020000000
0!
0'
#745030000000
1!
b110 %
1'
b110 +
#745040000000
0!
0'
#745050000000
1!
b111 %
1'
b111 +
#745060000000
0!
0'
#745070000000
1!
0$
b1000 %
1'
0*
b1000 +
#745080000000
0!
0'
#745090000000
1!
b1001 %
1'
b1001 +
#745100000000
0!
0'
#745110000000
1!
b0 %
1'
b0 +
#745120000000
0!
0'
#745130000000
1!
1$
b1 %
1'
1*
b1 +
#745140000000
0!
0'
#745150000000
1!
b10 %
1'
b10 +
#745160000000
0!
0'
#745170000000
1!
b11 %
1'
b11 +
#745180000000
0!
0'
#745190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#745200000000
0!
0'
#745210000000
1!
b101 %
1'
b101 +
#745220000000
0!
0'
#745230000000
1!
0$
b110 %
1'
0*
b110 +
#745240000000
0!
0'
#745250000000
1!
b111 %
1'
b111 +
#745260000000
0!
0'
#745270000000
1!
b1000 %
1'
b1000 +
#745280000000
0!
0'
#745290000000
1!
b1001 %
1'
b1001 +
#745300000000
0!
0'
#745310000000
1!
b0 %
1'
b0 +
#745320000000
0!
0'
#745330000000
1!
1$
b1 %
1'
1*
b1 +
#745340000000
0!
0'
#745350000000
1!
b10 %
1'
b10 +
#745360000000
0!
0'
#745370000000
1!
b11 %
1'
b11 +
#745380000000
0!
0'
#745390000000
1!
b100 %
1'
b100 +
#745400000000
1"
1(
#745410000000
0!
0"
b100 &
0'
0(
b100 ,
#745420000000
1!
b101 %
1'
b101 +
#745430000000
0!
0'
#745440000000
1!
b110 %
1'
b110 +
#745450000000
0!
0'
#745460000000
1!
b111 %
1'
b111 +
#745470000000
0!
0'
#745480000000
1!
0$
b1000 %
1'
0*
b1000 +
#745490000000
0!
0'
#745500000000
1!
b1001 %
1'
b1001 +
#745510000000
0!
0'
#745520000000
1!
b0 %
1'
b0 +
#745530000000
0!
0'
#745540000000
1!
1$
b1 %
1'
1*
b1 +
#745550000000
0!
0'
#745560000000
1!
b10 %
1'
b10 +
#745570000000
0!
0'
#745580000000
1!
b11 %
1'
b11 +
#745590000000
0!
0'
#745600000000
1!
b100 %
1'
b100 +
#745610000000
0!
0'
#745620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#745630000000
0!
0'
#745640000000
1!
0$
b110 %
1'
0*
b110 +
#745650000000
0!
0'
#745660000000
1!
b111 %
1'
b111 +
#745670000000
0!
0'
#745680000000
1!
b1000 %
1'
b1000 +
#745690000000
0!
0'
#745700000000
1!
b1001 %
1'
b1001 +
#745710000000
0!
0'
#745720000000
1!
b0 %
1'
b0 +
#745730000000
0!
0'
#745740000000
1!
1$
b1 %
1'
1*
b1 +
#745750000000
0!
0'
#745760000000
1!
b10 %
1'
b10 +
#745770000000
0!
0'
#745780000000
1!
b11 %
1'
b11 +
#745790000000
0!
0'
#745800000000
1!
b100 %
1'
b100 +
#745810000000
0!
0'
#745820000000
1!
b101 %
1'
b101 +
#745830000000
1"
1(
#745840000000
0!
0"
b100 &
0'
0(
b100 ,
#745850000000
1!
b110 %
1'
b110 +
#745860000000
0!
0'
#745870000000
1!
b111 %
1'
b111 +
#745880000000
0!
0'
#745890000000
1!
0$
b1000 %
1'
0*
b1000 +
#745900000000
0!
0'
#745910000000
1!
b1001 %
1'
b1001 +
#745920000000
0!
0'
#745930000000
1!
b0 %
1'
b0 +
#745940000000
0!
0'
#745950000000
1!
1$
b1 %
1'
1*
b1 +
#745960000000
0!
0'
#745970000000
1!
b10 %
1'
b10 +
#745980000000
0!
0'
#745990000000
1!
b11 %
1'
b11 +
#746000000000
0!
0'
#746010000000
1!
b100 %
1'
b100 +
#746020000000
0!
0'
#746030000000
1!
b101 %
1'
b101 +
#746040000000
0!
0'
#746050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#746060000000
0!
0'
#746070000000
1!
b111 %
1'
b111 +
#746080000000
0!
0'
#746090000000
1!
b1000 %
1'
b1000 +
#746100000000
0!
0'
#746110000000
1!
b1001 %
1'
b1001 +
#746120000000
0!
0'
#746130000000
1!
b0 %
1'
b0 +
#746140000000
0!
0'
#746150000000
1!
1$
b1 %
1'
1*
b1 +
#746160000000
0!
0'
#746170000000
1!
b10 %
1'
b10 +
#746180000000
0!
0'
#746190000000
1!
b11 %
1'
b11 +
#746200000000
0!
0'
#746210000000
1!
b100 %
1'
b100 +
#746220000000
0!
0'
#746230000000
1!
b101 %
1'
b101 +
#746240000000
0!
0'
#746250000000
1!
0$
b110 %
1'
0*
b110 +
#746260000000
1"
1(
#746270000000
0!
0"
b100 &
0'
0(
b100 ,
#746280000000
1!
1$
b111 %
1'
1*
b111 +
#746290000000
0!
0'
#746300000000
1!
0$
b1000 %
1'
0*
b1000 +
#746310000000
0!
0'
#746320000000
1!
b1001 %
1'
b1001 +
#746330000000
0!
0'
#746340000000
1!
b0 %
1'
b0 +
#746350000000
0!
0'
#746360000000
1!
1$
b1 %
1'
1*
b1 +
#746370000000
0!
0'
#746380000000
1!
b10 %
1'
b10 +
#746390000000
0!
0'
#746400000000
1!
b11 %
1'
b11 +
#746410000000
0!
0'
#746420000000
1!
b100 %
1'
b100 +
#746430000000
0!
0'
#746440000000
1!
b101 %
1'
b101 +
#746450000000
0!
0'
#746460000000
1!
b110 %
1'
b110 +
#746470000000
0!
0'
#746480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#746490000000
0!
0'
#746500000000
1!
b1000 %
1'
b1000 +
#746510000000
0!
0'
#746520000000
1!
b1001 %
1'
b1001 +
#746530000000
0!
0'
#746540000000
1!
b0 %
1'
b0 +
#746550000000
0!
0'
#746560000000
1!
1$
b1 %
1'
1*
b1 +
#746570000000
0!
0'
#746580000000
1!
b10 %
1'
b10 +
#746590000000
0!
0'
#746600000000
1!
b11 %
1'
b11 +
#746610000000
0!
0'
#746620000000
1!
b100 %
1'
b100 +
#746630000000
0!
0'
#746640000000
1!
b101 %
1'
b101 +
#746650000000
0!
0'
#746660000000
1!
0$
b110 %
1'
0*
b110 +
#746670000000
0!
0'
#746680000000
1!
b111 %
1'
b111 +
#746690000000
1"
1(
#746700000000
0!
0"
b100 &
0'
0(
b100 ,
#746710000000
1!
b1000 %
1'
b1000 +
#746720000000
0!
0'
#746730000000
1!
b1001 %
1'
b1001 +
#746740000000
0!
0'
#746750000000
1!
b0 %
1'
b0 +
#746760000000
0!
0'
#746770000000
1!
1$
b1 %
1'
1*
b1 +
#746780000000
0!
0'
#746790000000
1!
b10 %
1'
b10 +
#746800000000
0!
0'
#746810000000
1!
b11 %
1'
b11 +
#746820000000
0!
0'
#746830000000
1!
b100 %
1'
b100 +
#746840000000
0!
0'
#746850000000
1!
b101 %
1'
b101 +
#746860000000
0!
0'
#746870000000
1!
b110 %
1'
b110 +
#746880000000
0!
0'
#746890000000
1!
b111 %
1'
b111 +
#746900000000
0!
0'
#746910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#746920000000
0!
0'
#746930000000
1!
b1001 %
1'
b1001 +
#746940000000
0!
0'
#746950000000
1!
b0 %
1'
b0 +
#746960000000
0!
0'
#746970000000
1!
1$
b1 %
1'
1*
b1 +
#746980000000
0!
0'
#746990000000
1!
b10 %
1'
b10 +
#747000000000
0!
0'
#747010000000
1!
b11 %
1'
b11 +
#747020000000
0!
0'
#747030000000
1!
b100 %
1'
b100 +
#747040000000
0!
0'
#747050000000
1!
b101 %
1'
b101 +
#747060000000
0!
0'
#747070000000
1!
0$
b110 %
1'
0*
b110 +
#747080000000
0!
0'
#747090000000
1!
b111 %
1'
b111 +
#747100000000
0!
0'
#747110000000
1!
b1000 %
1'
b1000 +
#747120000000
1"
1(
#747130000000
0!
0"
b100 &
0'
0(
b100 ,
#747140000000
1!
b1001 %
1'
b1001 +
#747150000000
0!
0'
#747160000000
1!
b0 %
1'
b0 +
#747170000000
0!
0'
#747180000000
1!
1$
b1 %
1'
1*
b1 +
#747190000000
0!
0'
#747200000000
1!
b10 %
1'
b10 +
#747210000000
0!
0'
#747220000000
1!
b11 %
1'
b11 +
#747230000000
0!
0'
#747240000000
1!
b100 %
1'
b100 +
#747250000000
0!
0'
#747260000000
1!
b101 %
1'
b101 +
#747270000000
0!
0'
#747280000000
1!
b110 %
1'
b110 +
#747290000000
0!
0'
#747300000000
1!
b111 %
1'
b111 +
#747310000000
0!
0'
#747320000000
1!
0$
b1000 %
1'
0*
b1000 +
#747330000000
0!
0'
#747340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#747350000000
0!
0'
#747360000000
1!
b0 %
1'
b0 +
#747370000000
0!
0'
#747380000000
1!
1$
b1 %
1'
1*
b1 +
#747390000000
0!
0'
#747400000000
1!
b10 %
1'
b10 +
#747410000000
0!
0'
#747420000000
1!
b11 %
1'
b11 +
#747430000000
0!
0'
#747440000000
1!
b100 %
1'
b100 +
#747450000000
0!
0'
#747460000000
1!
b101 %
1'
b101 +
#747470000000
0!
0'
#747480000000
1!
0$
b110 %
1'
0*
b110 +
#747490000000
0!
0'
#747500000000
1!
b111 %
1'
b111 +
#747510000000
0!
0'
#747520000000
1!
b1000 %
1'
b1000 +
#747530000000
0!
0'
#747540000000
1!
b1001 %
1'
b1001 +
#747550000000
1"
1(
#747560000000
0!
0"
b100 &
0'
0(
b100 ,
#747570000000
1!
b0 %
1'
b0 +
#747580000000
0!
0'
#747590000000
1!
1$
b1 %
1'
1*
b1 +
#747600000000
0!
0'
#747610000000
1!
b10 %
1'
b10 +
#747620000000
0!
0'
#747630000000
1!
b11 %
1'
b11 +
#747640000000
0!
0'
#747650000000
1!
b100 %
1'
b100 +
#747660000000
0!
0'
#747670000000
1!
b101 %
1'
b101 +
#747680000000
0!
0'
#747690000000
1!
b110 %
1'
b110 +
#747700000000
0!
0'
#747710000000
1!
b111 %
1'
b111 +
#747720000000
0!
0'
#747730000000
1!
0$
b1000 %
1'
0*
b1000 +
#747740000000
0!
0'
#747750000000
1!
b1001 %
1'
b1001 +
#747760000000
0!
0'
#747770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#747780000000
0!
0'
#747790000000
1!
1$
b1 %
1'
1*
b1 +
#747800000000
0!
0'
#747810000000
1!
b10 %
1'
b10 +
#747820000000
0!
0'
#747830000000
1!
b11 %
1'
b11 +
#747840000000
0!
0'
#747850000000
1!
b100 %
1'
b100 +
#747860000000
0!
0'
#747870000000
1!
b101 %
1'
b101 +
#747880000000
0!
0'
#747890000000
1!
0$
b110 %
1'
0*
b110 +
#747900000000
0!
0'
#747910000000
1!
b111 %
1'
b111 +
#747920000000
0!
0'
#747930000000
1!
b1000 %
1'
b1000 +
#747940000000
0!
0'
#747950000000
1!
b1001 %
1'
b1001 +
#747960000000
0!
0'
#747970000000
1!
b0 %
1'
b0 +
#747980000000
1"
1(
#747990000000
0!
0"
b100 &
0'
0(
b100 ,
#748000000000
1!
1$
b1 %
1'
1*
b1 +
#748010000000
0!
0'
#748020000000
1!
b10 %
1'
b10 +
#748030000000
0!
0'
#748040000000
1!
b11 %
1'
b11 +
#748050000000
0!
0'
#748060000000
1!
b100 %
1'
b100 +
#748070000000
0!
0'
#748080000000
1!
b101 %
1'
b101 +
#748090000000
0!
0'
#748100000000
1!
b110 %
1'
b110 +
#748110000000
0!
0'
#748120000000
1!
b111 %
1'
b111 +
#748130000000
0!
0'
#748140000000
1!
0$
b1000 %
1'
0*
b1000 +
#748150000000
0!
0'
#748160000000
1!
b1001 %
1'
b1001 +
#748170000000
0!
0'
#748180000000
1!
b0 %
1'
b0 +
#748190000000
0!
0'
#748200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#748210000000
0!
0'
#748220000000
1!
b10 %
1'
b10 +
#748230000000
0!
0'
#748240000000
1!
b11 %
1'
b11 +
#748250000000
0!
0'
#748260000000
1!
b100 %
1'
b100 +
#748270000000
0!
0'
#748280000000
1!
b101 %
1'
b101 +
#748290000000
0!
0'
#748300000000
1!
0$
b110 %
1'
0*
b110 +
#748310000000
0!
0'
#748320000000
1!
b111 %
1'
b111 +
#748330000000
0!
0'
#748340000000
1!
b1000 %
1'
b1000 +
#748350000000
0!
0'
#748360000000
1!
b1001 %
1'
b1001 +
#748370000000
0!
0'
#748380000000
1!
b0 %
1'
b0 +
#748390000000
0!
0'
#748400000000
1!
1$
b1 %
1'
1*
b1 +
#748410000000
1"
1(
#748420000000
0!
0"
b100 &
0'
0(
b100 ,
#748430000000
1!
b10 %
1'
b10 +
#748440000000
0!
0'
#748450000000
1!
b11 %
1'
b11 +
#748460000000
0!
0'
#748470000000
1!
b100 %
1'
b100 +
#748480000000
0!
0'
#748490000000
1!
b101 %
1'
b101 +
#748500000000
0!
0'
#748510000000
1!
b110 %
1'
b110 +
#748520000000
0!
0'
#748530000000
1!
b111 %
1'
b111 +
#748540000000
0!
0'
#748550000000
1!
0$
b1000 %
1'
0*
b1000 +
#748560000000
0!
0'
#748570000000
1!
b1001 %
1'
b1001 +
#748580000000
0!
0'
#748590000000
1!
b0 %
1'
b0 +
#748600000000
0!
0'
#748610000000
1!
1$
b1 %
1'
1*
b1 +
#748620000000
0!
0'
#748630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#748640000000
0!
0'
#748650000000
1!
b11 %
1'
b11 +
#748660000000
0!
0'
#748670000000
1!
b100 %
1'
b100 +
#748680000000
0!
0'
#748690000000
1!
b101 %
1'
b101 +
#748700000000
0!
0'
#748710000000
1!
0$
b110 %
1'
0*
b110 +
#748720000000
0!
0'
#748730000000
1!
b111 %
1'
b111 +
#748740000000
0!
0'
#748750000000
1!
b1000 %
1'
b1000 +
#748760000000
0!
0'
#748770000000
1!
b1001 %
1'
b1001 +
#748780000000
0!
0'
#748790000000
1!
b0 %
1'
b0 +
#748800000000
0!
0'
#748810000000
1!
1$
b1 %
1'
1*
b1 +
#748820000000
0!
0'
#748830000000
1!
b10 %
1'
b10 +
#748840000000
1"
1(
#748850000000
0!
0"
b100 &
0'
0(
b100 ,
#748860000000
1!
b11 %
1'
b11 +
#748870000000
0!
0'
#748880000000
1!
b100 %
1'
b100 +
#748890000000
0!
0'
#748900000000
1!
b101 %
1'
b101 +
#748910000000
0!
0'
#748920000000
1!
b110 %
1'
b110 +
#748930000000
0!
0'
#748940000000
1!
b111 %
1'
b111 +
#748950000000
0!
0'
#748960000000
1!
0$
b1000 %
1'
0*
b1000 +
#748970000000
0!
0'
#748980000000
1!
b1001 %
1'
b1001 +
#748990000000
0!
0'
#749000000000
1!
b0 %
1'
b0 +
#749010000000
0!
0'
#749020000000
1!
1$
b1 %
1'
1*
b1 +
#749030000000
0!
0'
#749040000000
1!
b10 %
1'
b10 +
#749050000000
0!
0'
#749060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#749070000000
0!
0'
#749080000000
1!
b100 %
1'
b100 +
#749090000000
0!
0'
#749100000000
1!
b101 %
1'
b101 +
#749110000000
0!
0'
#749120000000
1!
0$
b110 %
1'
0*
b110 +
#749130000000
0!
0'
#749140000000
1!
b111 %
1'
b111 +
#749150000000
0!
0'
#749160000000
1!
b1000 %
1'
b1000 +
#749170000000
0!
0'
#749180000000
1!
b1001 %
1'
b1001 +
#749190000000
0!
0'
#749200000000
1!
b0 %
1'
b0 +
#749210000000
0!
0'
#749220000000
1!
1$
b1 %
1'
1*
b1 +
#749230000000
0!
0'
#749240000000
1!
b10 %
1'
b10 +
#749250000000
0!
0'
#749260000000
1!
b11 %
1'
b11 +
#749270000000
1"
1(
#749280000000
0!
0"
b100 &
0'
0(
b100 ,
#749290000000
1!
b100 %
1'
b100 +
#749300000000
0!
0'
#749310000000
1!
b101 %
1'
b101 +
#749320000000
0!
0'
#749330000000
1!
b110 %
1'
b110 +
#749340000000
0!
0'
#749350000000
1!
b111 %
1'
b111 +
#749360000000
0!
0'
#749370000000
1!
0$
b1000 %
1'
0*
b1000 +
#749380000000
0!
0'
#749390000000
1!
b1001 %
1'
b1001 +
#749400000000
0!
0'
#749410000000
1!
b0 %
1'
b0 +
#749420000000
0!
0'
#749430000000
1!
1$
b1 %
1'
1*
b1 +
#749440000000
0!
0'
#749450000000
1!
b10 %
1'
b10 +
#749460000000
0!
0'
#749470000000
1!
b11 %
1'
b11 +
#749480000000
0!
0'
#749490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#749500000000
0!
0'
#749510000000
1!
b101 %
1'
b101 +
#749520000000
0!
0'
#749530000000
1!
0$
b110 %
1'
0*
b110 +
#749540000000
0!
0'
#749550000000
1!
b111 %
1'
b111 +
#749560000000
0!
0'
#749570000000
1!
b1000 %
1'
b1000 +
#749580000000
0!
0'
#749590000000
1!
b1001 %
1'
b1001 +
#749600000000
0!
0'
#749610000000
1!
b0 %
1'
b0 +
#749620000000
0!
0'
#749630000000
1!
1$
b1 %
1'
1*
b1 +
#749640000000
0!
0'
#749650000000
1!
b10 %
1'
b10 +
#749660000000
0!
0'
#749670000000
1!
b11 %
1'
b11 +
#749680000000
0!
0'
#749690000000
1!
b100 %
1'
b100 +
#749700000000
1"
1(
#749710000000
0!
0"
b100 &
0'
0(
b100 ,
#749720000000
1!
b101 %
1'
b101 +
#749730000000
0!
0'
#749740000000
1!
b110 %
1'
b110 +
#749750000000
0!
0'
#749760000000
1!
b111 %
1'
b111 +
#749770000000
0!
0'
#749780000000
1!
0$
b1000 %
1'
0*
b1000 +
#749790000000
0!
0'
#749800000000
1!
b1001 %
1'
b1001 +
#749810000000
0!
0'
#749820000000
1!
b0 %
1'
b0 +
#749830000000
0!
0'
#749840000000
1!
1$
b1 %
1'
1*
b1 +
#749850000000
0!
0'
#749860000000
1!
b10 %
1'
b10 +
#749870000000
0!
0'
#749880000000
1!
b11 %
1'
b11 +
#749890000000
0!
0'
#749900000000
1!
b100 %
1'
b100 +
#749910000000
0!
0'
#749920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#749930000000
0!
0'
#749940000000
1!
0$
b110 %
1'
0*
b110 +
#749950000000
0!
0'
#749960000000
1!
b111 %
1'
b111 +
#749970000000
0!
0'
#749980000000
1!
b1000 %
1'
b1000 +
#749990000000
0!
0'
#750000000000
1!
b1001 %
1'
b1001 +
#750010000000
0!
0'
#750020000000
1!
b0 %
1'
b0 +
#750030000000
0!
0'
#750040000000
1!
1$
b1 %
1'
1*
b1 +
#750050000000
0!
0'
#750060000000
1!
b10 %
1'
b10 +
#750070000000
0!
0'
#750080000000
1!
b11 %
1'
b11 +
#750090000000
0!
0'
#750100000000
1!
b100 %
1'
b100 +
#750110000000
0!
0'
#750120000000
1!
b101 %
1'
b101 +
#750130000000
1"
1(
#750140000000
0!
0"
b100 &
0'
0(
b100 ,
#750150000000
1!
b110 %
1'
b110 +
#750160000000
0!
0'
#750170000000
1!
b111 %
1'
b111 +
#750180000000
0!
0'
#750190000000
1!
0$
b1000 %
1'
0*
b1000 +
#750200000000
0!
0'
#750210000000
1!
b1001 %
1'
b1001 +
#750220000000
0!
0'
#750230000000
1!
b0 %
1'
b0 +
#750240000000
0!
0'
#750250000000
1!
1$
b1 %
1'
1*
b1 +
#750260000000
0!
0'
#750270000000
1!
b10 %
1'
b10 +
#750280000000
0!
0'
#750290000000
1!
b11 %
1'
b11 +
#750300000000
0!
0'
#750310000000
1!
b100 %
1'
b100 +
#750320000000
0!
0'
#750330000000
1!
b101 %
1'
b101 +
#750340000000
0!
0'
#750350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#750360000000
0!
0'
#750370000000
1!
b111 %
1'
b111 +
#750380000000
0!
0'
#750390000000
1!
b1000 %
1'
b1000 +
#750400000000
0!
0'
#750410000000
1!
b1001 %
1'
b1001 +
#750420000000
0!
0'
#750430000000
1!
b0 %
1'
b0 +
#750440000000
0!
0'
#750450000000
1!
1$
b1 %
1'
1*
b1 +
#750460000000
0!
0'
#750470000000
1!
b10 %
1'
b10 +
#750480000000
0!
0'
#750490000000
1!
b11 %
1'
b11 +
#750500000000
0!
0'
#750510000000
1!
b100 %
1'
b100 +
#750520000000
0!
0'
#750530000000
1!
b101 %
1'
b101 +
#750540000000
0!
0'
#750550000000
1!
0$
b110 %
1'
0*
b110 +
#750560000000
1"
1(
#750570000000
0!
0"
b100 &
0'
0(
b100 ,
#750580000000
1!
1$
b111 %
1'
1*
b111 +
#750590000000
0!
0'
#750600000000
1!
0$
b1000 %
1'
0*
b1000 +
#750610000000
0!
0'
#750620000000
1!
b1001 %
1'
b1001 +
#750630000000
0!
0'
#750640000000
1!
b0 %
1'
b0 +
#750650000000
0!
0'
#750660000000
1!
1$
b1 %
1'
1*
b1 +
#750670000000
0!
0'
#750680000000
1!
b10 %
1'
b10 +
#750690000000
0!
0'
#750700000000
1!
b11 %
1'
b11 +
#750710000000
0!
0'
#750720000000
1!
b100 %
1'
b100 +
#750730000000
0!
0'
#750740000000
1!
b101 %
1'
b101 +
#750750000000
0!
0'
#750760000000
1!
b110 %
1'
b110 +
#750770000000
0!
0'
#750780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#750790000000
0!
0'
#750800000000
1!
b1000 %
1'
b1000 +
#750810000000
0!
0'
#750820000000
1!
b1001 %
1'
b1001 +
#750830000000
0!
0'
#750840000000
1!
b0 %
1'
b0 +
#750850000000
0!
0'
#750860000000
1!
1$
b1 %
1'
1*
b1 +
#750870000000
0!
0'
#750880000000
1!
b10 %
1'
b10 +
#750890000000
0!
0'
#750900000000
1!
b11 %
1'
b11 +
#750910000000
0!
0'
#750920000000
1!
b100 %
1'
b100 +
#750930000000
0!
0'
#750940000000
1!
b101 %
1'
b101 +
#750950000000
0!
0'
#750960000000
1!
0$
b110 %
1'
0*
b110 +
#750970000000
0!
0'
#750980000000
1!
b111 %
1'
b111 +
#750990000000
1"
1(
#751000000000
0!
0"
b100 &
0'
0(
b100 ,
#751010000000
1!
b1000 %
1'
b1000 +
#751020000000
0!
0'
#751030000000
1!
b1001 %
1'
b1001 +
#751040000000
0!
0'
#751050000000
1!
b0 %
1'
b0 +
#751060000000
0!
0'
#751070000000
1!
1$
b1 %
1'
1*
b1 +
#751080000000
0!
0'
#751090000000
1!
b10 %
1'
b10 +
#751100000000
0!
0'
#751110000000
1!
b11 %
1'
b11 +
#751120000000
0!
0'
#751130000000
1!
b100 %
1'
b100 +
#751140000000
0!
0'
#751150000000
1!
b101 %
1'
b101 +
#751160000000
0!
0'
#751170000000
1!
b110 %
1'
b110 +
#751180000000
0!
0'
#751190000000
1!
b111 %
1'
b111 +
#751200000000
0!
0'
#751210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#751220000000
0!
0'
#751230000000
1!
b1001 %
1'
b1001 +
#751240000000
0!
0'
#751250000000
1!
b0 %
1'
b0 +
#751260000000
0!
0'
#751270000000
1!
1$
b1 %
1'
1*
b1 +
#751280000000
0!
0'
#751290000000
1!
b10 %
1'
b10 +
#751300000000
0!
0'
#751310000000
1!
b11 %
1'
b11 +
#751320000000
0!
0'
#751330000000
1!
b100 %
1'
b100 +
#751340000000
0!
0'
#751350000000
1!
b101 %
1'
b101 +
#751360000000
0!
0'
#751370000000
1!
0$
b110 %
1'
0*
b110 +
#751380000000
0!
0'
#751390000000
1!
b111 %
1'
b111 +
#751400000000
0!
0'
#751410000000
1!
b1000 %
1'
b1000 +
#751420000000
1"
1(
#751430000000
0!
0"
b100 &
0'
0(
b100 ,
#751440000000
1!
b1001 %
1'
b1001 +
#751450000000
0!
0'
#751460000000
1!
b0 %
1'
b0 +
#751470000000
0!
0'
#751480000000
1!
1$
b1 %
1'
1*
b1 +
#751490000000
0!
0'
#751500000000
1!
b10 %
1'
b10 +
#751510000000
0!
0'
#751520000000
1!
b11 %
1'
b11 +
#751530000000
0!
0'
#751540000000
1!
b100 %
1'
b100 +
#751550000000
0!
0'
#751560000000
1!
b101 %
1'
b101 +
#751570000000
0!
0'
#751580000000
1!
b110 %
1'
b110 +
#751590000000
0!
0'
#751600000000
1!
b111 %
1'
b111 +
#751610000000
0!
0'
#751620000000
1!
0$
b1000 %
1'
0*
b1000 +
#751630000000
0!
0'
#751640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#751650000000
0!
0'
#751660000000
1!
b0 %
1'
b0 +
#751670000000
0!
0'
#751680000000
1!
1$
b1 %
1'
1*
b1 +
#751690000000
0!
0'
#751700000000
1!
b10 %
1'
b10 +
#751710000000
0!
0'
#751720000000
1!
b11 %
1'
b11 +
#751730000000
0!
0'
#751740000000
1!
b100 %
1'
b100 +
#751750000000
0!
0'
#751760000000
1!
b101 %
1'
b101 +
#751770000000
0!
0'
#751780000000
1!
0$
b110 %
1'
0*
b110 +
#751790000000
0!
0'
#751800000000
1!
b111 %
1'
b111 +
#751810000000
0!
0'
#751820000000
1!
b1000 %
1'
b1000 +
#751830000000
0!
0'
#751840000000
1!
b1001 %
1'
b1001 +
#751850000000
1"
1(
#751860000000
0!
0"
b100 &
0'
0(
b100 ,
#751870000000
1!
b0 %
1'
b0 +
#751880000000
0!
0'
#751890000000
1!
1$
b1 %
1'
1*
b1 +
#751900000000
0!
0'
#751910000000
1!
b10 %
1'
b10 +
#751920000000
0!
0'
#751930000000
1!
b11 %
1'
b11 +
#751940000000
0!
0'
#751950000000
1!
b100 %
1'
b100 +
#751960000000
0!
0'
#751970000000
1!
b101 %
1'
b101 +
#751980000000
0!
0'
#751990000000
1!
b110 %
1'
b110 +
#752000000000
0!
0'
#752010000000
1!
b111 %
1'
b111 +
#752020000000
0!
0'
#752030000000
1!
0$
b1000 %
1'
0*
b1000 +
#752040000000
0!
0'
#752050000000
1!
b1001 %
1'
b1001 +
#752060000000
0!
0'
#752070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#752080000000
0!
0'
#752090000000
1!
1$
b1 %
1'
1*
b1 +
#752100000000
0!
0'
#752110000000
1!
b10 %
1'
b10 +
#752120000000
0!
0'
#752130000000
1!
b11 %
1'
b11 +
#752140000000
0!
0'
#752150000000
1!
b100 %
1'
b100 +
#752160000000
0!
0'
#752170000000
1!
b101 %
1'
b101 +
#752180000000
0!
0'
#752190000000
1!
0$
b110 %
1'
0*
b110 +
#752200000000
0!
0'
#752210000000
1!
b111 %
1'
b111 +
#752220000000
0!
0'
#752230000000
1!
b1000 %
1'
b1000 +
#752240000000
0!
0'
#752250000000
1!
b1001 %
1'
b1001 +
#752260000000
0!
0'
#752270000000
1!
b0 %
1'
b0 +
#752280000000
1"
1(
#752290000000
0!
0"
b100 &
0'
0(
b100 ,
#752300000000
1!
1$
b1 %
1'
1*
b1 +
#752310000000
0!
0'
#752320000000
1!
b10 %
1'
b10 +
#752330000000
0!
0'
#752340000000
1!
b11 %
1'
b11 +
#752350000000
0!
0'
#752360000000
1!
b100 %
1'
b100 +
#752370000000
0!
0'
#752380000000
1!
b101 %
1'
b101 +
#752390000000
0!
0'
#752400000000
1!
b110 %
1'
b110 +
#752410000000
0!
0'
#752420000000
1!
b111 %
1'
b111 +
#752430000000
0!
0'
#752440000000
1!
0$
b1000 %
1'
0*
b1000 +
#752450000000
0!
0'
#752460000000
1!
b1001 %
1'
b1001 +
#752470000000
0!
0'
#752480000000
1!
b0 %
1'
b0 +
#752490000000
0!
0'
#752500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#752510000000
0!
0'
#752520000000
1!
b10 %
1'
b10 +
#752530000000
0!
0'
#752540000000
1!
b11 %
1'
b11 +
#752550000000
0!
0'
#752560000000
1!
b100 %
1'
b100 +
#752570000000
0!
0'
#752580000000
1!
b101 %
1'
b101 +
#752590000000
0!
0'
#752600000000
1!
0$
b110 %
1'
0*
b110 +
#752610000000
0!
0'
#752620000000
1!
b111 %
1'
b111 +
#752630000000
0!
0'
#752640000000
1!
b1000 %
1'
b1000 +
#752650000000
0!
0'
#752660000000
1!
b1001 %
1'
b1001 +
#752670000000
0!
0'
#752680000000
1!
b0 %
1'
b0 +
#752690000000
0!
0'
#752700000000
1!
1$
b1 %
1'
1*
b1 +
#752710000000
1"
1(
#752720000000
0!
0"
b100 &
0'
0(
b100 ,
#752730000000
1!
b10 %
1'
b10 +
#752740000000
0!
0'
#752750000000
1!
b11 %
1'
b11 +
#752760000000
0!
0'
#752770000000
1!
b100 %
1'
b100 +
#752780000000
0!
0'
#752790000000
1!
b101 %
1'
b101 +
#752800000000
0!
0'
#752810000000
1!
b110 %
1'
b110 +
#752820000000
0!
0'
#752830000000
1!
b111 %
1'
b111 +
#752840000000
0!
0'
#752850000000
1!
0$
b1000 %
1'
0*
b1000 +
#752860000000
0!
0'
#752870000000
1!
b1001 %
1'
b1001 +
#752880000000
0!
0'
#752890000000
1!
b0 %
1'
b0 +
#752900000000
0!
0'
#752910000000
1!
1$
b1 %
1'
1*
b1 +
#752920000000
0!
0'
#752930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#752940000000
0!
0'
#752950000000
1!
b11 %
1'
b11 +
#752960000000
0!
0'
#752970000000
1!
b100 %
1'
b100 +
#752980000000
0!
0'
#752990000000
1!
b101 %
1'
b101 +
#753000000000
0!
0'
#753010000000
1!
0$
b110 %
1'
0*
b110 +
#753020000000
0!
0'
#753030000000
1!
b111 %
1'
b111 +
#753040000000
0!
0'
#753050000000
1!
b1000 %
1'
b1000 +
#753060000000
0!
0'
#753070000000
1!
b1001 %
1'
b1001 +
#753080000000
0!
0'
#753090000000
1!
b0 %
1'
b0 +
#753100000000
0!
0'
#753110000000
1!
1$
b1 %
1'
1*
b1 +
#753120000000
0!
0'
#753130000000
1!
b10 %
1'
b10 +
#753140000000
1"
1(
#753150000000
0!
0"
b100 &
0'
0(
b100 ,
#753160000000
1!
b11 %
1'
b11 +
#753170000000
0!
0'
#753180000000
1!
b100 %
1'
b100 +
#753190000000
0!
0'
#753200000000
1!
b101 %
1'
b101 +
#753210000000
0!
0'
#753220000000
1!
b110 %
1'
b110 +
#753230000000
0!
0'
#753240000000
1!
b111 %
1'
b111 +
#753250000000
0!
0'
#753260000000
1!
0$
b1000 %
1'
0*
b1000 +
#753270000000
0!
0'
#753280000000
1!
b1001 %
1'
b1001 +
#753290000000
0!
0'
#753300000000
1!
b0 %
1'
b0 +
#753310000000
0!
0'
#753320000000
1!
1$
b1 %
1'
1*
b1 +
#753330000000
0!
0'
#753340000000
1!
b10 %
1'
b10 +
#753350000000
0!
0'
#753360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#753370000000
0!
0'
#753380000000
1!
b100 %
1'
b100 +
#753390000000
0!
0'
#753400000000
1!
b101 %
1'
b101 +
#753410000000
0!
0'
#753420000000
1!
0$
b110 %
1'
0*
b110 +
#753430000000
0!
0'
#753440000000
1!
b111 %
1'
b111 +
#753450000000
0!
0'
#753460000000
1!
b1000 %
1'
b1000 +
#753470000000
0!
0'
#753480000000
1!
b1001 %
1'
b1001 +
#753490000000
0!
0'
#753500000000
1!
b0 %
1'
b0 +
#753510000000
0!
0'
#753520000000
1!
1$
b1 %
1'
1*
b1 +
#753530000000
0!
0'
#753540000000
1!
b10 %
1'
b10 +
#753550000000
0!
0'
#753560000000
1!
b11 %
1'
b11 +
#753570000000
1"
1(
#753580000000
0!
0"
b100 &
0'
0(
b100 ,
#753590000000
1!
b100 %
1'
b100 +
#753600000000
0!
0'
#753610000000
1!
b101 %
1'
b101 +
#753620000000
0!
0'
#753630000000
1!
b110 %
1'
b110 +
#753640000000
0!
0'
#753650000000
1!
b111 %
1'
b111 +
#753660000000
0!
0'
#753670000000
1!
0$
b1000 %
1'
0*
b1000 +
#753680000000
0!
0'
#753690000000
1!
b1001 %
1'
b1001 +
#753700000000
0!
0'
#753710000000
1!
b0 %
1'
b0 +
#753720000000
0!
0'
#753730000000
1!
1$
b1 %
1'
1*
b1 +
#753740000000
0!
0'
#753750000000
1!
b10 %
1'
b10 +
#753760000000
0!
0'
#753770000000
1!
b11 %
1'
b11 +
#753780000000
0!
0'
#753790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#753800000000
0!
0'
#753810000000
1!
b101 %
1'
b101 +
#753820000000
0!
0'
#753830000000
1!
0$
b110 %
1'
0*
b110 +
#753840000000
0!
0'
#753850000000
1!
b111 %
1'
b111 +
#753860000000
0!
0'
#753870000000
1!
b1000 %
1'
b1000 +
#753880000000
0!
0'
#753890000000
1!
b1001 %
1'
b1001 +
#753900000000
0!
0'
#753910000000
1!
b0 %
1'
b0 +
#753920000000
0!
0'
#753930000000
1!
1$
b1 %
1'
1*
b1 +
#753940000000
0!
0'
#753950000000
1!
b10 %
1'
b10 +
#753960000000
0!
0'
#753970000000
1!
b11 %
1'
b11 +
#753980000000
0!
0'
#753990000000
1!
b100 %
1'
b100 +
#754000000000
1"
1(
#754010000000
0!
0"
b100 &
0'
0(
b100 ,
#754020000000
1!
b101 %
1'
b101 +
#754030000000
0!
0'
#754040000000
1!
b110 %
1'
b110 +
#754050000000
0!
0'
#754060000000
1!
b111 %
1'
b111 +
#754070000000
0!
0'
#754080000000
1!
0$
b1000 %
1'
0*
b1000 +
#754090000000
0!
0'
#754100000000
1!
b1001 %
1'
b1001 +
#754110000000
0!
0'
#754120000000
1!
b0 %
1'
b0 +
#754130000000
0!
0'
#754140000000
1!
1$
b1 %
1'
1*
b1 +
#754150000000
0!
0'
#754160000000
1!
b10 %
1'
b10 +
#754170000000
0!
0'
#754180000000
1!
b11 %
1'
b11 +
#754190000000
0!
0'
#754200000000
1!
b100 %
1'
b100 +
#754210000000
0!
0'
#754220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#754230000000
0!
0'
#754240000000
1!
0$
b110 %
1'
0*
b110 +
#754250000000
0!
0'
#754260000000
1!
b111 %
1'
b111 +
#754270000000
0!
0'
#754280000000
1!
b1000 %
1'
b1000 +
#754290000000
0!
0'
#754300000000
1!
b1001 %
1'
b1001 +
#754310000000
0!
0'
#754320000000
1!
b0 %
1'
b0 +
#754330000000
0!
0'
#754340000000
1!
1$
b1 %
1'
1*
b1 +
#754350000000
0!
0'
#754360000000
1!
b10 %
1'
b10 +
#754370000000
0!
0'
#754380000000
1!
b11 %
1'
b11 +
#754390000000
0!
0'
#754400000000
1!
b100 %
1'
b100 +
#754410000000
0!
0'
#754420000000
1!
b101 %
1'
b101 +
#754430000000
1"
1(
#754440000000
0!
0"
b100 &
0'
0(
b100 ,
#754450000000
1!
b110 %
1'
b110 +
#754460000000
0!
0'
#754470000000
1!
b111 %
1'
b111 +
#754480000000
0!
0'
#754490000000
1!
0$
b1000 %
1'
0*
b1000 +
#754500000000
0!
0'
#754510000000
1!
b1001 %
1'
b1001 +
#754520000000
0!
0'
#754530000000
1!
b0 %
1'
b0 +
#754540000000
0!
0'
#754550000000
1!
1$
b1 %
1'
1*
b1 +
#754560000000
0!
0'
#754570000000
1!
b10 %
1'
b10 +
#754580000000
0!
0'
#754590000000
1!
b11 %
1'
b11 +
#754600000000
0!
0'
#754610000000
1!
b100 %
1'
b100 +
#754620000000
0!
0'
#754630000000
1!
b101 %
1'
b101 +
#754640000000
0!
0'
#754650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#754660000000
0!
0'
#754670000000
1!
b111 %
1'
b111 +
#754680000000
0!
0'
#754690000000
1!
b1000 %
1'
b1000 +
#754700000000
0!
0'
#754710000000
1!
b1001 %
1'
b1001 +
#754720000000
0!
0'
#754730000000
1!
b0 %
1'
b0 +
#754740000000
0!
0'
#754750000000
1!
1$
b1 %
1'
1*
b1 +
#754760000000
0!
0'
#754770000000
1!
b10 %
1'
b10 +
#754780000000
0!
0'
#754790000000
1!
b11 %
1'
b11 +
#754800000000
0!
0'
#754810000000
1!
b100 %
1'
b100 +
#754820000000
0!
0'
#754830000000
1!
b101 %
1'
b101 +
#754840000000
0!
0'
#754850000000
1!
0$
b110 %
1'
0*
b110 +
#754860000000
1"
1(
#754870000000
0!
0"
b100 &
0'
0(
b100 ,
#754880000000
1!
1$
b111 %
1'
1*
b111 +
#754890000000
0!
0'
#754900000000
1!
0$
b1000 %
1'
0*
b1000 +
#754910000000
0!
0'
#754920000000
1!
b1001 %
1'
b1001 +
#754930000000
0!
0'
#754940000000
1!
b0 %
1'
b0 +
#754950000000
0!
0'
#754960000000
1!
1$
b1 %
1'
1*
b1 +
#754970000000
0!
0'
#754980000000
1!
b10 %
1'
b10 +
#754990000000
0!
0'
#755000000000
1!
b11 %
1'
b11 +
#755010000000
0!
0'
#755020000000
1!
b100 %
1'
b100 +
#755030000000
0!
0'
#755040000000
1!
b101 %
1'
b101 +
#755050000000
0!
0'
#755060000000
1!
b110 %
1'
b110 +
#755070000000
0!
0'
#755080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#755090000000
0!
0'
#755100000000
1!
b1000 %
1'
b1000 +
#755110000000
0!
0'
#755120000000
1!
b1001 %
1'
b1001 +
#755130000000
0!
0'
#755140000000
1!
b0 %
1'
b0 +
#755150000000
0!
0'
#755160000000
1!
1$
b1 %
1'
1*
b1 +
#755170000000
0!
0'
#755180000000
1!
b10 %
1'
b10 +
#755190000000
0!
0'
#755200000000
1!
b11 %
1'
b11 +
#755210000000
0!
0'
#755220000000
1!
b100 %
1'
b100 +
#755230000000
0!
0'
#755240000000
1!
b101 %
1'
b101 +
#755250000000
0!
0'
#755260000000
1!
0$
b110 %
1'
0*
b110 +
#755270000000
0!
0'
#755280000000
1!
b111 %
1'
b111 +
#755290000000
1"
1(
#755300000000
0!
0"
b100 &
0'
0(
b100 ,
#755310000000
1!
b1000 %
1'
b1000 +
#755320000000
0!
0'
#755330000000
1!
b1001 %
1'
b1001 +
#755340000000
0!
0'
#755350000000
1!
b0 %
1'
b0 +
#755360000000
0!
0'
#755370000000
1!
1$
b1 %
1'
1*
b1 +
#755380000000
0!
0'
#755390000000
1!
b10 %
1'
b10 +
#755400000000
0!
0'
#755410000000
1!
b11 %
1'
b11 +
#755420000000
0!
0'
#755430000000
1!
b100 %
1'
b100 +
#755440000000
0!
0'
#755450000000
1!
b101 %
1'
b101 +
#755460000000
0!
0'
#755470000000
1!
b110 %
1'
b110 +
#755480000000
0!
0'
#755490000000
1!
b111 %
1'
b111 +
#755500000000
0!
0'
#755510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#755520000000
0!
0'
#755530000000
1!
b1001 %
1'
b1001 +
#755540000000
0!
0'
#755550000000
1!
b0 %
1'
b0 +
#755560000000
0!
0'
#755570000000
1!
1$
b1 %
1'
1*
b1 +
#755580000000
0!
0'
#755590000000
1!
b10 %
1'
b10 +
#755600000000
0!
0'
#755610000000
1!
b11 %
1'
b11 +
#755620000000
0!
0'
#755630000000
1!
b100 %
1'
b100 +
#755640000000
0!
0'
#755650000000
1!
b101 %
1'
b101 +
#755660000000
0!
0'
#755670000000
1!
0$
b110 %
1'
0*
b110 +
#755680000000
0!
0'
#755690000000
1!
b111 %
1'
b111 +
#755700000000
0!
0'
#755710000000
1!
b1000 %
1'
b1000 +
#755720000000
1"
1(
#755730000000
0!
0"
b100 &
0'
0(
b100 ,
#755740000000
1!
b1001 %
1'
b1001 +
#755750000000
0!
0'
#755760000000
1!
b0 %
1'
b0 +
#755770000000
0!
0'
#755780000000
1!
1$
b1 %
1'
1*
b1 +
#755790000000
0!
0'
#755800000000
1!
b10 %
1'
b10 +
#755810000000
0!
0'
#755820000000
1!
b11 %
1'
b11 +
#755830000000
0!
0'
#755840000000
1!
b100 %
1'
b100 +
#755850000000
0!
0'
#755860000000
1!
b101 %
1'
b101 +
#755870000000
0!
0'
#755880000000
1!
b110 %
1'
b110 +
#755890000000
0!
0'
#755900000000
1!
b111 %
1'
b111 +
#755910000000
0!
0'
#755920000000
1!
0$
b1000 %
1'
0*
b1000 +
#755930000000
0!
0'
#755940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#755950000000
0!
0'
#755960000000
1!
b0 %
1'
b0 +
#755970000000
0!
0'
#755980000000
1!
1$
b1 %
1'
1*
b1 +
#755990000000
0!
0'
#756000000000
1!
b10 %
1'
b10 +
#756010000000
0!
0'
#756020000000
1!
b11 %
1'
b11 +
#756030000000
0!
0'
#756040000000
1!
b100 %
1'
b100 +
#756050000000
0!
0'
#756060000000
1!
b101 %
1'
b101 +
#756070000000
0!
0'
#756080000000
1!
0$
b110 %
1'
0*
b110 +
#756090000000
0!
0'
#756100000000
1!
b111 %
1'
b111 +
#756110000000
0!
0'
#756120000000
1!
b1000 %
1'
b1000 +
#756130000000
0!
0'
#756140000000
1!
b1001 %
1'
b1001 +
#756150000000
1"
1(
#756160000000
0!
0"
b100 &
0'
0(
b100 ,
#756170000000
1!
b0 %
1'
b0 +
#756180000000
0!
0'
#756190000000
1!
1$
b1 %
1'
1*
b1 +
#756200000000
0!
0'
#756210000000
1!
b10 %
1'
b10 +
#756220000000
0!
0'
#756230000000
1!
b11 %
1'
b11 +
#756240000000
0!
0'
#756250000000
1!
b100 %
1'
b100 +
#756260000000
0!
0'
#756270000000
1!
b101 %
1'
b101 +
#756280000000
0!
0'
#756290000000
1!
b110 %
1'
b110 +
#756300000000
0!
0'
#756310000000
1!
b111 %
1'
b111 +
#756320000000
0!
0'
#756330000000
1!
0$
b1000 %
1'
0*
b1000 +
#756340000000
0!
0'
#756350000000
1!
b1001 %
1'
b1001 +
#756360000000
0!
0'
#756370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#756380000000
0!
0'
#756390000000
1!
1$
b1 %
1'
1*
b1 +
#756400000000
0!
0'
#756410000000
1!
b10 %
1'
b10 +
#756420000000
0!
0'
#756430000000
1!
b11 %
1'
b11 +
#756440000000
0!
0'
#756450000000
1!
b100 %
1'
b100 +
#756460000000
0!
0'
#756470000000
1!
b101 %
1'
b101 +
#756480000000
0!
0'
#756490000000
1!
0$
b110 %
1'
0*
b110 +
#756500000000
0!
0'
#756510000000
1!
b111 %
1'
b111 +
#756520000000
0!
0'
#756530000000
1!
b1000 %
1'
b1000 +
#756540000000
0!
0'
#756550000000
1!
b1001 %
1'
b1001 +
#756560000000
0!
0'
#756570000000
1!
b0 %
1'
b0 +
#756580000000
1"
1(
#756590000000
0!
0"
b100 &
0'
0(
b100 ,
#756600000000
1!
1$
b1 %
1'
1*
b1 +
#756610000000
0!
0'
#756620000000
1!
b10 %
1'
b10 +
#756630000000
0!
0'
#756640000000
1!
b11 %
1'
b11 +
#756650000000
0!
0'
#756660000000
1!
b100 %
1'
b100 +
#756670000000
0!
0'
#756680000000
1!
b101 %
1'
b101 +
#756690000000
0!
0'
#756700000000
1!
b110 %
1'
b110 +
#756710000000
0!
0'
#756720000000
1!
b111 %
1'
b111 +
#756730000000
0!
0'
#756740000000
1!
0$
b1000 %
1'
0*
b1000 +
#756750000000
0!
0'
#756760000000
1!
b1001 %
1'
b1001 +
#756770000000
0!
0'
#756780000000
1!
b0 %
1'
b0 +
#756790000000
0!
0'
#756800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#756810000000
0!
0'
#756820000000
1!
b10 %
1'
b10 +
#756830000000
0!
0'
#756840000000
1!
b11 %
1'
b11 +
#756850000000
0!
0'
#756860000000
1!
b100 %
1'
b100 +
#756870000000
0!
0'
#756880000000
1!
b101 %
1'
b101 +
#756890000000
0!
0'
#756900000000
1!
0$
b110 %
1'
0*
b110 +
#756910000000
0!
0'
#756920000000
1!
b111 %
1'
b111 +
#756930000000
0!
0'
#756940000000
1!
b1000 %
1'
b1000 +
#756950000000
0!
0'
#756960000000
1!
b1001 %
1'
b1001 +
#756970000000
0!
0'
#756980000000
1!
b0 %
1'
b0 +
#756990000000
0!
0'
#757000000000
1!
1$
b1 %
1'
1*
b1 +
#757010000000
1"
1(
#757020000000
0!
0"
b100 &
0'
0(
b100 ,
#757030000000
1!
b10 %
1'
b10 +
#757040000000
0!
0'
#757050000000
1!
b11 %
1'
b11 +
#757060000000
0!
0'
#757070000000
1!
b100 %
1'
b100 +
#757080000000
0!
0'
#757090000000
1!
b101 %
1'
b101 +
#757100000000
0!
0'
#757110000000
1!
b110 %
1'
b110 +
#757120000000
0!
0'
#757130000000
1!
b111 %
1'
b111 +
#757140000000
0!
0'
#757150000000
1!
0$
b1000 %
1'
0*
b1000 +
#757160000000
0!
0'
#757170000000
1!
b1001 %
1'
b1001 +
#757180000000
0!
0'
#757190000000
1!
b0 %
1'
b0 +
#757200000000
0!
0'
#757210000000
1!
1$
b1 %
1'
1*
b1 +
#757220000000
0!
0'
#757230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#757240000000
0!
0'
#757250000000
1!
b11 %
1'
b11 +
#757260000000
0!
0'
#757270000000
1!
b100 %
1'
b100 +
#757280000000
0!
0'
#757290000000
1!
b101 %
1'
b101 +
#757300000000
0!
0'
#757310000000
1!
0$
b110 %
1'
0*
b110 +
#757320000000
0!
0'
#757330000000
1!
b111 %
1'
b111 +
#757340000000
0!
0'
#757350000000
1!
b1000 %
1'
b1000 +
#757360000000
0!
0'
#757370000000
1!
b1001 %
1'
b1001 +
#757380000000
0!
0'
#757390000000
1!
b0 %
1'
b0 +
#757400000000
0!
0'
#757410000000
1!
1$
b1 %
1'
1*
b1 +
#757420000000
0!
0'
#757430000000
1!
b10 %
1'
b10 +
#757440000000
1"
1(
#757450000000
0!
0"
b100 &
0'
0(
b100 ,
#757460000000
1!
b11 %
1'
b11 +
#757470000000
0!
0'
#757480000000
1!
b100 %
1'
b100 +
#757490000000
0!
0'
#757500000000
1!
b101 %
1'
b101 +
#757510000000
0!
0'
#757520000000
1!
b110 %
1'
b110 +
#757530000000
0!
0'
#757540000000
1!
b111 %
1'
b111 +
#757550000000
0!
0'
#757560000000
1!
0$
b1000 %
1'
0*
b1000 +
#757570000000
0!
0'
#757580000000
1!
b1001 %
1'
b1001 +
#757590000000
0!
0'
#757600000000
1!
b0 %
1'
b0 +
#757610000000
0!
0'
#757620000000
1!
1$
b1 %
1'
1*
b1 +
#757630000000
0!
0'
#757640000000
1!
b10 %
1'
b10 +
#757650000000
0!
0'
#757660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#757670000000
0!
0'
#757680000000
1!
b100 %
1'
b100 +
#757690000000
0!
0'
#757700000000
1!
b101 %
1'
b101 +
#757710000000
0!
0'
#757720000000
1!
0$
b110 %
1'
0*
b110 +
#757730000000
0!
0'
#757740000000
1!
b111 %
1'
b111 +
#757750000000
0!
0'
#757760000000
1!
b1000 %
1'
b1000 +
#757770000000
0!
0'
#757780000000
1!
b1001 %
1'
b1001 +
#757790000000
0!
0'
#757800000000
1!
b0 %
1'
b0 +
#757810000000
0!
0'
#757820000000
1!
1$
b1 %
1'
1*
b1 +
#757830000000
0!
0'
#757840000000
1!
b10 %
1'
b10 +
#757850000000
0!
0'
#757860000000
1!
b11 %
1'
b11 +
#757870000000
1"
1(
#757880000000
0!
0"
b100 &
0'
0(
b100 ,
#757890000000
1!
b100 %
1'
b100 +
#757900000000
0!
0'
#757910000000
1!
b101 %
1'
b101 +
#757920000000
0!
0'
#757930000000
1!
b110 %
1'
b110 +
#757940000000
0!
0'
#757950000000
1!
b111 %
1'
b111 +
#757960000000
0!
0'
#757970000000
1!
0$
b1000 %
1'
0*
b1000 +
#757980000000
0!
0'
#757990000000
1!
b1001 %
1'
b1001 +
#758000000000
0!
0'
#758010000000
1!
b0 %
1'
b0 +
#758020000000
0!
0'
#758030000000
1!
1$
b1 %
1'
1*
b1 +
#758040000000
0!
0'
#758050000000
1!
b10 %
1'
b10 +
#758060000000
0!
0'
#758070000000
1!
b11 %
1'
b11 +
#758080000000
0!
0'
#758090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#758100000000
0!
0'
#758110000000
1!
b101 %
1'
b101 +
#758120000000
0!
0'
#758130000000
1!
0$
b110 %
1'
0*
b110 +
#758140000000
0!
0'
#758150000000
1!
b111 %
1'
b111 +
#758160000000
0!
0'
#758170000000
1!
b1000 %
1'
b1000 +
#758180000000
0!
0'
#758190000000
1!
b1001 %
1'
b1001 +
#758200000000
0!
0'
#758210000000
1!
b0 %
1'
b0 +
#758220000000
0!
0'
#758230000000
1!
1$
b1 %
1'
1*
b1 +
#758240000000
0!
0'
#758250000000
1!
b10 %
1'
b10 +
#758260000000
0!
0'
#758270000000
1!
b11 %
1'
b11 +
#758280000000
0!
0'
#758290000000
1!
b100 %
1'
b100 +
#758300000000
1"
1(
#758310000000
0!
0"
b100 &
0'
0(
b100 ,
#758320000000
1!
b101 %
1'
b101 +
#758330000000
0!
0'
#758340000000
1!
b110 %
1'
b110 +
#758350000000
0!
0'
#758360000000
1!
b111 %
1'
b111 +
#758370000000
0!
0'
#758380000000
1!
0$
b1000 %
1'
0*
b1000 +
#758390000000
0!
0'
#758400000000
1!
b1001 %
1'
b1001 +
#758410000000
0!
0'
#758420000000
1!
b0 %
1'
b0 +
#758430000000
0!
0'
#758440000000
1!
1$
b1 %
1'
1*
b1 +
#758450000000
0!
0'
#758460000000
1!
b10 %
1'
b10 +
#758470000000
0!
0'
#758480000000
1!
b11 %
1'
b11 +
#758490000000
0!
0'
#758500000000
1!
b100 %
1'
b100 +
#758510000000
0!
0'
#758520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#758530000000
0!
0'
#758540000000
1!
0$
b110 %
1'
0*
b110 +
#758550000000
0!
0'
#758560000000
1!
b111 %
1'
b111 +
#758570000000
0!
0'
#758580000000
1!
b1000 %
1'
b1000 +
#758590000000
0!
0'
#758600000000
1!
b1001 %
1'
b1001 +
#758610000000
0!
0'
#758620000000
1!
b0 %
1'
b0 +
#758630000000
0!
0'
#758640000000
1!
1$
b1 %
1'
1*
b1 +
#758650000000
0!
0'
#758660000000
1!
b10 %
1'
b10 +
#758670000000
0!
0'
#758680000000
1!
b11 %
1'
b11 +
#758690000000
0!
0'
#758700000000
1!
b100 %
1'
b100 +
#758710000000
0!
0'
#758720000000
1!
b101 %
1'
b101 +
#758730000000
1"
1(
#758740000000
0!
0"
b100 &
0'
0(
b100 ,
#758750000000
1!
b110 %
1'
b110 +
#758760000000
0!
0'
#758770000000
1!
b111 %
1'
b111 +
#758780000000
0!
0'
#758790000000
1!
0$
b1000 %
1'
0*
b1000 +
#758800000000
0!
0'
#758810000000
1!
b1001 %
1'
b1001 +
#758820000000
0!
0'
#758830000000
1!
b0 %
1'
b0 +
#758840000000
0!
0'
#758850000000
1!
1$
b1 %
1'
1*
b1 +
#758860000000
0!
0'
#758870000000
1!
b10 %
1'
b10 +
#758880000000
0!
0'
#758890000000
1!
b11 %
1'
b11 +
#758900000000
0!
0'
#758910000000
1!
b100 %
1'
b100 +
#758920000000
0!
0'
#758930000000
1!
b101 %
1'
b101 +
#758940000000
0!
0'
#758950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#758960000000
0!
0'
#758970000000
1!
b111 %
1'
b111 +
#758980000000
0!
0'
#758990000000
1!
b1000 %
1'
b1000 +
#759000000000
0!
0'
#759010000000
1!
b1001 %
1'
b1001 +
#759020000000
0!
0'
#759030000000
1!
b0 %
1'
b0 +
#759040000000
0!
0'
#759050000000
1!
1$
b1 %
1'
1*
b1 +
#759060000000
0!
0'
#759070000000
1!
b10 %
1'
b10 +
#759080000000
0!
0'
#759090000000
1!
b11 %
1'
b11 +
#759100000000
0!
0'
#759110000000
1!
b100 %
1'
b100 +
#759120000000
0!
0'
#759130000000
1!
b101 %
1'
b101 +
#759140000000
0!
0'
#759150000000
1!
0$
b110 %
1'
0*
b110 +
#759160000000
1"
1(
#759170000000
0!
0"
b100 &
0'
0(
b100 ,
#759180000000
1!
1$
b111 %
1'
1*
b111 +
#759190000000
0!
0'
#759200000000
1!
0$
b1000 %
1'
0*
b1000 +
#759210000000
0!
0'
#759220000000
1!
b1001 %
1'
b1001 +
#759230000000
0!
0'
#759240000000
1!
b0 %
1'
b0 +
#759250000000
0!
0'
#759260000000
1!
1$
b1 %
1'
1*
b1 +
#759270000000
0!
0'
#759280000000
1!
b10 %
1'
b10 +
#759290000000
0!
0'
#759300000000
1!
b11 %
1'
b11 +
#759310000000
0!
0'
#759320000000
1!
b100 %
1'
b100 +
#759330000000
0!
0'
#759340000000
1!
b101 %
1'
b101 +
#759350000000
0!
0'
#759360000000
1!
b110 %
1'
b110 +
#759370000000
0!
0'
#759380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#759390000000
0!
0'
#759400000000
1!
b1000 %
1'
b1000 +
#759410000000
0!
0'
#759420000000
1!
b1001 %
1'
b1001 +
#759430000000
0!
0'
#759440000000
1!
b0 %
1'
b0 +
#759450000000
0!
0'
#759460000000
1!
1$
b1 %
1'
1*
b1 +
#759470000000
0!
0'
#759480000000
1!
b10 %
1'
b10 +
#759490000000
0!
0'
#759500000000
1!
b11 %
1'
b11 +
#759510000000
0!
0'
#759520000000
1!
b100 %
1'
b100 +
#759530000000
0!
0'
#759540000000
1!
b101 %
1'
b101 +
#759550000000
0!
0'
#759560000000
1!
0$
b110 %
1'
0*
b110 +
#759570000000
0!
0'
#759580000000
1!
b111 %
1'
b111 +
#759590000000
1"
1(
#759600000000
0!
0"
b100 &
0'
0(
b100 ,
#759610000000
1!
b1000 %
1'
b1000 +
#759620000000
0!
0'
#759630000000
1!
b1001 %
1'
b1001 +
#759640000000
0!
0'
#759650000000
1!
b0 %
1'
b0 +
#759660000000
0!
0'
#759670000000
1!
1$
b1 %
1'
1*
b1 +
#759680000000
0!
0'
#759690000000
1!
b10 %
1'
b10 +
#759700000000
0!
0'
#759710000000
1!
b11 %
1'
b11 +
#759720000000
0!
0'
#759730000000
1!
b100 %
1'
b100 +
#759740000000
0!
0'
#759750000000
1!
b101 %
1'
b101 +
#759760000000
0!
0'
#759770000000
1!
b110 %
1'
b110 +
#759780000000
0!
0'
#759790000000
1!
b111 %
1'
b111 +
#759800000000
0!
0'
#759810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#759820000000
0!
0'
#759830000000
1!
b1001 %
1'
b1001 +
#759840000000
0!
0'
#759850000000
1!
b0 %
1'
b0 +
#759860000000
0!
0'
#759870000000
1!
1$
b1 %
1'
1*
b1 +
#759880000000
0!
0'
#759890000000
1!
b10 %
1'
b10 +
#759900000000
0!
0'
#759910000000
1!
b11 %
1'
b11 +
#759920000000
0!
0'
#759930000000
1!
b100 %
1'
b100 +
#759940000000
0!
0'
#759950000000
1!
b101 %
1'
b101 +
#759960000000
0!
0'
#759970000000
1!
0$
b110 %
1'
0*
b110 +
#759980000000
0!
0'
#759990000000
1!
b111 %
1'
b111 +
#760000000000
0!
0'
#760010000000
1!
b1000 %
1'
b1000 +
#760020000000
1"
1(
#760030000000
0!
0"
b100 &
0'
0(
b100 ,
#760040000000
1!
b1001 %
1'
b1001 +
#760050000000
0!
0'
#760060000000
1!
b0 %
1'
b0 +
#760070000000
0!
0'
#760080000000
1!
1$
b1 %
1'
1*
b1 +
#760090000000
0!
0'
#760100000000
1!
b10 %
1'
b10 +
#760110000000
0!
0'
#760120000000
1!
b11 %
1'
b11 +
#760130000000
0!
0'
#760140000000
1!
b100 %
1'
b100 +
#760150000000
0!
0'
#760160000000
1!
b101 %
1'
b101 +
#760170000000
0!
0'
#760180000000
1!
b110 %
1'
b110 +
#760190000000
0!
0'
#760200000000
1!
b111 %
1'
b111 +
#760210000000
0!
0'
#760220000000
1!
0$
b1000 %
1'
0*
b1000 +
#760230000000
0!
0'
#760240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#760250000000
0!
0'
#760260000000
1!
b0 %
1'
b0 +
#760270000000
0!
0'
#760280000000
1!
1$
b1 %
1'
1*
b1 +
#760290000000
0!
0'
#760300000000
1!
b10 %
1'
b10 +
#760310000000
0!
0'
#760320000000
1!
b11 %
1'
b11 +
#760330000000
0!
0'
#760340000000
1!
b100 %
1'
b100 +
#760350000000
0!
0'
#760360000000
1!
b101 %
1'
b101 +
#760370000000
0!
0'
#760380000000
1!
0$
b110 %
1'
0*
b110 +
#760390000000
0!
0'
#760400000000
1!
b111 %
1'
b111 +
#760410000000
0!
0'
#760420000000
1!
b1000 %
1'
b1000 +
#760430000000
0!
0'
#760440000000
1!
b1001 %
1'
b1001 +
#760450000000
1"
1(
#760460000000
0!
0"
b100 &
0'
0(
b100 ,
#760470000000
1!
b0 %
1'
b0 +
#760480000000
0!
0'
#760490000000
1!
1$
b1 %
1'
1*
b1 +
#760500000000
0!
0'
#760510000000
1!
b10 %
1'
b10 +
#760520000000
0!
0'
#760530000000
1!
b11 %
1'
b11 +
#760540000000
0!
0'
#760550000000
1!
b100 %
1'
b100 +
#760560000000
0!
0'
#760570000000
1!
b101 %
1'
b101 +
#760580000000
0!
0'
#760590000000
1!
b110 %
1'
b110 +
#760600000000
0!
0'
#760610000000
1!
b111 %
1'
b111 +
#760620000000
0!
0'
#760630000000
1!
0$
b1000 %
1'
0*
b1000 +
#760640000000
0!
0'
#760650000000
1!
b1001 %
1'
b1001 +
#760660000000
0!
0'
#760670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#760680000000
0!
0'
#760690000000
1!
1$
b1 %
1'
1*
b1 +
#760700000000
0!
0'
#760710000000
1!
b10 %
1'
b10 +
#760720000000
0!
0'
#760730000000
1!
b11 %
1'
b11 +
#760740000000
0!
0'
#760750000000
1!
b100 %
1'
b100 +
#760760000000
0!
0'
#760770000000
1!
b101 %
1'
b101 +
#760780000000
0!
0'
#760790000000
1!
0$
b110 %
1'
0*
b110 +
#760800000000
0!
0'
#760810000000
1!
b111 %
1'
b111 +
#760820000000
0!
0'
#760830000000
1!
b1000 %
1'
b1000 +
#760840000000
0!
0'
#760850000000
1!
b1001 %
1'
b1001 +
#760860000000
0!
0'
#760870000000
1!
b0 %
1'
b0 +
#760880000000
1"
1(
#760890000000
0!
0"
b100 &
0'
0(
b100 ,
#760900000000
1!
1$
b1 %
1'
1*
b1 +
#760910000000
0!
0'
#760920000000
1!
b10 %
1'
b10 +
#760930000000
0!
0'
#760940000000
1!
b11 %
1'
b11 +
#760950000000
0!
0'
#760960000000
1!
b100 %
1'
b100 +
#760970000000
0!
0'
#760980000000
1!
b101 %
1'
b101 +
#760990000000
0!
0'
#761000000000
1!
b110 %
1'
b110 +
#761010000000
0!
0'
#761020000000
1!
b111 %
1'
b111 +
#761030000000
0!
0'
#761040000000
1!
0$
b1000 %
1'
0*
b1000 +
#761050000000
0!
0'
#761060000000
1!
b1001 %
1'
b1001 +
#761070000000
0!
0'
#761080000000
1!
b0 %
1'
b0 +
#761090000000
0!
0'
#761100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#761110000000
0!
0'
#761120000000
1!
b10 %
1'
b10 +
#761130000000
0!
0'
#761140000000
1!
b11 %
1'
b11 +
#761150000000
0!
0'
#761160000000
1!
b100 %
1'
b100 +
#761170000000
0!
0'
#761180000000
1!
b101 %
1'
b101 +
#761190000000
0!
0'
#761200000000
1!
0$
b110 %
1'
0*
b110 +
#761210000000
0!
0'
#761220000000
1!
b111 %
1'
b111 +
#761230000000
0!
0'
#761240000000
1!
b1000 %
1'
b1000 +
#761250000000
0!
0'
#761260000000
1!
b1001 %
1'
b1001 +
#761270000000
0!
0'
#761280000000
1!
b0 %
1'
b0 +
#761290000000
0!
0'
#761300000000
1!
1$
b1 %
1'
1*
b1 +
#761310000000
1"
1(
#761320000000
0!
0"
b100 &
0'
0(
b100 ,
#761330000000
1!
b10 %
1'
b10 +
#761340000000
0!
0'
#761350000000
1!
b11 %
1'
b11 +
#761360000000
0!
0'
#761370000000
1!
b100 %
1'
b100 +
#761380000000
0!
0'
#761390000000
1!
b101 %
1'
b101 +
#761400000000
0!
0'
#761410000000
1!
b110 %
1'
b110 +
#761420000000
0!
0'
#761430000000
1!
b111 %
1'
b111 +
#761440000000
0!
0'
#761450000000
1!
0$
b1000 %
1'
0*
b1000 +
#761460000000
0!
0'
#761470000000
1!
b1001 %
1'
b1001 +
#761480000000
0!
0'
#761490000000
1!
b0 %
1'
b0 +
#761500000000
0!
0'
#761510000000
1!
1$
b1 %
1'
1*
b1 +
#761520000000
0!
0'
#761530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#761540000000
0!
0'
#761550000000
1!
b11 %
1'
b11 +
#761560000000
0!
0'
#761570000000
1!
b100 %
1'
b100 +
#761580000000
0!
0'
#761590000000
1!
b101 %
1'
b101 +
#761600000000
0!
0'
#761610000000
1!
0$
b110 %
1'
0*
b110 +
#761620000000
0!
0'
#761630000000
1!
b111 %
1'
b111 +
#761640000000
0!
0'
#761650000000
1!
b1000 %
1'
b1000 +
#761660000000
0!
0'
#761670000000
1!
b1001 %
1'
b1001 +
#761680000000
0!
0'
#761690000000
1!
b0 %
1'
b0 +
#761700000000
0!
0'
#761710000000
1!
1$
b1 %
1'
1*
b1 +
#761720000000
0!
0'
#761730000000
1!
b10 %
1'
b10 +
#761740000000
1"
1(
#761750000000
0!
0"
b100 &
0'
0(
b100 ,
#761760000000
1!
b11 %
1'
b11 +
#761770000000
0!
0'
#761780000000
1!
b100 %
1'
b100 +
#761790000000
0!
0'
#761800000000
1!
b101 %
1'
b101 +
#761810000000
0!
0'
#761820000000
1!
b110 %
1'
b110 +
#761830000000
0!
0'
#761840000000
1!
b111 %
1'
b111 +
#761850000000
0!
0'
#761860000000
1!
0$
b1000 %
1'
0*
b1000 +
#761870000000
0!
0'
#761880000000
1!
b1001 %
1'
b1001 +
#761890000000
0!
0'
#761900000000
1!
b0 %
1'
b0 +
#761910000000
0!
0'
#761920000000
1!
1$
b1 %
1'
1*
b1 +
#761930000000
0!
0'
#761940000000
1!
b10 %
1'
b10 +
#761950000000
0!
0'
#761960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#761970000000
0!
0'
#761980000000
1!
b100 %
1'
b100 +
#761990000000
0!
0'
#762000000000
1!
b101 %
1'
b101 +
#762010000000
0!
0'
#762020000000
1!
0$
b110 %
1'
0*
b110 +
#762030000000
0!
0'
#762040000000
1!
b111 %
1'
b111 +
#762050000000
0!
0'
#762060000000
1!
b1000 %
1'
b1000 +
#762070000000
0!
0'
#762080000000
1!
b1001 %
1'
b1001 +
#762090000000
0!
0'
#762100000000
1!
b0 %
1'
b0 +
#762110000000
0!
0'
#762120000000
1!
1$
b1 %
1'
1*
b1 +
#762130000000
0!
0'
#762140000000
1!
b10 %
1'
b10 +
#762150000000
0!
0'
#762160000000
1!
b11 %
1'
b11 +
#762170000000
1"
1(
#762180000000
0!
0"
b100 &
0'
0(
b100 ,
#762190000000
1!
b100 %
1'
b100 +
#762200000000
0!
0'
#762210000000
1!
b101 %
1'
b101 +
#762220000000
0!
0'
#762230000000
1!
b110 %
1'
b110 +
#762240000000
0!
0'
#762250000000
1!
b111 %
1'
b111 +
#762260000000
0!
0'
#762270000000
1!
0$
b1000 %
1'
0*
b1000 +
#762280000000
0!
0'
#762290000000
1!
b1001 %
1'
b1001 +
#762300000000
0!
0'
#762310000000
1!
b0 %
1'
b0 +
#762320000000
0!
0'
#762330000000
1!
1$
b1 %
1'
1*
b1 +
#762340000000
0!
0'
#762350000000
1!
b10 %
1'
b10 +
#762360000000
0!
0'
#762370000000
1!
b11 %
1'
b11 +
#762380000000
0!
0'
#762390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#762400000000
0!
0'
#762410000000
1!
b101 %
1'
b101 +
#762420000000
0!
0'
#762430000000
1!
0$
b110 %
1'
0*
b110 +
#762440000000
0!
0'
#762450000000
1!
b111 %
1'
b111 +
#762460000000
0!
0'
#762470000000
1!
b1000 %
1'
b1000 +
#762480000000
0!
0'
#762490000000
1!
b1001 %
1'
b1001 +
#762500000000
0!
0'
#762510000000
1!
b0 %
1'
b0 +
#762520000000
0!
0'
#762530000000
1!
1$
b1 %
1'
1*
b1 +
#762540000000
0!
0'
#762550000000
1!
b10 %
1'
b10 +
#762560000000
0!
0'
#762570000000
1!
b11 %
1'
b11 +
#762580000000
0!
0'
#762590000000
1!
b100 %
1'
b100 +
#762600000000
1"
1(
#762610000000
0!
0"
b100 &
0'
0(
b100 ,
#762620000000
1!
b101 %
1'
b101 +
#762630000000
0!
0'
#762640000000
1!
b110 %
1'
b110 +
#762650000000
0!
0'
#762660000000
1!
b111 %
1'
b111 +
#762670000000
0!
0'
#762680000000
1!
0$
b1000 %
1'
0*
b1000 +
#762690000000
0!
0'
#762700000000
1!
b1001 %
1'
b1001 +
#762710000000
0!
0'
#762720000000
1!
b0 %
1'
b0 +
#762730000000
0!
0'
#762740000000
1!
1$
b1 %
1'
1*
b1 +
#762750000000
0!
0'
#762760000000
1!
b10 %
1'
b10 +
#762770000000
0!
0'
#762780000000
1!
b11 %
1'
b11 +
#762790000000
0!
0'
#762800000000
1!
b100 %
1'
b100 +
#762810000000
0!
0'
#762820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#762830000000
0!
0'
#762840000000
1!
0$
b110 %
1'
0*
b110 +
#762850000000
0!
0'
#762860000000
1!
b111 %
1'
b111 +
#762870000000
0!
0'
#762880000000
1!
b1000 %
1'
b1000 +
#762890000000
0!
0'
#762900000000
1!
b1001 %
1'
b1001 +
#762910000000
0!
0'
#762920000000
1!
b0 %
1'
b0 +
#762930000000
0!
0'
#762940000000
1!
1$
b1 %
1'
1*
b1 +
#762950000000
0!
0'
#762960000000
1!
b10 %
1'
b10 +
#762970000000
0!
0'
#762980000000
1!
b11 %
1'
b11 +
#762990000000
0!
0'
#763000000000
1!
b100 %
1'
b100 +
#763010000000
0!
0'
#763020000000
1!
b101 %
1'
b101 +
#763030000000
1"
1(
#763040000000
0!
0"
b100 &
0'
0(
b100 ,
#763050000000
1!
b110 %
1'
b110 +
#763060000000
0!
0'
#763070000000
1!
b111 %
1'
b111 +
#763080000000
0!
0'
#763090000000
1!
0$
b1000 %
1'
0*
b1000 +
#763100000000
0!
0'
#763110000000
1!
b1001 %
1'
b1001 +
#763120000000
0!
0'
#763130000000
1!
b0 %
1'
b0 +
#763140000000
0!
0'
#763150000000
1!
1$
b1 %
1'
1*
b1 +
#763160000000
0!
0'
#763170000000
1!
b10 %
1'
b10 +
#763180000000
0!
0'
#763190000000
1!
b11 %
1'
b11 +
#763200000000
0!
0'
#763210000000
1!
b100 %
1'
b100 +
#763220000000
0!
0'
#763230000000
1!
b101 %
1'
b101 +
#763240000000
0!
0'
#763250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#763260000000
0!
0'
#763270000000
1!
b111 %
1'
b111 +
#763280000000
0!
0'
#763290000000
1!
b1000 %
1'
b1000 +
#763300000000
0!
0'
#763310000000
1!
b1001 %
1'
b1001 +
#763320000000
0!
0'
#763330000000
1!
b0 %
1'
b0 +
#763340000000
0!
0'
#763350000000
1!
1$
b1 %
1'
1*
b1 +
#763360000000
0!
0'
#763370000000
1!
b10 %
1'
b10 +
#763380000000
0!
0'
#763390000000
1!
b11 %
1'
b11 +
#763400000000
0!
0'
#763410000000
1!
b100 %
1'
b100 +
#763420000000
0!
0'
#763430000000
1!
b101 %
1'
b101 +
#763440000000
0!
0'
#763450000000
1!
0$
b110 %
1'
0*
b110 +
#763460000000
1"
1(
#763470000000
0!
0"
b100 &
0'
0(
b100 ,
#763480000000
1!
1$
b111 %
1'
1*
b111 +
#763490000000
0!
0'
#763500000000
1!
0$
b1000 %
1'
0*
b1000 +
#763510000000
0!
0'
#763520000000
1!
b1001 %
1'
b1001 +
#763530000000
0!
0'
#763540000000
1!
b0 %
1'
b0 +
#763550000000
0!
0'
#763560000000
1!
1$
b1 %
1'
1*
b1 +
#763570000000
0!
0'
#763580000000
1!
b10 %
1'
b10 +
#763590000000
0!
0'
#763600000000
1!
b11 %
1'
b11 +
#763610000000
0!
0'
#763620000000
1!
b100 %
1'
b100 +
#763630000000
0!
0'
#763640000000
1!
b101 %
1'
b101 +
#763650000000
0!
0'
#763660000000
1!
b110 %
1'
b110 +
#763670000000
0!
0'
#763680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#763690000000
0!
0'
#763700000000
1!
b1000 %
1'
b1000 +
#763710000000
0!
0'
#763720000000
1!
b1001 %
1'
b1001 +
#763730000000
0!
0'
#763740000000
1!
b0 %
1'
b0 +
#763750000000
0!
0'
#763760000000
1!
1$
b1 %
1'
1*
b1 +
#763770000000
0!
0'
#763780000000
1!
b10 %
1'
b10 +
#763790000000
0!
0'
#763800000000
1!
b11 %
1'
b11 +
#763810000000
0!
0'
#763820000000
1!
b100 %
1'
b100 +
#763830000000
0!
0'
#763840000000
1!
b101 %
1'
b101 +
#763850000000
0!
0'
#763860000000
1!
0$
b110 %
1'
0*
b110 +
#763870000000
0!
0'
#763880000000
1!
b111 %
1'
b111 +
#763890000000
1"
1(
#763900000000
0!
0"
b100 &
0'
0(
b100 ,
#763910000000
1!
b1000 %
1'
b1000 +
#763920000000
0!
0'
#763930000000
1!
b1001 %
1'
b1001 +
#763940000000
0!
0'
#763950000000
1!
b0 %
1'
b0 +
#763960000000
0!
0'
#763970000000
1!
1$
b1 %
1'
1*
b1 +
#763980000000
0!
0'
#763990000000
1!
b10 %
1'
b10 +
#764000000000
0!
0'
#764010000000
1!
b11 %
1'
b11 +
#764020000000
0!
0'
#764030000000
1!
b100 %
1'
b100 +
#764040000000
0!
0'
#764050000000
1!
b101 %
1'
b101 +
#764060000000
0!
0'
#764070000000
1!
b110 %
1'
b110 +
#764080000000
0!
0'
#764090000000
1!
b111 %
1'
b111 +
#764100000000
0!
0'
#764110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#764120000000
0!
0'
#764130000000
1!
b1001 %
1'
b1001 +
#764140000000
0!
0'
#764150000000
1!
b0 %
1'
b0 +
#764160000000
0!
0'
#764170000000
1!
1$
b1 %
1'
1*
b1 +
#764180000000
0!
0'
#764190000000
1!
b10 %
1'
b10 +
#764200000000
0!
0'
#764210000000
1!
b11 %
1'
b11 +
#764220000000
0!
0'
#764230000000
1!
b100 %
1'
b100 +
#764240000000
0!
0'
#764250000000
1!
b101 %
1'
b101 +
#764260000000
0!
0'
#764270000000
1!
0$
b110 %
1'
0*
b110 +
#764280000000
0!
0'
#764290000000
1!
b111 %
1'
b111 +
#764300000000
0!
0'
#764310000000
1!
b1000 %
1'
b1000 +
#764320000000
1"
1(
#764330000000
0!
0"
b100 &
0'
0(
b100 ,
#764340000000
1!
b1001 %
1'
b1001 +
#764350000000
0!
0'
#764360000000
1!
b0 %
1'
b0 +
#764370000000
0!
0'
#764380000000
1!
1$
b1 %
1'
1*
b1 +
#764390000000
0!
0'
#764400000000
1!
b10 %
1'
b10 +
#764410000000
0!
0'
#764420000000
1!
b11 %
1'
b11 +
#764430000000
0!
0'
#764440000000
1!
b100 %
1'
b100 +
#764450000000
0!
0'
#764460000000
1!
b101 %
1'
b101 +
#764470000000
0!
0'
#764480000000
1!
b110 %
1'
b110 +
#764490000000
0!
0'
#764500000000
1!
b111 %
1'
b111 +
#764510000000
0!
0'
#764520000000
1!
0$
b1000 %
1'
0*
b1000 +
#764530000000
0!
0'
#764540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#764550000000
0!
0'
#764560000000
1!
b0 %
1'
b0 +
#764570000000
0!
0'
#764580000000
1!
1$
b1 %
1'
1*
b1 +
#764590000000
0!
0'
#764600000000
1!
b10 %
1'
b10 +
#764610000000
0!
0'
#764620000000
1!
b11 %
1'
b11 +
#764630000000
0!
0'
#764640000000
1!
b100 %
1'
b100 +
#764650000000
0!
0'
#764660000000
1!
b101 %
1'
b101 +
#764670000000
0!
0'
#764680000000
1!
0$
b110 %
1'
0*
b110 +
#764690000000
0!
0'
#764700000000
1!
b111 %
1'
b111 +
#764710000000
0!
0'
#764720000000
1!
b1000 %
1'
b1000 +
#764730000000
0!
0'
#764740000000
1!
b1001 %
1'
b1001 +
#764750000000
1"
1(
#764760000000
0!
0"
b100 &
0'
0(
b100 ,
#764770000000
1!
b0 %
1'
b0 +
#764780000000
0!
0'
#764790000000
1!
1$
b1 %
1'
1*
b1 +
#764800000000
0!
0'
#764810000000
1!
b10 %
1'
b10 +
#764820000000
0!
0'
#764830000000
1!
b11 %
1'
b11 +
#764840000000
0!
0'
#764850000000
1!
b100 %
1'
b100 +
#764860000000
0!
0'
#764870000000
1!
b101 %
1'
b101 +
#764880000000
0!
0'
#764890000000
1!
b110 %
1'
b110 +
#764900000000
0!
0'
#764910000000
1!
b111 %
1'
b111 +
#764920000000
0!
0'
#764930000000
1!
0$
b1000 %
1'
0*
b1000 +
#764940000000
0!
0'
#764950000000
1!
b1001 %
1'
b1001 +
#764960000000
0!
0'
#764970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#764980000000
0!
0'
#764990000000
1!
1$
b1 %
1'
1*
b1 +
#765000000000
0!
0'
#765010000000
1!
b10 %
1'
b10 +
#765020000000
0!
0'
#765030000000
1!
b11 %
1'
b11 +
#765040000000
0!
0'
#765050000000
1!
b100 %
1'
b100 +
#765060000000
0!
0'
#765070000000
1!
b101 %
1'
b101 +
#765080000000
0!
0'
#765090000000
1!
0$
b110 %
1'
0*
b110 +
#765100000000
0!
0'
#765110000000
1!
b111 %
1'
b111 +
#765120000000
0!
0'
#765130000000
1!
b1000 %
1'
b1000 +
#765140000000
0!
0'
#765150000000
1!
b1001 %
1'
b1001 +
#765160000000
0!
0'
#765170000000
1!
b0 %
1'
b0 +
#765180000000
1"
1(
#765190000000
0!
0"
b100 &
0'
0(
b100 ,
#765200000000
1!
1$
b1 %
1'
1*
b1 +
#765210000000
0!
0'
#765220000000
1!
b10 %
1'
b10 +
#765230000000
0!
0'
#765240000000
1!
b11 %
1'
b11 +
#765250000000
0!
0'
#765260000000
1!
b100 %
1'
b100 +
#765270000000
0!
0'
#765280000000
1!
b101 %
1'
b101 +
#765290000000
0!
0'
#765300000000
1!
b110 %
1'
b110 +
#765310000000
0!
0'
#765320000000
1!
b111 %
1'
b111 +
#765330000000
0!
0'
#765340000000
1!
0$
b1000 %
1'
0*
b1000 +
#765350000000
0!
0'
#765360000000
1!
b1001 %
1'
b1001 +
#765370000000
0!
0'
#765380000000
1!
b0 %
1'
b0 +
#765390000000
0!
0'
#765400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#765410000000
0!
0'
#765420000000
1!
b10 %
1'
b10 +
#765430000000
0!
0'
#765440000000
1!
b11 %
1'
b11 +
#765450000000
0!
0'
#765460000000
1!
b100 %
1'
b100 +
#765470000000
0!
0'
#765480000000
1!
b101 %
1'
b101 +
#765490000000
0!
0'
#765500000000
1!
0$
b110 %
1'
0*
b110 +
#765510000000
0!
0'
#765520000000
1!
b111 %
1'
b111 +
#765530000000
0!
0'
#765540000000
1!
b1000 %
1'
b1000 +
#765550000000
0!
0'
#765560000000
1!
b1001 %
1'
b1001 +
#765570000000
0!
0'
#765580000000
1!
b0 %
1'
b0 +
#765590000000
0!
0'
#765600000000
1!
1$
b1 %
1'
1*
b1 +
#765610000000
1"
1(
#765620000000
0!
0"
b100 &
0'
0(
b100 ,
#765630000000
1!
b10 %
1'
b10 +
#765640000000
0!
0'
#765650000000
1!
b11 %
1'
b11 +
#765660000000
0!
0'
#765670000000
1!
b100 %
1'
b100 +
#765680000000
0!
0'
#765690000000
1!
b101 %
1'
b101 +
#765700000000
0!
0'
#765710000000
1!
b110 %
1'
b110 +
#765720000000
0!
0'
#765730000000
1!
b111 %
1'
b111 +
#765740000000
0!
0'
#765750000000
1!
0$
b1000 %
1'
0*
b1000 +
#765760000000
0!
0'
#765770000000
1!
b1001 %
1'
b1001 +
#765780000000
0!
0'
#765790000000
1!
b0 %
1'
b0 +
#765800000000
0!
0'
#765810000000
1!
1$
b1 %
1'
1*
b1 +
#765820000000
0!
0'
#765830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#765840000000
0!
0'
#765850000000
1!
b11 %
1'
b11 +
#765860000000
0!
0'
#765870000000
1!
b100 %
1'
b100 +
#765880000000
0!
0'
#765890000000
1!
b101 %
1'
b101 +
#765900000000
0!
0'
#765910000000
1!
0$
b110 %
1'
0*
b110 +
#765920000000
0!
0'
#765930000000
1!
b111 %
1'
b111 +
#765940000000
0!
0'
#765950000000
1!
b1000 %
1'
b1000 +
#765960000000
0!
0'
#765970000000
1!
b1001 %
1'
b1001 +
#765980000000
0!
0'
#765990000000
1!
b0 %
1'
b0 +
#766000000000
0!
0'
#766010000000
1!
1$
b1 %
1'
1*
b1 +
#766020000000
0!
0'
#766030000000
1!
b10 %
1'
b10 +
#766040000000
1"
1(
#766050000000
0!
0"
b100 &
0'
0(
b100 ,
#766060000000
1!
b11 %
1'
b11 +
#766070000000
0!
0'
#766080000000
1!
b100 %
1'
b100 +
#766090000000
0!
0'
#766100000000
1!
b101 %
1'
b101 +
#766110000000
0!
0'
#766120000000
1!
b110 %
1'
b110 +
#766130000000
0!
0'
#766140000000
1!
b111 %
1'
b111 +
#766150000000
0!
0'
#766160000000
1!
0$
b1000 %
1'
0*
b1000 +
#766170000000
0!
0'
#766180000000
1!
b1001 %
1'
b1001 +
#766190000000
0!
0'
#766200000000
1!
b0 %
1'
b0 +
#766210000000
0!
0'
#766220000000
1!
1$
b1 %
1'
1*
b1 +
#766230000000
0!
0'
#766240000000
1!
b10 %
1'
b10 +
#766250000000
0!
0'
#766260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#766270000000
0!
0'
#766280000000
1!
b100 %
1'
b100 +
#766290000000
0!
0'
#766300000000
1!
b101 %
1'
b101 +
#766310000000
0!
0'
#766320000000
1!
0$
b110 %
1'
0*
b110 +
#766330000000
0!
0'
#766340000000
1!
b111 %
1'
b111 +
#766350000000
0!
0'
#766360000000
1!
b1000 %
1'
b1000 +
#766370000000
0!
0'
#766380000000
1!
b1001 %
1'
b1001 +
#766390000000
0!
0'
#766400000000
1!
b0 %
1'
b0 +
#766410000000
0!
0'
#766420000000
1!
1$
b1 %
1'
1*
b1 +
#766430000000
0!
0'
#766440000000
1!
b10 %
1'
b10 +
#766450000000
0!
0'
#766460000000
1!
b11 %
1'
b11 +
#766470000000
1"
1(
#766480000000
0!
0"
b100 &
0'
0(
b100 ,
#766490000000
1!
b100 %
1'
b100 +
#766500000000
0!
0'
#766510000000
1!
b101 %
1'
b101 +
#766520000000
0!
0'
#766530000000
1!
b110 %
1'
b110 +
#766540000000
0!
0'
#766550000000
1!
b111 %
1'
b111 +
#766560000000
0!
0'
#766570000000
1!
0$
b1000 %
1'
0*
b1000 +
#766580000000
0!
0'
#766590000000
1!
b1001 %
1'
b1001 +
#766600000000
0!
0'
#766610000000
1!
b0 %
1'
b0 +
#766620000000
0!
0'
#766630000000
1!
1$
b1 %
1'
1*
b1 +
#766640000000
0!
0'
#766650000000
1!
b10 %
1'
b10 +
#766660000000
0!
0'
#766670000000
1!
b11 %
1'
b11 +
#766680000000
0!
0'
#766690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#766700000000
0!
0'
#766710000000
1!
b101 %
1'
b101 +
#766720000000
0!
0'
#766730000000
1!
0$
b110 %
1'
0*
b110 +
#766740000000
0!
0'
#766750000000
1!
b111 %
1'
b111 +
#766760000000
0!
0'
#766770000000
1!
b1000 %
1'
b1000 +
#766780000000
0!
0'
#766790000000
1!
b1001 %
1'
b1001 +
#766800000000
0!
0'
#766810000000
1!
b0 %
1'
b0 +
#766820000000
0!
0'
#766830000000
1!
1$
b1 %
1'
1*
b1 +
#766840000000
0!
0'
#766850000000
1!
b10 %
1'
b10 +
#766860000000
0!
0'
#766870000000
1!
b11 %
1'
b11 +
#766880000000
0!
0'
#766890000000
1!
b100 %
1'
b100 +
#766900000000
1"
1(
#766910000000
0!
0"
b100 &
0'
0(
b100 ,
#766920000000
1!
b101 %
1'
b101 +
#766930000000
0!
0'
#766940000000
1!
b110 %
1'
b110 +
#766950000000
0!
0'
#766960000000
1!
b111 %
1'
b111 +
#766970000000
0!
0'
#766980000000
1!
0$
b1000 %
1'
0*
b1000 +
#766990000000
0!
0'
#767000000000
1!
b1001 %
1'
b1001 +
#767010000000
0!
0'
#767020000000
1!
b0 %
1'
b0 +
#767030000000
0!
0'
#767040000000
1!
1$
b1 %
1'
1*
b1 +
#767050000000
0!
0'
#767060000000
1!
b10 %
1'
b10 +
#767070000000
0!
0'
#767080000000
1!
b11 %
1'
b11 +
#767090000000
0!
0'
#767100000000
1!
b100 %
1'
b100 +
#767110000000
0!
0'
#767120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#767130000000
0!
0'
#767140000000
1!
0$
b110 %
1'
0*
b110 +
#767150000000
0!
0'
#767160000000
1!
b111 %
1'
b111 +
#767170000000
0!
0'
#767180000000
1!
b1000 %
1'
b1000 +
#767190000000
0!
0'
#767200000000
1!
b1001 %
1'
b1001 +
#767210000000
0!
0'
#767220000000
1!
b0 %
1'
b0 +
#767230000000
0!
0'
#767240000000
1!
1$
b1 %
1'
1*
b1 +
#767250000000
0!
0'
#767260000000
1!
b10 %
1'
b10 +
#767270000000
0!
0'
#767280000000
1!
b11 %
1'
b11 +
#767290000000
0!
0'
#767300000000
1!
b100 %
1'
b100 +
#767310000000
0!
0'
#767320000000
1!
b101 %
1'
b101 +
#767330000000
1"
1(
#767340000000
0!
0"
b100 &
0'
0(
b100 ,
#767350000000
1!
b110 %
1'
b110 +
#767360000000
0!
0'
#767370000000
1!
b111 %
1'
b111 +
#767380000000
0!
0'
#767390000000
1!
0$
b1000 %
1'
0*
b1000 +
#767400000000
0!
0'
#767410000000
1!
b1001 %
1'
b1001 +
#767420000000
0!
0'
#767430000000
1!
b0 %
1'
b0 +
#767440000000
0!
0'
#767450000000
1!
1$
b1 %
1'
1*
b1 +
#767460000000
0!
0'
#767470000000
1!
b10 %
1'
b10 +
#767480000000
0!
0'
#767490000000
1!
b11 %
1'
b11 +
#767500000000
0!
0'
#767510000000
1!
b100 %
1'
b100 +
#767520000000
0!
0'
#767530000000
1!
b101 %
1'
b101 +
#767540000000
0!
0'
#767550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#767560000000
0!
0'
#767570000000
1!
b111 %
1'
b111 +
#767580000000
0!
0'
#767590000000
1!
b1000 %
1'
b1000 +
#767600000000
0!
0'
#767610000000
1!
b1001 %
1'
b1001 +
#767620000000
0!
0'
#767630000000
1!
b0 %
1'
b0 +
#767640000000
0!
0'
#767650000000
1!
1$
b1 %
1'
1*
b1 +
#767660000000
0!
0'
#767670000000
1!
b10 %
1'
b10 +
#767680000000
0!
0'
#767690000000
1!
b11 %
1'
b11 +
#767700000000
0!
0'
#767710000000
1!
b100 %
1'
b100 +
#767720000000
0!
0'
#767730000000
1!
b101 %
1'
b101 +
#767740000000
0!
0'
#767750000000
1!
0$
b110 %
1'
0*
b110 +
#767760000000
1"
1(
#767770000000
0!
0"
b100 &
0'
0(
b100 ,
#767780000000
1!
1$
b111 %
1'
1*
b111 +
#767790000000
0!
0'
#767800000000
1!
0$
b1000 %
1'
0*
b1000 +
#767810000000
0!
0'
#767820000000
1!
b1001 %
1'
b1001 +
#767830000000
0!
0'
#767840000000
1!
b0 %
1'
b0 +
#767850000000
0!
0'
#767860000000
1!
1$
b1 %
1'
1*
b1 +
#767870000000
0!
0'
#767880000000
1!
b10 %
1'
b10 +
#767890000000
0!
0'
#767900000000
1!
b11 %
1'
b11 +
#767910000000
0!
0'
#767920000000
1!
b100 %
1'
b100 +
#767930000000
0!
0'
#767940000000
1!
b101 %
1'
b101 +
#767950000000
0!
0'
#767960000000
1!
b110 %
1'
b110 +
#767970000000
0!
0'
#767980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#767990000000
0!
0'
#768000000000
1!
b1000 %
1'
b1000 +
#768010000000
0!
0'
#768020000000
1!
b1001 %
1'
b1001 +
#768030000000
0!
0'
#768040000000
1!
b0 %
1'
b0 +
#768050000000
0!
0'
#768060000000
1!
1$
b1 %
1'
1*
b1 +
#768070000000
0!
0'
#768080000000
1!
b10 %
1'
b10 +
#768090000000
0!
0'
#768100000000
1!
b11 %
1'
b11 +
#768110000000
0!
0'
#768120000000
1!
b100 %
1'
b100 +
#768130000000
0!
0'
#768140000000
1!
b101 %
1'
b101 +
#768150000000
0!
0'
#768160000000
1!
0$
b110 %
1'
0*
b110 +
#768170000000
0!
0'
#768180000000
1!
b111 %
1'
b111 +
#768190000000
1"
1(
#768200000000
0!
0"
b100 &
0'
0(
b100 ,
#768210000000
1!
b1000 %
1'
b1000 +
#768220000000
0!
0'
#768230000000
1!
b1001 %
1'
b1001 +
#768240000000
0!
0'
#768250000000
1!
b0 %
1'
b0 +
#768260000000
0!
0'
#768270000000
1!
1$
b1 %
1'
1*
b1 +
#768280000000
0!
0'
#768290000000
1!
b10 %
1'
b10 +
#768300000000
0!
0'
#768310000000
1!
b11 %
1'
b11 +
#768320000000
0!
0'
#768330000000
1!
b100 %
1'
b100 +
#768340000000
0!
0'
#768350000000
1!
b101 %
1'
b101 +
#768360000000
0!
0'
#768370000000
1!
b110 %
1'
b110 +
#768380000000
0!
0'
#768390000000
1!
b111 %
1'
b111 +
#768400000000
0!
0'
#768410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#768420000000
0!
0'
#768430000000
1!
b1001 %
1'
b1001 +
#768440000000
0!
0'
#768450000000
1!
b0 %
1'
b0 +
#768460000000
0!
0'
#768470000000
1!
1$
b1 %
1'
1*
b1 +
#768480000000
0!
0'
#768490000000
1!
b10 %
1'
b10 +
#768500000000
0!
0'
#768510000000
1!
b11 %
1'
b11 +
#768520000000
0!
0'
#768530000000
1!
b100 %
1'
b100 +
#768540000000
0!
0'
#768550000000
1!
b101 %
1'
b101 +
#768560000000
0!
0'
#768570000000
1!
0$
b110 %
1'
0*
b110 +
#768580000000
0!
0'
#768590000000
1!
b111 %
1'
b111 +
#768600000000
0!
0'
#768610000000
1!
b1000 %
1'
b1000 +
#768620000000
1"
1(
#768630000000
0!
0"
b100 &
0'
0(
b100 ,
#768640000000
1!
b1001 %
1'
b1001 +
#768650000000
0!
0'
#768660000000
1!
b0 %
1'
b0 +
#768670000000
0!
0'
#768680000000
1!
1$
b1 %
1'
1*
b1 +
#768690000000
0!
0'
#768700000000
1!
b10 %
1'
b10 +
#768710000000
0!
0'
#768720000000
1!
b11 %
1'
b11 +
#768730000000
0!
0'
#768740000000
1!
b100 %
1'
b100 +
#768750000000
0!
0'
#768760000000
1!
b101 %
1'
b101 +
#768770000000
0!
0'
#768780000000
1!
b110 %
1'
b110 +
#768790000000
0!
0'
#768800000000
1!
b111 %
1'
b111 +
#768810000000
0!
0'
#768820000000
1!
0$
b1000 %
1'
0*
b1000 +
#768830000000
0!
0'
#768840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#768850000000
0!
0'
#768860000000
1!
b0 %
1'
b0 +
#768870000000
0!
0'
#768880000000
1!
1$
b1 %
1'
1*
b1 +
#768890000000
0!
0'
#768900000000
1!
b10 %
1'
b10 +
#768910000000
0!
0'
#768920000000
1!
b11 %
1'
b11 +
#768930000000
0!
0'
#768940000000
1!
b100 %
1'
b100 +
#768950000000
0!
0'
#768960000000
1!
b101 %
1'
b101 +
#768970000000
0!
0'
#768980000000
1!
0$
b110 %
1'
0*
b110 +
#768990000000
0!
0'
#769000000000
1!
b111 %
1'
b111 +
#769010000000
0!
0'
#769020000000
1!
b1000 %
1'
b1000 +
#769030000000
0!
0'
#769040000000
1!
b1001 %
1'
b1001 +
#769050000000
1"
1(
#769060000000
0!
0"
b100 &
0'
0(
b100 ,
#769070000000
1!
b0 %
1'
b0 +
#769080000000
0!
0'
#769090000000
1!
1$
b1 %
1'
1*
b1 +
#769100000000
0!
0'
#769110000000
1!
b10 %
1'
b10 +
#769120000000
0!
0'
#769130000000
1!
b11 %
1'
b11 +
#769140000000
0!
0'
#769150000000
1!
b100 %
1'
b100 +
#769160000000
0!
0'
#769170000000
1!
b101 %
1'
b101 +
#769180000000
0!
0'
#769190000000
1!
b110 %
1'
b110 +
#769200000000
0!
0'
#769210000000
1!
b111 %
1'
b111 +
#769220000000
0!
0'
#769230000000
1!
0$
b1000 %
1'
0*
b1000 +
#769240000000
0!
0'
#769250000000
1!
b1001 %
1'
b1001 +
#769260000000
0!
0'
#769270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#769280000000
0!
0'
#769290000000
1!
1$
b1 %
1'
1*
b1 +
#769300000000
0!
0'
#769310000000
1!
b10 %
1'
b10 +
#769320000000
0!
0'
#769330000000
1!
b11 %
1'
b11 +
#769340000000
0!
0'
#769350000000
1!
b100 %
1'
b100 +
#769360000000
0!
0'
#769370000000
1!
b101 %
1'
b101 +
#769380000000
0!
0'
#769390000000
1!
0$
b110 %
1'
0*
b110 +
#769400000000
0!
0'
#769410000000
1!
b111 %
1'
b111 +
#769420000000
0!
0'
#769430000000
1!
b1000 %
1'
b1000 +
#769440000000
0!
0'
#769450000000
1!
b1001 %
1'
b1001 +
#769460000000
0!
0'
#769470000000
1!
b0 %
1'
b0 +
#769480000000
1"
1(
#769490000000
0!
0"
b100 &
0'
0(
b100 ,
#769500000000
1!
1$
b1 %
1'
1*
b1 +
#769510000000
0!
0'
#769520000000
1!
b10 %
1'
b10 +
#769530000000
0!
0'
#769540000000
1!
b11 %
1'
b11 +
#769550000000
0!
0'
#769560000000
1!
b100 %
1'
b100 +
#769570000000
0!
0'
#769580000000
1!
b101 %
1'
b101 +
#769590000000
0!
0'
#769600000000
1!
b110 %
1'
b110 +
#769610000000
0!
0'
#769620000000
1!
b111 %
1'
b111 +
#769630000000
0!
0'
#769640000000
1!
0$
b1000 %
1'
0*
b1000 +
#769650000000
0!
0'
#769660000000
1!
b1001 %
1'
b1001 +
#769670000000
0!
0'
#769680000000
1!
b0 %
1'
b0 +
#769690000000
0!
0'
#769700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#769710000000
0!
0'
#769720000000
1!
b10 %
1'
b10 +
#769730000000
0!
0'
#769740000000
1!
b11 %
1'
b11 +
#769750000000
0!
0'
#769760000000
1!
b100 %
1'
b100 +
#769770000000
0!
0'
#769780000000
1!
b101 %
1'
b101 +
#769790000000
0!
0'
#769800000000
1!
0$
b110 %
1'
0*
b110 +
#769810000000
0!
0'
#769820000000
1!
b111 %
1'
b111 +
#769830000000
0!
0'
#769840000000
1!
b1000 %
1'
b1000 +
#769850000000
0!
0'
#769860000000
1!
b1001 %
1'
b1001 +
#769870000000
0!
0'
#769880000000
1!
b0 %
1'
b0 +
#769890000000
0!
0'
#769900000000
1!
1$
b1 %
1'
1*
b1 +
#769910000000
1"
1(
#769920000000
0!
0"
b100 &
0'
0(
b100 ,
#769930000000
1!
b10 %
1'
b10 +
#769940000000
0!
0'
#769950000000
1!
b11 %
1'
b11 +
#769960000000
0!
0'
#769970000000
1!
b100 %
1'
b100 +
#769980000000
0!
0'
#769990000000
1!
b101 %
1'
b101 +
#770000000000
0!
0'
#770010000000
1!
b110 %
1'
b110 +
#770020000000
0!
0'
#770030000000
1!
b111 %
1'
b111 +
#770040000000
0!
0'
#770050000000
1!
0$
b1000 %
1'
0*
b1000 +
#770060000000
0!
0'
#770070000000
1!
b1001 %
1'
b1001 +
#770080000000
0!
0'
#770090000000
1!
b0 %
1'
b0 +
#770100000000
0!
0'
#770110000000
1!
1$
b1 %
1'
1*
b1 +
#770120000000
0!
0'
#770130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#770140000000
0!
0'
#770150000000
1!
b11 %
1'
b11 +
#770160000000
0!
0'
#770170000000
1!
b100 %
1'
b100 +
#770180000000
0!
0'
#770190000000
1!
b101 %
1'
b101 +
#770200000000
0!
0'
#770210000000
1!
0$
b110 %
1'
0*
b110 +
#770220000000
0!
0'
#770230000000
1!
b111 %
1'
b111 +
#770240000000
0!
0'
#770250000000
1!
b1000 %
1'
b1000 +
#770260000000
0!
0'
#770270000000
1!
b1001 %
1'
b1001 +
#770280000000
0!
0'
#770290000000
1!
b0 %
1'
b0 +
#770300000000
0!
0'
#770310000000
1!
1$
b1 %
1'
1*
b1 +
#770320000000
0!
0'
#770330000000
1!
b10 %
1'
b10 +
#770340000000
1"
1(
#770350000000
0!
0"
b100 &
0'
0(
b100 ,
#770360000000
1!
b11 %
1'
b11 +
#770370000000
0!
0'
#770380000000
1!
b100 %
1'
b100 +
#770390000000
0!
0'
#770400000000
1!
b101 %
1'
b101 +
#770410000000
0!
0'
#770420000000
1!
b110 %
1'
b110 +
#770430000000
0!
0'
#770440000000
1!
b111 %
1'
b111 +
#770450000000
0!
0'
#770460000000
1!
0$
b1000 %
1'
0*
b1000 +
#770470000000
0!
0'
#770480000000
1!
b1001 %
1'
b1001 +
#770490000000
0!
0'
#770500000000
1!
b0 %
1'
b0 +
#770510000000
0!
0'
#770520000000
1!
1$
b1 %
1'
1*
b1 +
#770530000000
0!
0'
#770540000000
1!
b10 %
1'
b10 +
#770550000000
0!
0'
#770560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#770570000000
0!
0'
#770580000000
1!
b100 %
1'
b100 +
#770590000000
0!
0'
#770600000000
1!
b101 %
1'
b101 +
#770610000000
0!
0'
#770620000000
1!
0$
b110 %
1'
0*
b110 +
#770630000000
0!
0'
#770640000000
1!
b111 %
1'
b111 +
#770650000000
0!
0'
#770660000000
1!
b1000 %
1'
b1000 +
#770670000000
0!
0'
#770680000000
1!
b1001 %
1'
b1001 +
#770690000000
0!
0'
#770700000000
1!
b0 %
1'
b0 +
#770710000000
0!
0'
#770720000000
1!
1$
b1 %
1'
1*
b1 +
#770730000000
0!
0'
#770740000000
1!
b10 %
1'
b10 +
#770750000000
0!
0'
#770760000000
1!
b11 %
1'
b11 +
#770770000000
1"
1(
#770780000000
0!
0"
b100 &
0'
0(
b100 ,
#770790000000
1!
b100 %
1'
b100 +
#770800000000
0!
0'
#770810000000
1!
b101 %
1'
b101 +
#770820000000
0!
0'
#770830000000
1!
b110 %
1'
b110 +
#770840000000
0!
0'
#770850000000
1!
b111 %
1'
b111 +
#770860000000
0!
0'
#770870000000
1!
0$
b1000 %
1'
0*
b1000 +
#770880000000
0!
0'
#770890000000
1!
b1001 %
1'
b1001 +
#770900000000
0!
0'
#770910000000
1!
b0 %
1'
b0 +
#770920000000
0!
0'
#770930000000
1!
1$
b1 %
1'
1*
b1 +
#770940000000
0!
0'
#770950000000
1!
b10 %
1'
b10 +
#770960000000
0!
0'
#770970000000
1!
b11 %
1'
b11 +
#770980000000
0!
0'
#770990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#771000000000
0!
0'
#771010000000
1!
b101 %
1'
b101 +
#771020000000
0!
0'
#771030000000
1!
0$
b110 %
1'
0*
b110 +
#771040000000
0!
0'
#771050000000
1!
b111 %
1'
b111 +
#771060000000
0!
0'
#771070000000
1!
b1000 %
1'
b1000 +
#771080000000
0!
0'
#771090000000
1!
b1001 %
1'
b1001 +
#771100000000
0!
0'
#771110000000
1!
b0 %
1'
b0 +
#771120000000
0!
0'
#771130000000
1!
1$
b1 %
1'
1*
b1 +
#771140000000
0!
0'
#771150000000
1!
b10 %
1'
b10 +
#771160000000
0!
0'
#771170000000
1!
b11 %
1'
b11 +
#771180000000
0!
0'
#771190000000
1!
b100 %
1'
b100 +
#771200000000
1"
1(
#771210000000
0!
0"
b100 &
0'
0(
b100 ,
#771220000000
1!
b101 %
1'
b101 +
#771230000000
0!
0'
#771240000000
1!
b110 %
1'
b110 +
#771250000000
0!
0'
#771260000000
1!
b111 %
1'
b111 +
#771270000000
0!
0'
#771280000000
1!
0$
b1000 %
1'
0*
b1000 +
#771290000000
0!
0'
#771300000000
1!
b1001 %
1'
b1001 +
#771310000000
0!
0'
#771320000000
1!
b0 %
1'
b0 +
#771330000000
0!
0'
#771340000000
1!
1$
b1 %
1'
1*
b1 +
#771350000000
0!
0'
#771360000000
1!
b10 %
1'
b10 +
#771370000000
0!
0'
#771380000000
1!
b11 %
1'
b11 +
#771390000000
0!
0'
#771400000000
1!
b100 %
1'
b100 +
#771410000000
0!
0'
#771420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#771430000000
0!
0'
#771440000000
1!
0$
b110 %
1'
0*
b110 +
#771450000000
0!
0'
#771460000000
1!
b111 %
1'
b111 +
#771470000000
0!
0'
#771480000000
1!
b1000 %
1'
b1000 +
#771490000000
0!
0'
#771500000000
1!
b1001 %
1'
b1001 +
#771510000000
0!
0'
#771520000000
1!
b0 %
1'
b0 +
#771530000000
0!
0'
#771540000000
1!
1$
b1 %
1'
1*
b1 +
#771550000000
0!
0'
#771560000000
1!
b10 %
1'
b10 +
#771570000000
0!
0'
#771580000000
1!
b11 %
1'
b11 +
#771590000000
0!
0'
#771600000000
1!
b100 %
1'
b100 +
#771610000000
0!
0'
#771620000000
1!
b101 %
1'
b101 +
#771630000000
1"
1(
#771640000000
0!
0"
b100 &
0'
0(
b100 ,
#771650000000
1!
b110 %
1'
b110 +
#771660000000
0!
0'
#771670000000
1!
b111 %
1'
b111 +
#771680000000
0!
0'
#771690000000
1!
0$
b1000 %
1'
0*
b1000 +
#771700000000
0!
0'
#771710000000
1!
b1001 %
1'
b1001 +
#771720000000
0!
0'
#771730000000
1!
b0 %
1'
b0 +
#771740000000
0!
0'
#771750000000
1!
1$
b1 %
1'
1*
b1 +
#771760000000
0!
0'
#771770000000
1!
b10 %
1'
b10 +
#771780000000
0!
0'
#771790000000
1!
b11 %
1'
b11 +
#771800000000
0!
0'
#771810000000
1!
b100 %
1'
b100 +
#771820000000
0!
0'
#771830000000
1!
b101 %
1'
b101 +
#771840000000
0!
0'
#771850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#771860000000
0!
0'
#771870000000
1!
b111 %
1'
b111 +
#771880000000
0!
0'
#771890000000
1!
b1000 %
1'
b1000 +
#771900000000
0!
0'
#771910000000
1!
b1001 %
1'
b1001 +
#771920000000
0!
0'
#771930000000
1!
b0 %
1'
b0 +
#771940000000
0!
0'
#771950000000
1!
1$
b1 %
1'
1*
b1 +
#771960000000
0!
0'
#771970000000
1!
b10 %
1'
b10 +
#771980000000
0!
0'
#771990000000
1!
b11 %
1'
b11 +
#772000000000
0!
0'
#772010000000
1!
b100 %
1'
b100 +
#772020000000
0!
0'
#772030000000
1!
b101 %
1'
b101 +
#772040000000
0!
0'
#772050000000
1!
0$
b110 %
1'
0*
b110 +
#772060000000
1"
1(
#772070000000
0!
0"
b100 &
0'
0(
b100 ,
#772080000000
1!
1$
b111 %
1'
1*
b111 +
#772090000000
0!
0'
#772100000000
1!
0$
b1000 %
1'
0*
b1000 +
#772110000000
0!
0'
#772120000000
1!
b1001 %
1'
b1001 +
#772130000000
0!
0'
#772140000000
1!
b0 %
1'
b0 +
#772150000000
0!
0'
#772160000000
1!
1$
b1 %
1'
1*
b1 +
#772170000000
0!
0'
#772180000000
1!
b10 %
1'
b10 +
#772190000000
0!
0'
#772200000000
1!
b11 %
1'
b11 +
#772210000000
0!
0'
#772220000000
1!
b100 %
1'
b100 +
#772230000000
0!
0'
#772240000000
1!
b101 %
1'
b101 +
#772250000000
0!
0'
#772260000000
1!
b110 %
1'
b110 +
#772270000000
0!
0'
#772280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#772290000000
0!
0'
#772300000000
1!
b1000 %
1'
b1000 +
#772310000000
0!
0'
#772320000000
1!
b1001 %
1'
b1001 +
#772330000000
0!
0'
#772340000000
1!
b0 %
1'
b0 +
#772350000000
0!
0'
#772360000000
1!
1$
b1 %
1'
1*
b1 +
#772370000000
0!
0'
#772380000000
1!
b10 %
1'
b10 +
#772390000000
0!
0'
#772400000000
1!
b11 %
1'
b11 +
#772410000000
0!
0'
#772420000000
1!
b100 %
1'
b100 +
#772430000000
0!
0'
#772440000000
1!
b101 %
1'
b101 +
#772450000000
0!
0'
#772460000000
1!
0$
b110 %
1'
0*
b110 +
#772470000000
0!
0'
#772480000000
1!
b111 %
1'
b111 +
#772490000000
1"
1(
#772500000000
0!
0"
b100 &
0'
0(
b100 ,
#772510000000
1!
b1000 %
1'
b1000 +
#772520000000
0!
0'
#772530000000
1!
b1001 %
1'
b1001 +
#772540000000
0!
0'
#772550000000
1!
b0 %
1'
b0 +
#772560000000
0!
0'
#772570000000
1!
1$
b1 %
1'
1*
b1 +
#772580000000
0!
0'
#772590000000
1!
b10 %
1'
b10 +
#772600000000
0!
0'
#772610000000
1!
b11 %
1'
b11 +
#772620000000
0!
0'
#772630000000
1!
b100 %
1'
b100 +
#772640000000
0!
0'
#772650000000
1!
b101 %
1'
b101 +
#772660000000
0!
0'
#772670000000
1!
b110 %
1'
b110 +
#772680000000
0!
0'
#772690000000
1!
b111 %
1'
b111 +
#772700000000
0!
0'
#772710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#772720000000
0!
0'
#772730000000
1!
b1001 %
1'
b1001 +
#772740000000
0!
0'
#772750000000
1!
b0 %
1'
b0 +
#772760000000
0!
0'
#772770000000
1!
1$
b1 %
1'
1*
b1 +
#772780000000
0!
0'
#772790000000
1!
b10 %
1'
b10 +
#772800000000
0!
0'
#772810000000
1!
b11 %
1'
b11 +
#772820000000
0!
0'
#772830000000
1!
b100 %
1'
b100 +
#772840000000
0!
0'
#772850000000
1!
b101 %
1'
b101 +
#772860000000
0!
0'
#772870000000
1!
0$
b110 %
1'
0*
b110 +
#772880000000
0!
0'
#772890000000
1!
b111 %
1'
b111 +
#772900000000
0!
0'
#772910000000
1!
b1000 %
1'
b1000 +
#772920000000
1"
1(
#772930000000
0!
0"
b100 &
0'
0(
b100 ,
#772940000000
1!
b1001 %
1'
b1001 +
#772950000000
0!
0'
#772960000000
1!
b0 %
1'
b0 +
#772970000000
0!
0'
#772980000000
1!
1$
b1 %
1'
1*
b1 +
#772990000000
0!
0'
#773000000000
1!
b10 %
1'
b10 +
#773010000000
0!
0'
#773020000000
1!
b11 %
1'
b11 +
#773030000000
0!
0'
#773040000000
1!
b100 %
1'
b100 +
#773050000000
0!
0'
#773060000000
1!
b101 %
1'
b101 +
#773070000000
0!
0'
#773080000000
1!
b110 %
1'
b110 +
#773090000000
0!
0'
#773100000000
1!
b111 %
1'
b111 +
#773110000000
0!
0'
#773120000000
1!
0$
b1000 %
1'
0*
b1000 +
#773130000000
0!
0'
#773140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#773150000000
0!
0'
#773160000000
1!
b0 %
1'
b0 +
#773170000000
0!
0'
#773180000000
1!
1$
b1 %
1'
1*
b1 +
#773190000000
0!
0'
#773200000000
1!
b10 %
1'
b10 +
#773210000000
0!
0'
#773220000000
1!
b11 %
1'
b11 +
#773230000000
0!
0'
#773240000000
1!
b100 %
1'
b100 +
#773250000000
0!
0'
#773260000000
1!
b101 %
1'
b101 +
#773270000000
0!
0'
#773280000000
1!
0$
b110 %
1'
0*
b110 +
#773290000000
0!
0'
#773300000000
1!
b111 %
1'
b111 +
#773310000000
0!
0'
#773320000000
1!
b1000 %
1'
b1000 +
#773330000000
0!
0'
#773340000000
1!
b1001 %
1'
b1001 +
#773350000000
1"
1(
#773360000000
0!
0"
b100 &
0'
0(
b100 ,
#773370000000
1!
b0 %
1'
b0 +
#773380000000
0!
0'
#773390000000
1!
1$
b1 %
1'
1*
b1 +
#773400000000
0!
0'
#773410000000
1!
b10 %
1'
b10 +
#773420000000
0!
0'
#773430000000
1!
b11 %
1'
b11 +
#773440000000
0!
0'
#773450000000
1!
b100 %
1'
b100 +
#773460000000
0!
0'
#773470000000
1!
b101 %
1'
b101 +
#773480000000
0!
0'
#773490000000
1!
b110 %
1'
b110 +
#773500000000
0!
0'
#773510000000
1!
b111 %
1'
b111 +
#773520000000
0!
0'
#773530000000
1!
0$
b1000 %
1'
0*
b1000 +
#773540000000
0!
0'
#773550000000
1!
b1001 %
1'
b1001 +
#773560000000
0!
0'
#773570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#773580000000
0!
0'
#773590000000
1!
1$
b1 %
1'
1*
b1 +
#773600000000
0!
0'
#773610000000
1!
b10 %
1'
b10 +
#773620000000
0!
0'
#773630000000
1!
b11 %
1'
b11 +
#773640000000
0!
0'
#773650000000
1!
b100 %
1'
b100 +
#773660000000
0!
0'
#773670000000
1!
b101 %
1'
b101 +
#773680000000
0!
0'
#773690000000
1!
0$
b110 %
1'
0*
b110 +
#773700000000
0!
0'
#773710000000
1!
b111 %
1'
b111 +
#773720000000
0!
0'
#773730000000
1!
b1000 %
1'
b1000 +
#773740000000
0!
0'
#773750000000
1!
b1001 %
1'
b1001 +
#773760000000
0!
0'
#773770000000
1!
b0 %
1'
b0 +
#773780000000
1"
1(
#773790000000
0!
0"
b100 &
0'
0(
b100 ,
#773800000000
1!
1$
b1 %
1'
1*
b1 +
#773810000000
0!
0'
#773820000000
1!
b10 %
1'
b10 +
#773830000000
0!
0'
#773840000000
1!
b11 %
1'
b11 +
#773850000000
0!
0'
#773860000000
1!
b100 %
1'
b100 +
#773870000000
0!
0'
#773880000000
1!
b101 %
1'
b101 +
#773890000000
0!
0'
#773900000000
1!
b110 %
1'
b110 +
#773910000000
0!
0'
#773920000000
1!
b111 %
1'
b111 +
#773930000000
0!
0'
#773940000000
1!
0$
b1000 %
1'
0*
b1000 +
#773950000000
0!
0'
#773960000000
1!
b1001 %
1'
b1001 +
#773970000000
0!
0'
#773980000000
1!
b0 %
1'
b0 +
#773990000000
0!
0'
#774000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#774010000000
0!
0'
#774020000000
1!
b10 %
1'
b10 +
#774030000000
0!
0'
#774040000000
1!
b11 %
1'
b11 +
#774050000000
0!
0'
#774060000000
1!
b100 %
1'
b100 +
#774070000000
0!
0'
#774080000000
1!
b101 %
1'
b101 +
#774090000000
0!
0'
#774100000000
1!
0$
b110 %
1'
0*
b110 +
#774110000000
0!
0'
#774120000000
1!
b111 %
1'
b111 +
#774130000000
0!
0'
#774140000000
1!
b1000 %
1'
b1000 +
#774150000000
0!
0'
#774160000000
1!
b1001 %
1'
b1001 +
#774170000000
0!
0'
#774180000000
1!
b0 %
1'
b0 +
#774190000000
0!
0'
#774200000000
1!
1$
b1 %
1'
1*
b1 +
#774210000000
1"
1(
#774220000000
0!
0"
b100 &
0'
0(
b100 ,
#774230000000
1!
b10 %
1'
b10 +
#774240000000
0!
0'
#774250000000
1!
b11 %
1'
b11 +
#774260000000
0!
0'
#774270000000
1!
b100 %
1'
b100 +
#774280000000
0!
0'
#774290000000
1!
b101 %
1'
b101 +
#774300000000
0!
0'
#774310000000
1!
b110 %
1'
b110 +
#774320000000
0!
0'
#774330000000
1!
b111 %
1'
b111 +
#774340000000
0!
0'
#774350000000
1!
0$
b1000 %
1'
0*
b1000 +
#774360000000
0!
0'
#774370000000
1!
b1001 %
1'
b1001 +
#774380000000
0!
0'
#774390000000
1!
b0 %
1'
b0 +
#774400000000
0!
0'
#774410000000
1!
1$
b1 %
1'
1*
b1 +
#774420000000
0!
0'
#774430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#774440000000
0!
0'
#774450000000
1!
b11 %
1'
b11 +
#774460000000
0!
0'
#774470000000
1!
b100 %
1'
b100 +
#774480000000
0!
0'
#774490000000
1!
b101 %
1'
b101 +
#774500000000
0!
0'
#774510000000
1!
0$
b110 %
1'
0*
b110 +
#774520000000
0!
0'
#774530000000
1!
b111 %
1'
b111 +
#774540000000
0!
0'
#774550000000
1!
b1000 %
1'
b1000 +
#774560000000
0!
0'
#774570000000
1!
b1001 %
1'
b1001 +
#774580000000
0!
0'
#774590000000
1!
b0 %
1'
b0 +
#774600000000
0!
0'
#774610000000
1!
1$
b1 %
1'
1*
b1 +
#774620000000
0!
0'
#774630000000
1!
b10 %
1'
b10 +
#774640000000
1"
1(
#774650000000
0!
0"
b100 &
0'
0(
b100 ,
#774660000000
1!
b11 %
1'
b11 +
#774670000000
0!
0'
#774680000000
1!
b100 %
1'
b100 +
#774690000000
0!
0'
#774700000000
1!
b101 %
1'
b101 +
#774710000000
0!
0'
#774720000000
1!
b110 %
1'
b110 +
#774730000000
0!
0'
#774740000000
1!
b111 %
1'
b111 +
#774750000000
0!
0'
#774760000000
1!
0$
b1000 %
1'
0*
b1000 +
#774770000000
0!
0'
#774780000000
1!
b1001 %
1'
b1001 +
#774790000000
0!
0'
#774800000000
1!
b0 %
1'
b0 +
#774810000000
0!
0'
#774820000000
1!
1$
b1 %
1'
1*
b1 +
#774830000000
0!
0'
#774840000000
1!
b10 %
1'
b10 +
#774850000000
0!
0'
#774860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#774870000000
0!
0'
#774880000000
1!
b100 %
1'
b100 +
#774890000000
0!
0'
#774900000000
1!
b101 %
1'
b101 +
#774910000000
0!
0'
#774920000000
1!
0$
b110 %
1'
0*
b110 +
#774930000000
0!
0'
#774940000000
1!
b111 %
1'
b111 +
#774950000000
0!
0'
#774960000000
1!
b1000 %
1'
b1000 +
#774970000000
0!
0'
#774980000000
1!
b1001 %
1'
b1001 +
#774990000000
0!
0'
#775000000000
1!
b0 %
1'
b0 +
#775010000000
0!
0'
#775020000000
1!
1$
b1 %
1'
1*
b1 +
#775030000000
0!
0'
#775040000000
1!
b10 %
1'
b10 +
#775050000000
0!
0'
#775060000000
1!
b11 %
1'
b11 +
#775070000000
1"
1(
#775080000000
0!
0"
b100 &
0'
0(
b100 ,
#775090000000
1!
b100 %
1'
b100 +
#775100000000
0!
0'
#775110000000
1!
b101 %
1'
b101 +
#775120000000
0!
0'
#775130000000
1!
b110 %
1'
b110 +
#775140000000
0!
0'
#775150000000
1!
b111 %
1'
b111 +
#775160000000
0!
0'
#775170000000
1!
0$
b1000 %
1'
0*
b1000 +
#775180000000
0!
0'
#775190000000
1!
b1001 %
1'
b1001 +
#775200000000
0!
0'
#775210000000
1!
b0 %
1'
b0 +
#775220000000
0!
0'
#775230000000
1!
1$
b1 %
1'
1*
b1 +
#775240000000
0!
0'
#775250000000
1!
b10 %
1'
b10 +
#775260000000
0!
0'
#775270000000
1!
b11 %
1'
b11 +
#775280000000
0!
0'
#775290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#775300000000
0!
0'
#775310000000
1!
b101 %
1'
b101 +
#775320000000
0!
0'
#775330000000
1!
0$
b110 %
1'
0*
b110 +
#775340000000
0!
0'
#775350000000
1!
b111 %
1'
b111 +
#775360000000
0!
0'
#775370000000
1!
b1000 %
1'
b1000 +
#775380000000
0!
0'
#775390000000
1!
b1001 %
1'
b1001 +
#775400000000
0!
0'
#775410000000
1!
b0 %
1'
b0 +
#775420000000
0!
0'
#775430000000
1!
1$
b1 %
1'
1*
b1 +
#775440000000
0!
0'
#775450000000
1!
b10 %
1'
b10 +
#775460000000
0!
0'
#775470000000
1!
b11 %
1'
b11 +
#775480000000
0!
0'
#775490000000
1!
b100 %
1'
b100 +
#775500000000
1"
1(
#775510000000
0!
0"
b100 &
0'
0(
b100 ,
#775520000000
1!
b101 %
1'
b101 +
#775530000000
0!
0'
#775540000000
1!
b110 %
1'
b110 +
#775550000000
0!
0'
#775560000000
1!
b111 %
1'
b111 +
#775570000000
0!
0'
#775580000000
1!
0$
b1000 %
1'
0*
b1000 +
#775590000000
0!
0'
#775600000000
1!
b1001 %
1'
b1001 +
#775610000000
0!
0'
#775620000000
1!
b0 %
1'
b0 +
#775630000000
0!
0'
#775640000000
1!
1$
b1 %
1'
1*
b1 +
#775650000000
0!
0'
#775660000000
1!
b10 %
1'
b10 +
#775670000000
0!
0'
#775680000000
1!
b11 %
1'
b11 +
#775690000000
0!
0'
#775700000000
1!
b100 %
1'
b100 +
#775710000000
0!
0'
#775720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#775730000000
0!
0'
#775740000000
1!
0$
b110 %
1'
0*
b110 +
#775750000000
0!
0'
#775760000000
1!
b111 %
1'
b111 +
#775770000000
0!
0'
#775780000000
1!
b1000 %
1'
b1000 +
#775790000000
0!
0'
#775800000000
1!
b1001 %
1'
b1001 +
#775810000000
0!
0'
#775820000000
1!
b0 %
1'
b0 +
#775830000000
0!
0'
#775840000000
1!
1$
b1 %
1'
1*
b1 +
#775850000000
0!
0'
#775860000000
1!
b10 %
1'
b10 +
#775870000000
0!
0'
#775880000000
1!
b11 %
1'
b11 +
#775890000000
0!
0'
#775900000000
1!
b100 %
1'
b100 +
#775910000000
0!
0'
#775920000000
1!
b101 %
1'
b101 +
#775930000000
1"
1(
#775940000000
0!
0"
b100 &
0'
0(
b100 ,
#775950000000
1!
b110 %
1'
b110 +
#775960000000
0!
0'
#775970000000
1!
b111 %
1'
b111 +
#775980000000
0!
0'
#775990000000
1!
0$
b1000 %
1'
0*
b1000 +
#776000000000
0!
0'
#776010000000
1!
b1001 %
1'
b1001 +
#776020000000
0!
0'
#776030000000
1!
b0 %
1'
b0 +
#776040000000
0!
0'
#776050000000
1!
1$
b1 %
1'
1*
b1 +
#776060000000
0!
0'
#776070000000
1!
b10 %
1'
b10 +
#776080000000
0!
0'
#776090000000
1!
b11 %
1'
b11 +
#776100000000
0!
0'
#776110000000
1!
b100 %
1'
b100 +
#776120000000
0!
0'
#776130000000
1!
b101 %
1'
b101 +
#776140000000
0!
0'
#776150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#776160000000
0!
0'
#776170000000
1!
b111 %
1'
b111 +
#776180000000
0!
0'
#776190000000
1!
b1000 %
1'
b1000 +
#776200000000
0!
0'
#776210000000
1!
b1001 %
1'
b1001 +
#776220000000
0!
0'
#776230000000
1!
b0 %
1'
b0 +
#776240000000
0!
0'
#776250000000
1!
1$
b1 %
1'
1*
b1 +
#776260000000
0!
0'
#776270000000
1!
b10 %
1'
b10 +
#776280000000
0!
0'
#776290000000
1!
b11 %
1'
b11 +
#776300000000
0!
0'
#776310000000
1!
b100 %
1'
b100 +
#776320000000
0!
0'
#776330000000
1!
b101 %
1'
b101 +
#776340000000
0!
0'
#776350000000
1!
0$
b110 %
1'
0*
b110 +
#776360000000
1"
1(
#776370000000
0!
0"
b100 &
0'
0(
b100 ,
#776380000000
1!
1$
b111 %
1'
1*
b111 +
#776390000000
0!
0'
#776400000000
1!
0$
b1000 %
1'
0*
b1000 +
#776410000000
0!
0'
#776420000000
1!
b1001 %
1'
b1001 +
#776430000000
0!
0'
#776440000000
1!
b0 %
1'
b0 +
#776450000000
0!
0'
#776460000000
1!
1$
b1 %
1'
1*
b1 +
#776470000000
0!
0'
#776480000000
1!
b10 %
1'
b10 +
#776490000000
0!
0'
#776500000000
1!
b11 %
1'
b11 +
#776510000000
0!
0'
#776520000000
1!
b100 %
1'
b100 +
#776530000000
0!
0'
#776540000000
1!
b101 %
1'
b101 +
#776550000000
0!
0'
#776560000000
1!
b110 %
1'
b110 +
#776570000000
0!
0'
#776580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#776590000000
0!
0'
#776600000000
1!
b1000 %
1'
b1000 +
#776610000000
0!
0'
#776620000000
1!
b1001 %
1'
b1001 +
#776630000000
0!
0'
#776640000000
1!
b0 %
1'
b0 +
#776650000000
0!
0'
#776660000000
1!
1$
b1 %
1'
1*
b1 +
#776670000000
0!
0'
#776680000000
1!
b10 %
1'
b10 +
#776690000000
0!
0'
#776700000000
1!
b11 %
1'
b11 +
#776710000000
0!
0'
#776720000000
1!
b100 %
1'
b100 +
#776730000000
0!
0'
#776740000000
1!
b101 %
1'
b101 +
#776750000000
0!
0'
#776760000000
1!
0$
b110 %
1'
0*
b110 +
#776770000000
0!
0'
#776780000000
1!
b111 %
1'
b111 +
#776790000000
1"
1(
#776800000000
0!
0"
b100 &
0'
0(
b100 ,
#776810000000
1!
b1000 %
1'
b1000 +
#776820000000
0!
0'
#776830000000
1!
b1001 %
1'
b1001 +
#776840000000
0!
0'
#776850000000
1!
b0 %
1'
b0 +
#776860000000
0!
0'
#776870000000
1!
1$
b1 %
1'
1*
b1 +
#776880000000
0!
0'
#776890000000
1!
b10 %
1'
b10 +
#776900000000
0!
0'
#776910000000
1!
b11 %
1'
b11 +
#776920000000
0!
0'
#776930000000
1!
b100 %
1'
b100 +
#776940000000
0!
0'
#776950000000
1!
b101 %
1'
b101 +
#776960000000
0!
0'
#776970000000
1!
b110 %
1'
b110 +
#776980000000
0!
0'
#776990000000
1!
b111 %
1'
b111 +
#777000000000
0!
0'
#777010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#777020000000
0!
0'
#777030000000
1!
b1001 %
1'
b1001 +
#777040000000
0!
0'
#777050000000
1!
b0 %
1'
b0 +
#777060000000
0!
0'
#777070000000
1!
1$
b1 %
1'
1*
b1 +
#777080000000
0!
0'
#777090000000
1!
b10 %
1'
b10 +
#777100000000
0!
0'
#777110000000
1!
b11 %
1'
b11 +
#777120000000
0!
0'
#777130000000
1!
b100 %
1'
b100 +
#777140000000
0!
0'
#777150000000
1!
b101 %
1'
b101 +
#777160000000
0!
0'
#777170000000
1!
0$
b110 %
1'
0*
b110 +
#777180000000
0!
0'
#777190000000
1!
b111 %
1'
b111 +
#777200000000
0!
0'
#777210000000
1!
b1000 %
1'
b1000 +
#777220000000
1"
1(
#777230000000
0!
0"
b100 &
0'
0(
b100 ,
#777240000000
1!
b1001 %
1'
b1001 +
#777250000000
0!
0'
#777260000000
1!
b0 %
1'
b0 +
#777270000000
0!
0'
#777280000000
1!
1$
b1 %
1'
1*
b1 +
#777290000000
0!
0'
#777300000000
1!
b10 %
1'
b10 +
#777310000000
0!
0'
#777320000000
1!
b11 %
1'
b11 +
#777330000000
0!
0'
#777340000000
1!
b100 %
1'
b100 +
#777350000000
0!
0'
#777360000000
1!
b101 %
1'
b101 +
#777370000000
0!
0'
#777380000000
1!
b110 %
1'
b110 +
#777390000000
0!
0'
#777400000000
1!
b111 %
1'
b111 +
#777410000000
0!
0'
#777420000000
1!
0$
b1000 %
1'
0*
b1000 +
#777430000000
0!
0'
#777440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#777450000000
0!
0'
#777460000000
1!
b0 %
1'
b0 +
#777470000000
0!
0'
#777480000000
1!
1$
b1 %
1'
1*
b1 +
#777490000000
0!
0'
#777500000000
1!
b10 %
1'
b10 +
#777510000000
0!
0'
#777520000000
1!
b11 %
1'
b11 +
#777530000000
0!
0'
#777540000000
1!
b100 %
1'
b100 +
#777550000000
0!
0'
#777560000000
1!
b101 %
1'
b101 +
#777570000000
0!
0'
#777580000000
1!
0$
b110 %
1'
0*
b110 +
#777590000000
0!
0'
#777600000000
1!
b111 %
1'
b111 +
#777610000000
0!
0'
#777620000000
1!
b1000 %
1'
b1000 +
#777630000000
0!
0'
#777640000000
1!
b1001 %
1'
b1001 +
#777650000000
1"
1(
#777660000000
0!
0"
b100 &
0'
0(
b100 ,
#777670000000
1!
b0 %
1'
b0 +
#777680000000
0!
0'
#777690000000
1!
1$
b1 %
1'
1*
b1 +
#777700000000
0!
0'
#777710000000
1!
b10 %
1'
b10 +
#777720000000
0!
0'
#777730000000
1!
b11 %
1'
b11 +
#777740000000
0!
0'
#777750000000
1!
b100 %
1'
b100 +
#777760000000
0!
0'
#777770000000
1!
b101 %
1'
b101 +
#777780000000
0!
0'
#777790000000
1!
b110 %
1'
b110 +
#777800000000
0!
0'
#777810000000
1!
b111 %
1'
b111 +
#777820000000
0!
0'
#777830000000
1!
0$
b1000 %
1'
0*
b1000 +
#777840000000
0!
0'
#777850000000
1!
b1001 %
1'
b1001 +
#777860000000
0!
0'
#777870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#777880000000
0!
0'
#777890000000
1!
1$
b1 %
1'
1*
b1 +
#777900000000
0!
0'
#777910000000
1!
b10 %
1'
b10 +
#777920000000
0!
0'
#777930000000
1!
b11 %
1'
b11 +
#777940000000
0!
0'
#777950000000
1!
b100 %
1'
b100 +
#777960000000
0!
0'
#777970000000
1!
b101 %
1'
b101 +
#777980000000
0!
0'
#777990000000
1!
0$
b110 %
1'
0*
b110 +
#778000000000
0!
0'
#778010000000
1!
b111 %
1'
b111 +
#778020000000
0!
0'
#778030000000
1!
b1000 %
1'
b1000 +
#778040000000
0!
0'
#778050000000
1!
b1001 %
1'
b1001 +
#778060000000
0!
0'
#778070000000
1!
b0 %
1'
b0 +
#778080000000
1"
1(
#778090000000
0!
0"
b100 &
0'
0(
b100 ,
#778100000000
1!
1$
b1 %
1'
1*
b1 +
#778110000000
0!
0'
#778120000000
1!
b10 %
1'
b10 +
#778130000000
0!
0'
#778140000000
1!
b11 %
1'
b11 +
#778150000000
0!
0'
#778160000000
1!
b100 %
1'
b100 +
#778170000000
0!
0'
#778180000000
1!
b101 %
1'
b101 +
#778190000000
0!
0'
#778200000000
1!
b110 %
1'
b110 +
#778210000000
0!
0'
#778220000000
1!
b111 %
1'
b111 +
#778230000000
0!
0'
#778240000000
1!
0$
b1000 %
1'
0*
b1000 +
#778250000000
0!
0'
#778260000000
1!
b1001 %
1'
b1001 +
#778270000000
0!
0'
#778280000000
1!
b0 %
1'
b0 +
#778290000000
0!
0'
#778300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#778310000000
0!
0'
#778320000000
1!
b10 %
1'
b10 +
#778330000000
0!
0'
#778340000000
1!
b11 %
1'
b11 +
#778350000000
0!
0'
#778360000000
1!
b100 %
1'
b100 +
#778370000000
0!
0'
#778380000000
1!
b101 %
1'
b101 +
#778390000000
0!
0'
#778400000000
1!
0$
b110 %
1'
0*
b110 +
#778410000000
0!
0'
#778420000000
1!
b111 %
1'
b111 +
#778430000000
0!
0'
#778440000000
1!
b1000 %
1'
b1000 +
#778450000000
0!
0'
#778460000000
1!
b1001 %
1'
b1001 +
#778470000000
0!
0'
#778480000000
1!
b0 %
1'
b0 +
#778490000000
0!
0'
#778500000000
1!
1$
b1 %
1'
1*
b1 +
#778510000000
1"
1(
#778520000000
0!
0"
b100 &
0'
0(
b100 ,
#778530000000
1!
b10 %
1'
b10 +
#778540000000
0!
0'
#778550000000
1!
b11 %
1'
b11 +
#778560000000
0!
0'
#778570000000
1!
b100 %
1'
b100 +
#778580000000
0!
0'
#778590000000
1!
b101 %
1'
b101 +
#778600000000
0!
0'
#778610000000
1!
b110 %
1'
b110 +
#778620000000
0!
0'
#778630000000
1!
b111 %
1'
b111 +
#778640000000
0!
0'
#778650000000
1!
0$
b1000 %
1'
0*
b1000 +
#778660000000
0!
0'
#778670000000
1!
b1001 %
1'
b1001 +
#778680000000
0!
0'
#778690000000
1!
b0 %
1'
b0 +
#778700000000
0!
0'
#778710000000
1!
1$
b1 %
1'
1*
b1 +
#778720000000
0!
0'
#778730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#778740000000
0!
0'
#778750000000
1!
b11 %
1'
b11 +
#778760000000
0!
0'
#778770000000
1!
b100 %
1'
b100 +
#778780000000
0!
0'
#778790000000
1!
b101 %
1'
b101 +
#778800000000
0!
0'
#778810000000
1!
0$
b110 %
1'
0*
b110 +
#778820000000
0!
0'
#778830000000
1!
b111 %
1'
b111 +
#778840000000
0!
0'
#778850000000
1!
b1000 %
1'
b1000 +
#778860000000
0!
0'
#778870000000
1!
b1001 %
1'
b1001 +
#778880000000
0!
0'
#778890000000
1!
b0 %
1'
b0 +
#778900000000
0!
0'
#778910000000
1!
1$
b1 %
1'
1*
b1 +
#778920000000
0!
0'
#778930000000
1!
b10 %
1'
b10 +
#778940000000
1"
1(
#778950000000
0!
0"
b100 &
0'
0(
b100 ,
#778960000000
1!
b11 %
1'
b11 +
#778970000000
0!
0'
#778980000000
1!
b100 %
1'
b100 +
#778990000000
0!
0'
#779000000000
1!
b101 %
1'
b101 +
#779010000000
0!
0'
#779020000000
1!
b110 %
1'
b110 +
#779030000000
0!
0'
#779040000000
1!
b111 %
1'
b111 +
#779050000000
0!
0'
#779060000000
1!
0$
b1000 %
1'
0*
b1000 +
#779070000000
0!
0'
#779080000000
1!
b1001 %
1'
b1001 +
#779090000000
0!
0'
#779100000000
1!
b0 %
1'
b0 +
#779110000000
0!
0'
#779120000000
1!
1$
b1 %
1'
1*
b1 +
#779130000000
0!
0'
#779140000000
1!
b10 %
1'
b10 +
#779150000000
0!
0'
#779160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#779170000000
0!
0'
#779180000000
1!
b100 %
1'
b100 +
#779190000000
0!
0'
#779200000000
1!
b101 %
1'
b101 +
#779210000000
0!
0'
#779220000000
1!
0$
b110 %
1'
0*
b110 +
#779230000000
0!
0'
#779240000000
1!
b111 %
1'
b111 +
#779250000000
0!
0'
#779260000000
1!
b1000 %
1'
b1000 +
#779270000000
0!
0'
#779280000000
1!
b1001 %
1'
b1001 +
#779290000000
0!
0'
#779300000000
1!
b0 %
1'
b0 +
#779310000000
0!
0'
#779320000000
1!
1$
b1 %
1'
1*
b1 +
#779330000000
0!
0'
#779340000000
1!
b10 %
1'
b10 +
#779350000000
0!
0'
#779360000000
1!
b11 %
1'
b11 +
#779370000000
1"
1(
#779380000000
0!
0"
b100 &
0'
0(
b100 ,
#779390000000
1!
b100 %
1'
b100 +
#779400000000
0!
0'
#779410000000
1!
b101 %
1'
b101 +
#779420000000
0!
0'
#779430000000
1!
b110 %
1'
b110 +
#779440000000
0!
0'
#779450000000
1!
b111 %
1'
b111 +
#779460000000
0!
0'
#779470000000
1!
0$
b1000 %
1'
0*
b1000 +
#779480000000
0!
0'
#779490000000
1!
b1001 %
1'
b1001 +
#779500000000
0!
0'
#779510000000
1!
b0 %
1'
b0 +
#779520000000
0!
0'
#779530000000
1!
1$
b1 %
1'
1*
b1 +
#779540000000
0!
0'
#779550000000
1!
b10 %
1'
b10 +
#779560000000
0!
0'
#779570000000
1!
b11 %
1'
b11 +
#779580000000
0!
0'
#779590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#779600000000
0!
0'
#779610000000
1!
b101 %
1'
b101 +
#779620000000
0!
0'
#779630000000
1!
0$
b110 %
1'
0*
b110 +
#779640000000
0!
0'
#779650000000
1!
b111 %
1'
b111 +
#779660000000
0!
0'
#779670000000
1!
b1000 %
1'
b1000 +
#779680000000
0!
0'
#779690000000
1!
b1001 %
1'
b1001 +
#779700000000
0!
0'
#779710000000
1!
b0 %
1'
b0 +
#779720000000
0!
0'
#779730000000
1!
1$
b1 %
1'
1*
b1 +
#779740000000
0!
0'
#779750000000
1!
b10 %
1'
b10 +
#779760000000
0!
0'
#779770000000
1!
b11 %
1'
b11 +
#779780000000
0!
0'
#779790000000
1!
b100 %
1'
b100 +
#779800000000
1"
1(
#779810000000
0!
0"
b100 &
0'
0(
b100 ,
#779820000000
1!
b101 %
1'
b101 +
#779830000000
0!
0'
#779840000000
1!
b110 %
1'
b110 +
#779850000000
0!
0'
#779860000000
1!
b111 %
1'
b111 +
#779870000000
0!
0'
#779880000000
1!
0$
b1000 %
1'
0*
b1000 +
#779890000000
0!
0'
#779900000000
1!
b1001 %
1'
b1001 +
#779910000000
0!
0'
#779920000000
1!
b0 %
1'
b0 +
#779930000000
0!
0'
#779940000000
1!
1$
b1 %
1'
1*
b1 +
#779950000000
0!
0'
#779960000000
1!
b10 %
1'
b10 +
#779970000000
0!
0'
#779980000000
1!
b11 %
1'
b11 +
#779990000000
0!
0'
#780000000000
1!
b100 %
1'
b100 +
#780010000000
0!
0'
#780020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#780030000000
0!
0'
#780040000000
1!
0$
b110 %
1'
0*
b110 +
#780050000000
0!
0'
#780060000000
1!
b111 %
1'
b111 +
#780070000000
0!
0'
#780080000000
1!
b1000 %
1'
b1000 +
#780090000000
0!
0'
#780100000000
1!
b1001 %
1'
b1001 +
#780110000000
0!
0'
#780120000000
1!
b0 %
1'
b0 +
#780130000000
0!
0'
#780140000000
1!
1$
b1 %
1'
1*
b1 +
#780150000000
0!
0'
#780160000000
1!
b10 %
1'
b10 +
#780170000000
0!
0'
#780180000000
1!
b11 %
1'
b11 +
#780190000000
0!
0'
#780200000000
1!
b100 %
1'
b100 +
#780210000000
0!
0'
#780220000000
1!
b101 %
1'
b101 +
#780230000000
1"
1(
#780240000000
0!
0"
b100 &
0'
0(
b100 ,
#780250000000
1!
b110 %
1'
b110 +
#780260000000
0!
0'
#780270000000
1!
b111 %
1'
b111 +
#780280000000
0!
0'
#780290000000
1!
0$
b1000 %
1'
0*
b1000 +
#780300000000
0!
0'
#780310000000
1!
b1001 %
1'
b1001 +
#780320000000
0!
0'
#780330000000
1!
b0 %
1'
b0 +
#780340000000
0!
0'
#780350000000
1!
1$
b1 %
1'
1*
b1 +
#780360000000
0!
0'
#780370000000
1!
b10 %
1'
b10 +
#780380000000
0!
0'
#780390000000
1!
b11 %
1'
b11 +
#780400000000
0!
0'
#780410000000
1!
b100 %
1'
b100 +
#780420000000
0!
0'
#780430000000
1!
b101 %
1'
b101 +
#780440000000
0!
0'
#780450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#780460000000
0!
0'
#780470000000
1!
b111 %
1'
b111 +
#780480000000
0!
0'
#780490000000
1!
b1000 %
1'
b1000 +
#780500000000
0!
0'
#780510000000
1!
b1001 %
1'
b1001 +
#780520000000
0!
0'
#780530000000
1!
b0 %
1'
b0 +
#780540000000
0!
0'
#780550000000
1!
1$
b1 %
1'
1*
b1 +
#780560000000
0!
0'
#780570000000
1!
b10 %
1'
b10 +
#780580000000
0!
0'
#780590000000
1!
b11 %
1'
b11 +
#780600000000
0!
0'
#780610000000
1!
b100 %
1'
b100 +
#780620000000
0!
0'
#780630000000
1!
b101 %
1'
b101 +
#780640000000
0!
0'
#780650000000
1!
0$
b110 %
1'
0*
b110 +
#780660000000
1"
1(
#780670000000
0!
0"
b100 &
0'
0(
b100 ,
#780680000000
1!
1$
b111 %
1'
1*
b111 +
#780690000000
0!
0'
#780700000000
1!
0$
b1000 %
1'
0*
b1000 +
#780710000000
0!
0'
#780720000000
1!
b1001 %
1'
b1001 +
#780730000000
0!
0'
#780740000000
1!
b0 %
1'
b0 +
#780750000000
0!
0'
#780760000000
1!
1$
b1 %
1'
1*
b1 +
#780770000000
0!
0'
#780780000000
1!
b10 %
1'
b10 +
#780790000000
0!
0'
#780800000000
1!
b11 %
1'
b11 +
#780810000000
0!
0'
#780820000000
1!
b100 %
1'
b100 +
#780830000000
0!
0'
#780840000000
1!
b101 %
1'
b101 +
#780850000000
0!
0'
#780860000000
1!
b110 %
1'
b110 +
#780870000000
0!
0'
#780880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#780890000000
0!
0'
#780900000000
1!
b1000 %
1'
b1000 +
#780910000000
0!
0'
#780920000000
1!
b1001 %
1'
b1001 +
#780930000000
0!
0'
#780940000000
1!
b0 %
1'
b0 +
#780950000000
0!
0'
#780960000000
1!
1$
b1 %
1'
1*
b1 +
#780970000000
0!
0'
#780980000000
1!
b10 %
1'
b10 +
#780990000000
0!
0'
#781000000000
1!
b11 %
1'
b11 +
#781010000000
0!
0'
#781020000000
1!
b100 %
1'
b100 +
#781030000000
0!
0'
#781040000000
1!
b101 %
1'
b101 +
#781050000000
0!
0'
#781060000000
1!
0$
b110 %
1'
0*
b110 +
#781070000000
0!
0'
#781080000000
1!
b111 %
1'
b111 +
#781090000000
1"
1(
#781100000000
0!
0"
b100 &
0'
0(
b100 ,
#781110000000
1!
b1000 %
1'
b1000 +
#781120000000
0!
0'
#781130000000
1!
b1001 %
1'
b1001 +
#781140000000
0!
0'
#781150000000
1!
b0 %
1'
b0 +
#781160000000
0!
0'
#781170000000
1!
1$
b1 %
1'
1*
b1 +
#781180000000
0!
0'
#781190000000
1!
b10 %
1'
b10 +
#781200000000
0!
0'
#781210000000
1!
b11 %
1'
b11 +
#781220000000
0!
0'
#781230000000
1!
b100 %
1'
b100 +
#781240000000
0!
0'
#781250000000
1!
b101 %
1'
b101 +
#781260000000
0!
0'
#781270000000
1!
b110 %
1'
b110 +
#781280000000
0!
0'
#781290000000
1!
b111 %
1'
b111 +
#781300000000
0!
0'
#781310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#781320000000
0!
0'
#781330000000
1!
b1001 %
1'
b1001 +
#781340000000
0!
0'
#781350000000
1!
b0 %
1'
b0 +
#781360000000
0!
0'
#781370000000
1!
1$
b1 %
1'
1*
b1 +
#781380000000
0!
0'
#781390000000
1!
b10 %
1'
b10 +
#781400000000
0!
0'
#781410000000
1!
b11 %
1'
b11 +
#781420000000
0!
0'
#781430000000
1!
b100 %
1'
b100 +
#781440000000
0!
0'
#781450000000
1!
b101 %
1'
b101 +
#781460000000
0!
0'
#781470000000
1!
0$
b110 %
1'
0*
b110 +
#781480000000
0!
0'
#781490000000
1!
b111 %
1'
b111 +
#781500000000
0!
0'
#781510000000
1!
b1000 %
1'
b1000 +
#781520000000
1"
1(
#781530000000
0!
0"
b100 &
0'
0(
b100 ,
#781540000000
1!
b1001 %
1'
b1001 +
#781550000000
0!
0'
#781560000000
1!
b0 %
1'
b0 +
#781570000000
0!
0'
#781580000000
1!
1$
b1 %
1'
1*
b1 +
#781590000000
0!
0'
#781600000000
1!
b10 %
1'
b10 +
#781610000000
0!
0'
#781620000000
1!
b11 %
1'
b11 +
#781630000000
0!
0'
#781640000000
1!
b100 %
1'
b100 +
#781650000000
0!
0'
#781660000000
1!
b101 %
1'
b101 +
#781670000000
0!
0'
#781680000000
1!
b110 %
1'
b110 +
#781690000000
0!
0'
#781700000000
1!
b111 %
1'
b111 +
#781710000000
0!
0'
#781720000000
1!
0$
b1000 %
1'
0*
b1000 +
#781730000000
0!
0'
#781740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#781750000000
0!
0'
#781760000000
1!
b0 %
1'
b0 +
#781770000000
0!
0'
#781780000000
1!
1$
b1 %
1'
1*
b1 +
#781790000000
0!
0'
#781800000000
1!
b10 %
1'
b10 +
#781810000000
0!
0'
#781820000000
1!
b11 %
1'
b11 +
#781830000000
0!
0'
#781840000000
1!
b100 %
1'
b100 +
#781850000000
0!
0'
#781860000000
1!
b101 %
1'
b101 +
#781870000000
0!
0'
#781880000000
1!
0$
b110 %
1'
0*
b110 +
#781890000000
0!
0'
#781900000000
1!
b111 %
1'
b111 +
#781910000000
0!
0'
#781920000000
1!
b1000 %
1'
b1000 +
#781930000000
0!
0'
#781940000000
1!
b1001 %
1'
b1001 +
#781950000000
1"
1(
#781960000000
0!
0"
b100 &
0'
0(
b100 ,
#781970000000
1!
b0 %
1'
b0 +
#781980000000
0!
0'
#781990000000
1!
1$
b1 %
1'
1*
b1 +
#782000000000
0!
0'
#782010000000
1!
b10 %
1'
b10 +
#782020000000
0!
0'
#782030000000
1!
b11 %
1'
b11 +
#782040000000
0!
0'
#782050000000
1!
b100 %
1'
b100 +
#782060000000
0!
0'
#782070000000
1!
b101 %
1'
b101 +
#782080000000
0!
0'
#782090000000
1!
b110 %
1'
b110 +
#782100000000
0!
0'
#782110000000
1!
b111 %
1'
b111 +
#782120000000
0!
0'
#782130000000
1!
0$
b1000 %
1'
0*
b1000 +
#782140000000
0!
0'
#782150000000
1!
b1001 %
1'
b1001 +
#782160000000
0!
0'
#782170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#782180000000
0!
0'
#782190000000
1!
1$
b1 %
1'
1*
b1 +
#782200000000
0!
0'
#782210000000
1!
b10 %
1'
b10 +
#782220000000
0!
0'
#782230000000
1!
b11 %
1'
b11 +
#782240000000
0!
0'
#782250000000
1!
b100 %
1'
b100 +
#782260000000
0!
0'
#782270000000
1!
b101 %
1'
b101 +
#782280000000
0!
0'
#782290000000
1!
0$
b110 %
1'
0*
b110 +
#782300000000
0!
0'
#782310000000
1!
b111 %
1'
b111 +
#782320000000
0!
0'
#782330000000
1!
b1000 %
1'
b1000 +
#782340000000
0!
0'
#782350000000
1!
b1001 %
1'
b1001 +
#782360000000
0!
0'
#782370000000
1!
b0 %
1'
b0 +
#782380000000
1"
1(
#782390000000
0!
0"
b100 &
0'
0(
b100 ,
#782400000000
1!
1$
b1 %
1'
1*
b1 +
#782410000000
0!
0'
#782420000000
1!
b10 %
1'
b10 +
#782430000000
0!
0'
#782440000000
1!
b11 %
1'
b11 +
#782450000000
0!
0'
#782460000000
1!
b100 %
1'
b100 +
#782470000000
0!
0'
#782480000000
1!
b101 %
1'
b101 +
#782490000000
0!
0'
#782500000000
1!
b110 %
1'
b110 +
#782510000000
0!
0'
#782520000000
1!
b111 %
1'
b111 +
#782530000000
0!
0'
#782540000000
1!
0$
b1000 %
1'
0*
b1000 +
#782550000000
0!
0'
#782560000000
1!
b1001 %
1'
b1001 +
#782570000000
0!
0'
#782580000000
1!
b0 %
1'
b0 +
#782590000000
0!
0'
#782600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#782610000000
0!
0'
#782620000000
1!
b10 %
1'
b10 +
#782630000000
0!
0'
#782640000000
1!
b11 %
1'
b11 +
#782650000000
0!
0'
#782660000000
1!
b100 %
1'
b100 +
#782670000000
0!
0'
#782680000000
1!
b101 %
1'
b101 +
#782690000000
0!
0'
#782700000000
1!
0$
b110 %
1'
0*
b110 +
#782710000000
0!
0'
#782720000000
1!
b111 %
1'
b111 +
#782730000000
0!
0'
#782740000000
1!
b1000 %
1'
b1000 +
#782750000000
0!
0'
#782760000000
1!
b1001 %
1'
b1001 +
#782770000000
0!
0'
#782780000000
1!
b0 %
1'
b0 +
#782790000000
0!
0'
#782800000000
1!
1$
b1 %
1'
1*
b1 +
#782810000000
1"
1(
#782820000000
0!
0"
b100 &
0'
0(
b100 ,
#782830000000
1!
b10 %
1'
b10 +
#782840000000
0!
0'
#782850000000
1!
b11 %
1'
b11 +
#782860000000
0!
0'
#782870000000
1!
b100 %
1'
b100 +
#782880000000
0!
0'
#782890000000
1!
b101 %
1'
b101 +
#782900000000
0!
0'
#782910000000
1!
b110 %
1'
b110 +
#782920000000
0!
0'
#782930000000
1!
b111 %
1'
b111 +
#782940000000
0!
0'
#782950000000
1!
0$
b1000 %
1'
0*
b1000 +
#782960000000
0!
0'
#782970000000
1!
b1001 %
1'
b1001 +
#782980000000
0!
0'
#782990000000
1!
b0 %
1'
b0 +
#783000000000
0!
0'
#783010000000
1!
1$
b1 %
1'
1*
b1 +
#783020000000
0!
0'
#783030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#783040000000
0!
0'
#783050000000
1!
b11 %
1'
b11 +
#783060000000
0!
0'
#783070000000
1!
b100 %
1'
b100 +
#783080000000
0!
0'
#783090000000
1!
b101 %
1'
b101 +
#783100000000
0!
0'
#783110000000
1!
0$
b110 %
1'
0*
b110 +
#783120000000
0!
0'
#783130000000
1!
b111 %
1'
b111 +
#783140000000
0!
0'
#783150000000
1!
b1000 %
1'
b1000 +
#783160000000
0!
0'
#783170000000
1!
b1001 %
1'
b1001 +
#783180000000
0!
0'
#783190000000
1!
b0 %
1'
b0 +
#783200000000
0!
0'
#783210000000
1!
1$
b1 %
1'
1*
b1 +
#783220000000
0!
0'
#783230000000
1!
b10 %
1'
b10 +
#783240000000
1"
1(
#783250000000
0!
0"
b100 &
0'
0(
b100 ,
#783260000000
1!
b11 %
1'
b11 +
#783270000000
0!
0'
#783280000000
1!
b100 %
1'
b100 +
#783290000000
0!
0'
#783300000000
1!
b101 %
1'
b101 +
#783310000000
0!
0'
#783320000000
1!
b110 %
1'
b110 +
#783330000000
0!
0'
#783340000000
1!
b111 %
1'
b111 +
#783350000000
0!
0'
#783360000000
1!
0$
b1000 %
1'
0*
b1000 +
#783370000000
0!
0'
#783380000000
1!
b1001 %
1'
b1001 +
#783390000000
0!
0'
#783400000000
1!
b0 %
1'
b0 +
#783410000000
0!
0'
#783420000000
1!
1$
b1 %
1'
1*
b1 +
#783430000000
0!
0'
#783440000000
1!
b10 %
1'
b10 +
#783450000000
0!
0'
#783460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#783470000000
0!
0'
#783480000000
1!
b100 %
1'
b100 +
#783490000000
0!
0'
#783500000000
1!
b101 %
1'
b101 +
#783510000000
0!
0'
#783520000000
1!
0$
b110 %
1'
0*
b110 +
#783530000000
0!
0'
#783540000000
1!
b111 %
1'
b111 +
#783550000000
0!
0'
#783560000000
1!
b1000 %
1'
b1000 +
#783570000000
0!
0'
#783580000000
1!
b1001 %
1'
b1001 +
#783590000000
0!
0'
#783600000000
1!
b0 %
1'
b0 +
#783610000000
0!
0'
#783620000000
1!
1$
b1 %
1'
1*
b1 +
#783630000000
0!
0'
#783640000000
1!
b10 %
1'
b10 +
#783650000000
0!
0'
#783660000000
1!
b11 %
1'
b11 +
#783670000000
1"
1(
#783680000000
0!
0"
b100 &
0'
0(
b100 ,
#783690000000
1!
b100 %
1'
b100 +
#783700000000
0!
0'
#783710000000
1!
b101 %
1'
b101 +
#783720000000
0!
0'
#783730000000
1!
b110 %
1'
b110 +
#783740000000
0!
0'
#783750000000
1!
b111 %
1'
b111 +
#783760000000
0!
0'
#783770000000
1!
0$
b1000 %
1'
0*
b1000 +
#783780000000
0!
0'
#783790000000
1!
b1001 %
1'
b1001 +
#783800000000
0!
0'
#783810000000
1!
b0 %
1'
b0 +
#783820000000
0!
0'
#783830000000
1!
1$
b1 %
1'
1*
b1 +
#783840000000
0!
0'
#783850000000
1!
b10 %
1'
b10 +
#783860000000
0!
0'
#783870000000
1!
b11 %
1'
b11 +
#783880000000
0!
0'
#783890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#783900000000
0!
0'
#783910000000
1!
b101 %
1'
b101 +
#783920000000
0!
0'
#783930000000
1!
0$
b110 %
1'
0*
b110 +
#783940000000
0!
0'
#783950000000
1!
b111 %
1'
b111 +
#783960000000
0!
0'
#783970000000
1!
b1000 %
1'
b1000 +
#783980000000
0!
0'
#783990000000
1!
b1001 %
1'
b1001 +
#784000000000
0!
0'
#784010000000
1!
b0 %
1'
b0 +
#784020000000
0!
0'
#784030000000
1!
1$
b1 %
1'
1*
b1 +
#784040000000
0!
0'
#784050000000
1!
b10 %
1'
b10 +
#784060000000
0!
0'
#784070000000
1!
b11 %
1'
b11 +
#784080000000
0!
0'
#784090000000
1!
b100 %
1'
b100 +
#784100000000
1"
1(
#784110000000
0!
0"
b100 &
0'
0(
b100 ,
#784120000000
1!
b101 %
1'
b101 +
#784130000000
0!
0'
#784140000000
1!
b110 %
1'
b110 +
#784150000000
0!
0'
#784160000000
1!
b111 %
1'
b111 +
#784170000000
0!
0'
#784180000000
1!
0$
b1000 %
1'
0*
b1000 +
#784190000000
0!
0'
#784200000000
1!
b1001 %
1'
b1001 +
#784210000000
0!
0'
#784220000000
1!
b0 %
1'
b0 +
#784230000000
0!
0'
#784240000000
1!
1$
b1 %
1'
1*
b1 +
#784250000000
0!
0'
#784260000000
1!
b10 %
1'
b10 +
#784270000000
0!
0'
#784280000000
1!
b11 %
1'
b11 +
#784290000000
0!
0'
#784300000000
1!
b100 %
1'
b100 +
#784310000000
0!
0'
#784320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#784330000000
0!
0'
#784340000000
1!
0$
b110 %
1'
0*
b110 +
#784350000000
0!
0'
#784360000000
1!
b111 %
1'
b111 +
#784370000000
0!
0'
#784380000000
1!
b1000 %
1'
b1000 +
#784390000000
0!
0'
#784400000000
1!
b1001 %
1'
b1001 +
#784410000000
0!
0'
#784420000000
1!
b0 %
1'
b0 +
#784430000000
0!
0'
#784440000000
1!
1$
b1 %
1'
1*
b1 +
#784450000000
0!
0'
#784460000000
1!
b10 %
1'
b10 +
#784470000000
0!
0'
#784480000000
1!
b11 %
1'
b11 +
#784490000000
0!
0'
#784500000000
1!
b100 %
1'
b100 +
#784510000000
0!
0'
#784520000000
1!
b101 %
1'
b101 +
#784530000000
1"
1(
#784540000000
0!
0"
b100 &
0'
0(
b100 ,
#784550000000
1!
b110 %
1'
b110 +
#784560000000
0!
0'
#784570000000
1!
b111 %
1'
b111 +
#784580000000
0!
0'
#784590000000
1!
0$
b1000 %
1'
0*
b1000 +
#784600000000
0!
0'
#784610000000
1!
b1001 %
1'
b1001 +
#784620000000
0!
0'
#784630000000
1!
b0 %
1'
b0 +
#784640000000
0!
0'
#784650000000
1!
1$
b1 %
1'
1*
b1 +
#784660000000
0!
0'
#784670000000
1!
b10 %
1'
b10 +
#784680000000
0!
0'
#784690000000
1!
b11 %
1'
b11 +
#784700000000
0!
0'
#784710000000
1!
b100 %
1'
b100 +
#784720000000
0!
0'
#784730000000
1!
b101 %
1'
b101 +
#784740000000
0!
0'
#784750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#784760000000
0!
0'
#784770000000
1!
b111 %
1'
b111 +
#784780000000
0!
0'
#784790000000
1!
b1000 %
1'
b1000 +
#784800000000
0!
0'
#784810000000
1!
b1001 %
1'
b1001 +
#784820000000
0!
0'
#784830000000
1!
b0 %
1'
b0 +
#784840000000
0!
0'
#784850000000
1!
1$
b1 %
1'
1*
b1 +
#784860000000
0!
0'
#784870000000
1!
b10 %
1'
b10 +
#784880000000
0!
0'
#784890000000
1!
b11 %
1'
b11 +
#784900000000
0!
0'
#784910000000
1!
b100 %
1'
b100 +
#784920000000
0!
0'
#784930000000
1!
b101 %
1'
b101 +
#784940000000
0!
0'
#784950000000
1!
0$
b110 %
1'
0*
b110 +
#784960000000
1"
1(
#784970000000
0!
0"
b100 &
0'
0(
b100 ,
#784980000000
1!
1$
b111 %
1'
1*
b111 +
#784990000000
0!
0'
#785000000000
1!
0$
b1000 %
1'
0*
b1000 +
#785010000000
0!
0'
#785020000000
1!
b1001 %
1'
b1001 +
#785030000000
0!
0'
#785040000000
1!
b0 %
1'
b0 +
#785050000000
0!
0'
#785060000000
1!
1$
b1 %
1'
1*
b1 +
#785070000000
0!
0'
#785080000000
1!
b10 %
1'
b10 +
#785090000000
0!
0'
#785100000000
1!
b11 %
1'
b11 +
#785110000000
0!
0'
#785120000000
1!
b100 %
1'
b100 +
#785130000000
0!
0'
#785140000000
1!
b101 %
1'
b101 +
#785150000000
0!
0'
#785160000000
1!
b110 %
1'
b110 +
#785170000000
0!
0'
#785180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#785190000000
0!
0'
#785200000000
1!
b1000 %
1'
b1000 +
#785210000000
0!
0'
#785220000000
1!
b1001 %
1'
b1001 +
#785230000000
0!
0'
#785240000000
1!
b0 %
1'
b0 +
#785250000000
0!
0'
#785260000000
1!
1$
b1 %
1'
1*
b1 +
#785270000000
0!
0'
#785280000000
1!
b10 %
1'
b10 +
#785290000000
0!
0'
#785300000000
1!
b11 %
1'
b11 +
#785310000000
0!
0'
#785320000000
1!
b100 %
1'
b100 +
#785330000000
0!
0'
#785340000000
1!
b101 %
1'
b101 +
#785350000000
0!
0'
#785360000000
1!
0$
b110 %
1'
0*
b110 +
#785370000000
0!
0'
#785380000000
1!
b111 %
1'
b111 +
#785390000000
1"
1(
#785400000000
0!
0"
b100 &
0'
0(
b100 ,
#785410000000
1!
b1000 %
1'
b1000 +
#785420000000
0!
0'
#785430000000
1!
b1001 %
1'
b1001 +
#785440000000
0!
0'
#785450000000
1!
b0 %
1'
b0 +
#785460000000
0!
0'
#785470000000
1!
1$
b1 %
1'
1*
b1 +
#785480000000
0!
0'
#785490000000
1!
b10 %
1'
b10 +
#785500000000
0!
0'
#785510000000
1!
b11 %
1'
b11 +
#785520000000
0!
0'
#785530000000
1!
b100 %
1'
b100 +
#785540000000
0!
0'
#785550000000
1!
b101 %
1'
b101 +
#785560000000
0!
0'
#785570000000
1!
b110 %
1'
b110 +
#785580000000
0!
0'
#785590000000
1!
b111 %
1'
b111 +
#785600000000
0!
0'
#785610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#785620000000
0!
0'
#785630000000
1!
b1001 %
1'
b1001 +
#785640000000
0!
0'
#785650000000
1!
b0 %
1'
b0 +
#785660000000
0!
0'
#785670000000
1!
1$
b1 %
1'
1*
b1 +
#785680000000
0!
0'
#785690000000
1!
b10 %
1'
b10 +
#785700000000
0!
0'
#785710000000
1!
b11 %
1'
b11 +
#785720000000
0!
0'
#785730000000
1!
b100 %
1'
b100 +
#785740000000
0!
0'
#785750000000
1!
b101 %
1'
b101 +
#785760000000
0!
0'
#785770000000
1!
0$
b110 %
1'
0*
b110 +
#785780000000
0!
0'
#785790000000
1!
b111 %
1'
b111 +
#785800000000
0!
0'
#785810000000
1!
b1000 %
1'
b1000 +
#785820000000
1"
1(
#785830000000
0!
0"
b100 &
0'
0(
b100 ,
#785840000000
1!
b1001 %
1'
b1001 +
#785850000000
0!
0'
#785860000000
1!
b0 %
1'
b0 +
#785870000000
0!
0'
#785880000000
1!
1$
b1 %
1'
1*
b1 +
#785890000000
0!
0'
#785900000000
1!
b10 %
1'
b10 +
#785910000000
0!
0'
#785920000000
1!
b11 %
1'
b11 +
#785930000000
0!
0'
#785940000000
1!
b100 %
1'
b100 +
#785950000000
0!
0'
#785960000000
1!
b101 %
1'
b101 +
#785970000000
0!
0'
#785980000000
1!
b110 %
1'
b110 +
#785990000000
0!
0'
#786000000000
1!
b111 %
1'
b111 +
#786010000000
0!
0'
#786020000000
1!
0$
b1000 %
1'
0*
b1000 +
#786030000000
0!
0'
#786040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#786050000000
0!
0'
#786060000000
1!
b0 %
1'
b0 +
#786070000000
0!
0'
#786080000000
1!
1$
b1 %
1'
1*
b1 +
#786090000000
0!
0'
#786100000000
1!
b10 %
1'
b10 +
#786110000000
0!
0'
#786120000000
1!
b11 %
1'
b11 +
#786130000000
0!
0'
#786140000000
1!
b100 %
1'
b100 +
#786150000000
0!
0'
#786160000000
1!
b101 %
1'
b101 +
#786170000000
0!
0'
#786180000000
1!
0$
b110 %
1'
0*
b110 +
#786190000000
0!
0'
#786200000000
1!
b111 %
1'
b111 +
#786210000000
0!
0'
#786220000000
1!
b1000 %
1'
b1000 +
#786230000000
0!
0'
#786240000000
1!
b1001 %
1'
b1001 +
#786250000000
1"
1(
#786260000000
0!
0"
b100 &
0'
0(
b100 ,
#786270000000
1!
b0 %
1'
b0 +
#786280000000
0!
0'
#786290000000
1!
1$
b1 %
1'
1*
b1 +
#786300000000
0!
0'
#786310000000
1!
b10 %
1'
b10 +
#786320000000
0!
0'
#786330000000
1!
b11 %
1'
b11 +
#786340000000
0!
0'
#786350000000
1!
b100 %
1'
b100 +
#786360000000
0!
0'
#786370000000
1!
b101 %
1'
b101 +
#786380000000
0!
0'
#786390000000
1!
b110 %
1'
b110 +
#786400000000
0!
0'
#786410000000
1!
b111 %
1'
b111 +
#786420000000
0!
0'
#786430000000
1!
0$
b1000 %
1'
0*
b1000 +
#786440000000
0!
0'
#786450000000
1!
b1001 %
1'
b1001 +
#786460000000
0!
0'
#786470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#786480000000
0!
0'
#786490000000
1!
1$
b1 %
1'
1*
b1 +
#786500000000
0!
0'
#786510000000
1!
b10 %
1'
b10 +
#786520000000
0!
0'
#786530000000
1!
b11 %
1'
b11 +
#786540000000
0!
0'
#786550000000
1!
b100 %
1'
b100 +
#786560000000
0!
0'
#786570000000
1!
b101 %
1'
b101 +
#786580000000
0!
0'
#786590000000
1!
0$
b110 %
1'
0*
b110 +
#786600000000
0!
0'
#786610000000
1!
b111 %
1'
b111 +
#786620000000
0!
0'
#786630000000
1!
b1000 %
1'
b1000 +
#786640000000
0!
0'
#786650000000
1!
b1001 %
1'
b1001 +
#786660000000
0!
0'
#786670000000
1!
b0 %
1'
b0 +
#786680000000
1"
1(
#786690000000
0!
0"
b100 &
0'
0(
b100 ,
#786700000000
1!
1$
b1 %
1'
1*
b1 +
#786710000000
0!
0'
#786720000000
1!
b10 %
1'
b10 +
#786730000000
0!
0'
#786740000000
1!
b11 %
1'
b11 +
#786750000000
0!
0'
#786760000000
1!
b100 %
1'
b100 +
#786770000000
0!
0'
#786780000000
1!
b101 %
1'
b101 +
#786790000000
0!
0'
#786800000000
1!
b110 %
1'
b110 +
#786810000000
0!
0'
#786820000000
1!
b111 %
1'
b111 +
#786830000000
0!
0'
#786840000000
1!
0$
b1000 %
1'
0*
b1000 +
#786850000000
0!
0'
#786860000000
1!
b1001 %
1'
b1001 +
#786870000000
0!
0'
#786880000000
1!
b0 %
1'
b0 +
#786890000000
0!
0'
#786900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#786910000000
0!
0'
#786920000000
1!
b10 %
1'
b10 +
#786930000000
0!
0'
#786940000000
1!
b11 %
1'
b11 +
#786950000000
0!
0'
#786960000000
1!
b100 %
1'
b100 +
#786970000000
0!
0'
#786980000000
1!
b101 %
1'
b101 +
#786990000000
0!
0'
#787000000000
1!
0$
b110 %
1'
0*
b110 +
#787010000000
0!
0'
#787020000000
1!
b111 %
1'
b111 +
#787030000000
0!
0'
#787040000000
1!
b1000 %
1'
b1000 +
#787050000000
0!
0'
#787060000000
1!
b1001 %
1'
b1001 +
#787070000000
0!
0'
#787080000000
1!
b0 %
1'
b0 +
#787090000000
0!
0'
#787100000000
1!
1$
b1 %
1'
1*
b1 +
#787110000000
1"
1(
#787120000000
0!
0"
b100 &
0'
0(
b100 ,
#787130000000
1!
b10 %
1'
b10 +
#787140000000
0!
0'
#787150000000
1!
b11 %
1'
b11 +
#787160000000
0!
0'
#787170000000
1!
b100 %
1'
b100 +
#787180000000
0!
0'
#787190000000
1!
b101 %
1'
b101 +
#787200000000
0!
0'
#787210000000
1!
b110 %
1'
b110 +
#787220000000
0!
0'
#787230000000
1!
b111 %
1'
b111 +
#787240000000
0!
0'
#787250000000
1!
0$
b1000 %
1'
0*
b1000 +
#787260000000
0!
0'
#787270000000
1!
b1001 %
1'
b1001 +
#787280000000
0!
0'
#787290000000
1!
b0 %
1'
b0 +
#787300000000
0!
0'
#787310000000
1!
1$
b1 %
1'
1*
b1 +
#787320000000
0!
0'
#787330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#787340000000
0!
0'
#787350000000
1!
b11 %
1'
b11 +
#787360000000
0!
0'
#787370000000
1!
b100 %
1'
b100 +
#787380000000
0!
0'
#787390000000
1!
b101 %
1'
b101 +
#787400000000
0!
0'
#787410000000
1!
0$
b110 %
1'
0*
b110 +
#787420000000
0!
0'
#787430000000
1!
b111 %
1'
b111 +
#787440000000
0!
0'
#787450000000
1!
b1000 %
1'
b1000 +
#787460000000
0!
0'
#787470000000
1!
b1001 %
1'
b1001 +
#787480000000
0!
0'
#787490000000
1!
b0 %
1'
b0 +
#787500000000
0!
0'
#787510000000
1!
1$
b1 %
1'
1*
b1 +
#787520000000
0!
0'
#787530000000
1!
b10 %
1'
b10 +
#787540000000
1"
1(
#787550000000
0!
0"
b100 &
0'
0(
b100 ,
#787560000000
1!
b11 %
1'
b11 +
#787570000000
0!
0'
#787580000000
1!
b100 %
1'
b100 +
#787590000000
0!
0'
#787600000000
1!
b101 %
1'
b101 +
#787610000000
0!
0'
#787620000000
1!
b110 %
1'
b110 +
#787630000000
0!
0'
#787640000000
1!
b111 %
1'
b111 +
#787650000000
0!
0'
#787660000000
1!
0$
b1000 %
1'
0*
b1000 +
#787670000000
0!
0'
#787680000000
1!
b1001 %
1'
b1001 +
#787690000000
0!
0'
#787700000000
1!
b0 %
1'
b0 +
#787710000000
0!
0'
#787720000000
1!
1$
b1 %
1'
1*
b1 +
#787730000000
0!
0'
#787740000000
1!
b10 %
1'
b10 +
#787750000000
0!
0'
#787760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#787770000000
0!
0'
#787780000000
1!
b100 %
1'
b100 +
#787790000000
0!
0'
#787800000000
1!
b101 %
1'
b101 +
#787810000000
0!
0'
#787820000000
1!
0$
b110 %
1'
0*
b110 +
#787830000000
0!
0'
#787840000000
1!
b111 %
1'
b111 +
#787850000000
0!
0'
#787860000000
1!
b1000 %
1'
b1000 +
#787870000000
0!
0'
#787880000000
1!
b1001 %
1'
b1001 +
#787890000000
0!
0'
#787900000000
1!
b0 %
1'
b0 +
#787910000000
0!
0'
#787920000000
1!
1$
b1 %
1'
1*
b1 +
#787930000000
0!
0'
#787940000000
1!
b10 %
1'
b10 +
#787950000000
0!
0'
#787960000000
1!
b11 %
1'
b11 +
#787970000000
1"
1(
#787980000000
0!
0"
b100 &
0'
0(
b100 ,
#787990000000
1!
b100 %
1'
b100 +
#788000000000
0!
0'
#788010000000
1!
b101 %
1'
b101 +
#788020000000
0!
0'
#788030000000
1!
b110 %
1'
b110 +
#788040000000
0!
0'
#788050000000
1!
b111 %
1'
b111 +
#788060000000
0!
0'
#788070000000
1!
0$
b1000 %
1'
0*
b1000 +
#788080000000
0!
0'
#788090000000
1!
b1001 %
1'
b1001 +
#788100000000
0!
0'
#788110000000
1!
b0 %
1'
b0 +
#788120000000
0!
0'
#788130000000
1!
1$
b1 %
1'
1*
b1 +
#788140000000
0!
0'
#788150000000
1!
b10 %
1'
b10 +
#788160000000
0!
0'
#788170000000
1!
b11 %
1'
b11 +
#788180000000
0!
0'
#788190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#788200000000
0!
0'
#788210000000
1!
b101 %
1'
b101 +
#788220000000
0!
0'
#788230000000
1!
0$
b110 %
1'
0*
b110 +
#788240000000
0!
0'
#788250000000
1!
b111 %
1'
b111 +
#788260000000
0!
0'
#788270000000
1!
b1000 %
1'
b1000 +
#788280000000
0!
0'
#788290000000
1!
b1001 %
1'
b1001 +
#788300000000
0!
0'
#788310000000
1!
b0 %
1'
b0 +
#788320000000
0!
0'
#788330000000
1!
1$
b1 %
1'
1*
b1 +
#788340000000
0!
0'
#788350000000
1!
b10 %
1'
b10 +
#788360000000
0!
0'
#788370000000
1!
b11 %
1'
b11 +
#788380000000
0!
0'
#788390000000
1!
b100 %
1'
b100 +
#788400000000
1"
1(
#788410000000
0!
0"
b100 &
0'
0(
b100 ,
#788420000000
1!
b101 %
1'
b101 +
#788430000000
0!
0'
#788440000000
1!
b110 %
1'
b110 +
#788450000000
0!
0'
#788460000000
1!
b111 %
1'
b111 +
#788470000000
0!
0'
#788480000000
1!
0$
b1000 %
1'
0*
b1000 +
#788490000000
0!
0'
#788500000000
1!
b1001 %
1'
b1001 +
#788510000000
0!
0'
#788520000000
1!
b0 %
1'
b0 +
#788530000000
0!
0'
#788540000000
1!
1$
b1 %
1'
1*
b1 +
#788550000000
0!
0'
#788560000000
1!
b10 %
1'
b10 +
#788570000000
0!
0'
#788580000000
1!
b11 %
1'
b11 +
#788590000000
0!
0'
#788600000000
1!
b100 %
1'
b100 +
#788610000000
0!
0'
#788620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#788630000000
0!
0'
#788640000000
1!
0$
b110 %
1'
0*
b110 +
#788650000000
0!
0'
#788660000000
1!
b111 %
1'
b111 +
#788670000000
0!
0'
#788680000000
1!
b1000 %
1'
b1000 +
#788690000000
0!
0'
#788700000000
1!
b1001 %
1'
b1001 +
#788710000000
0!
0'
#788720000000
1!
b0 %
1'
b0 +
#788730000000
0!
0'
#788740000000
1!
1$
b1 %
1'
1*
b1 +
#788750000000
0!
0'
#788760000000
1!
b10 %
1'
b10 +
#788770000000
0!
0'
#788780000000
1!
b11 %
1'
b11 +
#788790000000
0!
0'
#788800000000
1!
b100 %
1'
b100 +
#788810000000
0!
0'
#788820000000
1!
b101 %
1'
b101 +
#788830000000
1"
1(
#788840000000
0!
0"
b100 &
0'
0(
b100 ,
#788850000000
1!
b110 %
1'
b110 +
#788860000000
0!
0'
#788870000000
1!
b111 %
1'
b111 +
#788880000000
0!
0'
#788890000000
1!
0$
b1000 %
1'
0*
b1000 +
#788900000000
0!
0'
#788910000000
1!
b1001 %
1'
b1001 +
#788920000000
0!
0'
#788930000000
1!
b0 %
1'
b0 +
#788940000000
0!
0'
#788950000000
1!
1$
b1 %
1'
1*
b1 +
#788960000000
0!
0'
#788970000000
1!
b10 %
1'
b10 +
#788980000000
0!
0'
#788990000000
1!
b11 %
1'
b11 +
#789000000000
0!
0'
#789010000000
1!
b100 %
1'
b100 +
#789020000000
0!
0'
#789030000000
1!
b101 %
1'
b101 +
#789040000000
0!
0'
#789050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#789060000000
0!
0'
#789070000000
1!
b111 %
1'
b111 +
#789080000000
0!
0'
#789090000000
1!
b1000 %
1'
b1000 +
#789100000000
0!
0'
#789110000000
1!
b1001 %
1'
b1001 +
#789120000000
0!
0'
#789130000000
1!
b0 %
1'
b0 +
#789140000000
0!
0'
#789150000000
1!
1$
b1 %
1'
1*
b1 +
#789160000000
0!
0'
#789170000000
1!
b10 %
1'
b10 +
#789180000000
0!
0'
#789190000000
1!
b11 %
1'
b11 +
#789200000000
0!
0'
#789210000000
1!
b100 %
1'
b100 +
#789220000000
0!
0'
#789230000000
1!
b101 %
1'
b101 +
#789240000000
0!
0'
#789250000000
1!
0$
b110 %
1'
0*
b110 +
#789260000000
1"
1(
#789270000000
0!
0"
b100 &
0'
0(
b100 ,
#789280000000
1!
1$
b111 %
1'
1*
b111 +
#789290000000
0!
0'
#789300000000
1!
0$
b1000 %
1'
0*
b1000 +
#789310000000
0!
0'
#789320000000
1!
b1001 %
1'
b1001 +
#789330000000
0!
0'
#789340000000
1!
b0 %
1'
b0 +
#789350000000
0!
0'
#789360000000
1!
1$
b1 %
1'
1*
b1 +
#789370000000
0!
0'
#789380000000
1!
b10 %
1'
b10 +
#789390000000
0!
0'
#789400000000
1!
b11 %
1'
b11 +
#789410000000
0!
0'
#789420000000
1!
b100 %
1'
b100 +
#789430000000
0!
0'
#789440000000
1!
b101 %
1'
b101 +
#789450000000
0!
0'
#789460000000
1!
b110 %
1'
b110 +
#789470000000
0!
0'
#789480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#789490000000
0!
0'
#789500000000
1!
b1000 %
1'
b1000 +
#789510000000
0!
0'
#789520000000
1!
b1001 %
1'
b1001 +
#789530000000
0!
0'
#789540000000
1!
b0 %
1'
b0 +
#789550000000
0!
0'
#789560000000
1!
1$
b1 %
1'
1*
b1 +
#789570000000
0!
0'
#789580000000
1!
b10 %
1'
b10 +
#789590000000
0!
0'
#789600000000
1!
b11 %
1'
b11 +
#789610000000
0!
0'
#789620000000
1!
b100 %
1'
b100 +
#789630000000
0!
0'
#789640000000
1!
b101 %
1'
b101 +
#789650000000
0!
0'
#789660000000
1!
0$
b110 %
1'
0*
b110 +
#789670000000
0!
0'
#789680000000
1!
b111 %
1'
b111 +
#789690000000
1"
1(
#789700000000
0!
0"
b100 &
0'
0(
b100 ,
#789710000000
1!
b1000 %
1'
b1000 +
#789720000000
0!
0'
#789730000000
1!
b1001 %
1'
b1001 +
#789740000000
0!
0'
#789750000000
1!
b0 %
1'
b0 +
#789760000000
0!
0'
#789770000000
1!
1$
b1 %
1'
1*
b1 +
#789780000000
0!
0'
#789790000000
1!
b10 %
1'
b10 +
#789800000000
0!
0'
#789810000000
1!
b11 %
1'
b11 +
#789820000000
0!
0'
#789830000000
1!
b100 %
1'
b100 +
#789840000000
0!
0'
#789850000000
1!
b101 %
1'
b101 +
#789860000000
0!
0'
#789870000000
1!
b110 %
1'
b110 +
#789880000000
0!
0'
#789890000000
1!
b111 %
1'
b111 +
#789900000000
0!
0'
#789910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#789920000000
0!
0'
#789930000000
1!
b1001 %
1'
b1001 +
#789940000000
0!
0'
#789950000000
1!
b0 %
1'
b0 +
#789960000000
0!
0'
#789970000000
1!
1$
b1 %
1'
1*
b1 +
#789980000000
0!
0'
#789990000000
1!
b10 %
1'
b10 +
#790000000000
0!
0'
#790010000000
1!
b11 %
1'
b11 +
#790020000000
0!
0'
#790030000000
1!
b100 %
1'
b100 +
#790040000000
0!
0'
#790050000000
1!
b101 %
1'
b101 +
#790060000000
0!
0'
#790070000000
1!
0$
b110 %
1'
0*
b110 +
#790080000000
0!
0'
#790090000000
1!
b111 %
1'
b111 +
#790100000000
0!
0'
#790110000000
1!
b1000 %
1'
b1000 +
#790120000000
1"
1(
#790130000000
0!
0"
b100 &
0'
0(
b100 ,
#790140000000
1!
b1001 %
1'
b1001 +
#790150000000
0!
0'
#790160000000
1!
b0 %
1'
b0 +
#790170000000
0!
0'
#790180000000
1!
1$
b1 %
1'
1*
b1 +
#790190000000
0!
0'
#790200000000
1!
b10 %
1'
b10 +
#790210000000
0!
0'
#790220000000
1!
b11 %
1'
b11 +
#790230000000
0!
0'
#790240000000
1!
b100 %
1'
b100 +
#790250000000
0!
0'
#790260000000
1!
b101 %
1'
b101 +
#790270000000
0!
0'
#790280000000
1!
b110 %
1'
b110 +
#790290000000
0!
0'
#790300000000
1!
b111 %
1'
b111 +
#790310000000
0!
0'
#790320000000
1!
0$
b1000 %
1'
0*
b1000 +
#790330000000
0!
0'
#790340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#790350000000
0!
0'
#790360000000
1!
b0 %
1'
b0 +
#790370000000
0!
0'
#790380000000
1!
1$
b1 %
1'
1*
b1 +
#790390000000
0!
0'
#790400000000
1!
b10 %
1'
b10 +
#790410000000
0!
0'
#790420000000
1!
b11 %
1'
b11 +
#790430000000
0!
0'
#790440000000
1!
b100 %
1'
b100 +
#790450000000
0!
0'
#790460000000
1!
b101 %
1'
b101 +
#790470000000
0!
0'
#790480000000
1!
0$
b110 %
1'
0*
b110 +
#790490000000
0!
0'
#790500000000
1!
b111 %
1'
b111 +
#790510000000
0!
0'
#790520000000
1!
b1000 %
1'
b1000 +
#790530000000
0!
0'
#790540000000
1!
b1001 %
1'
b1001 +
#790550000000
1"
1(
#790560000000
0!
0"
b100 &
0'
0(
b100 ,
#790570000000
1!
b0 %
1'
b0 +
#790580000000
0!
0'
#790590000000
1!
1$
b1 %
1'
1*
b1 +
#790600000000
0!
0'
#790610000000
1!
b10 %
1'
b10 +
#790620000000
0!
0'
#790630000000
1!
b11 %
1'
b11 +
#790640000000
0!
0'
#790650000000
1!
b100 %
1'
b100 +
#790660000000
0!
0'
#790670000000
1!
b101 %
1'
b101 +
#790680000000
0!
0'
#790690000000
1!
b110 %
1'
b110 +
#790700000000
0!
0'
#790710000000
1!
b111 %
1'
b111 +
#790720000000
0!
0'
#790730000000
1!
0$
b1000 %
1'
0*
b1000 +
#790740000000
0!
0'
#790750000000
1!
b1001 %
1'
b1001 +
#790760000000
0!
0'
#790770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#790780000000
0!
0'
#790790000000
1!
1$
b1 %
1'
1*
b1 +
#790800000000
0!
0'
#790810000000
1!
b10 %
1'
b10 +
#790820000000
0!
0'
#790830000000
1!
b11 %
1'
b11 +
#790840000000
0!
0'
#790850000000
1!
b100 %
1'
b100 +
#790860000000
0!
0'
#790870000000
1!
b101 %
1'
b101 +
#790880000000
0!
0'
#790890000000
1!
0$
b110 %
1'
0*
b110 +
#790900000000
0!
0'
#790910000000
1!
b111 %
1'
b111 +
#790920000000
0!
0'
#790930000000
1!
b1000 %
1'
b1000 +
#790940000000
0!
0'
#790950000000
1!
b1001 %
1'
b1001 +
#790960000000
0!
0'
#790970000000
1!
b0 %
1'
b0 +
#790980000000
1"
1(
#790990000000
0!
0"
b100 &
0'
0(
b100 ,
#791000000000
1!
1$
b1 %
1'
1*
b1 +
#791010000000
0!
0'
#791020000000
1!
b10 %
1'
b10 +
#791030000000
0!
0'
#791040000000
1!
b11 %
1'
b11 +
#791050000000
0!
0'
#791060000000
1!
b100 %
1'
b100 +
#791070000000
0!
0'
#791080000000
1!
b101 %
1'
b101 +
#791090000000
0!
0'
#791100000000
1!
b110 %
1'
b110 +
#791110000000
0!
0'
#791120000000
1!
b111 %
1'
b111 +
#791130000000
0!
0'
#791140000000
1!
0$
b1000 %
1'
0*
b1000 +
#791150000000
0!
0'
#791160000000
1!
b1001 %
1'
b1001 +
#791170000000
0!
0'
#791180000000
1!
b0 %
1'
b0 +
#791190000000
0!
0'
#791200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#791210000000
0!
0'
#791220000000
1!
b10 %
1'
b10 +
#791230000000
0!
0'
#791240000000
1!
b11 %
1'
b11 +
#791250000000
0!
0'
#791260000000
1!
b100 %
1'
b100 +
#791270000000
0!
0'
#791280000000
1!
b101 %
1'
b101 +
#791290000000
0!
0'
#791300000000
1!
0$
b110 %
1'
0*
b110 +
#791310000000
0!
0'
#791320000000
1!
b111 %
1'
b111 +
#791330000000
0!
0'
#791340000000
1!
b1000 %
1'
b1000 +
#791350000000
0!
0'
#791360000000
1!
b1001 %
1'
b1001 +
#791370000000
0!
0'
#791380000000
1!
b0 %
1'
b0 +
#791390000000
0!
0'
#791400000000
1!
1$
b1 %
1'
1*
b1 +
#791410000000
1"
1(
#791420000000
0!
0"
b100 &
0'
0(
b100 ,
#791430000000
1!
b10 %
1'
b10 +
#791440000000
0!
0'
#791450000000
1!
b11 %
1'
b11 +
#791460000000
0!
0'
#791470000000
1!
b100 %
1'
b100 +
#791480000000
0!
0'
#791490000000
1!
b101 %
1'
b101 +
#791500000000
0!
0'
#791510000000
1!
b110 %
1'
b110 +
#791520000000
0!
0'
#791530000000
1!
b111 %
1'
b111 +
#791540000000
0!
0'
#791550000000
1!
0$
b1000 %
1'
0*
b1000 +
#791560000000
0!
0'
#791570000000
1!
b1001 %
1'
b1001 +
#791580000000
0!
0'
#791590000000
1!
b0 %
1'
b0 +
#791600000000
0!
0'
#791610000000
1!
1$
b1 %
1'
1*
b1 +
#791620000000
0!
0'
#791630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#791640000000
0!
0'
#791650000000
1!
b11 %
1'
b11 +
#791660000000
0!
0'
#791670000000
1!
b100 %
1'
b100 +
#791680000000
0!
0'
#791690000000
1!
b101 %
1'
b101 +
#791700000000
0!
0'
#791710000000
1!
0$
b110 %
1'
0*
b110 +
#791720000000
0!
0'
#791730000000
1!
b111 %
1'
b111 +
#791740000000
0!
0'
#791750000000
1!
b1000 %
1'
b1000 +
#791760000000
0!
0'
#791770000000
1!
b1001 %
1'
b1001 +
#791780000000
0!
0'
#791790000000
1!
b0 %
1'
b0 +
#791800000000
0!
0'
#791810000000
1!
1$
b1 %
1'
1*
b1 +
#791820000000
0!
0'
#791830000000
1!
b10 %
1'
b10 +
#791840000000
1"
1(
#791850000000
0!
0"
b100 &
0'
0(
b100 ,
#791860000000
1!
b11 %
1'
b11 +
#791870000000
0!
0'
#791880000000
1!
b100 %
1'
b100 +
#791890000000
0!
0'
#791900000000
1!
b101 %
1'
b101 +
#791910000000
0!
0'
#791920000000
1!
b110 %
1'
b110 +
#791930000000
0!
0'
#791940000000
1!
b111 %
1'
b111 +
#791950000000
0!
0'
#791960000000
1!
0$
b1000 %
1'
0*
b1000 +
#791970000000
0!
0'
#791980000000
1!
b1001 %
1'
b1001 +
#791990000000
0!
0'
#792000000000
1!
b0 %
1'
b0 +
#792010000000
0!
0'
#792020000000
1!
1$
b1 %
1'
1*
b1 +
#792030000000
0!
0'
#792040000000
1!
b10 %
1'
b10 +
#792050000000
0!
0'
#792060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#792070000000
0!
0'
#792080000000
1!
b100 %
1'
b100 +
#792090000000
0!
0'
#792100000000
1!
b101 %
1'
b101 +
#792110000000
0!
0'
#792120000000
1!
0$
b110 %
1'
0*
b110 +
#792130000000
0!
0'
#792140000000
1!
b111 %
1'
b111 +
#792150000000
0!
0'
#792160000000
1!
b1000 %
1'
b1000 +
#792170000000
0!
0'
#792180000000
1!
b1001 %
1'
b1001 +
#792190000000
0!
0'
#792200000000
1!
b0 %
1'
b0 +
#792210000000
0!
0'
#792220000000
1!
1$
b1 %
1'
1*
b1 +
#792230000000
0!
0'
#792240000000
1!
b10 %
1'
b10 +
#792250000000
0!
0'
#792260000000
1!
b11 %
1'
b11 +
#792270000000
1"
1(
#792280000000
0!
0"
b100 &
0'
0(
b100 ,
#792290000000
1!
b100 %
1'
b100 +
#792300000000
0!
0'
#792310000000
1!
b101 %
1'
b101 +
#792320000000
0!
0'
#792330000000
1!
b110 %
1'
b110 +
#792340000000
0!
0'
#792350000000
1!
b111 %
1'
b111 +
#792360000000
0!
0'
#792370000000
1!
0$
b1000 %
1'
0*
b1000 +
#792380000000
0!
0'
#792390000000
1!
b1001 %
1'
b1001 +
#792400000000
0!
0'
#792410000000
1!
b0 %
1'
b0 +
#792420000000
0!
0'
#792430000000
1!
1$
b1 %
1'
1*
b1 +
#792440000000
0!
0'
#792450000000
1!
b10 %
1'
b10 +
#792460000000
0!
0'
#792470000000
1!
b11 %
1'
b11 +
#792480000000
0!
0'
#792490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#792500000000
0!
0'
#792510000000
1!
b101 %
1'
b101 +
#792520000000
0!
0'
#792530000000
1!
0$
b110 %
1'
0*
b110 +
#792540000000
0!
0'
#792550000000
1!
b111 %
1'
b111 +
#792560000000
0!
0'
#792570000000
1!
b1000 %
1'
b1000 +
#792580000000
0!
0'
#792590000000
1!
b1001 %
1'
b1001 +
#792600000000
0!
0'
#792610000000
1!
b0 %
1'
b0 +
#792620000000
0!
0'
#792630000000
1!
1$
b1 %
1'
1*
b1 +
#792640000000
0!
0'
#792650000000
1!
b10 %
1'
b10 +
#792660000000
0!
0'
#792670000000
1!
b11 %
1'
b11 +
#792680000000
0!
0'
#792690000000
1!
b100 %
1'
b100 +
#792700000000
1"
1(
#792710000000
0!
0"
b100 &
0'
0(
b100 ,
#792720000000
1!
b101 %
1'
b101 +
#792730000000
0!
0'
#792740000000
1!
b110 %
1'
b110 +
#792750000000
0!
0'
#792760000000
1!
b111 %
1'
b111 +
#792770000000
0!
0'
#792780000000
1!
0$
b1000 %
1'
0*
b1000 +
#792790000000
0!
0'
#792800000000
1!
b1001 %
1'
b1001 +
#792810000000
0!
0'
#792820000000
1!
b0 %
1'
b0 +
#792830000000
0!
0'
#792840000000
1!
1$
b1 %
1'
1*
b1 +
#792850000000
0!
0'
#792860000000
1!
b10 %
1'
b10 +
#792870000000
0!
0'
#792880000000
1!
b11 %
1'
b11 +
#792890000000
0!
0'
#792900000000
1!
b100 %
1'
b100 +
#792910000000
0!
0'
#792920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#792930000000
0!
0'
#792940000000
1!
0$
b110 %
1'
0*
b110 +
#792950000000
0!
0'
#792960000000
1!
b111 %
1'
b111 +
#792970000000
0!
0'
#792980000000
1!
b1000 %
1'
b1000 +
#792990000000
0!
0'
#793000000000
1!
b1001 %
1'
b1001 +
#793010000000
0!
0'
#793020000000
1!
b0 %
1'
b0 +
#793030000000
0!
0'
#793040000000
1!
1$
b1 %
1'
1*
b1 +
#793050000000
0!
0'
#793060000000
1!
b10 %
1'
b10 +
#793070000000
0!
0'
#793080000000
1!
b11 %
1'
b11 +
#793090000000
0!
0'
#793100000000
1!
b100 %
1'
b100 +
#793110000000
0!
0'
#793120000000
1!
b101 %
1'
b101 +
#793130000000
1"
1(
#793140000000
0!
0"
b100 &
0'
0(
b100 ,
#793150000000
1!
b110 %
1'
b110 +
#793160000000
0!
0'
#793170000000
1!
b111 %
1'
b111 +
#793180000000
0!
0'
#793190000000
1!
0$
b1000 %
1'
0*
b1000 +
#793200000000
0!
0'
#793210000000
1!
b1001 %
1'
b1001 +
#793220000000
0!
0'
#793230000000
1!
b0 %
1'
b0 +
#793240000000
0!
0'
#793250000000
1!
1$
b1 %
1'
1*
b1 +
#793260000000
0!
0'
#793270000000
1!
b10 %
1'
b10 +
#793280000000
0!
0'
#793290000000
1!
b11 %
1'
b11 +
#793300000000
0!
0'
#793310000000
1!
b100 %
1'
b100 +
#793320000000
0!
0'
#793330000000
1!
b101 %
1'
b101 +
#793340000000
0!
0'
#793350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#793360000000
0!
0'
#793370000000
1!
b111 %
1'
b111 +
#793380000000
0!
0'
#793390000000
1!
b1000 %
1'
b1000 +
#793400000000
0!
0'
#793410000000
1!
b1001 %
1'
b1001 +
#793420000000
0!
0'
#793430000000
1!
b0 %
1'
b0 +
#793440000000
0!
0'
#793450000000
1!
1$
b1 %
1'
1*
b1 +
#793460000000
0!
0'
#793470000000
1!
b10 %
1'
b10 +
#793480000000
0!
0'
#793490000000
1!
b11 %
1'
b11 +
#793500000000
0!
0'
#793510000000
1!
b100 %
1'
b100 +
#793520000000
0!
0'
#793530000000
1!
b101 %
1'
b101 +
#793540000000
0!
0'
#793550000000
1!
0$
b110 %
1'
0*
b110 +
#793560000000
1"
1(
#793570000000
0!
0"
b100 &
0'
0(
b100 ,
#793580000000
1!
1$
b111 %
1'
1*
b111 +
#793590000000
0!
0'
#793600000000
1!
0$
b1000 %
1'
0*
b1000 +
#793610000000
0!
0'
#793620000000
1!
b1001 %
1'
b1001 +
#793630000000
0!
0'
#793640000000
1!
b0 %
1'
b0 +
#793650000000
0!
0'
#793660000000
1!
1$
b1 %
1'
1*
b1 +
#793670000000
0!
0'
#793680000000
1!
b10 %
1'
b10 +
#793690000000
0!
0'
#793700000000
1!
b11 %
1'
b11 +
#793710000000
0!
0'
#793720000000
1!
b100 %
1'
b100 +
#793730000000
0!
0'
#793740000000
1!
b101 %
1'
b101 +
#793750000000
0!
0'
#793760000000
1!
b110 %
1'
b110 +
#793770000000
0!
0'
#793780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#793790000000
0!
0'
#793800000000
1!
b1000 %
1'
b1000 +
#793810000000
0!
0'
#793820000000
1!
b1001 %
1'
b1001 +
#793830000000
0!
0'
#793840000000
1!
b0 %
1'
b0 +
#793850000000
0!
0'
#793860000000
1!
1$
b1 %
1'
1*
b1 +
#793870000000
0!
0'
#793880000000
1!
b10 %
1'
b10 +
#793890000000
0!
0'
#793900000000
1!
b11 %
1'
b11 +
#793910000000
0!
0'
#793920000000
1!
b100 %
1'
b100 +
#793930000000
0!
0'
#793940000000
1!
b101 %
1'
b101 +
#793950000000
0!
0'
#793960000000
1!
0$
b110 %
1'
0*
b110 +
#793970000000
0!
0'
#793980000000
1!
b111 %
1'
b111 +
#793990000000
1"
1(
#794000000000
0!
0"
b100 &
0'
0(
b100 ,
#794010000000
1!
b1000 %
1'
b1000 +
#794020000000
0!
0'
#794030000000
1!
b1001 %
1'
b1001 +
#794040000000
0!
0'
#794050000000
1!
b0 %
1'
b0 +
#794060000000
0!
0'
#794070000000
1!
1$
b1 %
1'
1*
b1 +
#794080000000
0!
0'
#794090000000
1!
b10 %
1'
b10 +
#794100000000
0!
0'
#794110000000
1!
b11 %
1'
b11 +
#794120000000
0!
0'
#794130000000
1!
b100 %
1'
b100 +
#794140000000
0!
0'
#794150000000
1!
b101 %
1'
b101 +
#794160000000
0!
0'
#794170000000
1!
b110 %
1'
b110 +
#794180000000
0!
0'
#794190000000
1!
b111 %
1'
b111 +
#794200000000
0!
0'
#794210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#794220000000
0!
0'
#794230000000
1!
b1001 %
1'
b1001 +
#794240000000
0!
0'
#794250000000
1!
b0 %
1'
b0 +
#794260000000
0!
0'
#794270000000
1!
1$
b1 %
1'
1*
b1 +
#794280000000
0!
0'
#794290000000
1!
b10 %
1'
b10 +
#794300000000
0!
0'
#794310000000
1!
b11 %
1'
b11 +
#794320000000
0!
0'
#794330000000
1!
b100 %
1'
b100 +
#794340000000
0!
0'
#794350000000
1!
b101 %
1'
b101 +
#794360000000
0!
0'
#794370000000
1!
0$
b110 %
1'
0*
b110 +
#794380000000
0!
0'
#794390000000
1!
b111 %
1'
b111 +
#794400000000
0!
0'
#794410000000
1!
b1000 %
1'
b1000 +
#794420000000
1"
1(
#794430000000
0!
0"
b100 &
0'
0(
b100 ,
#794440000000
1!
b1001 %
1'
b1001 +
#794450000000
0!
0'
#794460000000
1!
b0 %
1'
b0 +
#794470000000
0!
0'
#794480000000
1!
1$
b1 %
1'
1*
b1 +
#794490000000
0!
0'
#794500000000
1!
b10 %
1'
b10 +
#794510000000
0!
0'
#794520000000
1!
b11 %
1'
b11 +
#794530000000
0!
0'
#794540000000
1!
b100 %
1'
b100 +
#794550000000
0!
0'
#794560000000
1!
b101 %
1'
b101 +
#794570000000
0!
0'
#794580000000
1!
b110 %
1'
b110 +
#794590000000
0!
0'
#794600000000
1!
b111 %
1'
b111 +
#794610000000
0!
0'
#794620000000
1!
0$
b1000 %
1'
0*
b1000 +
#794630000000
0!
0'
#794640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#794650000000
0!
0'
#794660000000
1!
b0 %
1'
b0 +
#794670000000
0!
0'
#794680000000
1!
1$
b1 %
1'
1*
b1 +
#794690000000
0!
0'
#794700000000
1!
b10 %
1'
b10 +
#794710000000
0!
0'
#794720000000
1!
b11 %
1'
b11 +
#794730000000
0!
0'
#794740000000
1!
b100 %
1'
b100 +
#794750000000
0!
0'
#794760000000
1!
b101 %
1'
b101 +
#794770000000
0!
0'
#794780000000
1!
0$
b110 %
1'
0*
b110 +
#794790000000
0!
0'
#794800000000
1!
b111 %
1'
b111 +
#794810000000
0!
0'
#794820000000
1!
b1000 %
1'
b1000 +
#794830000000
0!
0'
#794840000000
1!
b1001 %
1'
b1001 +
#794850000000
1"
1(
#794860000000
0!
0"
b100 &
0'
0(
b100 ,
#794870000000
1!
b0 %
1'
b0 +
#794880000000
0!
0'
#794890000000
1!
1$
b1 %
1'
1*
b1 +
#794900000000
0!
0'
#794910000000
1!
b10 %
1'
b10 +
#794920000000
0!
0'
#794930000000
1!
b11 %
1'
b11 +
#794940000000
0!
0'
#794950000000
1!
b100 %
1'
b100 +
#794960000000
0!
0'
#794970000000
1!
b101 %
1'
b101 +
#794980000000
0!
0'
#794990000000
1!
b110 %
1'
b110 +
#795000000000
0!
0'
#795010000000
1!
b111 %
1'
b111 +
#795020000000
0!
0'
#795030000000
1!
0$
b1000 %
1'
0*
b1000 +
#795040000000
0!
0'
#795050000000
1!
b1001 %
1'
b1001 +
#795060000000
0!
0'
#795070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#795080000000
0!
0'
#795090000000
1!
1$
b1 %
1'
1*
b1 +
#795100000000
0!
0'
#795110000000
1!
b10 %
1'
b10 +
#795120000000
0!
0'
#795130000000
1!
b11 %
1'
b11 +
#795140000000
0!
0'
#795150000000
1!
b100 %
1'
b100 +
#795160000000
0!
0'
#795170000000
1!
b101 %
1'
b101 +
#795180000000
0!
0'
#795190000000
1!
0$
b110 %
1'
0*
b110 +
#795200000000
0!
0'
#795210000000
1!
b111 %
1'
b111 +
#795220000000
0!
0'
#795230000000
1!
b1000 %
1'
b1000 +
#795240000000
0!
0'
#795250000000
1!
b1001 %
1'
b1001 +
#795260000000
0!
0'
#795270000000
1!
b0 %
1'
b0 +
#795280000000
1"
1(
#795290000000
0!
0"
b100 &
0'
0(
b100 ,
#795300000000
1!
1$
b1 %
1'
1*
b1 +
#795310000000
0!
0'
#795320000000
1!
b10 %
1'
b10 +
#795330000000
0!
0'
#795340000000
1!
b11 %
1'
b11 +
#795350000000
0!
0'
#795360000000
1!
b100 %
1'
b100 +
#795370000000
0!
0'
#795380000000
1!
b101 %
1'
b101 +
#795390000000
0!
0'
#795400000000
1!
b110 %
1'
b110 +
#795410000000
0!
0'
#795420000000
1!
b111 %
1'
b111 +
#795430000000
0!
0'
#795440000000
1!
0$
b1000 %
1'
0*
b1000 +
#795450000000
0!
0'
#795460000000
1!
b1001 %
1'
b1001 +
#795470000000
0!
0'
#795480000000
1!
b0 %
1'
b0 +
#795490000000
0!
0'
#795500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#795510000000
0!
0'
#795520000000
1!
b10 %
1'
b10 +
#795530000000
0!
0'
#795540000000
1!
b11 %
1'
b11 +
#795550000000
0!
0'
#795560000000
1!
b100 %
1'
b100 +
#795570000000
0!
0'
#795580000000
1!
b101 %
1'
b101 +
#795590000000
0!
0'
#795600000000
1!
0$
b110 %
1'
0*
b110 +
#795610000000
0!
0'
#795620000000
1!
b111 %
1'
b111 +
#795630000000
0!
0'
#795640000000
1!
b1000 %
1'
b1000 +
#795650000000
0!
0'
#795660000000
1!
b1001 %
1'
b1001 +
#795670000000
0!
0'
#795680000000
1!
b0 %
1'
b0 +
#795690000000
0!
0'
#795700000000
1!
1$
b1 %
1'
1*
b1 +
#795710000000
1"
1(
#795720000000
0!
0"
b100 &
0'
0(
b100 ,
#795730000000
1!
b10 %
1'
b10 +
#795740000000
0!
0'
#795750000000
1!
b11 %
1'
b11 +
#795760000000
0!
0'
#795770000000
1!
b100 %
1'
b100 +
#795780000000
0!
0'
#795790000000
1!
b101 %
1'
b101 +
#795800000000
0!
0'
#795810000000
1!
b110 %
1'
b110 +
#795820000000
0!
0'
#795830000000
1!
b111 %
1'
b111 +
#795840000000
0!
0'
#795850000000
1!
0$
b1000 %
1'
0*
b1000 +
#795860000000
0!
0'
#795870000000
1!
b1001 %
1'
b1001 +
#795880000000
0!
0'
#795890000000
1!
b0 %
1'
b0 +
#795900000000
0!
0'
#795910000000
1!
1$
b1 %
1'
1*
b1 +
#795920000000
0!
0'
#795930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#795940000000
0!
0'
#795950000000
1!
b11 %
1'
b11 +
#795960000000
0!
0'
#795970000000
1!
b100 %
1'
b100 +
#795980000000
0!
0'
#795990000000
1!
b101 %
1'
b101 +
#796000000000
0!
0'
#796010000000
1!
0$
b110 %
1'
0*
b110 +
#796020000000
0!
0'
#796030000000
1!
b111 %
1'
b111 +
#796040000000
0!
0'
#796050000000
1!
b1000 %
1'
b1000 +
#796060000000
0!
0'
#796070000000
1!
b1001 %
1'
b1001 +
#796080000000
0!
0'
#796090000000
1!
b0 %
1'
b0 +
#796100000000
0!
0'
#796110000000
1!
1$
b1 %
1'
1*
b1 +
#796120000000
0!
0'
#796130000000
1!
b10 %
1'
b10 +
#796140000000
1"
1(
#796150000000
0!
0"
b100 &
0'
0(
b100 ,
#796160000000
1!
b11 %
1'
b11 +
#796170000000
0!
0'
#796180000000
1!
b100 %
1'
b100 +
#796190000000
0!
0'
#796200000000
1!
b101 %
1'
b101 +
#796210000000
0!
0'
#796220000000
1!
b110 %
1'
b110 +
#796230000000
0!
0'
#796240000000
1!
b111 %
1'
b111 +
#796250000000
0!
0'
#796260000000
1!
0$
b1000 %
1'
0*
b1000 +
#796270000000
0!
0'
#796280000000
1!
b1001 %
1'
b1001 +
#796290000000
0!
0'
#796300000000
1!
b0 %
1'
b0 +
#796310000000
0!
0'
#796320000000
1!
1$
b1 %
1'
1*
b1 +
#796330000000
0!
0'
#796340000000
1!
b10 %
1'
b10 +
#796350000000
0!
0'
#796360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#796370000000
0!
0'
#796380000000
1!
b100 %
1'
b100 +
#796390000000
0!
0'
#796400000000
1!
b101 %
1'
b101 +
#796410000000
0!
0'
#796420000000
1!
0$
b110 %
1'
0*
b110 +
#796430000000
0!
0'
#796440000000
1!
b111 %
1'
b111 +
#796450000000
0!
0'
#796460000000
1!
b1000 %
1'
b1000 +
#796470000000
0!
0'
#796480000000
1!
b1001 %
1'
b1001 +
#796490000000
0!
0'
#796500000000
1!
b0 %
1'
b0 +
#796510000000
0!
0'
#796520000000
1!
1$
b1 %
1'
1*
b1 +
#796530000000
0!
0'
#796540000000
1!
b10 %
1'
b10 +
#796550000000
0!
0'
#796560000000
1!
b11 %
1'
b11 +
#796570000000
1"
1(
#796580000000
0!
0"
b100 &
0'
0(
b100 ,
#796590000000
1!
b100 %
1'
b100 +
#796600000000
0!
0'
#796610000000
1!
b101 %
1'
b101 +
#796620000000
0!
0'
#796630000000
1!
b110 %
1'
b110 +
#796640000000
0!
0'
#796650000000
1!
b111 %
1'
b111 +
#796660000000
0!
0'
#796670000000
1!
0$
b1000 %
1'
0*
b1000 +
#796680000000
0!
0'
#796690000000
1!
b1001 %
1'
b1001 +
#796700000000
0!
0'
#796710000000
1!
b0 %
1'
b0 +
#796720000000
0!
0'
#796730000000
1!
1$
b1 %
1'
1*
b1 +
#796740000000
0!
0'
#796750000000
1!
b10 %
1'
b10 +
#796760000000
0!
0'
#796770000000
1!
b11 %
1'
b11 +
#796780000000
0!
0'
#796790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#796800000000
0!
0'
#796810000000
1!
b101 %
1'
b101 +
#796820000000
0!
0'
#796830000000
1!
0$
b110 %
1'
0*
b110 +
#796840000000
0!
0'
#796850000000
1!
b111 %
1'
b111 +
#796860000000
0!
0'
#796870000000
1!
b1000 %
1'
b1000 +
#796880000000
0!
0'
#796890000000
1!
b1001 %
1'
b1001 +
#796900000000
0!
0'
#796910000000
1!
b0 %
1'
b0 +
#796920000000
0!
0'
#796930000000
1!
1$
b1 %
1'
1*
b1 +
#796940000000
0!
0'
#796950000000
1!
b10 %
1'
b10 +
#796960000000
0!
0'
#796970000000
1!
b11 %
1'
b11 +
#796980000000
0!
0'
#796990000000
1!
b100 %
1'
b100 +
#797000000000
1"
1(
#797010000000
0!
0"
b100 &
0'
0(
b100 ,
#797020000000
1!
b101 %
1'
b101 +
#797030000000
0!
0'
#797040000000
1!
b110 %
1'
b110 +
#797050000000
0!
0'
#797060000000
1!
b111 %
1'
b111 +
#797070000000
0!
0'
#797080000000
1!
0$
b1000 %
1'
0*
b1000 +
#797090000000
0!
0'
#797100000000
1!
b1001 %
1'
b1001 +
#797110000000
0!
0'
#797120000000
1!
b0 %
1'
b0 +
#797130000000
0!
0'
#797140000000
1!
1$
b1 %
1'
1*
b1 +
#797150000000
0!
0'
#797160000000
1!
b10 %
1'
b10 +
#797170000000
0!
0'
#797180000000
1!
b11 %
1'
b11 +
#797190000000
0!
0'
#797200000000
1!
b100 %
1'
b100 +
#797210000000
0!
0'
#797220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#797230000000
0!
0'
#797240000000
1!
0$
b110 %
1'
0*
b110 +
#797250000000
0!
0'
#797260000000
1!
b111 %
1'
b111 +
#797270000000
0!
0'
#797280000000
1!
b1000 %
1'
b1000 +
#797290000000
0!
0'
#797300000000
1!
b1001 %
1'
b1001 +
#797310000000
0!
0'
#797320000000
1!
b0 %
1'
b0 +
#797330000000
0!
0'
#797340000000
1!
1$
b1 %
1'
1*
b1 +
#797350000000
0!
0'
#797360000000
1!
b10 %
1'
b10 +
#797370000000
0!
0'
#797380000000
1!
b11 %
1'
b11 +
#797390000000
0!
0'
#797400000000
1!
b100 %
1'
b100 +
#797410000000
0!
0'
#797420000000
1!
b101 %
1'
b101 +
#797430000000
1"
1(
#797440000000
0!
0"
b100 &
0'
0(
b100 ,
#797450000000
1!
b110 %
1'
b110 +
#797460000000
0!
0'
#797470000000
1!
b111 %
1'
b111 +
#797480000000
0!
0'
#797490000000
1!
0$
b1000 %
1'
0*
b1000 +
#797500000000
0!
0'
#797510000000
1!
b1001 %
1'
b1001 +
#797520000000
0!
0'
#797530000000
1!
b0 %
1'
b0 +
#797540000000
0!
0'
#797550000000
1!
1$
b1 %
1'
1*
b1 +
#797560000000
0!
0'
#797570000000
1!
b10 %
1'
b10 +
#797580000000
0!
0'
#797590000000
1!
b11 %
1'
b11 +
#797600000000
0!
0'
#797610000000
1!
b100 %
1'
b100 +
#797620000000
0!
0'
#797630000000
1!
b101 %
1'
b101 +
#797640000000
0!
0'
#797650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#797660000000
0!
0'
#797670000000
1!
b111 %
1'
b111 +
#797680000000
0!
0'
#797690000000
1!
b1000 %
1'
b1000 +
#797700000000
0!
0'
#797710000000
1!
b1001 %
1'
b1001 +
#797720000000
0!
0'
#797730000000
1!
b0 %
1'
b0 +
#797740000000
0!
0'
#797750000000
1!
1$
b1 %
1'
1*
b1 +
#797760000000
0!
0'
#797770000000
1!
b10 %
1'
b10 +
#797780000000
0!
0'
#797790000000
1!
b11 %
1'
b11 +
#797800000000
0!
0'
#797810000000
1!
b100 %
1'
b100 +
#797820000000
0!
0'
#797830000000
1!
b101 %
1'
b101 +
#797840000000
0!
0'
#797850000000
1!
0$
b110 %
1'
0*
b110 +
#797860000000
1"
1(
#797870000000
0!
0"
b100 &
0'
0(
b100 ,
#797880000000
1!
1$
b111 %
1'
1*
b111 +
#797890000000
0!
0'
#797900000000
1!
0$
b1000 %
1'
0*
b1000 +
#797910000000
0!
0'
#797920000000
1!
b1001 %
1'
b1001 +
#797930000000
0!
0'
#797940000000
1!
b0 %
1'
b0 +
#797950000000
0!
0'
#797960000000
1!
1$
b1 %
1'
1*
b1 +
#797970000000
0!
0'
#797980000000
1!
b10 %
1'
b10 +
#797990000000
0!
0'
#798000000000
1!
b11 %
1'
b11 +
#798010000000
0!
0'
#798020000000
1!
b100 %
1'
b100 +
#798030000000
0!
0'
#798040000000
1!
b101 %
1'
b101 +
#798050000000
0!
0'
#798060000000
1!
b110 %
1'
b110 +
#798070000000
0!
0'
#798080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#798090000000
0!
0'
#798100000000
1!
b1000 %
1'
b1000 +
#798110000000
0!
0'
#798120000000
1!
b1001 %
1'
b1001 +
#798130000000
0!
0'
#798140000000
1!
b0 %
1'
b0 +
#798150000000
0!
0'
#798160000000
1!
1$
b1 %
1'
1*
b1 +
#798170000000
0!
0'
#798180000000
1!
b10 %
1'
b10 +
#798190000000
0!
0'
#798200000000
1!
b11 %
1'
b11 +
#798210000000
0!
0'
#798220000000
1!
b100 %
1'
b100 +
#798230000000
0!
0'
#798240000000
1!
b101 %
1'
b101 +
#798250000000
0!
0'
#798260000000
1!
0$
b110 %
1'
0*
b110 +
#798270000000
0!
0'
#798280000000
1!
b111 %
1'
b111 +
#798290000000
1"
1(
#798300000000
0!
0"
b100 &
0'
0(
b100 ,
#798310000000
1!
b1000 %
1'
b1000 +
#798320000000
0!
0'
#798330000000
1!
b1001 %
1'
b1001 +
#798340000000
0!
0'
#798350000000
1!
b0 %
1'
b0 +
#798360000000
0!
0'
#798370000000
1!
1$
b1 %
1'
1*
b1 +
#798380000000
0!
0'
#798390000000
1!
b10 %
1'
b10 +
#798400000000
0!
0'
#798410000000
1!
b11 %
1'
b11 +
#798420000000
0!
0'
#798430000000
1!
b100 %
1'
b100 +
#798440000000
0!
0'
#798450000000
1!
b101 %
1'
b101 +
#798460000000
0!
0'
#798470000000
1!
b110 %
1'
b110 +
#798480000000
0!
0'
#798490000000
1!
b111 %
1'
b111 +
#798500000000
0!
0'
#798510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#798520000000
0!
0'
#798530000000
1!
b1001 %
1'
b1001 +
#798540000000
0!
0'
#798550000000
1!
b0 %
1'
b0 +
#798560000000
0!
0'
#798570000000
1!
1$
b1 %
1'
1*
b1 +
#798580000000
0!
0'
#798590000000
1!
b10 %
1'
b10 +
#798600000000
0!
0'
#798610000000
1!
b11 %
1'
b11 +
#798620000000
0!
0'
#798630000000
1!
b100 %
1'
b100 +
#798640000000
0!
0'
#798650000000
1!
b101 %
1'
b101 +
#798660000000
0!
0'
#798670000000
1!
0$
b110 %
1'
0*
b110 +
#798680000000
0!
0'
#798690000000
1!
b111 %
1'
b111 +
#798700000000
0!
0'
#798710000000
1!
b1000 %
1'
b1000 +
#798720000000
1"
1(
#798730000000
0!
0"
b100 &
0'
0(
b100 ,
#798740000000
1!
b1001 %
1'
b1001 +
#798750000000
0!
0'
#798760000000
1!
b0 %
1'
b0 +
#798770000000
0!
0'
#798780000000
1!
1$
b1 %
1'
1*
b1 +
#798790000000
0!
0'
#798800000000
1!
b10 %
1'
b10 +
#798810000000
0!
0'
#798820000000
1!
b11 %
1'
b11 +
#798830000000
0!
0'
#798840000000
1!
b100 %
1'
b100 +
#798850000000
0!
0'
#798860000000
1!
b101 %
1'
b101 +
#798870000000
0!
0'
#798880000000
1!
b110 %
1'
b110 +
#798890000000
0!
0'
#798900000000
1!
b111 %
1'
b111 +
#798910000000
0!
0'
#798920000000
1!
0$
b1000 %
1'
0*
b1000 +
#798930000000
0!
0'
#798940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#798950000000
0!
0'
#798960000000
1!
b0 %
1'
b0 +
#798970000000
0!
0'
#798980000000
1!
1$
b1 %
1'
1*
b1 +
#798990000000
0!
0'
#799000000000
1!
b10 %
1'
b10 +
#799010000000
0!
0'
#799020000000
1!
b11 %
1'
b11 +
#799030000000
0!
0'
#799040000000
1!
b100 %
1'
b100 +
#799050000000
0!
0'
#799060000000
1!
b101 %
1'
b101 +
#799070000000
0!
0'
#799080000000
1!
0$
b110 %
1'
0*
b110 +
#799090000000
0!
0'
#799100000000
1!
b111 %
1'
b111 +
#799110000000
0!
0'
#799120000000
1!
b1000 %
1'
b1000 +
#799130000000
0!
0'
#799140000000
1!
b1001 %
1'
b1001 +
#799150000000
1"
1(
#799160000000
0!
0"
b100 &
0'
0(
b100 ,
#799170000000
1!
b0 %
1'
b0 +
#799180000000
0!
0'
#799190000000
1!
1$
b1 %
1'
1*
b1 +
#799200000000
0!
0'
#799210000000
1!
b10 %
1'
b10 +
#799220000000
0!
0'
#799230000000
1!
b11 %
1'
b11 +
#799240000000
0!
0'
#799250000000
1!
b100 %
1'
b100 +
#799260000000
0!
0'
#799270000000
1!
b101 %
1'
b101 +
#799280000000
0!
0'
#799290000000
1!
b110 %
1'
b110 +
#799300000000
0!
0'
#799310000000
1!
b111 %
1'
b111 +
#799320000000
0!
0'
#799330000000
1!
0$
b1000 %
1'
0*
b1000 +
#799340000000
0!
0'
#799350000000
1!
b1001 %
1'
b1001 +
#799360000000
0!
0'
#799370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#799380000000
0!
0'
#799390000000
1!
1$
b1 %
1'
1*
b1 +
#799400000000
0!
0'
#799410000000
1!
b10 %
1'
b10 +
#799420000000
0!
0'
#799430000000
1!
b11 %
1'
b11 +
#799440000000
0!
0'
#799450000000
1!
b100 %
1'
b100 +
#799460000000
0!
0'
#799470000000
1!
b101 %
1'
b101 +
#799480000000
0!
0'
#799490000000
1!
0$
b110 %
1'
0*
b110 +
#799500000000
0!
0'
#799510000000
1!
b111 %
1'
b111 +
#799520000000
0!
0'
#799530000000
1!
b1000 %
1'
b1000 +
#799540000000
0!
0'
#799550000000
1!
b1001 %
1'
b1001 +
#799560000000
0!
0'
#799570000000
1!
b0 %
1'
b0 +
#799580000000
1"
1(
#799590000000
0!
0"
b100 &
0'
0(
b100 ,
#799600000000
1!
1$
b1 %
1'
1*
b1 +
#799610000000
0!
0'
#799620000000
1!
b10 %
1'
b10 +
#799630000000
0!
0'
#799640000000
1!
b11 %
1'
b11 +
#799650000000
0!
0'
#799660000000
1!
b100 %
1'
b100 +
#799670000000
0!
0'
#799680000000
1!
b101 %
1'
b101 +
#799690000000
0!
0'
#799700000000
1!
b110 %
1'
b110 +
#799710000000
0!
0'
#799720000000
1!
b111 %
1'
b111 +
#799730000000
0!
0'
#799740000000
1!
0$
b1000 %
1'
0*
b1000 +
#799750000000
0!
0'
#799760000000
1!
b1001 %
1'
b1001 +
#799770000000
0!
0'
#799780000000
1!
b0 %
1'
b0 +
#799790000000
0!
0'
#799800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#799810000000
0!
0'
#799820000000
1!
b10 %
1'
b10 +
#799830000000
0!
0'
#799840000000
1!
b11 %
1'
b11 +
#799850000000
0!
0'
#799860000000
1!
b100 %
1'
b100 +
#799870000000
0!
0'
#799880000000
1!
b101 %
1'
b101 +
#799890000000
0!
0'
#799900000000
1!
0$
b110 %
1'
0*
b110 +
#799910000000
0!
0'
#799920000000
1!
b111 %
1'
b111 +
#799930000000
0!
0'
#799940000000
1!
b1000 %
1'
b1000 +
#799950000000
0!
0'
#799960000000
1!
b1001 %
1'
b1001 +
#799970000000
0!
0'
#799980000000
1!
b0 %
1'
b0 +
#799990000000
0!
0'
#800000000000
1!
1$
b1 %
1'
1*
b1 +
#800010000000
1"
1(
#800020000000
0!
0"
b100 &
0'
0(
b100 ,
#800030000000
1!
b10 %
1'
b10 +
#800040000000
0!
0'
#800050000000
1!
b11 %
1'
b11 +
#800060000000
0!
0'
#800070000000
1!
b100 %
1'
b100 +
#800080000000
0!
0'
#800090000000
1!
b101 %
1'
b101 +
#800100000000
0!
0'
#800110000000
1!
b110 %
1'
b110 +
#800120000000
0!
0'
#800130000000
1!
b111 %
1'
b111 +
#800140000000
0!
0'
#800150000000
1!
0$
b1000 %
1'
0*
b1000 +
#800160000000
0!
0'
#800170000000
1!
b1001 %
1'
b1001 +
#800180000000
0!
0'
#800190000000
1!
b0 %
1'
b0 +
#800200000000
0!
0'
#800210000000
1!
1$
b1 %
1'
1*
b1 +
#800220000000
0!
0'
#800230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#800240000000
0!
0'
#800250000000
1!
b11 %
1'
b11 +
#800260000000
0!
0'
#800270000000
1!
b100 %
1'
b100 +
#800280000000
0!
0'
#800290000000
1!
b101 %
1'
b101 +
#800300000000
0!
0'
#800310000000
1!
0$
b110 %
1'
0*
b110 +
#800320000000
0!
0'
#800330000000
1!
b111 %
1'
b111 +
#800340000000
0!
0'
#800350000000
1!
b1000 %
1'
b1000 +
#800360000000
0!
0'
#800370000000
1!
b1001 %
1'
b1001 +
#800380000000
0!
0'
#800390000000
1!
b0 %
1'
b0 +
#800400000000
0!
0'
#800410000000
1!
1$
b1 %
1'
1*
b1 +
#800420000000
0!
0'
#800430000000
1!
b10 %
1'
b10 +
#800440000000
1"
1(
#800450000000
0!
0"
b100 &
0'
0(
b100 ,
#800460000000
1!
b11 %
1'
b11 +
#800470000000
0!
0'
#800480000000
1!
b100 %
1'
b100 +
#800490000000
0!
0'
#800500000000
1!
b101 %
1'
b101 +
#800510000000
0!
0'
#800520000000
1!
b110 %
1'
b110 +
#800530000000
0!
0'
#800540000000
1!
b111 %
1'
b111 +
#800550000000
0!
0'
#800560000000
1!
0$
b1000 %
1'
0*
b1000 +
#800570000000
0!
0'
#800580000000
1!
b1001 %
1'
b1001 +
#800590000000
0!
0'
#800600000000
1!
b0 %
1'
b0 +
#800610000000
0!
0'
#800620000000
1!
1$
b1 %
1'
1*
b1 +
#800630000000
0!
0'
#800640000000
1!
b10 %
1'
b10 +
#800650000000
0!
0'
#800660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#800670000000
0!
0'
#800680000000
1!
b100 %
1'
b100 +
#800690000000
0!
0'
#800700000000
1!
b101 %
1'
b101 +
#800710000000
0!
0'
#800720000000
1!
0$
b110 %
1'
0*
b110 +
#800730000000
0!
0'
#800740000000
1!
b111 %
1'
b111 +
#800750000000
0!
0'
#800760000000
1!
b1000 %
1'
b1000 +
#800770000000
0!
0'
#800780000000
1!
b1001 %
1'
b1001 +
#800790000000
0!
0'
#800800000000
1!
b0 %
1'
b0 +
#800810000000
0!
0'
#800820000000
1!
1$
b1 %
1'
1*
b1 +
#800830000000
0!
0'
#800840000000
1!
b10 %
1'
b10 +
#800850000000
0!
0'
#800860000000
1!
b11 %
1'
b11 +
#800870000000
1"
1(
#800880000000
0!
0"
b100 &
0'
0(
b100 ,
#800890000000
1!
b100 %
1'
b100 +
#800900000000
0!
0'
#800910000000
1!
b101 %
1'
b101 +
#800920000000
0!
0'
#800930000000
1!
b110 %
1'
b110 +
#800940000000
0!
0'
#800950000000
1!
b111 %
1'
b111 +
#800960000000
0!
0'
#800970000000
1!
0$
b1000 %
1'
0*
b1000 +
#800980000000
0!
0'
#800990000000
1!
b1001 %
1'
b1001 +
#801000000000
0!
0'
#801010000000
1!
b0 %
1'
b0 +
#801020000000
0!
0'
#801030000000
1!
1$
b1 %
1'
1*
b1 +
#801040000000
0!
0'
#801050000000
1!
b10 %
1'
b10 +
#801060000000
0!
0'
#801070000000
1!
b11 %
1'
b11 +
#801080000000
0!
0'
#801090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#801100000000
0!
0'
#801110000000
1!
b101 %
1'
b101 +
#801120000000
0!
0'
#801130000000
1!
0$
b110 %
1'
0*
b110 +
#801140000000
0!
0'
#801150000000
1!
b111 %
1'
b111 +
#801160000000
0!
0'
#801170000000
1!
b1000 %
1'
b1000 +
#801180000000
0!
0'
#801190000000
1!
b1001 %
1'
b1001 +
#801200000000
0!
0'
#801210000000
1!
b0 %
1'
b0 +
#801220000000
0!
0'
#801230000000
1!
1$
b1 %
1'
1*
b1 +
#801240000000
0!
0'
#801250000000
1!
b10 %
1'
b10 +
#801260000000
0!
0'
#801270000000
1!
b11 %
1'
b11 +
#801280000000
0!
0'
#801290000000
1!
b100 %
1'
b100 +
#801300000000
1"
1(
#801310000000
0!
0"
b100 &
0'
0(
b100 ,
#801320000000
1!
b101 %
1'
b101 +
#801330000000
0!
0'
#801340000000
1!
b110 %
1'
b110 +
#801350000000
0!
0'
#801360000000
1!
b111 %
1'
b111 +
#801370000000
0!
0'
#801380000000
1!
0$
b1000 %
1'
0*
b1000 +
#801390000000
0!
0'
#801400000000
1!
b1001 %
1'
b1001 +
#801410000000
0!
0'
#801420000000
1!
b0 %
1'
b0 +
#801430000000
0!
0'
#801440000000
1!
1$
b1 %
1'
1*
b1 +
#801450000000
0!
0'
#801460000000
1!
b10 %
1'
b10 +
#801470000000
0!
0'
#801480000000
1!
b11 %
1'
b11 +
#801490000000
0!
0'
#801500000000
1!
b100 %
1'
b100 +
#801510000000
0!
0'
#801520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#801530000000
0!
0'
#801540000000
1!
0$
b110 %
1'
0*
b110 +
#801550000000
0!
0'
#801560000000
1!
b111 %
1'
b111 +
#801570000000
0!
0'
#801580000000
1!
b1000 %
1'
b1000 +
#801590000000
0!
0'
#801600000000
1!
b1001 %
1'
b1001 +
#801610000000
0!
0'
#801620000000
1!
b0 %
1'
b0 +
#801630000000
0!
0'
#801640000000
1!
1$
b1 %
1'
1*
b1 +
#801650000000
0!
0'
#801660000000
1!
b10 %
1'
b10 +
#801670000000
0!
0'
#801680000000
1!
b11 %
1'
b11 +
#801690000000
0!
0'
#801700000000
1!
b100 %
1'
b100 +
#801710000000
0!
0'
#801720000000
1!
b101 %
1'
b101 +
#801730000000
1"
1(
#801740000000
0!
0"
b100 &
0'
0(
b100 ,
#801750000000
1!
b110 %
1'
b110 +
#801760000000
0!
0'
#801770000000
1!
b111 %
1'
b111 +
#801780000000
0!
0'
#801790000000
1!
0$
b1000 %
1'
0*
b1000 +
#801800000000
0!
0'
#801810000000
1!
b1001 %
1'
b1001 +
#801820000000
0!
0'
#801830000000
1!
b0 %
1'
b0 +
#801840000000
0!
0'
#801850000000
1!
1$
b1 %
1'
1*
b1 +
#801860000000
0!
0'
#801870000000
1!
b10 %
1'
b10 +
#801880000000
0!
0'
#801890000000
1!
b11 %
1'
b11 +
#801900000000
0!
0'
#801910000000
1!
b100 %
1'
b100 +
#801920000000
0!
0'
#801930000000
1!
b101 %
1'
b101 +
#801940000000
0!
0'
#801950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#801960000000
0!
0'
#801970000000
1!
b111 %
1'
b111 +
#801980000000
0!
0'
#801990000000
1!
b1000 %
1'
b1000 +
#802000000000
0!
0'
#802010000000
1!
b1001 %
1'
b1001 +
#802020000000
0!
0'
#802030000000
1!
b0 %
1'
b0 +
#802040000000
0!
0'
#802050000000
1!
1$
b1 %
1'
1*
b1 +
#802060000000
0!
0'
#802070000000
1!
b10 %
1'
b10 +
#802080000000
0!
0'
#802090000000
1!
b11 %
1'
b11 +
#802100000000
0!
0'
#802110000000
1!
b100 %
1'
b100 +
#802120000000
0!
0'
#802130000000
1!
b101 %
1'
b101 +
#802140000000
0!
0'
#802150000000
1!
0$
b110 %
1'
0*
b110 +
#802160000000
1"
1(
#802170000000
0!
0"
b100 &
0'
0(
b100 ,
#802180000000
1!
1$
b111 %
1'
1*
b111 +
#802190000000
0!
0'
#802200000000
1!
0$
b1000 %
1'
0*
b1000 +
#802210000000
0!
0'
#802220000000
1!
b1001 %
1'
b1001 +
#802230000000
0!
0'
#802240000000
1!
b0 %
1'
b0 +
#802250000000
0!
0'
#802260000000
1!
1$
b1 %
1'
1*
b1 +
#802270000000
0!
0'
#802280000000
1!
b10 %
1'
b10 +
#802290000000
0!
0'
#802300000000
1!
b11 %
1'
b11 +
#802310000000
0!
0'
#802320000000
1!
b100 %
1'
b100 +
#802330000000
0!
0'
#802340000000
1!
b101 %
1'
b101 +
#802350000000
0!
0'
#802360000000
1!
b110 %
1'
b110 +
#802370000000
0!
0'
#802380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#802390000000
0!
0'
#802400000000
1!
b1000 %
1'
b1000 +
#802410000000
0!
0'
#802420000000
1!
b1001 %
1'
b1001 +
#802430000000
0!
0'
#802440000000
1!
b0 %
1'
b0 +
#802450000000
0!
0'
#802460000000
1!
1$
b1 %
1'
1*
b1 +
#802470000000
0!
0'
#802480000000
1!
b10 %
1'
b10 +
#802490000000
0!
0'
#802500000000
1!
b11 %
1'
b11 +
#802510000000
0!
0'
#802520000000
1!
b100 %
1'
b100 +
#802530000000
0!
0'
#802540000000
1!
b101 %
1'
b101 +
#802550000000
0!
0'
#802560000000
1!
0$
b110 %
1'
0*
b110 +
#802570000000
0!
0'
#802580000000
1!
b111 %
1'
b111 +
#802590000000
1"
1(
#802600000000
0!
0"
b100 &
0'
0(
b100 ,
#802610000000
1!
b1000 %
1'
b1000 +
#802620000000
0!
0'
#802630000000
1!
b1001 %
1'
b1001 +
#802640000000
0!
0'
#802650000000
1!
b0 %
1'
b0 +
#802660000000
0!
0'
#802670000000
1!
1$
b1 %
1'
1*
b1 +
#802680000000
0!
0'
#802690000000
1!
b10 %
1'
b10 +
#802700000000
0!
0'
#802710000000
1!
b11 %
1'
b11 +
#802720000000
0!
0'
#802730000000
1!
b100 %
1'
b100 +
#802740000000
0!
0'
#802750000000
1!
b101 %
1'
b101 +
#802760000000
0!
0'
#802770000000
1!
b110 %
1'
b110 +
#802780000000
0!
0'
#802790000000
1!
b111 %
1'
b111 +
#802800000000
0!
0'
#802810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#802820000000
0!
0'
#802830000000
1!
b1001 %
1'
b1001 +
#802840000000
0!
0'
#802850000000
1!
b0 %
1'
b0 +
#802860000000
0!
0'
#802870000000
1!
1$
b1 %
1'
1*
b1 +
#802880000000
0!
0'
#802890000000
1!
b10 %
1'
b10 +
#802900000000
0!
0'
#802910000000
1!
b11 %
1'
b11 +
#802920000000
0!
0'
#802930000000
1!
b100 %
1'
b100 +
#802940000000
0!
0'
#802950000000
1!
b101 %
1'
b101 +
#802960000000
0!
0'
#802970000000
1!
0$
b110 %
1'
0*
b110 +
#802980000000
0!
0'
#802990000000
1!
b111 %
1'
b111 +
#803000000000
0!
0'
#803010000000
1!
b1000 %
1'
b1000 +
#803020000000
1"
1(
#803030000000
0!
0"
b100 &
0'
0(
b100 ,
#803040000000
1!
b1001 %
1'
b1001 +
#803050000000
0!
0'
#803060000000
1!
b0 %
1'
b0 +
#803070000000
0!
0'
#803080000000
1!
1$
b1 %
1'
1*
b1 +
#803090000000
0!
0'
#803100000000
1!
b10 %
1'
b10 +
#803110000000
0!
0'
#803120000000
1!
b11 %
1'
b11 +
#803130000000
0!
0'
#803140000000
1!
b100 %
1'
b100 +
#803150000000
0!
0'
#803160000000
1!
b101 %
1'
b101 +
#803170000000
0!
0'
#803180000000
1!
b110 %
1'
b110 +
#803190000000
0!
0'
#803200000000
1!
b111 %
1'
b111 +
#803210000000
0!
0'
#803220000000
1!
0$
b1000 %
1'
0*
b1000 +
#803230000000
0!
0'
#803240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#803250000000
0!
0'
#803260000000
1!
b0 %
1'
b0 +
#803270000000
0!
0'
#803280000000
1!
1$
b1 %
1'
1*
b1 +
#803290000000
0!
0'
#803300000000
1!
b10 %
1'
b10 +
#803310000000
0!
0'
#803320000000
1!
b11 %
1'
b11 +
#803330000000
0!
0'
#803340000000
1!
b100 %
1'
b100 +
#803350000000
0!
0'
#803360000000
1!
b101 %
1'
b101 +
#803370000000
0!
0'
#803380000000
1!
0$
b110 %
1'
0*
b110 +
#803390000000
0!
0'
#803400000000
1!
b111 %
1'
b111 +
#803410000000
0!
0'
#803420000000
1!
b1000 %
1'
b1000 +
#803430000000
0!
0'
#803440000000
1!
b1001 %
1'
b1001 +
#803450000000
1"
1(
#803460000000
0!
0"
b100 &
0'
0(
b100 ,
#803470000000
1!
b0 %
1'
b0 +
#803480000000
0!
0'
#803490000000
1!
1$
b1 %
1'
1*
b1 +
#803500000000
0!
0'
#803510000000
1!
b10 %
1'
b10 +
#803520000000
0!
0'
#803530000000
1!
b11 %
1'
b11 +
#803540000000
0!
0'
#803550000000
1!
b100 %
1'
b100 +
#803560000000
0!
0'
#803570000000
1!
b101 %
1'
b101 +
#803580000000
0!
0'
#803590000000
1!
b110 %
1'
b110 +
#803600000000
0!
0'
#803610000000
1!
b111 %
1'
b111 +
#803620000000
0!
0'
#803630000000
1!
0$
b1000 %
1'
0*
b1000 +
#803640000000
0!
0'
#803650000000
1!
b1001 %
1'
b1001 +
#803660000000
0!
0'
#803670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#803680000000
0!
0'
#803690000000
1!
1$
b1 %
1'
1*
b1 +
#803700000000
0!
0'
#803710000000
1!
b10 %
1'
b10 +
#803720000000
0!
0'
#803730000000
1!
b11 %
1'
b11 +
#803740000000
0!
0'
#803750000000
1!
b100 %
1'
b100 +
#803760000000
0!
0'
#803770000000
1!
b101 %
1'
b101 +
#803780000000
0!
0'
#803790000000
1!
0$
b110 %
1'
0*
b110 +
#803800000000
0!
0'
#803810000000
1!
b111 %
1'
b111 +
#803820000000
0!
0'
#803830000000
1!
b1000 %
1'
b1000 +
#803840000000
0!
0'
#803850000000
1!
b1001 %
1'
b1001 +
#803860000000
0!
0'
#803870000000
1!
b0 %
1'
b0 +
#803880000000
1"
1(
#803890000000
0!
0"
b100 &
0'
0(
b100 ,
#803900000000
1!
1$
b1 %
1'
1*
b1 +
#803910000000
0!
0'
#803920000000
1!
b10 %
1'
b10 +
#803930000000
0!
0'
#803940000000
1!
b11 %
1'
b11 +
#803950000000
0!
0'
#803960000000
1!
b100 %
1'
b100 +
#803970000000
0!
0'
#803980000000
1!
b101 %
1'
b101 +
#803990000000
0!
0'
#804000000000
1!
b110 %
1'
b110 +
#804010000000
0!
0'
#804020000000
1!
b111 %
1'
b111 +
#804030000000
0!
0'
#804040000000
1!
0$
b1000 %
1'
0*
b1000 +
#804050000000
0!
0'
#804060000000
1!
b1001 %
1'
b1001 +
#804070000000
0!
0'
#804080000000
1!
b0 %
1'
b0 +
#804090000000
0!
0'
#804100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#804110000000
0!
0'
#804120000000
1!
b10 %
1'
b10 +
#804130000000
0!
0'
#804140000000
1!
b11 %
1'
b11 +
#804150000000
0!
0'
#804160000000
1!
b100 %
1'
b100 +
#804170000000
0!
0'
#804180000000
1!
b101 %
1'
b101 +
#804190000000
0!
0'
#804200000000
1!
0$
b110 %
1'
0*
b110 +
#804210000000
0!
0'
#804220000000
1!
b111 %
1'
b111 +
#804230000000
0!
0'
#804240000000
1!
b1000 %
1'
b1000 +
#804250000000
0!
0'
#804260000000
1!
b1001 %
1'
b1001 +
#804270000000
0!
0'
#804280000000
1!
b0 %
1'
b0 +
#804290000000
0!
0'
#804300000000
1!
1$
b1 %
1'
1*
b1 +
#804310000000
1"
1(
#804320000000
0!
0"
b100 &
0'
0(
b100 ,
#804330000000
1!
b10 %
1'
b10 +
#804340000000
0!
0'
#804350000000
1!
b11 %
1'
b11 +
#804360000000
0!
0'
#804370000000
1!
b100 %
1'
b100 +
#804380000000
0!
0'
#804390000000
1!
b101 %
1'
b101 +
#804400000000
0!
0'
#804410000000
1!
b110 %
1'
b110 +
#804420000000
0!
0'
#804430000000
1!
b111 %
1'
b111 +
#804440000000
0!
0'
#804450000000
1!
0$
b1000 %
1'
0*
b1000 +
#804460000000
0!
0'
#804470000000
1!
b1001 %
1'
b1001 +
#804480000000
0!
0'
#804490000000
1!
b0 %
1'
b0 +
#804500000000
0!
0'
#804510000000
1!
1$
b1 %
1'
1*
b1 +
#804520000000
0!
0'
#804530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#804540000000
0!
0'
#804550000000
1!
b11 %
1'
b11 +
#804560000000
0!
0'
#804570000000
1!
b100 %
1'
b100 +
#804580000000
0!
0'
#804590000000
1!
b101 %
1'
b101 +
#804600000000
0!
0'
#804610000000
1!
0$
b110 %
1'
0*
b110 +
#804620000000
0!
0'
#804630000000
1!
b111 %
1'
b111 +
#804640000000
0!
0'
#804650000000
1!
b1000 %
1'
b1000 +
#804660000000
0!
0'
#804670000000
1!
b1001 %
1'
b1001 +
#804680000000
0!
0'
#804690000000
1!
b0 %
1'
b0 +
#804700000000
0!
0'
#804710000000
1!
1$
b1 %
1'
1*
b1 +
#804720000000
0!
0'
#804730000000
1!
b10 %
1'
b10 +
#804740000000
1"
1(
#804750000000
0!
0"
b100 &
0'
0(
b100 ,
#804760000000
1!
b11 %
1'
b11 +
#804770000000
0!
0'
#804780000000
1!
b100 %
1'
b100 +
#804790000000
0!
0'
#804800000000
1!
b101 %
1'
b101 +
#804810000000
0!
0'
#804820000000
1!
b110 %
1'
b110 +
#804830000000
0!
0'
#804840000000
1!
b111 %
1'
b111 +
#804850000000
0!
0'
#804860000000
1!
0$
b1000 %
1'
0*
b1000 +
#804870000000
0!
0'
#804880000000
1!
b1001 %
1'
b1001 +
#804890000000
0!
0'
#804900000000
1!
b0 %
1'
b0 +
#804910000000
0!
0'
#804920000000
1!
1$
b1 %
1'
1*
b1 +
#804930000000
0!
0'
#804940000000
1!
b10 %
1'
b10 +
#804950000000
0!
0'
#804960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#804970000000
0!
0'
#804980000000
1!
b100 %
1'
b100 +
#804990000000
0!
0'
#805000000000
1!
b101 %
1'
b101 +
#805010000000
0!
0'
#805020000000
1!
0$
b110 %
1'
0*
b110 +
#805030000000
0!
0'
#805040000000
1!
b111 %
1'
b111 +
#805050000000
0!
0'
#805060000000
1!
b1000 %
1'
b1000 +
#805070000000
0!
0'
#805080000000
1!
b1001 %
1'
b1001 +
#805090000000
0!
0'
#805100000000
1!
b0 %
1'
b0 +
#805110000000
0!
0'
#805120000000
1!
1$
b1 %
1'
1*
b1 +
#805130000000
0!
0'
#805140000000
1!
b10 %
1'
b10 +
#805150000000
0!
0'
#805160000000
1!
b11 %
1'
b11 +
#805170000000
1"
1(
#805180000000
0!
0"
b100 &
0'
0(
b100 ,
#805190000000
1!
b100 %
1'
b100 +
#805200000000
0!
0'
#805210000000
1!
b101 %
1'
b101 +
#805220000000
0!
0'
#805230000000
1!
b110 %
1'
b110 +
#805240000000
0!
0'
#805250000000
1!
b111 %
1'
b111 +
#805260000000
0!
0'
#805270000000
1!
0$
b1000 %
1'
0*
b1000 +
#805280000000
0!
0'
#805290000000
1!
b1001 %
1'
b1001 +
#805300000000
0!
0'
#805310000000
1!
b0 %
1'
b0 +
#805320000000
0!
0'
#805330000000
1!
1$
b1 %
1'
1*
b1 +
#805340000000
0!
0'
#805350000000
1!
b10 %
1'
b10 +
#805360000000
0!
0'
#805370000000
1!
b11 %
1'
b11 +
#805380000000
0!
0'
#805390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#805400000000
0!
0'
#805410000000
1!
b101 %
1'
b101 +
#805420000000
0!
0'
#805430000000
1!
0$
b110 %
1'
0*
b110 +
#805440000000
0!
0'
#805450000000
1!
b111 %
1'
b111 +
#805460000000
0!
0'
#805470000000
1!
b1000 %
1'
b1000 +
#805480000000
0!
0'
#805490000000
1!
b1001 %
1'
b1001 +
#805500000000
0!
0'
#805510000000
1!
b0 %
1'
b0 +
#805520000000
0!
0'
#805530000000
1!
1$
b1 %
1'
1*
b1 +
#805540000000
0!
0'
#805550000000
1!
b10 %
1'
b10 +
#805560000000
0!
0'
#805570000000
1!
b11 %
1'
b11 +
#805580000000
0!
0'
#805590000000
1!
b100 %
1'
b100 +
#805600000000
1"
1(
#805610000000
0!
0"
b100 &
0'
0(
b100 ,
#805620000000
1!
b101 %
1'
b101 +
#805630000000
0!
0'
#805640000000
1!
b110 %
1'
b110 +
#805650000000
0!
0'
#805660000000
1!
b111 %
1'
b111 +
#805670000000
0!
0'
#805680000000
1!
0$
b1000 %
1'
0*
b1000 +
#805690000000
0!
0'
#805700000000
1!
b1001 %
1'
b1001 +
#805710000000
0!
0'
#805720000000
1!
b0 %
1'
b0 +
#805730000000
0!
0'
#805740000000
1!
1$
b1 %
1'
1*
b1 +
#805750000000
0!
0'
#805760000000
1!
b10 %
1'
b10 +
#805770000000
0!
0'
#805780000000
1!
b11 %
1'
b11 +
#805790000000
0!
0'
#805800000000
1!
b100 %
1'
b100 +
#805810000000
0!
0'
#805820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#805830000000
0!
0'
#805840000000
1!
0$
b110 %
1'
0*
b110 +
#805850000000
0!
0'
#805860000000
1!
b111 %
1'
b111 +
#805870000000
0!
0'
#805880000000
1!
b1000 %
1'
b1000 +
#805890000000
0!
0'
#805900000000
1!
b1001 %
1'
b1001 +
#805910000000
0!
0'
#805920000000
1!
b0 %
1'
b0 +
#805930000000
0!
0'
#805940000000
1!
1$
b1 %
1'
1*
b1 +
#805950000000
0!
0'
#805960000000
1!
b10 %
1'
b10 +
#805970000000
0!
0'
#805980000000
1!
b11 %
1'
b11 +
#805990000000
0!
0'
#806000000000
1!
b100 %
1'
b100 +
#806010000000
0!
0'
#806020000000
1!
b101 %
1'
b101 +
#806030000000
1"
1(
#806040000000
0!
0"
b100 &
0'
0(
b100 ,
#806050000000
1!
b110 %
1'
b110 +
#806060000000
0!
0'
#806070000000
1!
b111 %
1'
b111 +
#806080000000
0!
0'
#806090000000
1!
0$
b1000 %
1'
0*
b1000 +
#806100000000
0!
0'
#806110000000
1!
b1001 %
1'
b1001 +
#806120000000
0!
0'
#806130000000
1!
b0 %
1'
b0 +
#806140000000
0!
0'
#806150000000
1!
1$
b1 %
1'
1*
b1 +
#806160000000
0!
0'
#806170000000
1!
b10 %
1'
b10 +
#806180000000
0!
0'
#806190000000
1!
b11 %
1'
b11 +
#806200000000
0!
0'
#806210000000
1!
b100 %
1'
b100 +
#806220000000
0!
0'
#806230000000
1!
b101 %
1'
b101 +
#806240000000
0!
0'
#806250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#806260000000
0!
0'
#806270000000
1!
b111 %
1'
b111 +
#806280000000
0!
0'
#806290000000
1!
b1000 %
1'
b1000 +
#806300000000
0!
0'
#806310000000
1!
b1001 %
1'
b1001 +
#806320000000
0!
0'
#806330000000
1!
b0 %
1'
b0 +
#806340000000
0!
0'
#806350000000
1!
1$
b1 %
1'
1*
b1 +
#806360000000
0!
0'
#806370000000
1!
b10 %
1'
b10 +
#806380000000
0!
0'
#806390000000
1!
b11 %
1'
b11 +
#806400000000
0!
0'
#806410000000
1!
b100 %
1'
b100 +
#806420000000
0!
0'
#806430000000
1!
b101 %
1'
b101 +
#806440000000
0!
0'
#806450000000
1!
0$
b110 %
1'
0*
b110 +
#806460000000
1"
1(
#806470000000
0!
0"
b100 &
0'
0(
b100 ,
#806480000000
1!
1$
b111 %
1'
1*
b111 +
#806490000000
0!
0'
#806500000000
1!
0$
b1000 %
1'
0*
b1000 +
#806510000000
0!
0'
#806520000000
1!
b1001 %
1'
b1001 +
#806530000000
0!
0'
#806540000000
1!
b0 %
1'
b0 +
#806550000000
0!
0'
#806560000000
1!
1$
b1 %
1'
1*
b1 +
#806570000000
0!
0'
#806580000000
1!
b10 %
1'
b10 +
#806590000000
0!
0'
#806600000000
1!
b11 %
1'
b11 +
#806610000000
0!
0'
#806620000000
1!
b100 %
1'
b100 +
#806630000000
0!
0'
#806640000000
1!
b101 %
1'
b101 +
#806650000000
0!
0'
#806660000000
1!
b110 %
1'
b110 +
#806670000000
0!
0'
#806680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#806690000000
0!
0'
#806700000000
1!
b1000 %
1'
b1000 +
#806710000000
0!
0'
#806720000000
1!
b1001 %
1'
b1001 +
#806730000000
0!
0'
#806740000000
1!
b0 %
1'
b0 +
#806750000000
0!
0'
#806760000000
1!
1$
b1 %
1'
1*
b1 +
#806770000000
0!
0'
#806780000000
1!
b10 %
1'
b10 +
#806790000000
0!
0'
#806800000000
1!
b11 %
1'
b11 +
#806810000000
0!
0'
#806820000000
1!
b100 %
1'
b100 +
#806830000000
0!
0'
#806840000000
1!
b101 %
1'
b101 +
#806850000000
0!
0'
#806860000000
1!
0$
b110 %
1'
0*
b110 +
#806870000000
0!
0'
#806880000000
1!
b111 %
1'
b111 +
#806890000000
1"
1(
#806900000000
0!
0"
b100 &
0'
0(
b100 ,
#806910000000
1!
b1000 %
1'
b1000 +
#806920000000
0!
0'
#806930000000
1!
b1001 %
1'
b1001 +
#806940000000
0!
0'
#806950000000
1!
b0 %
1'
b0 +
#806960000000
0!
0'
#806970000000
1!
1$
b1 %
1'
1*
b1 +
#806980000000
0!
0'
#806990000000
1!
b10 %
1'
b10 +
#807000000000
0!
0'
#807010000000
1!
b11 %
1'
b11 +
#807020000000
0!
0'
#807030000000
1!
b100 %
1'
b100 +
#807040000000
0!
0'
#807050000000
1!
b101 %
1'
b101 +
#807060000000
0!
0'
#807070000000
1!
b110 %
1'
b110 +
#807080000000
0!
0'
#807090000000
1!
b111 %
1'
b111 +
#807100000000
0!
0'
#807110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#807120000000
0!
0'
#807130000000
1!
b1001 %
1'
b1001 +
#807140000000
0!
0'
#807150000000
1!
b0 %
1'
b0 +
#807160000000
0!
0'
#807170000000
1!
1$
b1 %
1'
1*
b1 +
#807180000000
0!
0'
#807190000000
1!
b10 %
1'
b10 +
#807200000000
0!
0'
#807210000000
1!
b11 %
1'
b11 +
#807220000000
0!
0'
#807230000000
1!
b100 %
1'
b100 +
#807240000000
0!
0'
#807250000000
1!
b101 %
1'
b101 +
#807260000000
0!
0'
#807270000000
1!
0$
b110 %
1'
0*
b110 +
#807280000000
0!
0'
#807290000000
1!
b111 %
1'
b111 +
#807300000000
0!
0'
#807310000000
1!
b1000 %
1'
b1000 +
#807320000000
1"
1(
#807330000000
0!
0"
b100 &
0'
0(
b100 ,
#807340000000
1!
b1001 %
1'
b1001 +
#807350000000
0!
0'
#807360000000
1!
b0 %
1'
b0 +
#807370000000
0!
0'
#807380000000
1!
1$
b1 %
1'
1*
b1 +
#807390000000
0!
0'
#807400000000
1!
b10 %
1'
b10 +
#807410000000
0!
0'
#807420000000
1!
b11 %
1'
b11 +
#807430000000
0!
0'
#807440000000
1!
b100 %
1'
b100 +
#807450000000
0!
0'
#807460000000
1!
b101 %
1'
b101 +
#807470000000
0!
0'
#807480000000
1!
b110 %
1'
b110 +
#807490000000
0!
0'
#807500000000
1!
b111 %
1'
b111 +
#807510000000
0!
0'
#807520000000
1!
0$
b1000 %
1'
0*
b1000 +
#807530000000
0!
0'
#807540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#807550000000
0!
0'
#807560000000
1!
b0 %
1'
b0 +
#807570000000
0!
0'
#807580000000
1!
1$
b1 %
1'
1*
b1 +
#807590000000
0!
0'
#807600000000
1!
b10 %
1'
b10 +
#807610000000
0!
0'
#807620000000
1!
b11 %
1'
b11 +
#807630000000
0!
0'
#807640000000
1!
b100 %
1'
b100 +
#807650000000
0!
0'
#807660000000
1!
b101 %
1'
b101 +
#807670000000
0!
0'
#807680000000
1!
0$
b110 %
1'
0*
b110 +
#807690000000
0!
0'
#807700000000
1!
b111 %
1'
b111 +
#807710000000
0!
0'
#807720000000
1!
b1000 %
1'
b1000 +
#807730000000
0!
0'
#807740000000
1!
b1001 %
1'
b1001 +
#807750000000
1"
1(
#807760000000
0!
0"
b100 &
0'
0(
b100 ,
#807770000000
1!
b0 %
1'
b0 +
#807780000000
0!
0'
#807790000000
1!
1$
b1 %
1'
1*
b1 +
#807800000000
0!
0'
#807810000000
1!
b10 %
1'
b10 +
#807820000000
0!
0'
#807830000000
1!
b11 %
1'
b11 +
#807840000000
0!
0'
#807850000000
1!
b100 %
1'
b100 +
#807860000000
0!
0'
#807870000000
1!
b101 %
1'
b101 +
#807880000000
0!
0'
#807890000000
1!
b110 %
1'
b110 +
#807900000000
0!
0'
#807910000000
1!
b111 %
1'
b111 +
#807920000000
0!
0'
#807930000000
1!
0$
b1000 %
1'
0*
b1000 +
#807940000000
0!
0'
#807950000000
1!
b1001 %
1'
b1001 +
#807960000000
0!
0'
#807970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#807980000000
0!
0'
#807990000000
1!
1$
b1 %
1'
1*
b1 +
#808000000000
0!
0'
#808010000000
1!
b10 %
1'
b10 +
#808020000000
0!
0'
#808030000000
1!
b11 %
1'
b11 +
#808040000000
0!
0'
#808050000000
1!
b100 %
1'
b100 +
#808060000000
0!
0'
#808070000000
1!
b101 %
1'
b101 +
#808080000000
0!
0'
#808090000000
1!
0$
b110 %
1'
0*
b110 +
#808100000000
0!
0'
#808110000000
1!
b111 %
1'
b111 +
#808120000000
0!
0'
#808130000000
1!
b1000 %
1'
b1000 +
#808140000000
0!
0'
#808150000000
1!
b1001 %
1'
b1001 +
#808160000000
0!
0'
#808170000000
1!
b0 %
1'
b0 +
#808180000000
1"
1(
#808190000000
0!
0"
b100 &
0'
0(
b100 ,
#808200000000
1!
1$
b1 %
1'
1*
b1 +
#808210000000
0!
0'
#808220000000
1!
b10 %
1'
b10 +
#808230000000
0!
0'
#808240000000
1!
b11 %
1'
b11 +
#808250000000
0!
0'
#808260000000
1!
b100 %
1'
b100 +
#808270000000
0!
0'
#808280000000
1!
b101 %
1'
b101 +
#808290000000
0!
0'
#808300000000
1!
b110 %
1'
b110 +
#808310000000
0!
0'
#808320000000
1!
b111 %
1'
b111 +
#808330000000
0!
0'
#808340000000
1!
0$
b1000 %
1'
0*
b1000 +
#808350000000
0!
0'
#808360000000
1!
b1001 %
1'
b1001 +
#808370000000
0!
0'
#808380000000
1!
b0 %
1'
b0 +
#808390000000
0!
0'
#808400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#808410000000
0!
0'
#808420000000
1!
b10 %
1'
b10 +
#808430000000
0!
0'
#808440000000
1!
b11 %
1'
b11 +
#808450000000
0!
0'
#808460000000
1!
b100 %
1'
b100 +
#808470000000
0!
0'
#808480000000
1!
b101 %
1'
b101 +
#808490000000
0!
0'
#808500000000
1!
0$
b110 %
1'
0*
b110 +
#808510000000
0!
0'
#808520000000
1!
b111 %
1'
b111 +
#808530000000
0!
0'
#808540000000
1!
b1000 %
1'
b1000 +
#808550000000
0!
0'
#808560000000
1!
b1001 %
1'
b1001 +
#808570000000
0!
0'
#808580000000
1!
b0 %
1'
b0 +
#808590000000
0!
0'
#808600000000
1!
1$
b1 %
1'
1*
b1 +
#808610000000
1"
1(
#808620000000
0!
0"
b100 &
0'
0(
b100 ,
#808630000000
1!
b10 %
1'
b10 +
#808640000000
0!
0'
#808650000000
1!
b11 %
1'
b11 +
#808660000000
0!
0'
#808670000000
1!
b100 %
1'
b100 +
#808680000000
0!
0'
#808690000000
1!
b101 %
1'
b101 +
#808700000000
0!
0'
#808710000000
1!
b110 %
1'
b110 +
#808720000000
0!
0'
#808730000000
1!
b111 %
1'
b111 +
#808740000000
0!
0'
#808750000000
1!
0$
b1000 %
1'
0*
b1000 +
#808760000000
0!
0'
#808770000000
1!
b1001 %
1'
b1001 +
#808780000000
0!
0'
#808790000000
1!
b0 %
1'
b0 +
#808800000000
0!
0'
#808810000000
1!
1$
b1 %
1'
1*
b1 +
#808820000000
0!
0'
#808830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#808840000000
0!
0'
#808850000000
1!
b11 %
1'
b11 +
#808860000000
0!
0'
#808870000000
1!
b100 %
1'
b100 +
#808880000000
0!
0'
#808890000000
1!
b101 %
1'
b101 +
#808900000000
0!
0'
#808910000000
1!
0$
b110 %
1'
0*
b110 +
#808920000000
0!
0'
#808930000000
1!
b111 %
1'
b111 +
#808940000000
0!
0'
#808950000000
1!
b1000 %
1'
b1000 +
#808960000000
0!
0'
#808970000000
1!
b1001 %
1'
b1001 +
#808980000000
0!
0'
#808990000000
1!
b0 %
1'
b0 +
#809000000000
0!
0'
#809010000000
1!
1$
b1 %
1'
1*
b1 +
#809020000000
0!
0'
#809030000000
1!
b10 %
1'
b10 +
#809040000000
1"
1(
#809050000000
0!
0"
b100 &
0'
0(
b100 ,
#809060000000
1!
b11 %
1'
b11 +
#809070000000
0!
0'
#809080000000
1!
b100 %
1'
b100 +
#809090000000
0!
0'
#809100000000
1!
b101 %
1'
b101 +
#809110000000
0!
0'
#809120000000
1!
b110 %
1'
b110 +
#809130000000
0!
0'
#809140000000
1!
b111 %
1'
b111 +
#809150000000
0!
0'
#809160000000
1!
0$
b1000 %
1'
0*
b1000 +
#809170000000
0!
0'
#809180000000
1!
b1001 %
1'
b1001 +
#809190000000
0!
0'
#809200000000
1!
b0 %
1'
b0 +
#809210000000
0!
0'
#809220000000
1!
1$
b1 %
1'
1*
b1 +
#809230000000
0!
0'
#809240000000
1!
b10 %
1'
b10 +
#809250000000
0!
0'
#809260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#809270000000
0!
0'
#809280000000
1!
b100 %
1'
b100 +
#809290000000
0!
0'
#809300000000
1!
b101 %
1'
b101 +
#809310000000
0!
0'
#809320000000
1!
0$
b110 %
1'
0*
b110 +
#809330000000
0!
0'
#809340000000
1!
b111 %
1'
b111 +
#809350000000
0!
0'
#809360000000
1!
b1000 %
1'
b1000 +
#809370000000
0!
0'
#809380000000
1!
b1001 %
1'
b1001 +
#809390000000
0!
0'
#809400000000
1!
b0 %
1'
b0 +
#809410000000
0!
0'
#809420000000
1!
1$
b1 %
1'
1*
b1 +
#809430000000
0!
0'
#809440000000
1!
b10 %
1'
b10 +
#809450000000
0!
0'
#809460000000
1!
b11 %
1'
b11 +
#809470000000
1"
1(
#809480000000
0!
0"
b100 &
0'
0(
b100 ,
#809490000000
1!
b100 %
1'
b100 +
#809500000000
0!
0'
#809510000000
1!
b101 %
1'
b101 +
#809520000000
0!
0'
#809530000000
1!
b110 %
1'
b110 +
#809540000000
0!
0'
#809550000000
1!
b111 %
1'
b111 +
#809560000000
0!
0'
#809570000000
1!
0$
b1000 %
1'
0*
b1000 +
#809580000000
0!
0'
#809590000000
1!
b1001 %
1'
b1001 +
#809600000000
0!
0'
#809610000000
1!
b0 %
1'
b0 +
#809620000000
0!
0'
#809630000000
1!
1$
b1 %
1'
1*
b1 +
#809640000000
0!
0'
#809650000000
1!
b10 %
1'
b10 +
#809660000000
0!
0'
#809670000000
1!
b11 %
1'
b11 +
#809680000000
0!
0'
#809690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#809700000000
0!
0'
#809710000000
1!
b101 %
1'
b101 +
#809720000000
0!
0'
#809730000000
1!
0$
b110 %
1'
0*
b110 +
#809740000000
0!
0'
#809750000000
1!
b111 %
1'
b111 +
#809760000000
0!
0'
#809770000000
1!
b1000 %
1'
b1000 +
#809780000000
0!
0'
#809790000000
1!
b1001 %
1'
b1001 +
#809800000000
0!
0'
#809810000000
1!
b0 %
1'
b0 +
#809820000000
0!
0'
#809830000000
1!
1$
b1 %
1'
1*
b1 +
#809840000000
0!
0'
#809850000000
1!
b10 %
1'
b10 +
#809860000000
0!
0'
#809870000000
1!
b11 %
1'
b11 +
#809880000000
0!
0'
#809890000000
1!
b100 %
1'
b100 +
#809900000000
1"
1(
#809910000000
0!
0"
b100 &
0'
0(
b100 ,
#809920000000
1!
b101 %
1'
b101 +
#809930000000
0!
0'
#809940000000
1!
b110 %
1'
b110 +
#809950000000
0!
0'
#809960000000
1!
b111 %
1'
b111 +
#809970000000
0!
0'
#809980000000
1!
0$
b1000 %
1'
0*
b1000 +
#809990000000
0!
0'
#810000000000
1!
b1001 %
1'
b1001 +
#810010000000
0!
0'
#810020000000
1!
b0 %
1'
b0 +
#810030000000
0!
0'
#810040000000
1!
1$
b1 %
1'
1*
b1 +
#810050000000
0!
0'
#810060000000
1!
b10 %
1'
b10 +
#810070000000
0!
0'
#810080000000
1!
b11 %
1'
b11 +
#810090000000
0!
0'
#810100000000
1!
b100 %
1'
b100 +
#810110000000
0!
0'
#810120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#810130000000
0!
0'
#810140000000
1!
0$
b110 %
1'
0*
b110 +
#810150000000
0!
0'
#810160000000
1!
b111 %
1'
b111 +
#810170000000
0!
0'
#810180000000
1!
b1000 %
1'
b1000 +
#810190000000
0!
0'
#810200000000
1!
b1001 %
1'
b1001 +
#810210000000
0!
0'
#810220000000
1!
b0 %
1'
b0 +
#810230000000
0!
0'
#810240000000
1!
1$
b1 %
1'
1*
b1 +
#810250000000
0!
0'
#810260000000
1!
b10 %
1'
b10 +
#810270000000
0!
0'
#810280000000
1!
b11 %
1'
b11 +
#810290000000
0!
0'
#810300000000
1!
b100 %
1'
b100 +
#810310000000
0!
0'
#810320000000
1!
b101 %
1'
b101 +
#810330000000
1"
1(
#810340000000
0!
0"
b100 &
0'
0(
b100 ,
#810350000000
1!
b110 %
1'
b110 +
#810360000000
0!
0'
#810370000000
1!
b111 %
1'
b111 +
#810380000000
0!
0'
#810390000000
1!
0$
b1000 %
1'
0*
b1000 +
#810400000000
0!
0'
#810410000000
1!
b1001 %
1'
b1001 +
#810420000000
0!
0'
#810430000000
1!
b0 %
1'
b0 +
#810440000000
0!
0'
#810450000000
1!
1$
b1 %
1'
1*
b1 +
#810460000000
0!
0'
#810470000000
1!
b10 %
1'
b10 +
#810480000000
0!
0'
#810490000000
1!
b11 %
1'
b11 +
#810500000000
0!
0'
#810510000000
1!
b100 %
1'
b100 +
#810520000000
0!
0'
#810530000000
1!
b101 %
1'
b101 +
#810540000000
0!
0'
#810550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#810560000000
0!
0'
#810570000000
1!
b111 %
1'
b111 +
#810580000000
0!
0'
#810590000000
1!
b1000 %
1'
b1000 +
#810600000000
0!
0'
#810610000000
1!
b1001 %
1'
b1001 +
#810620000000
0!
0'
#810630000000
1!
b0 %
1'
b0 +
#810640000000
0!
0'
#810650000000
1!
1$
b1 %
1'
1*
b1 +
#810660000000
0!
0'
#810670000000
1!
b10 %
1'
b10 +
#810680000000
0!
0'
#810690000000
1!
b11 %
1'
b11 +
#810700000000
0!
0'
#810710000000
1!
b100 %
1'
b100 +
#810720000000
0!
0'
#810730000000
1!
b101 %
1'
b101 +
#810740000000
0!
0'
#810750000000
1!
0$
b110 %
1'
0*
b110 +
#810760000000
1"
1(
#810770000000
0!
0"
b100 &
0'
0(
b100 ,
#810780000000
1!
1$
b111 %
1'
1*
b111 +
#810790000000
0!
0'
#810800000000
1!
0$
b1000 %
1'
0*
b1000 +
#810810000000
0!
0'
#810820000000
1!
b1001 %
1'
b1001 +
#810830000000
0!
0'
#810840000000
1!
b0 %
1'
b0 +
#810850000000
0!
0'
#810860000000
1!
1$
b1 %
1'
1*
b1 +
#810870000000
0!
0'
#810880000000
1!
b10 %
1'
b10 +
#810890000000
0!
0'
#810900000000
1!
b11 %
1'
b11 +
#810910000000
0!
0'
#810920000000
1!
b100 %
1'
b100 +
#810930000000
0!
0'
#810940000000
1!
b101 %
1'
b101 +
#810950000000
0!
0'
#810960000000
1!
b110 %
1'
b110 +
#810970000000
0!
0'
#810980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#810990000000
0!
0'
#811000000000
1!
b1000 %
1'
b1000 +
#811010000000
0!
0'
#811020000000
1!
b1001 %
1'
b1001 +
#811030000000
0!
0'
#811040000000
1!
b0 %
1'
b0 +
#811050000000
0!
0'
#811060000000
1!
1$
b1 %
1'
1*
b1 +
#811070000000
0!
0'
#811080000000
1!
b10 %
1'
b10 +
#811090000000
0!
0'
#811100000000
1!
b11 %
1'
b11 +
#811110000000
0!
0'
#811120000000
1!
b100 %
1'
b100 +
#811130000000
0!
0'
#811140000000
1!
b101 %
1'
b101 +
#811150000000
0!
0'
#811160000000
1!
0$
b110 %
1'
0*
b110 +
#811170000000
0!
0'
#811180000000
1!
b111 %
1'
b111 +
#811190000000
1"
1(
#811200000000
0!
0"
b100 &
0'
0(
b100 ,
#811210000000
1!
b1000 %
1'
b1000 +
#811220000000
0!
0'
#811230000000
1!
b1001 %
1'
b1001 +
#811240000000
0!
0'
#811250000000
1!
b0 %
1'
b0 +
#811260000000
0!
0'
#811270000000
1!
1$
b1 %
1'
1*
b1 +
#811280000000
0!
0'
#811290000000
1!
b10 %
1'
b10 +
#811300000000
0!
0'
#811310000000
1!
b11 %
1'
b11 +
#811320000000
0!
0'
#811330000000
1!
b100 %
1'
b100 +
#811340000000
0!
0'
#811350000000
1!
b101 %
1'
b101 +
#811360000000
0!
0'
#811370000000
1!
b110 %
1'
b110 +
#811380000000
0!
0'
#811390000000
1!
b111 %
1'
b111 +
#811400000000
0!
0'
#811410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#811420000000
0!
0'
#811430000000
1!
b1001 %
1'
b1001 +
#811440000000
0!
0'
#811450000000
1!
b0 %
1'
b0 +
#811460000000
0!
0'
#811470000000
1!
1$
b1 %
1'
1*
b1 +
#811480000000
0!
0'
#811490000000
1!
b10 %
1'
b10 +
#811500000000
0!
0'
#811510000000
1!
b11 %
1'
b11 +
#811520000000
0!
0'
#811530000000
1!
b100 %
1'
b100 +
#811540000000
0!
0'
#811550000000
1!
b101 %
1'
b101 +
#811560000000
0!
0'
#811570000000
1!
0$
b110 %
1'
0*
b110 +
#811580000000
0!
0'
#811590000000
1!
b111 %
1'
b111 +
#811600000000
0!
0'
#811610000000
1!
b1000 %
1'
b1000 +
#811620000000
1"
1(
#811630000000
0!
0"
b100 &
0'
0(
b100 ,
#811640000000
1!
b1001 %
1'
b1001 +
#811650000000
0!
0'
#811660000000
1!
b0 %
1'
b0 +
#811670000000
0!
0'
#811680000000
1!
1$
b1 %
1'
1*
b1 +
#811690000000
0!
0'
#811700000000
1!
b10 %
1'
b10 +
#811710000000
0!
0'
#811720000000
1!
b11 %
1'
b11 +
#811730000000
0!
0'
#811740000000
1!
b100 %
1'
b100 +
#811750000000
0!
0'
#811760000000
1!
b101 %
1'
b101 +
#811770000000
0!
0'
#811780000000
1!
b110 %
1'
b110 +
#811790000000
0!
0'
#811800000000
1!
b111 %
1'
b111 +
#811810000000
0!
0'
#811820000000
1!
0$
b1000 %
1'
0*
b1000 +
#811830000000
0!
0'
#811840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#811850000000
0!
0'
#811860000000
1!
b0 %
1'
b0 +
#811870000000
0!
0'
#811880000000
1!
1$
b1 %
1'
1*
b1 +
#811890000000
0!
0'
#811900000000
1!
b10 %
1'
b10 +
#811910000000
0!
0'
#811920000000
1!
b11 %
1'
b11 +
#811930000000
0!
0'
#811940000000
1!
b100 %
1'
b100 +
#811950000000
0!
0'
#811960000000
1!
b101 %
1'
b101 +
#811970000000
0!
0'
#811980000000
1!
0$
b110 %
1'
0*
b110 +
#811990000000
0!
0'
#812000000000
1!
b111 %
1'
b111 +
#812010000000
0!
0'
#812020000000
1!
b1000 %
1'
b1000 +
#812030000000
0!
0'
#812040000000
1!
b1001 %
1'
b1001 +
#812050000000
1"
1(
#812060000000
0!
0"
b100 &
0'
0(
b100 ,
#812070000000
1!
b0 %
1'
b0 +
#812080000000
0!
0'
#812090000000
1!
1$
b1 %
1'
1*
b1 +
#812100000000
0!
0'
#812110000000
1!
b10 %
1'
b10 +
#812120000000
0!
0'
#812130000000
1!
b11 %
1'
b11 +
#812140000000
0!
0'
#812150000000
1!
b100 %
1'
b100 +
#812160000000
0!
0'
#812170000000
1!
b101 %
1'
b101 +
#812180000000
0!
0'
#812190000000
1!
b110 %
1'
b110 +
#812200000000
0!
0'
#812210000000
1!
b111 %
1'
b111 +
#812220000000
0!
0'
#812230000000
1!
0$
b1000 %
1'
0*
b1000 +
#812240000000
0!
0'
#812250000000
1!
b1001 %
1'
b1001 +
#812260000000
0!
0'
#812270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#812280000000
0!
0'
#812290000000
1!
1$
b1 %
1'
1*
b1 +
#812300000000
0!
0'
#812310000000
1!
b10 %
1'
b10 +
#812320000000
0!
0'
#812330000000
1!
b11 %
1'
b11 +
#812340000000
0!
0'
#812350000000
1!
b100 %
1'
b100 +
#812360000000
0!
0'
#812370000000
1!
b101 %
1'
b101 +
#812380000000
0!
0'
#812390000000
1!
0$
b110 %
1'
0*
b110 +
#812400000000
0!
0'
#812410000000
1!
b111 %
1'
b111 +
#812420000000
0!
0'
#812430000000
1!
b1000 %
1'
b1000 +
#812440000000
0!
0'
#812450000000
1!
b1001 %
1'
b1001 +
#812460000000
0!
0'
#812470000000
1!
b0 %
1'
b0 +
#812480000000
1"
1(
#812490000000
0!
0"
b100 &
0'
0(
b100 ,
#812500000000
1!
1$
b1 %
1'
1*
b1 +
#812510000000
0!
0'
#812520000000
1!
b10 %
1'
b10 +
#812530000000
0!
0'
#812540000000
1!
b11 %
1'
b11 +
#812550000000
0!
0'
#812560000000
1!
b100 %
1'
b100 +
#812570000000
0!
0'
#812580000000
1!
b101 %
1'
b101 +
#812590000000
0!
0'
#812600000000
1!
b110 %
1'
b110 +
#812610000000
0!
0'
#812620000000
1!
b111 %
1'
b111 +
#812630000000
0!
0'
#812640000000
1!
0$
b1000 %
1'
0*
b1000 +
#812650000000
0!
0'
#812660000000
1!
b1001 %
1'
b1001 +
#812670000000
0!
0'
#812680000000
1!
b0 %
1'
b0 +
#812690000000
0!
0'
#812700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#812710000000
0!
0'
#812720000000
1!
b10 %
1'
b10 +
#812730000000
0!
0'
#812740000000
1!
b11 %
1'
b11 +
#812750000000
0!
0'
#812760000000
1!
b100 %
1'
b100 +
#812770000000
0!
0'
#812780000000
1!
b101 %
1'
b101 +
#812790000000
0!
0'
#812800000000
1!
0$
b110 %
1'
0*
b110 +
#812810000000
0!
0'
#812820000000
1!
b111 %
1'
b111 +
#812830000000
0!
0'
#812840000000
1!
b1000 %
1'
b1000 +
#812850000000
0!
0'
#812860000000
1!
b1001 %
1'
b1001 +
#812870000000
0!
0'
#812880000000
1!
b0 %
1'
b0 +
#812890000000
0!
0'
#812900000000
1!
1$
b1 %
1'
1*
b1 +
#812910000000
1"
1(
#812920000000
0!
0"
b100 &
0'
0(
b100 ,
#812930000000
1!
b10 %
1'
b10 +
#812940000000
0!
0'
#812950000000
1!
b11 %
1'
b11 +
#812960000000
0!
0'
#812970000000
1!
b100 %
1'
b100 +
#812980000000
0!
0'
#812990000000
1!
b101 %
1'
b101 +
#813000000000
0!
0'
#813010000000
1!
b110 %
1'
b110 +
#813020000000
0!
0'
#813030000000
1!
b111 %
1'
b111 +
#813040000000
0!
0'
#813050000000
1!
0$
b1000 %
1'
0*
b1000 +
#813060000000
0!
0'
#813070000000
1!
b1001 %
1'
b1001 +
#813080000000
0!
0'
#813090000000
1!
b0 %
1'
b0 +
#813100000000
0!
0'
#813110000000
1!
1$
b1 %
1'
1*
b1 +
#813120000000
0!
0'
#813130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#813140000000
0!
0'
#813150000000
1!
b11 %
1'
b11 +
#813160000000
0!
0'
#813170000000
1!
b100 %
1'
b100 +
#813180000000
0!
0'
#813190000000
1!
b101 %
1'
b101 +
#813200000000
0!
0'
#813210000000
1!
0$
b110 %
1'
0*
b110 +
#813220000000
0!
0'
#813230000000
1!
b111 %
1'
b111 +
#813240000000
0!
0'
#813250000000
1!
b1000 %
1'
b1000 +
#813260000000
0!
0'
#813270000000
1!
b1001 %
1'
b1001 +
#813280000000
0!
0'
#813290000000
1!
b0 %
1'
b0 +
#813300000000
0!
0'
#813310000000
1!
1$
b1 %
1'
1*
b1 +
#813320000000
0!
0'
#813330000000
1!
b10 %
1'
b10 +
#813340000000
1"
1(
#813350000000
0!
0"
b100 &
0'
0(
b100 ,
#813360000000
1!
b11 %
1'
b11 +
#813370000000
0!
0'
#813380000000
1!
b100 %
1'
b100 +
#813390000000
0!
0'
#813400000000
1!
b101 %
1'
b101 +
#813410000000
0!
0'
#813420000000
1!
b110 %
1'
b110 +
#813430000000
0!
0'
#813440000000
1!
b111 %
1'
b111 +
#813450000000
0!
0'
#813460000000
1!
0$
b1000 %
1'
0*
b1000 +
#813470000000
0!
0'
#813480000000
1!
b1001 %
1'
b1001 +
#813490000000
0!
0'
#813500000000
1!
b0 %
1'
b0 +
#813510000000
0!
0'
#813520000000
1!
1$
b1 %
1'
1*
b1 +
#813530000000
0!
0'
#813540000000
1!
b10 %
1'
b10 +
#813550000000
0!
0'
#813560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#813570000000
0!
0'
#813580000000
1!
b100 %
1'
b100 +
#813590000000
0!
0'
#813600000000
1!
b101 %
1'
b101 +
#813610000000
0!
0'
#813620000000
1!
0$
b110 %
1'
0*
b110 +
#813630000000
0!
0'
#813640000000
1!
b111 %
1'
b111 +
#813650000000
0!
0'
#813660000000
1!
b1000 %
1'
b1000 +
#813670000000
0!
0'
#813680000000
1!
b1001 %
1'
b1001 +
#813690000000
0!
0'
#813700000000
1!
b0 %
1'
b0 +
#813710000000
0!
0'
#813720000000
1!
1$
b1 %
1'
1*
b1 +
#813730000000
0!
0'
#813740000000
1!
b10 %
1'
b10 +
#813750000000
0!
0'
#813760000000
1!
b11 %
1'
b11 +
#813770000000
1"
1(
#813780000000
0!
0"
b100 &
0'
0(
b100 ,
#813790000000
1!
b100 %
1'
b100 +
#813800000000
0!
0'
#813810000000
1!
b101 %
1'
b101 +
#813820000000
0!
0'
#813830000000
1!
b110 %
1'
b110 +
#813840000000
0!
0'
#813850000000
1!
b111 %
1'
b111 +
#813860000000
0!
0'
#813870000000
1!
0$
b1000 %
1'
0*
b1000 +
#813880000000
0!
0'
#813890000000
1!
b1001 %
1'
b1001 +
#813900000000
0!
0'
#813910000000
1!
b0 %
1'
b0 +
#813920000000
0!
0'
#813930000000
1!
1$
b1 %
1'
1*
b1 +
#813940000000
0!
0'
#813950000000
1!
b10 %
1'
b10 +
#813960000000
0!
0'
#813970000000
1!
b11 %
1'
b11 +
#813980000000
0!
0'
#813990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#814000000000
0!
0'
#814010000000
1!
b101 %
1'
b101 +
#814020000000
0!
0'
#814030000000
1!
0$
b110 %
1'
0*
b110 +
#814040000000
0!
0'
#814050000000
1!
b111 %
1'
b111 +
#814060000000
0!
0'
#814070000000
1!
b1000 %
1'
b1000 +
#814080000000
0!
0'
#814090000000
1!
b1001 %
1'
b1001 +
#814100000000
0!
0'
#814110000000
1!
b0 %
1'
b0 +
#814120000000
0!
0'
#814130000000
1!
1$
b1 %
1'
1*
b1 +
#814140000000
0!
0'
#814150000000
1!
b10 %
1'
b10 +
#814160000000
0!
0'
#814170000000
1!
b11 %
1'
b11 +
#814180000000
0!
0'
#814190000000
1!
b100 %
1'
b100 +
#814200000000
1"
1(
#814210000000
0!
0"
b100 &
0'
0(
b100 ,
#814220000000
1!
b101 %
1'
b101 +
#814230000000
0!
0'
#814240000000
1!
b110 %
1'
b110 +
#814250000000
0!
0'
#814260000000
1!
b111 %
1'
b111 +
#814270000000
0!
0'
#814280000000
1!
0$
b1000 %
1'
0*
b1000 +
#814290000000
0!
0'
#814300000000
1!
b1001 %
1'
b1001 +
#814310000000
0!
0'
#814320000000
1!
b0 %
1'
b0 +
#814330000000
0!
0'
#814340000000
1!
1$
b1 %
1'
1*
b1 +
#814350000000
0!
0'
#814360000000
1!
b10 %
1'
b10 +
#814370000000
0!
0'
#814380000000
1!
b11 %
1'
b11 +
#814390000000
0!
0'
#814400000000
1!
b100 %
1'
b100 +
#814410000000
0!
0'
#814420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#814430000000
0!
0'
#814440000000
1!
0$
b110 %
1'
0*
b110 +
#814450000000
0!
0'
#814460000000
1!
b111 %
1'
b111 +
#814470000000
0!
0'
#814480000000
1!
b1000 %
1'
b1000 +
#814490000000
0!
0'
#814500000000
1!
b1001 %
1'
b1001 +
#814510000000
0!
0'
#814520000000
1!
b0 %
1'
b0 +
#814530000000
0!
0'
#814540000000
1!
1$
b1 %
1'
1*
b1 +
#814550000000
0!
0'
#814560000000
1!
b10 %
1'
b10 +
#814570000000
0!
0'
#814580000000
1!
b11 %
1'
b11 +
#814590000000
0!
0'
#814600000000
1!
b100 %
1'
b100 +
#814610000000
0!
0'
#814620000000
1!
b101 %
1'
b101 +
#814630000000
1"
1(
#814640000000
0!
0"
b100 &
0'
0(
b100 ,
#814650000000
1!
b110 %
1'
b110 +
#814660000000
0!
0'
#814670000000
1!
b111 %
1'
b111 +
#814680000000
0!
0'
#814690000000
1!
0$
b1000 %
1'
0*
b1000 +
#814700000000
0!
0'
#814710000000
1!
b1001 %
1'
b1001 +
#814720000000
0!
0'
#814730000000
1!
b0 %
1'
b0 +
#814740000000
0!
0'
#814750000000
1!
1$
b1 %
1'
1*
b1 +
#814760000000
0!
0'
#814770000000
1!
b10 %
1'
b10 +
#814780000000
0!
0'
#814790000000
1!
b11 %
1'
b11 +
#814800000000
0!
0'
#814810000000
1!
b100 %
1'
b100 +
#814820000000
0!
0'
#814830000000
1!
b101 %
1'
b101 +
#814840000000
0!
0'
#814850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#814860000000
0!
0'
#814870000000
1!
b111 %
1'
b111 +
#814880000000
0!
0'
#814890000000
1!
b1000 %
1'
b1000 +
#814900000000
0!
0'
#814910000000
1!
b1001 %
1'
b1001 +
#814920000000
0!
0'
#814930000000
1!
b0 %
1'
b0 +
#814940000000
0!
0'
#814950000000
1!
1$
b1 %
1'
1*
b1 +
#814960000000
0!
0'
#814970000000
1!
b10 %
1'
b10 +
#814980000000
0!
0'
#814990000000
1!
b11 %
1'
b11 +
#815000000000
0!
0'
#815010000000
1!
b100 %
1'
b100 +
#815020000000
0!
0'
#815030000000
1!
b101 %
1'
b101 +
#815040000000
0!
0'
#815050000000
1!
0$
b110 %
1'
0*
b110 +
#815060000000
1"
1(
#815070000000
0!
0"
b100 &
0'
0(
b100 ,
#815080000000
1!
1$
b111 %
1'
1*
b111 +
#815090000000
0!
0'
#815100000000
1!
0$
b1000 %
1'
0*
b1000 +
#815110000000
0!
0'
#815120000000
1!
b1001 %
1'
b1001 +
#815130000000
0!
0'
#815140000000
1!
b0 %
1'
b0 +
#815150000000
0!
0'
#815160000000
1!
1$
b1 %
1'
1*
b1 +
#815170000000
0!
0'
#815180000000
1!
b10 %
1'
b10 +
#815190000000
0!
0'
#815200000000
1!
b11 %
1'
b11 +
#815210000000
0!
0'
#815220000000
1!
b100 %
1'
b100 +
#815230000000
0!
0'
#815240000000
1!
b101 %
1'
b101 +
#815250000000
0!
0'
#815260000000
1!
b110 %
1'
b110 +
#815270000000
0!
0'
#815280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#815290000000
0!
0'
#815300000000
1!
b1000 %
1'
b1000 +
#815310000000
0!
0'
#815320000000
1!
b1001 %
1'
b1001 +
#815330000000
0!
0'
#815340000000
1!
b0 %
1'
b0 +
#815350000000
0!
0'
#815360000000
1!
1$
b1 %
1'
1*
b1 +
#815370000000
0!
0'
#815380000000
1!
b10 %
1'
b10 +
#815390000000
0!
0'
#815400000000
1!
b11 %
1'
b11 +
#815410000000
0!
0'
#815420000000
1!
b100 %
1'
b100 +
#815430000000
0!
0'
#815440000000
1!
b101 %
1'
b101 +
#815450000000
0!
0'
#815460000000
1!
0$
b110 %
1'
0*
b110 +
#815470000000
0!
0'
#815480000000
1!
b111 %
1'
b111 +
#815490000000
1"
1(
#815500000000
0!
0"
b100 &
0'
0(
b100 ,
#815510000000
1!
b1000 %
1'
b1000 +
#815520000000
0!
0'
#815530000000
1!
b1001 %
1'
b1001 +
#815540000000
0!
0'
#815550000000
1!
b0 %
1'
b0 +
#815560000000
0!
0'
#815570000000
1!
1$
b1 %
1'
1*
b1 +
#815580000000
0!
0'
#815590000000
1!
b10 %
1'
b10 +
#815600000000
0!
0'
#815610000000
1!
b11 %
1'
b11 +
#815620000000
0!
0'
#815630000000
1!
b100 %
1'
b100 +
#815640000000
0!
0'
#815650000000
1!
b101 %
1'
b101 +
#815660000000
0!
0'
#815670000000
1!
b110 %
1'
b110 +
#815680000000
0!
0'
#815690000000
1!
b111 %
1'
b111 +
#815700000000
0!
0'
#815710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#815720000000
0!
0'
#815730000000
1!
b1001 %
1'
b1001 +
#815740000000
0!
0'
#815750000000
1!
b0 %
1'
b0 +
#815760000000
0!
0'
#815770000000
1!
1$
b1 %
1'
1*
b1 +
#815780000000
0!
0'
#815790000000
1!
b10 %
1'
b10 +
#815800000000
0!
0'
#815810000000
1!
b11 %
1'
b11 +
#815820000000
0!
0'
#815830000000
1!
b100 %
1'
b100 +
#815840000000
0!
0'
#815850000000
1!
b101 %
1'
b101 +
#815860000000
0!
0'
#815870000000
1!
0$
b110 %
1'
0*
b110 +
#815880000000
0!
0'
#815890000000
1!
b111 %
1'
b111 +
#815900000000
0!
0'
#815910000000
1!
b1000 %
1'
b1000 +
#815920000000
1"
1(
#815930000000
0!
0"
b100 &
0'
0(
b100 ,
#815940000000
1!
b1001 %
1'
b1001 +
#815950000000
0!
0'
#815960000000
1!
b0 %
1'
b0 +
#815970000000
0!
0'
#815980000000
1!
1$
b1 %
1'
1*
b1 +
#815990000000
0!
0'
#816000000000
1!
b10 %
1'
b10 +
#816010000000
0!
0'
#816020000000
1!
b11 %
1'
b11 +
#816030000000
0!
0'
#816040000000
1!
b100 %
1'
b100 +
#816050000000
0!
0'
#816060000000
1!
b101 %
1'
b101 +
#816070000000
0!
0'
#816080000000
1!
b110 %
1'
b110 +
#816090000000
0!
0'
#816100000000
1!
b111 %
1'
b111 +
#816110000000
0!
0'
#816120000000
1!
0$
b1000 %
1'
0*
b1000 +
#816130000000
0!
0'
#816140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#816150000000
0!
0'
#816160000000
1!
b0 %
1'
b0 +
#816170000000
0!
0'
#816180000000
1!
1$
b1 %
1'
1*
b1 +
#816190000000
0!
0'
#816200000000
1!
b10 %
1'
b10 +
#816210000000
0!
0'
#816220000000
1!
b11 %
1'
b11 +
#816230000000
0!
0'
#816240000000
1!
b100 %
1'
b100 +
#816250000000
0!
0'
#816260000000
1!
b101 %
1'
b101 +
#816270000000
0!
0'
#816280000000
1!
0$
b110 %
1'
0*
b110 +
#816290000000
0!
0'
#816300000000
1!
b111 %
1'
b111 +
#816310000000
0!
0'
#816320000000
1!
b1000 %
1'
b1000 +
#816330000000
0!
0'
#816340000000
1!
b1001 %
1'
b1001 +
#816350000000
1"
1(
#816360000000
0!
0"
b100 &
0'
0(
b100 ,
#816370000000
1!
b0 %
1'
b0 +
#816380000000
0!
0'
#816390000000
1!
1$
b1 %
1'
1*
b1 +
#816400000000
0!
0'
#816410000000
1!
b10 %
1'
b10 +
#816420000000
0!
0'
#816430000000
1!
b11 %
1'
b11 +
#816440000000
0!
0'
#816450000000
1!
b100 %
1'
b100 +
#816460000000
0!
0'
#816470000000
1!
b101 %
1'
b101 +
#816480000000
0!
0'
#816490000000
1!
b110 %
1'
b110 +
#816500000000
0!
0'
#816510000000
1!
b111 %
1'
b111 +
#816520000000
0!
0'
#816530000000
1!
0$
b1000 %
1'
0*
b1000 +
#816540000000
0!
0'
#816550000000
1!
b1001 %
1'
b1001 +
#816560000000
0!
0'
#816570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#816580000000
0!
0'
#816590000000
1!
1$
b1 %
1'
1*
b1 +
#816600000000
0!
0'
#816610000000
1!
b10 %
1'
b10 +
#816620000000
0!
0'
#816630000000
1!
b11 %
1'
b11 +
#816640000000
0!
0'
#816650000000
1!
b100 %
1'
b100 +
#816660000000
0!
0'
#816670000000
1!
b101 %
1'
b101 +
#816680000000
0!
0'
#816690000000
1!
0$
b110 %
1'
0*
b110 +
#816700000000
0!
0'
#816710000000
1!
b111 %
1'
b111 +
#816720000000
0!
0'
#816730000000
1!
b1000 %
1'
b1000 +
#816740000000
0!
0'
#816750000000
1!
b1001 %
1'
b1001 +
#816760000000
0!
0'
#816770000000
1!
b0 %
1'
b0 +
#816780000000
1"
1(
#816790000000
0!
0"
b100 &
0'
0(
b100 ,
#816800000000
1!
1$
b1 %
1'
1*
b1 +
#816810000000
0!
0'
#816820000000
1!
b10 %
1'
b10 +
#816830000000
0!
0'
#816840000000
1!
b11 %
1'
b11 +
#816850000000
0!
0'
#816860000000
1!
b100 %
1'
b100 +
#816870000000
0!
0'
#816880000000
1!
b101 %
1'
b101 +
#816890000000
0!
0'
#816900000000
1!
b110 %
1'
b110 +
#816910000000
0!
0'
#816920000000
1!
b111 %
1'
b111 +
#816930000000
0!
0'
#816940000000
1!
0$
b1000 %
1'
0*
b1000 +
#816950000000
0!
0'
#816960000000
1!
b1001 %
1'
b1001 +
#816970000000
0!
0'
#816980000000
1!
b0 %
1'
b0 +
#816990000000
0!
0'
#817000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#817010000000
0!
0'
#817020000000
1!
b10 %
1'
b10 +
#817030000000
0!
0'
#817040000000
1!
b11 %
1'
b11 +
#817050000000
0!
0'
#817060000000
1!
b100 %
1'
b100 +
#817070000000
0!
0'
#817080000000
1!
b101 %
1'
b101 +
#817090000000
0!
0'
#817100000000
1!
0$
b110 %
1'
0*
b110 +
#817110000000
0!
0'
#817120000000
1!
b111 %
1'
b111 +
#817130000000
0!
0'
#817140000000
1!
b1000 %
1'
b1000 +
#817150000000
0!
0'
#817160000000
1!
b1001 %
1'
b1001 +
#817170000000
0!
0'
#817180000000
1!
b0 %
1'
b0 +
#817190000000
0!
0'
#817200000000
1!
1$
b1 %
1'
1*
b1 +
#817210000000
1"
1(
#817220000000
0!
0"
b100 &
0'
0(
b100 ,
#817230000000
1!
b10 %
1'
b10 +
#817240000000
0!
0'
#817250000000
1!
b11 %
1'
b11 +
#817260000000
0!
0'
#817270000000
1!
b100 %
1'
b100 +
#817280000000
0!
0'
#817290000000
1!
b101 %
1'
b101 +
#817300000000
0!
0'
#817310000000
1!
b110 %
1'
b110 +
#817320000000
0!
0'
#817330000000
1!
b111 %
1'
b111 +
#817340000000
0!
0'
#817350000000
1!
0$
b1000 %
1'
0*
b1000 +
#817360000000
0!
0'
#817370000000
1!
b1001 %
1'
b1001 +
#817380000000
0!
0'
#817390000000
1!
b0 %
1'
b0 +
#817400000000
0!
0'
#817410000000
1!
1$
b1 %
1'
1*
b1 +
#817420000000
0!
0'
#817430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#817440000000
0!
0'
#817450000000
1!
b11 %
1'
b11 +
#817460000000
0!
0'
#817470000000
1!
b100 %
1'
b100 +
#817480000000
0!
0'
#817490000000
1!
b101 %
1'
b101 +
#817500000000
0!
0'
#817510000000
1!
0$
b110 %
1'
0*
b110 +
#817520000000
0!
0'
#817530000000
1!
b111 %
1'
b111 +
#817540000000
0!
0'
#817550000000
1!
b1000 %
1'
b1000 +
#817560000000
0!
0'
#817570000000
1!
b1001 %
1'
b1001 +
#817580000000
0!
0'
#817590000000
1!
b0 %
1'
b0 +
#817600000000
0!
0'
#817610000000
1!
1$
b1 %
1'
1*
b1 +
#817620000000
0!
0'
#817630000000
1!
b10 %
1'
b10 +
#817640000000
1"
1(
#817650000000
0!
0"
b100 &
0'
0(
b100 ,
#817660000000
1!
b11 %
1'
b11 +
#817670000000
0!
0'
#817680000000
1!
b100 %
1'
b100 +
#817690000000
0!
0'
#817700000000
1!
b101 %
1'
b101 +
#817710000000
0!
0'
#817720000000
1!
b110 %
1'
b110 +
#817730000000
0!
0'
#817740000000
1!
b111 %
1'
b111 +
#817750000000
0!
0'
#817760000000
1!
0$
b1000 %
1'
0*
b1000 +
#817770000000
0!
0'
#817780000000
1!
b1001 %
1'
b1001 +
#817790000000
0!
0'
#817800000000
1!
b0 %
1'
b0 +
#817810000000
0!
0'
#817820000000
1!
1$
b1 %
1'
1*
b1 +
#817830000000
0!
0'
#817840000000
1!
b10 %
1'
b10 +
#817850000000
0!
0'
#817860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#817870000000
0!
0'
#817880000000
1!
b100 %
1'
b100 +
#817890000000
0!
0'
#817900000000
1!
b101 %
1'
b101 +
#817910000000
0!
0'
#817920000000
1!
0$
b110 %
1'
0*
b110 +
#817930000000
0!
0'
#817940000000
1!
b111 %
1'
b111 +
#817950000000
0!
0'
#817960000000
1!
b1000 %
1'
b1000 +
#817970000000
0!
0'
#817980000000
1!
b1001 %
1'
b1001 +
#817990000000
0!
0'
#818000000000
1!
b0 %
1'
b0 +
#818010000000
0!
0'
#818020000000
1!
1$
b1 %
1'
1*
b1 +
#818030000000
0!
0'
#818040000000
1!
b10 %
1'
b10 +
#818050000000
0!
0'
#818060000000
1!
b11 %
1'
b11 +
#818070000000
1"
1(
#818080000000
0!
0"
b100 &
0'
0(
b100 ,
#818090000000
1!
b100 %
1'
b100 +
#818100000000
0!
0'
#818110000000
1!
b101 %
1'
b101 +
#818120000000
0!
0'
#818130000000
1!
b110 %
1'
b110 +
#818140000000
0!
0'
#818150000000
1!
b111 %
1'
b111 +
#818160000000
0!
0'
#818170000000
1!
0$
b1000 %
1'
0*
b1000 +
#818180000000
0!
0'
#818190000000
1!
b1001 %
1'
b1001 +
#818200000000
0!
0'
#818210000000
1!
b0 %
1'
b0 +
#818220000000
0!
0'
#818230000000
1!
1$
b1 %
1'
1*
b1 +
#818240000000
0!
0'
#818250000000
1!
b10 %
1'
b10 +
#818260000000
0!
0'
#818270000000
1!
b11 %
1'
b11 +
#818280000000
0!
0'
#818290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#818300000000
0!
0'
#818310000000
1!
b101 %
1'
b101 +
#818320000000
0!
0'
#818330000000
1!
0$
b110 %
1'
0*
b110 +
#818340000000
0!
0'
#818350000000
1!
b111 %
1'
b111 +
#818360000000
0!
0'
#818370000000
1!
b1000 %
1'
b1000 +
#818380000000
0!
0'
#818390000000
1!
b1001 %
1'
b1001 +
#818400000000
0!
0'
#818410000000
1!
b0 %
1'
b0 +
#818420000000
0!
0'
#818430000000
1!
1$
b1 %
1'
1*
b1 +
#818440000000
0!
0'
#818450000000
1!
b10 %
1'
b10 +
#818460000000
0!
0'
#818470000000
1!
b11 %
1'
b11 +
#818480000000
0!
0'
#818490000000
1!
b100 %
1'
b100 +
#818500000000
1"
1(
#818510000000
0!
0"
b100 &
0'
0(
b100 ,
#818520000000
1!
b101 %
1'
b101 +
#818530000000
0!
0'
#818540000000
1!
b110 %
1'
b110 +
#818550000000
0!
0'
#818560000000
1!
b111 %
1'
b111 +
#818570000000
0!
0'
#818580000000
1!
0$
b1000 %
1'
0*
b1000 +
#818590000000
0!
0'
#818600000000
1!
b1001 %
1'
b1001 +
#818610000000
0!
0'
#818620000000
1!
b0 %
1'
b0 +
#818630000000
0!
0'
#818640000000
1!
1$
b1 %
1'
1*
b1 +
#818650000000
0!
0'
#818660000000
1!
b10 %
1'
b10 +
#818670000000
0!
0'
#818680000000
1!
b11 %
1'
b11 +
#818690000000
0!
0'
#818700000000
1!
b100 %
1'
b100 +
#818710000000
0!
0'
#818720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#818730000000
0!
0'
#818740000000
1!
0$
b110 %
1'
0*
b110 +
#818750000000
0!
0'
#818760000000
1!
b111 %
1'
b111 +
#818770000000
0!
0'
#818780000000
1!
b1000 %
1'
b1000 +
#818790000000
0!
0'
#818800000000
1!
b1001 %
1'
b1001 +
#818810000000
0!
0'
#818820000000
1!
b0 %
1'
b0 +
#818830000000
0!
0'
#818840000000
1!
1$
b1 %
1'
1*
b1 +
#818850000000
0!
0'
#818860000000
1!
b10 %
1'
b10 +
#818870000000
0!
0'
#818880000000
1!
b11 %
1'
b11 +
#818890000000
0!
0'
#818900000000
1!
b100 %
1'
b100 +
#818910000000
0!
0'
#818920000000
1!
b101 %
1'
b101 +
#818930000000
1"
1(
#818940000000
0!
0"
b100 &
0'
0(
b100 ,
#818950000000
1!
b110 %
1'
b110 +
#818960000000
0!
0'
#818970000000
1!
b111 %
1'
b111 +
#818980000000
0!
0'
#818990000000
1!
0$
b1000 %
1'
0*
b1000 +
#819000000000
0!
0'
#819010000000
1!
b1001 %
1'
b1001 +
#819020000000
0!
0'
#819030000000
1!
b0 %
1'
b0 +
#819040000000
0!
0'
#819050000000
1!
1$
b1 %
1'
1*
b1 +
#819060000000
0!
0'
#819070000000
1!
b10 %
1'
b10 +
#819080000000
0!
0'
#819090000000
1!
b11 %
1'
b11 +
#819100000000
0!
0'
#819110000000
1!
b100 %
1'
b100 +
#819120000000
0!
0'
#819130000000
1!
b101 %
1'
b101 +
#819140000000
0!
0'
#819150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#819160000000
0!
0'
#819170000000
1!
b111 %
1'
b111 +
#819180000000
0!
0'
#819190000000
1!
b1000 %
1'
b1000 +
#819200000000
0!
0'
#819210000000
1!
b1001 %
1'
b1001 +
#819220000000
0!
0'
#819230000000
1!
b0 %
1'
b0 +
#819240000000
0!
0'
#819250000000
1!
1$
b1 %
1'
1*
b1 +
#819260000000
0!
0'
#819270000000
1!
b10 %
1'
b10 +
#819280000000
0!
0'
#819290000000
1!
b11 %
1'
b11 +
#819300000000
0!
0'
#819310000000
1!
b100 %
1'
b100 +
#819320000000
0!
0'
#819330000000
1!
b101 %
1'
b101 +
#819340000000
0!
0'
#819350000000
1!
0$
b110 %
1'
0*
b110 +
#819360000000
1"
1(
#819370000000
0!
0"
b100 &
0'
0(
b100 ,
#819380000000
1!
1$
b111 %
1'
1*
b111 +
#819390000000
0!
0'
#819400000000
1!
0$
b1000 %
1'
0*
b1000 +
#819410000000
0!
0'
#819420000000
1!
b1001 %
1'
b1001 +
#819430000000
0!
0'
#819440000000
1!
b0 %
1'
b0 +
#819450000000
0!
0'
#819460000000
1!
1$
b1 %
1'
1*
b1 +
#819470000000
0!
0'
#819480000000
1!
b10 %
1'
b10 +
#819490000000
0!
0'
#819500000000
1!
b11 %
1'
b11 +
#819510000000
0!
0'
#819520000000
1!
b100 %
1'
b100 +
#819530000000
0!
0'
#819540000000
1!
b101 %
1'
b101 +
#819550000000
0!
0'
#819560000000
1!
b110 %
1'
b110 +
#819570000000
0!
0'
#819580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#819590000000
0!
0'
#819600000000
1!
b1000 %
1'
b1000 +
#819610000000
0!
0'
#819620000000
1!
b1001 %
1'
b1001 +
#819630000000
0!
0'
#819640000000
1!
b0 %
1'
b0 +
#819650000000
0!
0'
#819660000000
1!
1$
b1 %
1'
1*
b1 +
#819670000000
0!
0'
#819680000000
1!
b10 %
1'
b10 +
#819690000000
0!
0'
#819700000000
1!
b11 %
1'
b11 +
#819710000000
0!
0'
#819720000000
1!
b100 %
1'
b100 +
#819730000000
0!
0'
#819740000000
1!
b101 %
1'
b101 +
#819750000000
0!
0'
#819760000000
1!
0$
b110 %
1'
0*
b110 +
#819770000000
0!
0'
#819780000000
1!
b111 %
1'
b111 +
#819790000000
1"
1(
#819800000000
0!
0"
b100 &
0'
0(
b100 ,
#819810000000
1!
b1000 %
1'
b1000 +
#819820000000
0!
0'
#819830000000
1!
b1001 %
1'
b1001 +
#819840000000
0!
0'
#819850000000
1!
b0 %
1'
b0 +
#819860000000
0!
0'
#819870000000
1!
1$
b1 %
1'
1*
b1 +
#819880000000
0!
0'
#819890000000
1!
b10 %
1'
b10 +
#819900000000
0!
0'
#819910000000
1!
b11 %
1'
b11 +
#819920000000
0!
0'
#819930000000
1!
b100 %
1'
b100 +
#819940000000
0!
0'
#819950000000
1!
b101 %
1'
b101 +
#819960000000
0!
0'
#819970000000
1!
b110 %
1'
b110 +
#819980000000
0!
0'
#819990000000
1!
b111 %
1'
b111 +
#820000000000
0!
0'
#820010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#820020000000
0!
0'
#820030000000
1!
b1001 %
1'
b1001 +
#820040000000
0!
0'
#820050000000
1!
b0 %
1'
b0 +
#820060000000
0!
0'
#820070000000
1!
1$
b1 %
1'
1*
b1 +
#820080000000
0!
0'
#820090000000
1!
b10 %
1'
b10 +
#820100000000
0!
0'
#820110000000
1!
b11 %
1'
b11 +
#820120000000
0!
0'
#820130000000
1!
b100 %
1'
b100 +
#820140000000
0!
0'
#820150000000
1!
b101 %
1'
b101 +
#820160000000
0!
0'
#820170000000
1!
0$
b110 %
1'
0*
b110 +
#820180000000
0!
0'
#820190000000
1!
b111 %
1'
b111 +
#820200000000
0!
0'
#820210000000
1!
b1000 %
1'
b1000 +
#820220000000
1"
1(
#820230000000
0!
0"
b100 &
0'
0(
b100 ,
#820240000000
1!
b1001 %
1'
b1001 +
#820250000000
0!
0'
#820260000000
1!
b0 %
1'
b0 +
#820270000000
0!
0'
#820280000000
1!
1$
b1 %
1'
1*
b1 +
#820290000000
0!
0'
#820300000000
1!
b10 %
1'
b10 +
#820310000000
0!
0'
#820320000000
1!
b11 %
1'
b11 +
#820330000000
0!
0'
#820340000000
1!
b100 %
1'
b100 +
#820350000000
0!
0'
#820360000000
1!
b101 %
1'
b101 +
#820370000000
0!
0'
#820380000000
1!
b110 %
1'
b110 +
#820390000000
0!
0'
#820400000000
1!
b111 %
1'
b111 +
#820410000000
0!
0'
#820420000000
1!
0$
b1000 %
1'
0*
b1000 +
#820430000000
0!
0'
#820440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#820450000000
0!
0'
#820460000000
1!
b0 %
1'
b0 +
#820470000000
0!
0'
#820480000000
1!
1$
b1 %
1'
1*
b1 +
#820490000000
0!
0'
#820500000000
1!
b10 %
1'
b10 +
#820510000000
0!
0'
#820520000000
1!
b11 %
1'
b11 +
#820530000000
0!
0'
#820540000000
1!
b100 %
1'
b100 +
#820550000000
0!
0'
#820560000000
1!
b101 %
1'
b101 +
#820570000000
0!
0'
#820580000000
1!
0$
b110 %
1'
0*
b110 +
#820590000000
0!
0'
#820600000000
1!
b111 %
1'
b111 +
#820610000000
0!
0'
#820620000000
1!
b1000 %
1'
b1000 +
#820630000000
0!
0'
#820640000000
1!
b1001 %
1'
b1001 +
#820650000000
1"
1(
#820660000000
0!
0"
b100 &
0'
0(
b100 ,
#820670000000
1!
b0 %
1'
b0 +
#820680000000
0!
0'
#820690000000
1!
1$
b1 %
1'
1*
b1 +
#820700000000
0!
0'
#820710000000
1!
b10 %
1'
b10 +
#820720000000
0!
0'
#820730000000
1!
b11 %
1'
b11 +
#820740000000
0!
0'
#820750000000
1!
b100 %
1'
b100 +
#820760000000
0!
0'
#820770000000
1!
b101 %
1'
b101 +
#820780000000
0!
0'
#820790000000
1!
b110 %
1'
b110 +
#820800000000
0!
0'
#820810000000
1!
b111 %
1'
b111 +
#820820000000
0!
0'
#820830000000
1!
0$
b1000 %
1'
0*
b1000 +
#820840000000
0!
0'
#820850000000
1!
b1001 %
1'
b1001 +
#820860000000
0!
0'
#820870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#820880000000
0!
0'
#820890000000
1!
1$
b1 %
1'
1*
b1 +
#820900000000
0!
0'
#820910000000
1!
b10 %
1'
b10 +
#820920000000
0!
0'
#820930000000
1!
b11 %
1'
b11 +
#820940000000
0!
0'
#820950000000
1!
b100 %
1'
b100 +
#820960000000
0!
0'
#820970000000
1!
b101 %
1'
b101 +
#820980000000
0!
0'
#820990000000
1!
0$
b110 %
1'
0*
b110 +
#821000000000
0!
0'
#821010000000
1!
b111 %
1'
b111 +
#821020000000
0!
0'
#821030000000
1!
b1000 %
1'
b1000 +
#821040000000
0!
0'
#821050000000
1!
b1001 %
1'
b1001 +
#821060000000
0!
0'
#821070000000
1!
b0 %
1'
b0 +
#821080000000
1"
1(
#821090000000
0!
0"
b100 &
0'
0(
b100 ,
#821100000000
1!
1$
b1 %
1'
1*
b1 +
#821110000000
0!
0'
#821120000000
1!
b10 %
1'
b10 +
#821130000000
0!
0'
#821140000000
1!
b11 %
1'
b11 +
#821150000000
0!
0'
#821160000000
1!
b100 %
1'
b100 +
#821170000000
0!
0'
#821180000000
1!
b101 %
1'
b101 +
#821190000000
0!
0'
#821200000000
1!
b110 %
1'
b110 +
#821210000000
0!
0'
#821220000000
1!
b111 %
1'
b111 +
#821230000000
0!
0'
#821240000000
1!
0$
b1000 %
1'
0*
b1000 +
#821250000000
0!
0'
#821260000000
1!
b1001 %
1'
b1001 +
#821270000000
0!
0'
#821280000000
1!
b0 %
1'
b0 +
#821290000000
0!
0'
#821300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#821310000000
0!
0'
#821320000000
1!
b10 %
1'
b10 +
#821330000000
0!
0'
#821340000000
1!
b11 %
1'
b11 +
#821350000000
0!
0'
#821360000000
1!
b100 %
1'
b100 +
#821370000000
0!
0'
#821380000000
1!
b101 %
1'
b101 +
#821390000000
0!
0'
#821400000000
1!
0$
b110 %
1'
0*
b110 +
#821410000000
0!
0'
#821420000000
1!
b111 %
1'
b111 +
#821430000000
0!
0'
#821440000000
1!
b1000 %
1'
b1000 +
#821450000000
0!
0'
#821460000000
1!
b1001 %
1'
b1001 +
#821470000000
0!
0'
#821480000000
1!
b0 %
1'
b0 +
#821490000000
0!
0'
#821500000000
1!
1$
b1 %
1'
1*
b1 +
#821510000000
1"
1(
#821520000000
0!
0"
b100 &
0'
0(
b100 ,
#821530000000
1!
b10 %
1'
b10 +
#821540000000
0!
0'
#821550000000
1!
b11 %
1'
b11 +
#821560000000
0!
0'
#821570000000
1!
b100 %
1'
b100 +
#821580000000
0!
0'
#821590000000
1!
b101 %
1'
b101 +
#821600000000
0!
0'
#821610000000
1!
b110 %
1'
b110 +
#821620000000
0!
0'
#821630000000
1!
b111 %
1'
b111 +
#821640000000
0!
0'
#821650000000
1!
0$
b1000 %
1'
0*
b1000 +
#821660000000
0!
0'
#821670000000
1!
b1001 %
1'
b1001 +
#821680000000
0!
0'
#821690000000
1!
b0 %
1'
b0 +
#821700000000
0!
0'
#821710000000
1!
1$
b1 %
1'
1*
b1 +
#821720000000
0!
0'
#821730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#821740000000
0!
0'
#821750000000
1!
b11 %
1'
b11 +
#821760000000
0!
0'
#821770000000
1!
b100 %
1'
b100 +
#821780000000
0!
0'
#821790000000
1!
b101 %
1'
b101 +
#821800000000
0!
0'
#821810000000
1!
0$
b110 %
1'
0*
b110 +
#821820000000
0!
0'
#821830000000
1!
b111 %
1'
b111 +
#821840000000
0!
0'
#821850000000
1!
b1000 %
1'
b1000 +
#821860000000
0!
0'
#821870000000
1!
b1001 %
1'
b1001 +
#821880000000
0!
0'
#821890000000
1!
b0 %
1'
b0 +
#821900000000
0!
0'
#821910000000
1!
1$
b1 %
1'
1*
b1 +
#821920000000
0!
0'
#821930000000
1!
b10 %
1'
b10 +
#821940000000
1"
1(
#821950000000
0!
0"
b100 &
0'
0(
b100 ,
#821960000000
1!
b11 %
1'
b11 +
#821970000000
0!
0'
#821980000000
1!
b100 %
1'
b100 +
#821990000000
0!
0'
#822000000000
1!
b101 %
1'
b101 +
#822010000000
0!
0'
#822020000000
1!
b110 %
1'
b110 +
#822030000000
0!
0'
#822040000000
1!
b111 %
1'
b111 +
#822050000000
0!
0'
#822060000000
1!
0$
b1000 %
1'
0*
b1000 +
#822070000000
0!
0'
#822080000000
1!
b1001 %
1'
b1001 +
#822090000000
0!
0'
#822100000000
1!
b0 %
1'
b0 +
#822110000000
0!
0'
#822120000000
1!
1$
b1 %
1'
1*
b1 +
#822130000000
0!
0'
#822140000000
1!
b10 %
1'
b10 +
#822150000000
0!
0'
#822160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#822170000000
0!
0'
#822180000000
1!
b100 %
1'
b100 +
#822190000000
0!
0'
#822200000000
1!
b101 %
1'
b101 +
#822210000000
0!
0'
#822220000000
1!
0$
b110 %
1'
0*
b110 +
#822230000000
0!
0'
#822240000000
1!
b111 %
1'
b111 +
#822250000000
0!
0'
#822260000000
1!
b1000 %
1'
b1000 +
#822270000000
0!
0'
#822280000000
1!
b1001 %
1'
b1001 +
#822290000000
0!
0'
#822300000000
1!
b0 %
1'
b0 +
#822310000000
0!
0'
#822320000000
1!
1$
b1 %
1'
1*
b1 +
#822330000000
0!
0'
#822340000000
1!
b10 %
1'
b10 +
#822350000000
0!
0'
#822360000000
1!
b11 %
1'
b11 +
#822370000000
1"
1(
#822380000000
0!
0"
b100 &
0'
0(
b100 ,
#822390000000
1!
b100 %
1'
b100 +
#822400000000
0!
0'
#822410000000
1!
b101 %
1'
b101 +
#822420000000
0!
0'
#822430000000
1!
b110 %
1'
b110 +
#822440000000
0!
0'
#822450000000
1!
b111 %
1'
b111 +
#822460000000
0!
0'
#822470000000
1!
0$
b1000 %
1'
0*
b1000 +
#822480000000
0!
0'
#822490000000
1!
b1001 %
1'
b1001 +
#822500000000
0!
0'
#822510000000
1!
b0 %
1'
b0 +
#822520000000
0!
0'
#822530000000
1!
1$
b1 %
1'
1*
b1 +
#822540000000
0!
0'
#822550000000
1!
b10 %
1'
b10 +
#822560000000
0!
0'
#822570000000
1!
b11 %
1'
b11 +
#822580000000
0!
0'
#822590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#822600000000
0!
0'
#822610000000
1!
b101 %
1'
b101 +
#822620000000
0!
0'
#822630000000
1!
0$
b110 %
1'
0*
b110 +
#822640000000
0!
0'
#822650000000
1!
b111 %
1'
b111 +
#822660000000
0!
0'
#822670000000
1!
b1000 %
1'
b1000 +
#822680000000
0!
0'
#822690000000
1!
b1001 %
1'
b1001 +
#822700000000
0!
0'
#822710000000
1!
b0 %
1'
b0 +
#822720000000
0!
0'
#822730000000
1!
1$
b1 %
1'
1*
b1 +
#822740000000
0!
0'
#822750000000
1!
b10 %
1'
b10 +
#822760000000
0!
0'
#822770000000
1!
b11 %
1'
b11 +
#822780000000
0!
0'
#822790000000
1!
b100 %
1'
b100 +
#822800000000
1"
1(
#822810000000
0!
0"
b100 &
0'
0(
b100 ,
#822820000000
1!
b101 %
1'
b101 +
#822830000000
0!
0'
#822840000000
1!
b110 %
1'
b110 +
#822850000000
0!
0'
#822860000000
1!
b111 %
1'
b111 +
#822870000000
0!
0'
#822880000000
1!
0$
b1000 %
1'
0*
b1000 +
#822890000000
0!
0'
#822900000000
1!
b1001 %
1'
b1001 +
#822910000000
0!
0'
#822920000000
1!
b0 %
1'
b0 +
#822930000000
0!
0'
#822940000000
1!
1$
b1 %
1'
1*
b1 +
#822950000000
0!
0'
#822960000000
1!
b10 %
1'
b10 +
#822970000000
0!
0'
#822980000000
1!
b11 %
1'
b11 +
#822990000000
0!
0'
#823000000000
1!
b100 %
1'
b100 +
#823010000000
0!
0'
#823020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#823030000000
0!
0'
#823040000000
1!
0$
b110 %
1'
0*
b110 +
#823050000000
0!
0'
#823060000000
1!
b111 %
1'
b111 +
#823070000000
0!
0'
#823080000000
1!
b1000 %
1'
b1000 +
#823090000000
0!
0'
#823100000000
1!
b1001 %
1'
b1001 +
#823110000000
0!
0'
#823120000000
1!
b0 %
1'
b0 +
#823130000000
0!
0'
#823140000000
1!
1$
b1 %
1'
1*
b1 +
#823150000000
0!
0'
#823160000000
1!
b10 %
1'
b10 +
#823170000000
0!
0'
#823180000000
1!
b11 %
1'
b11 +
#823190000000
0!
0'
#823200000000
1!
b100 %
1'
b100 +
#823210000000
0!
0'
#823220000000
1!
b101 %
1'
b101 +
#823230000000
1"
1(
#823240000000
0!
0"
b100 &
0'
0(
b100 ,
#823250000000
1!
b110 %
1'
b110 +
#823260000000
0!
0'
#823270000000
1!
b111 %
1'
b111 +
#823280000000
0!
0'
#823290000000
1!
0$
b1000 %
1'
0*
b1000 +
#823300000000
0!
0'
#823310000000
1!
b1001 %
1'
b1001 +
#823320000000
0!
0'
#823330000000
1!
b0 %
1'
b0 +
#823340000000
0!
0'
#823350000000
1!
1$
b1 %
1'
1*
b1 +
#823360000000
0!
0'
#823370000000
1!
b10 %
1'
b10 +
#823380000000
0!
0'
#823390000000
1!
b11 %
1'
b11 +
#823400000000
0!
0'
#823410000000
1!
b100 %
1'
b100 +
#823420000000
0!
0'
#823430000000
1!
b101 %
1'
b101 +
#823440000000
0!
0'
#823450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#823460000000
0!
0'
#823470000000
1!
b111 %
1'
b111 +
#823480000000
0!
0'
#823490000000
1!
b1000 %
1'
b1000 +
#823500000000
0!
0'
#823510000000
1!
b1001 %
1'
b1001 +
#823520000000
0!
0'
#823530000000
1!
b0 %
1'
b0 +
#823540000000
0!
0'
#823550000000
1!
1$
b1 %
1'
1*
b1 +
#823560000000
0!
0'
#823570000000
1!
b10 %
1'
b10 +
#823580000000
0!
0'
#823590000000
1!
b11 %
1'
b11 +
#823600000000
0!
0'
#823610000000
1!
b100 %
1'
b100 +
#823620000000
0!
0'
#823630000000
1!
b101 %
1'
b101 +
#823640000000
0!
0'
#823650000000
1!
0$
b110 %
1'
0*
b110 +
#823660000000
1"
1(
#823670000000
0!
0"
b100 &
0'
0(
b100 ,
#823680000000
1!
1$
b111 %
1'
1*
b111 +
#823690000000
0!
0'
#823700000000
1!
0$
b1000 %
1'
0*
b1000 +
#823710000000
0!
0'
#823720000000
1!
b1001 %
1'
b1001 +
#823730000000
0!
0'
#823740000000
1!
b0 %
1'
b0 +
#823750000000
0!
0'
#823760000000
1!
1$
b1 %
1'
1*
b1 +
#823770000000
0!
0'
#823780000000
1!
b10 %
1'
b10 +
#823790000000
0!
0'
#823800000000
1!
b11 %
1'
b11 +
#823810000000
0!
0'
#823820000000
1!
b100 %
1'
b100 +
#823830000000
0!
0'
#823840000000
1!
b101 %
1'
b101 +
#823850000000
0!
0'
#823860000000
1!
b110 %
1'
b110 +
#823870000000
0!
0'
#823880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#823890000000
0!
0'
#823900000000
1!
b1000 %
1'
b1000 +
#823910000000
0!
0'
#823920000000
1!
b1001 %
1'
b1001 +
#823930000000
0!
0'
#823940000000
1!
b0 %
1'
b0 +
#823950000000
0!
0'
#823960000000
1!
1$
b1 %
1'
1*
b1 +
#823970000000
0!
0'
#823980000000
1!
b10 %
1'
b10 +
#823990000000
0!
0'
#824000000000
1!
b11 %
1'
b11 +
#824010000000
0!
0'
#824020000000
1!
b100 %
1'
b100 +
#824030000000
0!
0'
#824040000000
1!
b101 %
1'
b101 +
#824050000000
0!
0'
#824060000000
1!
0$
b110 %
1'
0*
b110 +
#824070000000
0!
0'
#824080000000
1!
b111 %
1'
b111 +
#824090000000
1"
1(
#824100000000
0!
0"
b100 &
0'
0(
b100 ,
#824110000000
1!
b1000 %
1'
b1000 +
#824120000000
0!
0'
#824130000000
1!
b1001 %
1'
b1001 +
#824140000000
0!
0'
#824150000000
1!
b0 %
1'
b0 +
#824160000000
0!
0'
#824170000000
1!
1$
b1 %
1'
1*
b1 +
#824180000000
0!
0'
#824190000000
1!
b10 %
1'
b10 +
#824200000000
0!
0'
#824210000000
1!
b11 %
1'
b11 +
#824220000000
0!
0'
#824230000000
1!
b100 %
1'
b100 +
#824240000000
0!
0'
#824250000000
1!
b101 %
1'
b101 +
#824260000000
0!
0'
#824270000000
1!
b110 %
1'
b110 +
#824280000000
0!
0'
#824290000000
1!
b111 %
1'
b111 +
#824300000000
0!
0'
#824310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#824320000000
0!
0'
#824330000000
1!
b1001 %
1'
b1001 +
#824340000000
0!
0'
#824350000000
1!
b0 %
1'
b0 +
#824360000000
0!
0'
#824370000000
1!
1$
b1 %
1'
1*
b1 +
#824380000000
0!
0'
#824390000000
1!
b10 %
1'
b10 +
#824400000000
0!
0'
#824410000000
1!
b11 %
1'
b11 +
#824420000000
0!
0'
#824430000000
1!
b100 %
1'
b100 +
#824440000000
0!
0'
#824450000000
1!
b101 %
1'
b101 +
#824460000000
0!
0'
#824470000000
1!
0$
b110 %
1'
0*
b110 +
#824480000000
0!
0'
#824490000000
1!
b111 %
1'
b111 +
#824500000000
0!
0'
#824510000000
1!
b1000 %
1'
b1000 +
#824520000000
1"
1(
#824530000000
0!
0"
b100 &
0'
0(
b100 ,
#824540000000
1!
b1001 %
1'
b1001 +
#824550000000
0!
0'
#824560000000
1!
b0 %
1'
b0 +
#824570000000
0!
0'
#824580000000
1!
1$
b1 %
1'
1*
b1 +
#824590000000
0!
0'
#824600000000
1!
b10 %
1'
b10 +
#824610000000
0!
0'
#824620000000
1!
b11 %
1'
b11 +
#824630000000
0!
0'
#824640000000
1!
b100 %
1'
b100 +
#824650000000
0!
0'
#824660000000
1!
b101 %
1'
b101 +
#824670000000
0!
0'
#824680000000
1!
b110 %
1'
b110 +
#824690000000
0!
0'
#824700000000
1!
b111 %
1'
b111 +
#824710000000
0!
0'
#824720000000
1!
0$
b1000 %
1'
0*
b1000 +
#824730000000
0!
0'
#824740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#824750000000
0!
0'
#824760000000
1!
b0 %
1'
b0 +
#824770000000
0!
0'
#824780000000
1!
1$
b1 %
1'
1*
b1 +
#824790000000
0!
0'
#824800000000
1!
b10 %
1'
b10 +
#824810000000
0!
0'
#824820000000
1!
b11 %
1'
b11 +
#824830000000
0!
0'
#824840000000
1!
b100 %
1'
b100 +
#824850000000
0!
0'
#824860000000
1!
b101 %
1'
b101 +
#824870000000
0!
0'
#824880000000
1!
0$
b110 %
1'
0*
b110 +
#824890000000
0!
0'
#824900000000
1!
b111 %
1'
b111 +
#824910000000
0!
0'
#824920000000
1!
b1000 %
1'
b1000 +
#824930000000
0!
0'
#824940000000
1!
b1001 %
1'
b1001 +
#824950000000
1"
1(
#824960000000
0!
0"
b100 &
0'
0(
b100 ,
#824970000000
1!
b0 %
1'
b0 +
#824980000000
0!
0'
#824990000000
1!
1$
b1 %
1'
1*
b1 +
#825000000000
0!
0'
#825010000000
1!
b10 %
1'
b10 +
#825020000000
0!
0'
#825030000000
1!
b11 %
1'
b11 +
#825040000000
0!
0'
#825050000000
1!
b100 %
1'
b100 +
#825060000000
0!
0'
#825070000000
1!
b101 %
1'
b101 +
#825080000000
0!
0'
#825090000000
1!
b110 %
1'
b110 +
#825100000000
0!
0'
#825110000000
1!
b111 %
1'
b111 +
#825120000000
0!
0'
#825130000000
1!
0$
b1000 %
1'
0*
b1000 +
#825140000000
0!
0'
#825150000000
1!
b1001 %
1'
b1001 +
#825160000000
0!
0'
#825170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#825180000000
0!
0'
#825190000000
1!
1$
b1 %
1'
1*
b1 +
#825200000000
0!
0'
#825210000000
1!
b10 %
1'
b10 +
#825220000000
0!
0'
#825230000000
1!
b11 %
1'
b11 +
#825240000000
0!
0'
#825250000000
1!
b100 %
1'
b100 +
#825260000000
0!
0'
#825270000000
1!
b101 %
1'
b101 +
#825280000000
0!
0'
#825290000000
1!
0$
b110 %
1'
0*
b110 +
#825300000000
0!
0'
#825310000000
1!
b111 %
1'
b111 +
#825320000000
0!
0'
#825330000000
1!
b1000 %
1'
b1000 +
#825340000000
0!
0'
#825350000000
1!
b1001 %
1'
b1001 +
#825360000000
0!
0'
#825370000000
1!
b0 %
1'
b0 +
#825380000000
1"
1(
#825390000000
0!
0"
b100 &
0'
0(
b100 ,
#825400000000
1!
1$
b1 %
1'
1*
b1 +
#825410000000
0!
0'
#825420000000
1!
b10 %
1'
b10 +
#825430000000
0!
0'
#825440000000
1!
b11 %
1'
b11 +
#825450000000
0!
0'
#825460000000
1!
b100 %
1'
b100 +
#825470000000
0!
0'
#825480000000
1!
b101 %
1'
b101 +
#825490000000
0!
0'
#825500000000
1!
b110 %
1'
b110 +
#825510000000
0!
0'
#825520000000
1!
b111 %
1'
b111 +
#825530000000
0!
0'
#825540000000
1!
0$
b1000 %
1'
0*
b1000 +
#825550000000
0!
0'
#825560000000
1!
b1001 %
1'
b1001 +
#825570000000
0!
0'
#825580000000
1!
b0 %
1'
b0 +
#825590000000
0!
0'
#825600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#825610000000
0!
0'
#825620000000
1!
b10 %
1'
b10 +
#825630000000
0!
0'
#825640000000
1!
b11 %
1'
b11 +
#825650000000
0!
0'
#825660000000
1!
b100 %
1'
b100 +
#825670000000
0!
0'
#825680000000
1!
b101 %
1'
b101 +
#825690000000
0!
0'
#825700000000
1!
0$
b110 %
1'
0*
b110 +
#825710000000
0!
0'
#825720000000
1!
b111 %
1'
b111 +
#825730000000
0!
0'
#825740000000
1!
b1000 %
1'
b1000 +
#825750000000
0!
0'
#825760000000
1!
b1001 %
1'
b1001 +
#825770000000
0!
0'
#825780000000
1!
b0 %
1'
b0 +
#825790000000
0!
0'
#825800000000
1!
1$
b1 %
1'
1*
b1 +
#825810000000
1"
1(
#825820000000
0!
0"
b100 &
0'
0(
b100 ,
#825830000000
1!
b10 %
1'
b10 +
#825840000000
0!
0'
#825850000000
1!
b11 %
1'
b11 +
#825860000000
0!
0'
#825870000000
1!
b100 %
1'
b100 +
#825880000000
0!
0'
#825890000000
1!
b101 %
1'
b101 +
#825900000000
0!
0'
#825910000000
1!
b110 %
1'
b110 +
#825920000000
0!
0'
#825930000000
1!
b111 %
1'
b111 +
#825940000000
0!
0'
#825950000000
1!
0$
b1000 %
1'
0*
b1000 +
#825960000000
0!
0'
#825970000000
1!
b1001 %
1'
b1001 +
#825980000000
0!
0'
#825990000000
1!
b0 %
1'
b0 +
#826000000000
0!
0'
#826010000000
1!
1$
b1 %
1'
1*
b1 +
#826020000000
0!
0'
#826030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#826040000000
0!
0'
#826050000000
1!
b11 %
1'
b11 +
#826060000000
0!
0'
#826070000000
1!
b100 %
1'
b100 +
#826080000000
0!
0'
#826090000000
1!
b101 %
1'
b101 +
#826100000000
0!
0'
#826110000000
1!
0$
b110 %
1'
0*
b110 +
#826120000000
0!
0'
#826130000000
1!
b111 %
1'
b111 +
#826140000000
0!
0'
#826150000000
1!
b1000 %
1'
b1000 +
#826160000000
0!
0'
#826170000000
1!
b1001 %
1'
b1001 +
#826180000000
0!
0'
#826190000000
1!
b0 %
1'
b0 +
#826200000000
0!
0'
#826210000000
1!
1$
b1 %
1'
1*
b1 +
#826220000000
0!
0'
#826230000000
1!
b10 %
1'
b10 +
#826240000000
1"
1(
#826250000000
0!
0"
b100 &
0'
0(
b100 ,
#826260000000
1!
b11 %
1'
b11 +
#826270000000
0!
0'
#826280000000
1!
b100 %
1'
b100 +
#826290000000
0!
0'
#826300000000
1!
b101 %
1'
b101 +
#826310000000
0!
0'
#826320000000
1!
b110 %
1'
b110 +
#826330000000
0!
0'
#826340000000
1!
b111 %
1'
b111 +
#826350000000
0!
0'
#826360000000
1!
0$
b1000 %
1'
0*
b1000 +
#826370000000
0!
0'
#826380000000
1!
b1001 %
1'
b1001 +
#826390000000
0!
0'
#826400000000
1!
b0 %
1'
b0 +
#826410000000
0!
0'
#826420000000
1!
1$
b1 %
1'
1*
b1 +
#826430000000
0!
0'
#826440000000
1!
b10 %
1'
b10 +
#826450000000
0!
0'
#826460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#826470000000
0!
0'
#826480000000
1!
b100 %
1'
b100 +
#826490000000
0!
0'
#826500000000
1!
b101 %
1'
b101 +
#826510000000
0!
0'
#826520000000
1!
0$
b110 %
1'
0*
b110 +
#826530000000
0!
0'
#826540000000
1!
b111 %
1'
b111 +
#826550000000
0!
0'
#826560000000
1!
b1000 %
1'
b1000 +
#826570000000
0!
0'
#826580000000
1!
b1001 %
1'
b1001 +
#826590000000
0!
0'
#826600000000
1!
b0 %
1'
b0 +
#826610000000
0!
0'
#826620000000
1!
1$
b1 %
1'
1*
b1 +
#826630000000
0!
0'
#826640000000
1!
b10 %
1'
b10 +
#826650000000
0!
0'
#826660000000
1!
b11 %
1'
b11 +
#826670000000
1"
1(
#826680000000
0!
0"
b100 &
0'
0(
b100 ,
#826690000000
1!
b100 %
1'
b100 +
#826700000000
0!
0'
#826710000000
1!
b101 %
1'
b101 +
#826720000000
0!
0'
#826730000000
1!
b110 %
1'
b110 +
#826740000000
0!
0'
#826750000000
1!
b111 %
1'
b111 +
#826760000000
0!
0'
#826770000000
1!
0$
b1000 %
1'
0*
b1000 +
#826780000000
0!
0'
#826790000000
1!
b1001 %
1'
b1001 +
#826800000000
0!
0'
#826810000000
1!
b0 %
1'
b0 +
#826820000000
0!
0'
#826830000000
1!
1$
b1 %
1'
1*
b1 +
#826840000000
0!
0'
#826850000000
1!
b10 %
1'
b10 +
#826860000000
0!
0'
#826870000000
1!
b11 %
1'
b11 +
#826880000000
0!
0'
#826890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#826900000000
0!
0'
#826910000000
1!
b101 %
1'
b101 +
#826920000000
0!
0'
#826930000000
1!
0$
b110 %
1'
0*
b110 +
#826940000000
0!
0'
#826950000000
1!
b111 %
1'
b111 +
#826960000000
0!
0'
#826970000000
1!
b1000 %
1'
b1000 +
#826980000000
0!
0'
#826990000000
1!
b1001 %
1'
b1001 +
#827000000000
0!
0'
#827010000000
1!
b0 %
1'
b0 +
#827020000000
0!
0'
#827030000000
1!
1$
b1 %
1'
1*
b1 +
#827040000000
0!
0'
#827050000000
1!
b10 %
1'
b10 +
#827060000000
0!
0'
#827070000000
1!
b11 %
1'
b11 +
#827080000000
0!
0'
#827090000000
1!
b100 %
1'
b100 +
#827100000000
1"
1(
#827110000000
0!
0"
b100 &
0'
0(
b100 ,
#827120000000
1!
b101 %
1'
b101 +
#827130000000
0!
0'
#827140000000
1!
b110 %
1'
b110 +
#827150000000
0!
0'
#827160000000
1!
b111 %
1'
b111 +
#827170000000
0!
0'
#827180000000
1!
0$
b1000 %
1'
0*
b1000 +
#827190000000
0!
0'
#827200000000
1!
b1001 %
1'
b1001 +
#827210000000
0!
0'
#827220000000
1!
b0 %
1'
b0 +
#827230000000
0!
0'
#827240000000
1!
1$
b1 %
1'
1*
b1 +
#827250000000
0!
0'
#827260000000
1!
b10 %
1'
b10 +
#827270000000
0!
0'
#827280000000
1!
b11 %
1'
b11 +
#827290000000
0!
0'
#827300000000
1!
b100 %
1'
b100 +
#827310000000
0!
0'
#827320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#827330000000
0!
0'
#827340000000
1!
0$
b110 %
1'
0*
b110 +
#827350000000
0!
0'
#827360000000
1!
b111 %
1'
b111 +
#827370000000
0!
0'
#827380000000
1!
b1000 %
1'
b1000 +
#827390000000
0!
0'
#827400000000
1!
b1001 %
1'
b1001 +
#827410000000
0!
0'
#827420000000
1!
b0 %
1'
b0 +
#827430000000
0!
0'
#827440000000
1!
1$
b1 %
1'
1*
b1 +
#827450000000
0!
0'
#827460000000
1!
b10 %
1'
b10 +
#827470000000
0!
0'
#827480000000
1!
b11 %
1'
b11 +
#827490000000
0!
0'
#827500000000
1!
b100 %
1'
b100 +
#827510000000
0!
0'
#827520000000
1!
b101 %
1'
b101 +
#827530000000
1"
1(
#827540000000
0!
0"
b100 &
0'
0(
b100 ,
#827550000000
1!
b110 %
1'
b110 +
#827560000000
0!
0'
#827570000000
1!
b111 %
1'
b111 +
#827580000000
0!
0'
#827590000000
1!
0$
b1000 %
1'
0*
b1000 +
#827600000000
0!
0'
#827610000000
1!
b1001 %
1'
b1001 +
#827620000000
0!
0'
#827630000000
1!
b0 %
1'
b0 +
#827640000000
0!
0'
#827650000000
1!
1$
b1 %
1'
1*
b1 +
#827660000000
0!
0'
#827670000000
1!
b10 %
1'
b10 +
#827680000000
0!
0'
#827690000000
1!
b11 %
1'
b11 +
#827700000000
0!
0'
#827710000000
1!
b100 %
1'
b100 +
#827720000000
0!
0'
#827730000000
1!
b101 %
1'
b101 +
#827740000000
0!
0'
#827750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#827760000000
0!
0'
#827770000000
1!
b111 %
1'
b111 +
#827780000000
0!
0'
#827790000000
1!
b1000 %
1'
b1000 +
#827800000000
0!
0'
#827810000000
1!
b1001 %
1'
b1001 +
#827820000000
0!
0'
#827830000000
1!
b0 %
1'
b0 +
#827840000000
0!
0'
#827850000000
1!
1$
b1 %
1'
1*
b1 +
#827860000000
0!
0'
#827870000000
1!
b10 %
1'
b10 +
#827880000000
0!
0'
#827890000000
1!
b11 %
1'
b11 +
#827900000000
0!
0'
#827910000000
1!
b100 %
1'
b100 +
#827920000000
0!
0'
#827930000000
1!
b101 %
1'
b101 +
#827940000000
0!
0'
#827950000000
1!
0$
b110 %
1'
0*
b110 +
#827960000000
1"
1(
#827970000000
0!
0"
b100 &
0'
0(
b100 ,
#827980000000
1!
1$
b111 %
1'
1*
b111 +
#827990000000
0!
0'
#828000000000
1!
0$
b1000 %
1'
0*
b1000 +
#828010000000
0!
0'
#828020000000
1!
b1001 %
1'
b1001 +
#828030000000
0!
0'
#828040000000
1!
b0 %
1'
b0 +
#828050000000
0!
0'
#828060000000
1!
1$
b1 %
1'
1*
b1 +
#828070000000
0!
0'
#828080000000
1!
b10 %
1'
b10 +
#828090000000
0!
0'
#828100000000
1!
b11 %
1'
b11 +
#828110000000
0!
0'
#828120000000
1!
b100 %
1'
b100 +
#828130000000
0!
0'
#828140000000
1!
b101 %
1'
b101 +
#828150000000
0!
0'
#828160000000
1!
b110 %
1'
b110 +
#828170000000
0!
0'
#828180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#828190000000
0!
0'
#828200000000
1!
b1000 %
1'
b1000 +
#828210000000
0!
0'
#828220000000
1!
b1001 %
1'
b1001 +
#828230000000
0!
0'
#828240000000
1!
b0 %
1'
b0 +
#828250000000
0!
0'
#828260000000
1!
1$
b1 %
1'
1*
b1 +
#828270000000
0!
0'
#828280000000
1!
b10 %
1'
b10 +
#828290000000
0!
0'
#828300000000
1!
b11 %
1'
b11 +
#828310000000
0!
0'
#828320000000
1!
b100 %
1'
b100 +
#828330000000
0!
0'
#828340000000
1!
b101 %
1'
b101 +
#828350000000
0!
0'
#828360000000
1!
0$
b110 %
1'
0*
b110 +
#828370000000
0!
0'
#828380000000
1!
b111 %
1'
b111 +
#828390000000
1"
1(
#828400000000
0!
0"
b100 &
0'
0(
b100 ,
#828410000000
1!
b1000 %
1'
b1000 +
#828420000000
0!
0'
#828430000000
1!
b1001 %
1'
b1001 +
#828440000000
0!
0'
#828450000000
1!
b0 %
1'
b0 +
#828460000000
0!
0'
#828470000000
1!
1$
b1 %
1'
1*
b1 +
#828480000000
0!
0'
#828490000000
1!
b10 %
1'
b10 +
#828500000000
0!
0'
#828510000000
1!
b11 %
1'
b11 +
#828520000000
0!
0'
#828530000000
1!
b100 %
1'
b100 +
#828540000000
0!
0'
#828550000000
1!
b101 %
1'
b101 +
#828560000000
0!
0'
#828570000000
1!
b110 %
1'
b110 +
#828580000000
0!
0'
#828590000000
1!
b111 %
1'
b111 +
#828600000000
0!
0'
#828610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#828620000000
0!
0'
#828630000000
1!
b1001 %
1'
b1001 +
#828640000000
0!
0'
#828650000000
1!
b0 %
1'
b0 +
#828660000000
0!
0'
#828670000000
1!
1$
b1 %
1'
1*
b1 +
#828680000000
0!
0'
#828690000000
1!
b10 %
1'
b10 +
#828700000000
0!
0'
#828710000000
1!
b11 %
1'
b11 +
#828720000000
0!
0'
#828730000000
1!
b100 %
1'
b100 +
#828740000000
0!
0'
#828750000000
1!
b101 %
1'
b101 +
#828760000000
0!
0'
#828770000000
1!
0$
b110 %
1'
0*
b110 +
#828780000000
0!
0'
#828790000000
1!
b111 %
1'
b111 +
#828800000000
0!
0'
#828810000000
1!
b1000 %
1'
b1000 +
#828820000000
1"
1(
#828830000000
0!
0"
b100 &
0'
0(
b100 ,
#828840000000
1!
b1001 %
1'
b1001 +
#828850000000
0!
0'
#828860000000
1!
b0 %
1'
b0 +
#828870000000
0!
0'
#828880000000
1!
1$
b1 %
1'
1*
b1 +
#828890000000
0!
0'
#828900000000
1!
b10 %
1'
b10 +
#828910000000
0!
0'
#828920000000
1!
b11 %
1'
b11 +
#828930000000
0!
0'
#828940000000
1!
b100 %
1'
b100 +
#828950000000
0!
0'
#828960000000
1!
b101 %
1'
b101 +
#828970000000
0!
0'
#828980000000
1!
b110 %
1'
b110 +
#828990000000
0!
0'
#829000000000
1!
b111 %
1'
b111 +
#829010000000
0!
0'
#829020000000
1!
0$
b1000 %
1'
0*
b1000 +
#829030000000
0!
0'
#829040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#829050000000
0!
0'
#829060000000
1!
b0 %
1'
b0 +
#829070000000
0!
0'
#829080000000
1!
1$
b1 %
1'
1*
b1 +
#829090000000
0!
0'
#829100000000
1!
b10 %
1'
b10 +
#829110000000
0!
0'
#829120000000
1!
b11 %
1'
b11 +
#829130000000
0!
0'
#829140000000
1!
b100 %
1'
b100 +
#829150000000
0!
0'
#829160000000
1!
b101 %
1'
b101 +
#829170000000
0!
0'
#829180000000
1!
0$
b110 %
1'
0*
b110 +
#829190000000
0!
0'
#829200000000
1!
b111 %
1'
b111 +
#829210000000
0!
0'
#829220000000
1!
b1000 %
1'
b1000 +
#829230000000
0!
0'
#829240000000
1!
b1001 %
1'
b1001 +
#829250000000
1"
1(
#829260000000
0!
0"
b100 &
0'
0(
b100 ,
#829270000000
1!
b0 %
1'
b0 +
#829280000000
0!
0'
#829290000000
1!
1$
b1 %
1'
1*
b1 +
#829300000000
0!
0'
#829310000000
1!
b10 %
1'
b10 +
#829320000000
0!
0'
#829330000000
1!
b11 %
1'
b11 +
#829340000000
0!
0'
#829350000000
1!
b100 %
1'
b100 +
#829360000000
0!
0'
#829370000000
1!
b101 %
1'
b101 +
#829380000000
0!
0'
#829390000000
1!
b110 %
1'
b110 +
#829400000000
0!
0'
#829410000000
1!
b111 %
1'
b111 +
#829420000000
0!
0'
#829430000000
1!
0$
b1000 %
1'
0*
b1000 +
#829440000000
0!
0'
#829450000000
1!
b1001 %
1'
b1001 +
#829460000000
0!
0'
#829470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#829480000000
0!
0'
#829490000000
1!
1$
b1 %
1'
1*
b1 +
#829500000000
0!
0'
#829510000000
1!
b10 %
1'
b10 +
#829520000000
0!
0'
#829530000000
1!
b11 %
1'
b11 +
#829540000000
0!
0'
#829550000000
1!
b100 %
1'
b100 +
#829560000000
0!
0'
#829570000000
1!
b101 %
1'
b101 +
#829580000000
0!
0'
#829590000000
1!
0$
b110 %
1'
0*
b110 +
#829600000000
0!
0'
#829610000000
1!
b111 %
1'
b111 +
#829620000000
0!
0'
#829630000000
1!
b1000 %
1'
b1000 +
#829640000000
0!
0'
#829650000000
1!
b1001 %
1'
b1001 +
#829660000000
0!
0'
#829670000000
1!
b0 %
1'
b0 +
#829680000000
1"
1(
#829690000000
0!
0"
b100 &
0'
0(
b100 ,
#829700000000
1!
1$
b1 %
1'
1*
b1 +
#829710000000
0!
0'
#829720000000
1!
b10 %
1'
b10 +
#829730000000
0!
0'
#829740000000
1!
b11 %
1'
b11 +
#829750000000
0!
0'
#829760000000
1!
b100 %
1'
b100 +
#829770000000
0!
0'
#829780000000
1!
b101 %
1'
b101 +
#829790000000
0!
0'
#829800000000
1!
b110 %
1'
b110 +
#829810000000
0!
0'
#829820000000
1!
b111 %
1'
b111 +
#829830000000
0!
0'
#829840000000
1!
0$
b1000 %
1'
0*
b1000 +
#829850000000
0!
0'
#829860000000
1!
b1001 %
1'
b1001 +
#829870000000
0!
0'
#829880000000
1!
b0 %
1'
b0 +
#829890000000
0!
0'
#829900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#829910000000
0!
0'
#829920000000
1!
b10 %
1'
b10 +
#829930000000
0!
0'
#829940000000
1!
b11 %
1'
b11 +
#829950000000
0!
0'
#829960000000
1!
b100 %
1'
b100 +
#829970000000
0!
0'
#829980000000
1!
b101 %
1'
b101 +
#829990000000
0!
0'
#830000000000
1!
0$
b110 %
1'
0*
b110 +
#830010000000
0!
0'
#830020000000
1!
b111 %
1'
b111 +
#830030000000
0!
0'
#830040000000
1!
b1000 %
1'
b1000 +
#830050000000
0!
0'
#830060000000
1!
b1001 %
1'
b1001 +
#830070000000
0!
0'
#830080000000
1!
b0 %
1'
b0 +
#830090000000
0!
0'
#830100000000
1!
1$
b1 %
1'
1*
b1 +
#830110000000
1"
1(
#830120000000
0!
0"
b100 &
0'
0(
b100 ,
#830130000000
1!
b10 %
1'
b10 +
#830140000000
0!
0'
#830150000000
1!
b11 %
1'
b11 +
#830160000000
0!
0'
#830170000000
1!
b100 %
1'
b100 +
#830180000000
0!
0'
#830190000000
1!
b101 %
1'
b101 +
#830200000000
0!
0'
#830210000000
1!
b110 %
1'
b110 +
#830220000000
0!
0'
#830230000000
1!
b111 %
1'
b111 +
#830240000000
0!
0'
#830250000000
1!
0$
b1000 %
1'
0*
b1000 +
#830260000000
0!
0'
#830270000000
1!
b1001 %
1'
b1001 +
#830280000000
0!
0'
#830290000000
1!
b0 %
1'
b0 +
#830300000000
0!
0'
#830310000000
1!
1$
b1 %
1'
1*
b1 +
#830320000000
0!
0'
#830330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#830340000000
0!
0'
#830350000000
1!
b11 %
1'
b11 +
#830360000000
0!
0'
#830370000000
1!
b100 %
1'
b100 +
#830380000000
0!
0'
#830390000000
1!
b101 %
1'
b101 +
#830400000000
0!
0'
#830410000000
1!
0$
b110 %
1'
0*
b110 +
#830420000000
0!
0'
#830430000000
1!
b111 %
1'
b111 +
#830440000000
0!
0'
#830450000000
1!
b1000 %
1'
b1000 +
#830460000000
0!
0'
#830470000000
1!
b1001 %
1'
b1001 +
#830480000000
0!
0'
#830490000000
1!
b0 %
1'
b0 +
#830500000000
0!
0'
#830510000000
1!
1$
b1 %
1'
1*
b1 +
#830520000000
0!
0'
#830530000000
1!
b10 %
1'
b10 +
#830540000000
1"
1(
#830550000000
0!
0"
b100 &
0'
0(
b100 ,
#830560000000
1!
b11 %
1'
b11 +
#830570000000
0!
0'
#830580000000
1!
b100 %
1'
b100 +
#830590000000
0!
0'
#830600000000
1!
b101 %
1'
b101 +
#830610000000
0!
0'
#830620000000
1!
b110 %
1'
b110 +
#830630000000
0!
0'
#830640000000
1!
b111 %
1'
b111 +
#830650000000
0!
0'
#830660000000
1!
0$
b1000 %
1'
0*
b1000 +
#830670000000
0!
0'
#830680000000
1!
b1001 %
1'
b1001 +
#830690000000
0!
0'
#830700000000
1!
b0 %
1'
b0 +
#830710000000
0!
0'
#830720000000
1!
1$
b1 %
1'
1*
b1 +
#830730000000
0!
0'
#830740000000
1!
b10 %
1'
b10 +
#830750000000
0!
0'
#830760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#830770000000
0!
0'
#830780000000
1!
b100 %
1'
b100 +
#830790000000
0!
0'
#830800000000
1!
b101 %
1'
b101 +
#830810000000
0!
0'
#830820000000
1!
0$
b110 %
1'
0*
b110 +
#830830000000
0!
0'
#830840000000
1!
b111 %
1'
b111 +
#830850000000
0!
0'
#830860000000
1!
b1000 %
1'
b1000 +
#830870000000
0!
0'
#830880000000
1!
b1001 %
1'
b1001 +
#830890000000
0!
0'
#830900000000
1!
b0 %
1'
b0 +
#830910000000
0!
0'
#830920000000
1!
1$
b1 %
1'
1*
b1 +
#830930000000
0!
0'
#830940000000
1!
b10 %
1'
b10 +
#830950000000
0!
0'
#830960000000
1!
b11 %
1'
b11 +
#830970000000
1"
1(
#830980000000
0!
0"
b100 &
0'
0(
b100 ,
#830990000000
1!
b100 %
1'
b100 +
#831000000000
0!
0'
#831010000000
1!
b101 %
1'
b101 +
#831020000000
0!
0'
#831030000000
1!
b110 %
1'
b110 +
#831040000000
0!
0'
#831050000000
1!
b111 %
1'
b111 +
#831060000000
0!
0'
#831070000000
1!
0$
b1000 %
1'
0*
b1000 +
#831080000000
0!
0'
#831090000000
1!
b1001 %
1'
b1001 +
#831100000000
0!
0'
#831110000000
1!
b0 %
1'
b0 +
#831120000000
0!
0'
#831130000000
1!
1$
b1 %
1'
1*
b1 +
#831140000000
0!
0'
#831150000000
1!
b10 %
1'
b10 +
#831160000000
0!
0'
#831170000000
1!
b11 %
1'
b11 +
#831180000000
0!
0'
#831190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#831200000000
0!
0'
#831210000000
1!
b101 %
1'
b101 +
#831220000000
0!
0'
#831230000000
1!
0$
b110 %
1'
0*
b110 +
#831240000000
0!
0'
#831250000000
1!
b111 %
1'
b111 +
#831260000000
0!
0'
#831270000000
1!
b1000 %
1'
b1000 +
#831280000000
0!
0'
#831290000000
1!
b1001 %
1'
b1001 +
#831300000000
0!
0'
#831310000000
1!
b0 %
1'
b0 +
#831320000000
0!
0'
#831330000000
1!
1$
b1 %
1'
1*
b1 +
#831340000000
0!
0'
#831350000000
1!
b10 %
1'
b10 +
#831360000000
0!
0'
#831370000000
1!
b11 %
1'
b11 +
#831380000000
0!
0'
#831390000000
1!
b100 %
1'
b100 +
#831400000000
1"
1(
#831410000000
0!
0"
b100 &
0'
0(
b100 ,
#831420000000
1!
b101 %
1'
b101 +
#831430000000
0!
0'
#831440000000
1!
b110 %
1'
b110 +
#831450000000
0!
0'
#831460000000
1!
b111 %
1'
b111 +
#831470000000
0!
0'
#831480000000
1!
0$
b1000 %
1'
0*
b1000 +
#831490000000
0!
0'
#831500000000
1!
b1001 %
1'
b1001 +
#831510000000
0!
0'
#831520000000
1!
b0 %
1'
b0 +
#831530000000
0!
0'
#831540000000
1!
1$
b1 %
1'
1*
b1 +
#831550000000
0!
0'
#831560000000
1!
b10 %
1'
b10 +
#831570000000
0!
0'
#831580000000
1!
b11 %
1'
b11 +
#831590000000
0!
0'
#831600000000
1!
b100 %
1'
b100 +
#831610000000
0!
0'
#831620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#831630000000
0!
0'
#831640000000
1!
0$
b110 %
1'
0*
b110 +
#831650000000
0!
0'
#831660000000
1!
b111 %
1'
b111 +
#831670000000
0!
0'
#831680000000
1!
b1000 %
1'
b1000 +
#831690000000
0!
0'
#831700000000
1!
b1001 %
1'
b1001 +
#831710000000
0!
0'
#831720000000
1!
b0 %
1'
b0 +
#831730000000
0!
0'
#831740000000
1!
1$
b1 %
1'
1*
b1 +
#831750000000
0!
0'
#831760000000
1!
b10 %
1'
b10 +
#831770000000
0!
0'
#831780000000
1!
b11 %
1'
b11 +
#831790000000
0!
0'
#831800000000
1!
b100 %
1'
b100 +
#831810000000
0!
0'
#831820000000
1!
b101 %
1'
b101 +
#831830000000
1"
1(
#831840000000
0!
0"
b100 &
0'
0(
b100 ,
#831850000000
1!
b110 %
1'
b110 +
#831860000000
0!
0'
#831870000000
1!
b111 %
1'
b111 +
#831880000000
0!
0'
#831890000000
1!
0$
b1000 %
1'
0*
b1000 +
#831900000000
0!
0'
#831910000000
1!
b1001 %
1'
b1001 +
#831920000000
0!
0'
#831930000000
1!
b0 %
1'
b0 +
#831940000000
0!
0'
#831950000000
1!
1$
b1 %
1'
1*
b1 +
#831960000000
0!
0'
#831970000000
1!
b10 %
1'
b10 +
#831980000000
0!
0'
#831990000000
1!
b11 %
1'
b11 +
#832000000000
0!
0'
#832010000000
1!
b100 %
1'
b100 +
#832020000000
0!
0'
#832030000000
1!
b101 %
1'
b101 +
#832040000000
0!
0'
#832050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#832060000000
0!
0'
#832070000000
1!
b111 %
1'
b111 +
#832080000000
0!
0'
#832090000000
1!
b1000 %
1'
b1000 +
#832100000000
0!
0'
#832110000000
1!
b1001 %
1'
b1001 +
#832120000000
0!
0'
#832130000000
1!
b0 %
1'
b0 +
#832140000000
0!
0'
#832150000000
1!
1$
b1 %
1'
1*
b1 +
#832160000000
0!
0'
#832170000000
1!
b10 %
1'
b10 +
#832180000000
0!
0'
#832190000000
1!
b11 %
1'
b11 +
#832200000000
0!
0'
#832210000000
1!
b100 %
1'
b100 +
#832220000000
0!
0'
#832230000000
1!
b101 %
1'
b101 +
#832240000000
0!
0'
#832250000000
1!
0$
b110 %
1'
0*
b110 +
#832260000000
1"
1(
#832270000000
0!
0"
b100 &
0'
0(
b100 ,
#832280000000
1!
1$
b111 %
1'
1*
b111 +
#832290000000
0!
0'
#832300000000
1!
0$
b1000 %
1'
0*
b1000 +
#832310000000
0!
0'
#832320000000
1!
b1001 %
1'
b1001 +
#832330000000
0!
0'
#832340000000
1!
b0 %
1'
b0 +
#832350000000
0!
0'
#832360000000
1!
1$
b1 %
1'
1*
b1 +
#832370000000
0!
0'
#832380000000
1!
b10 %
1'
b10 +
#832390000000
0!
0'
#832400000000
1!
b11 %
1'
b11 +
#832410000000
0!
0'
#832420000000
1!
b100 %
1'
b100 +
#832430000000
0!
0'
#832440000000
1!
b101 %
1'
b101 +
#832450000000
0!
0'
#832460000000
1!
b110 %
1'
b110 +
#832470000000
0!
0'
#832480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#832490000000
0!
0'
#832500000000
1!
b1000 %
1'
b1000 +
#832510000000
0!
0'
#832520000000
1!
b1001 %
1'
b1001 +
#832530000000
0!
0'
#832540000000
1!
b0 %
1'
b0 +
#832550000000
0!
0'
#832560000000
1!
1$
b1 %
1'
1*
b1 +
#832570000000
0!
0'
#832580000000
1!
b10 %
1'
b10 +
#832590000000
0!
0'
#832600000000
1!
b11 %
1'
b11 +
#832610000000
0!
0'
#832620000000
1!
b100 %
1'
b100 +
#832630000000
0!
0'
#832640000000
1!
b101 %
1'
b101 +
#832650000000
0!
0'
#832660000000
1!
0$
b110 %
1'
0*
b110 +
#832670000000
0!
0'
#832680000000
1!
b111 %
1'
b111 +
#832690000000
1"
1(
#832700000000
0!
0"
b100 &
0'
0(
b100 ,
#832710000000
1!
b1000 %
1'
b1000 +
#832720000000
0!
0'
#832730000000
1!
b1001 %
1'
b1001 +
#832740000000
0!
0'
#832750000000
1!
b0 %
1'
b0 +
#832760000000
0!
0'
#832770000000
1!
1$
b1 %
1'
1*
b1 +
#832780000000
0!
0'
#832790000000
1!
b10 %
1'
b10 +
#832800000000
0!
0'
#832810000000
1!
b11 %
1'
b11 +
#832820000000
0!
0'
#832830000000
1!
b100 %
1'
b100 +
#832840000000
0!
0'
#832850000000
1!
b101 %
1'
b101 +
#832860000000
0!
0'
#832870000000
1!
b110 %
1'
b110 +
#832880000000
0!
0'
#832890000000
1!
b111 %
1'
b111 +
#832900000000
0!
0'
#832910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#832920000000
0!
0'
#832930000000
1!
b1001 %
1'
b1001 +
#832940000000
0!
0'
#832950000000
1!
b0 %
1'
b0 +
#832960000000
0!
0'
#832970000000
1!
1$
b1 %
1'
1*
b1 +
#832980000000
0!
0'
#832990000000
1!
b10 %
1'
b10 +
#833000000000
0!
0'
#833010000000
1!
b11 %
1'
b11 +
#833020000000
0!
0'
#833030000000
1!
b100 %
1'
b100 +
#833040000000
0!
0'
#833050000000
1!
b101 %
1'
b101 +
#833060000000
0!
0'
#833070000000
1!
0$
b110 %
1'
0*
b110 +
#833080000000
0!
0'
#833090000000
1!
b111 %
1'
b111 +
#833100000000
0!
0'
#833110000000
1!
b1000 %
1'
b1000 +
#833120000000
1"
1(
#833130000000
0!
0"
b100 &
0'
0(
b100 ,
#833140000000
1!
b1001 %
1'
b1001 +
#833150000000
0!
0'
#833160000000
1!
b0 %
1'
b0 +
#833170000000
0!
0'
#833180000000
1!
1$
b1 %
1'
1*
b1 +
#833190000000
0!
0'
#833200000000
1!
b10 %
1'
b10 +
#833210000000
0!
0'
#833220000000
1!
b11 %
1'
b11 +
#833230000000
0!
0'
#833240000000
1!
b100 %
1'
b100 +
#833250000000
0!
0'
#833260000000
1!
b101 %
1'
b101 +
#833270000000
0!
0'
#833280000000
1!
b110 %
1'
b110 +
#833290000000
0!
0'
#833300000000
1!
b111 %
1'
b111 +
#833310000000
0!
0'
#833320000000
1!
0$
b1000 %
1'
0*
b1000 +
#833330000000
0!
0'
#833340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#833350000000
0!
0'
#833360000000
1!
b0 %
1'
b0 +
#833370000000
0!
0'
#833380000000
1!
1$
b1 %
1'
1*
b1 +
#833390000000
0!
0'
#833400000000
1!
b10 %
1'
b10 +
#833410000000
0!
0'
#833420000000
1!
b11 %
1'
b11 +
#833430000000
0!
0'
#833440000000
1!
b100 %
1'
b100 +
#833450000000
0!
0'
#833460000000
1!
b101 %
1'
b101 +
#833470000000
0!
0'
#833480000000
1!
0$
b110 %
1'
0*
b110 +
#833490000000
0!
0'
#833500000000
1!
b111 %
1'
b111 +
#833510000000
0!
0'
#833520000000
1!
b1000 %
1'
b1000 +
#833530000000
0!
0'
#833540000000
1!
b1001 %
1'
b1001 +
#833550000000
1"
1(
#833560000000
0!
0"
b100 &
0'
0(
b100 ,
#833570000000
1!
b0 %
1'
b0 +
#833580000000
0!
0'
#833590000000
1!
1$
b1 %
1'
1*
b1 +
#833600000000
0!
0'
#833610000000
1!
b10 %
1'
b10 +
#833620000000
0!
0'
#833630000000
1!
b11 %
1'
b11 +
#833640000000
0!
0'
#833650000000
1!
b100 %
1'
b100 +
#833660000000
0!
0'
#833670000000
1!
b101 %
1'
b101 +
#833680000000
0!
0'
#833690000000
1!
b110 %
1'
b110 +
#833700000000
0!
0'
#833710000000
1!
b111 %
1'
b111 +
#833720000000
0!
0'
#833730000000
1!
0$
b1000 %
1'
0*
b1000 +
#833740000000
0!
0'
#833750000000
1!
b1001 %
1'
b1001 +
#833760000000
0!
0'
#833770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#833780000000
0!
0'
#833790000000
1!
1$
b1 %
1'
1*
b1 +
#833800000000
0!
0'
#833810000000
1!
b10 %
1'
b10 +
#833820000000
0!
0'
#833830000000
1!
b11 %
1'
b11 +
#833840000000
0!
0'
#833850000000
1!
b100 %
1'
b100 +
#833860000000
0!
0'
#833870000000
1!
b101 %
1'
b101 +
#833880000000
0!
0'
#833890000000
1!
0$
b110 %
1'
0*
b110 +
#833900000000
0!
0'
#833910000000
1!
b111 %
1'
b111 +
#833920000000
0!
0'
#833930000000
1!
b1000 %
1'
b1000 +
#833940000000
0!
0'
#833950000000
1!
b1001 %
1'
b1001 +
#833960000000
0!
0'
#833970000000
1!
b0 %
1'
b0 +
#833980000000
1"
1(
#833990000000
0!
0"
b100 &
0'
0(
b100 ,
#834000000000
1!
1$
b1 %
1'
1*
b1 +
#834010000000
0!
0'
#834020000000
1!
b10 %
1'
b10 +
#834030000000
0!
0'
#834040000000
1!
b11 %
1'
b11 +
#834050000000
0!
0'
#834060000000
1!
b100 %
1'
b100 +
#834070000000
0!
0'
#834080000000
1!
b101 %
1'
b101 +
#834090000000
0!
0'
#834100000000
1!
b110 %
1'
b110 +
#834110000000
0!
0'
#834120000000
1!
b111 %
1'
b111 +
#834130000000
0!
0'
#834140000000
1!
0$
b1000 %
1'
0*
b1000 +
#834150000000
0!
0'
#834160000000
1!
b1001 %
1'
b1001 +
#834170000000
0!
0'
#834180000000
1!
b0 %
1'
b0 +
#834190000000
0!
0'
#834200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#834210000000
0!
0'
#834220000000
1!
b10 %
1'
b10 +
#834230000000
0!
0'
#834240000000
1!
b11 %
1'
b11 +
#834250000000
0!
0'
#834260000000
1!
b100 %
1'
b100 +
#834270000000
0!
0'
#834280000000
1!
b101 %
1'
b101 +
#834290000000
0!
0'
#834300000000
1!
0$
b110 %
1'
0*
b110 +
#834310000000
0!
0'
#834320000000
1!
b111 %
1'
b111 +
#834330000000
0!
0'
#834340000000
1!
b1000 %
1'
b1000 +
#834350000000
0!
0'
#834360000000
1!
b1001 %
1'
b1001 +
#834370000000
0!
0'
#834380000000
1!
b0 %
1'
b0 +
#834390000000
0!
0'
#834400000000
1!
1$
b1 %
1'
1*
b1 +
#834410000000
1"
1(
#834420000000
0!
0"
b100 &
0'
0(
b100 ,
#834430000000
1!
b10 %
1'
b10 +
#834440000000
0!
0'
#834450000000
1!
b11 %
1'
b11 +
#834460000000
0!
0'
#834470000000
1!
b100 %
1'
b100 +
#834480000000
0!
0'
#834490000000
1!
b101 %
1'
b101 +
#834500000000
0!
0'
#834510000000
1!
b110 %
1'
b110 +
#834520000000
0!
0'
#834530000000
1!
b111 %
1'
b111 +
#834540000000
0!
0'
#834550000000
1!
0$
b1000 %
1'
0*
b1000 +
#834560000000
0!
0'
#834570000000
1!
b1001 %
1'
b1001 +
#834580000000
0!
0'
#834590000000
1!
b0 %
1'
b0 +
#834600000000
0!
0'
#834610000000
1!
1$
b1 %
1'
1*
b1 +
#834620000000
0!
0'
#834630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#834640000000
0!
0'
#834650000000
1!
b11 %
1'
b11 +
#834660000000
0!
0'
#834670000000
1!
b100 %
1'
b100 +
#834680000000
0!
0'
#834690000000
1!
b101 %
1'
b101 +
#834700000000
0!
0'
#834710000000
1!
0$
b110 %
1'
0*
b110 +
#834720000000
0!
0'
#834730000000
1!
b111 %
1'
b111 +
#834740000000
0!
0'
#834750000000
1!
b1000 %
1'
b1000 +
#834760000000
0!
0'
#834770000000
1!
b1001 %
1'
b1001 +
#834780000000
0!
0'
#834790000000
1!
b0 %
1'
b0 +
#834800000000
0!
0'
#834810000000
1!
1$
b1 %
1'
1*
b1 +
#834820000000
0!
0'
#834830000000
1!
b10 %
1'
b10 +
#834840000000
1"
1(
#834850000000
0!
0"
b100 &
0'
0(
b100 ,
#834860000000
1!
b11 %
1'
b11 +
#834870000000
0!
0'
#834880000000
1!
b100 %
1'
b100 +
#834890000000
0!
0'
#834900000000
1!
b101 %
1'
b101 +
#834910000000
0!
0'
#834920000000
1!
b110 %
1'
b110 +
#834930000000
0!
0'
#834940000000
1!
b111 %
1'
b111 +
#834950000000
0!
0'
#834960000000
1!
0$
b1000 %
1'
0*
b1000 +
#834970000000
0!
0'
#834980000000
1!
b1001 %
1'
b1001 +
#834990000000
0!
0'
#835000000000
1!
b0 %
1'
b0 +
#835010000000
0!
0'
#835020000000
1!
1$
b1 %
1'
1*
b1 +
#835030000000
0!
0'
#835040000000
1!
b10 %
1'
b10 +
#835050000000
0!
0'
#835060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#835070000000
0!
0'
#835080000000
1!
b100 %
1'
b100 +
#835090000000
0!
0'
#835100000000
1!
b101 %
1'
b101 +
#835110000000
0!
0'
#835120000000
1!
0$
b110 %
1'
0*
b110 +
#835130000000
0!
0'
#835140000000
1!
b111 %
1'
b111 +
#835150000000
0!
0'
#835160000000
1!
b1000 %
1'
b1000 +
#835170000000
0!
0'
#835180000000
1!
b1001 %
1'
b1001 +
#835190000000
0!
0'
#835200000000
1!
b0 %
1'
b0 +
#835210000000
0!
0'
#835220000000
1!
1$
b1 %
1'
1*
b1 +
#835230000000
0!
0'
#835240000000
1!
b10 %
1'
b10 +
#835250000000
0!
0'
#835260000000
1!
b11 %
1'
b11 +
#835270000000
1"
1(
#835280000000
0!
0"
b100 &
0'
0(
b100 ,
#835290000000
1!
b100 %
1'
b100 +
#835300000000
0!
0'
#835310000000
1!
b101 %
1'
b101 +
#835320000000
0!
0'
#835330000000
1!
b110 %
1'
b110 +
#835340000000
0!
0'
#835350000000
1!
b111 %
1'
b111 +
#835360000000
0!
0'
#835370000000
1!
0$
b1000 %
1'
0*
b1000 +
#835380000000
0!
0'
#835390000000
1!
b1001 %
1'
b1001 +
#835400000000
0!
0'
#835410000000
1!
b0 %
1'
b0 +
#835420000000
0!
0'
#835430000000
1!
1$
b1 %
1'
1*
b1 +
#835440000000
0!
0'
#835450000000
1!
b10 %
1'
b10 +
#835460000000
0!
0'
#835470000000
1!
b11 %
1'
b11 +
#835480000000
0!
0'
#835490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#835500000000
0!
0'
#835510000000
1!
b101 %
1'
b101 +
#835520000000
0!
0'
#835530000000
1!
0$
b110 %
1'
0*
b110 +
#835540000000
0!
0'
#835550000000
1!
b111 %
1'
b111 +
#835560000000
0!
0'
#835570000000
1!
b1000 %
1'
b1000 +
#835580000000
0!
0'
#835590000000
1!
b1001 %
1'
b1001 +
#835600000000
0!
0'
#835610000000
1!
b0 %
1'
b0 +
#835620000000
0!
0'
#835630000000
1!
1$
b1 %
1'
1*
b1 +
#835640000000
0!
0'
#835650000000
1!
b10 %
1'
b10 +
#835660000000
0!
0'
#835670000000
1!
b11 %
1'
b11 +
#835680000000
0!
0'
#835690000000
1!
b100 %
1'
b100 +
#835700000000
1"
1(
#835710000000
0!
0"
b100 &
0'
0(
b100 ,
#835720000000
1!
b101 %
1'
b101 +
#835730000000
0!
0'
#835740000000
1!
b110 %
1'
b110 +
#835750000000
0!
0'
#835760000000
1!
b111 %
1'
b111 +
#835770000000
0!
0'
#835780000000
1!
0$
b1000 %
1'
0*
b1000 +
#835790000000
0!
0'
#835800000000
1!
b1001 %
1'
b1001 +
#835810000000
0!
0'
#835820000000
1!
b0 %
1'
b0 +
#835830000000
0!
0'
#835840000000
1!
1$
b1 %
1'
1*
b1 +
#835850000000
0!
0'
#835860000000
1!
b10 %
1'
b10 +
#835870000000
0!
0'
#835880000000
1!
b11 %
1'
b11 +
#835890000000
0!
0'
#835900000000
1!
b100 %
1'
b100 +
#835910000000
0!
0'
#835920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#835930000000
0!
0'
#835940000000
1!
0$
b110 %
1'
0*
b110 +
#835950000000
0!
0'
#835960000000
1!
b111 %
1'
b111 +
#835970000000
0!
0'
#835980000000
1!
b1000 %
1'
b1000 +
#835990000000
0!
0'
#836000000000
1!
b1001 %
1'
b1001 +
#836010000000
0!
0'
#836020000000
1!
b0 %
1'
b0 +
#836030000000
0!
0'
#836040000000
1!
1$
b1 %
1'
1*
b1 +
#836050000000
0!
0'
#836060000000
1!
b10 %
1'
b10 +
#836070000000
0!
0'
#836080000000
1!
b11 %
1'
b11 +
#836090000000
0!
0'
#836100000000
1!
b100 %
1'
b100 +
#836110000000
0!
0'
#836120000000
1!
b101 %
1'
b101 +
#836130000000
1"
1(
#836140000000
0!
0"
b100 &
0'
0(
b100 ,
#836150000000
1!
b110 %
1'
b110 +
#836160000000
0!
0'
#836170000000
1!
b111 %
1'
b111 +
#836180000000
0!
0'
#836190000000
1!
0$
b1000 %
1'
0*
b1000 +
#836200000000
0!
0'
#836210000000
1!
b1001 %
1'
b1001 +
#836220000000
0!
0'
#836230000000
1!
b0 %
1'
b0 +
#836240000000
0!
0'
#836250000000
1!
1$
b1 %
1'
1*
b1 +
#836260000000
0!
0'
#836270000000
1!
b10 %
1'
b10 +
#836280000000
0!
0'
#836290000000
1!
b11 %
1'
b11 +
#836300000000
0!
0'
#836310000000
1!
b100 %
1'
b100 +
#836320000000
0!
0'
#836330000000
1!
b101 %
1'
b101 +
#836340000000
0!
0'
#836350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#836360000000
0!
0'
#836370000000
1!
b111 %
1'
b111 +
#836380000000
0!
0'
#836390000000
1!
b1000 %
1'
b1000 +
#836400000000
0!
0'
#836410000000
1!
b1001 %
1'
b1001 +
#836420000000
0!
0'
#836430000000
1!
b0 %
1'
b0 +
#836440000000
0!
0'
#836450000000
1!
1$
b1 %
1'
1*
b1 +
#836460000000
0!
0'
#836470000000
1!
b10 %
1'
b10 +
#836480000000
0!
0'
#836490000000
1!
b11 %
1'
b11 +
#836500000000
0!
0'
#836510000000
1!
b100 %
1'
b100 +
#836520000000
0!
0'
#836530000000
1!
b101 %
1'
b101 +
#836540000000
0!
0'
#836550000000
1!
0$
b110 %
1'
0*
b110 +
#836560000000
1"
1(
#836570000000
0!
0"
b100 &
0'
0(
b100 ,
#836580000000
1!
1$
b111 %
1'
1*
b111 +
#836590000000
0!
0'
#836600000000
1!
0$
b1000 %
1'
0*
b1000 +
#836610000000
0!
0'
#836620000000
1!
b1001 %
1'
b1001 +
#836630000000
0!
0'
#836640000000
1!
b0 %
1'
b0 +
#836650000000
0!
0'
#836660000000
1!
1$
b1 %
1'
1*
b1 +
#836670000000
0!
0'
#836680000000
1!
b10 %
1'
b10 +
#836690000000
0!
0'
#836700000000
1!
b11 %
1'
b11 +
#836710000000
0!
0'
#836720000000
1!
b100 %
1'
b100 +
#836730000000
0!
0'
#836740000000
1!
b101 %
1'
b101 +
#836750000000
0!
0'
#836760000000
1!
b110 %
1'
b110 +
#836770000000
0!
0'
#836780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#836790000000
0!
0'
#836800000000
1!
b1000 %
1'
b1000 +
#836810000000
0!
0'
#836820000000
1!
b1001 %
1'
b1001 +
#836830000000
0!
0'
#836840000000
1!
b0 %
1'
b0 +
#836850000000
0!
0'
#836860000000
1!
1$
b1 %
1'
1*
b1 +
#836870000000
0!
0'
#836880000000
1!
b10 %
1'
b10 +
#836890000000
0!
0'
#836900000000
1!
b11 %
1'
b11 +
#836910000000
0!
0'
#836920000000
1!
b100 %
1'
b100 +
#836930000000
0!
0'
#836940000000
1!
b101 %
1'
b101 +
#836950000000
0!
0'
#836960000000
1!
0$
b110 %
1'
0*
b110 +
#836970000000
0!
0'
#836980000000
1!
b111 %
1'
b111 +
#836990000000
1"
1(
#837000000000
0!
0"
b100 &
0'
0(
b100 ,
#837010000000
1!
b1000 %
1'
b1000 +
#837020000000
0!
0'
#837030000000
1!
b1001 %
1'
b1001 +
#837040000000
0!
0'
#837050000000
1!
b0 %
1'
b0 +
#837060000000
0!
0'
#837070000000
1!
1$
b1 %
1'
1*
b1 +
#837080000000
0!
0'
#837090000000
1!
b10 %
1'
b10 +
#837100000000
0!
0'
#837110000000
1!
b11 %
1'
b11 +
#837120000000
0!
0'
#837130000000
1!
b100 %
1'
b100 +
#837140000000
0!
0'
#837150000000
1!
b101 %
1'
b101 +
#837160000000
0!
0'
#837170000000
1!
b110 %
1'
b110 +
#837180000000
0!
0'
#837190000000
1!
b111 %
1'
b111 +
#837200000000
0!
0'
#837210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#837220000000
0!
0'
#837230000000
1!
b1001 %
1'
b1001 +
#837240000000
0!
0'
#837250000000
1!
b0 %
1'
b0 +
#837260000000
0!
0'
#837270000000
1!
1$
b1 %
1'
1*
b1 +
#837280000000
0!
0'
#837290000000
1!
b10 %
1'
b10 +
#837300000000
0!
0'
#837310000000
1!
b11 %
1'
b11 +
#837320000000
0!
0'
#837330000000
1!
b100 %
1'
b100 +
#837340000000
0!
0'
#837350000000
1!
b101 %
1'
b101 +
#837360000000
0!
0'
#837370000000
1!
0$
b110 %
1'
0*
b110 +
#837380000000
0!
0'
#837390000000
1!
b111 %
1'
b111 +
#837400000000
0!
0'
#837410000000
1!
b1000 %
1'
b1000 +
#837420000000
1"
1(
#837430000000
0!
0"
b100 &
0'
0(
b100 ,
#837440000000
1!
b1001 %
1'
b1001 +
#837450000000
0!
0'
#837460000000
1!
b0 %
1'
b0 +
#837470000000
0!
0'
#837480000000
1!
1$
b1 %
1'
1*
b1 +
#837490000000
0!
0'
#837500000000
1!
b10 %
1'
b10 +
#837510000000
0!
0'
#837520000000
1!
b11 %
1'
b11 +
#837530000000
0!
0'
#837540000000
1!
b100 %
1'
b100 +
#837550000000
0!
0'
#837560000000
1!
b101 %
1'
b101 +
#837570000000
0!
0'
#837580000000
1!
b110 %
1'
b110 +
#837590000000
0!
0'
#837600000000
1!
b111 %
1'
b111 +
#837610000000
0!
0'
#837620000000
1!
0$
b1000 %
1'
0*
b1000 +
#837630000000
0!
0'
#837640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#837650000000
0!
0'
#837660000000
1!
b0 %
1'
b0 +
#837670000000
0!
0'
#837680000000
1!
1$
b1 %
1'
1*
b1 +
#837690000000
0!
0'
#837700000000
1!
b10 %
1'
b10 +
#837710000000
0!
0'
#837720000000
1!
b11 %
1'
b11 +
#837730000000
0!
0'
#837740000000
1!
b100 %
1'
b100 +
#837750000000
0!
0'
#837760000000
1!
b101 %
1'
b101 +
#837770000000
0!
0'
#837780000000
1!
0$
b110 %
1'
0*
b110 +
#837790000000
0!
0'
#837800000000
1!
b111 %
1'
b111 +
#837810000000
0!
0'
#837820000000
1!
b1000 %
1'
b1000 +
#837830000000
0!
0'
#837840000000
1!
b1001 %
1'
b1001 +
#837850000000
1"
1(
#837860000000
0!
0"
b100 &
0'
0(
b100 ,
#837870000000
1!
b0 %
1'
b0 +
#837880000000
0!
0'
#837890000000
1!
1$
b1 %
1'
1*
b1 +
#837900000000
0!
0'
#837910000000
1!
b10 %
1'
b10 +
#837920000000
0!
0'
#837930000000
1!
b11 %
1'
b11 +
#837940000000
0!
0'
#837950000000
1!
b100 %
1'
b100 +
#837960000000
0!
0'
#837970000000
1!
b101 %
1'
b101 +
#837980000000
0!
0'
#837990000000
1!
b110 %
1'
b110 +
#838000000000
0!
0'
#838010000000
1!
b111 %
1'
b111 +
#838020000000
0!
0'
#838030000000
1!
0$
b1000 %
1'
0*
b1000 +
#838040000000
0!
0'
#838050000000
1!
b1001 %
1'
b1001 +
#838060000000
0!
0'
#838070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#838080000000
0!
0'
#838090000000
1!
1$
b1 %
1'
1*
b1 +
#838100000000
0!
0'
#838110000000
1!
b10 %
1'
b10 +
#838120000000
0!
0'
#838130000000
1!
b11 %
1'
b11 +
#838140000000
0!
0'
#838150000000
1!
b100 %
1'
b100 +
#838160000000
0!
0'
#838170000000
1!
b101 %
1'
b101 +
#838180000000
0!
0'
#838190000000
1!
0$
b110 %
1'
0*
b110 +
#838200000000
0!
0'
#838210000000
1!
b111 %
1'
b111 +
#838220000000
0!
0'
#838230000000
1!
b1000 %
1'
b1000 +
#838240000000
0!
0'
#838250000000
1!
b1001 %
1'
b1001 +
#838260000000
0!
0'
#838270000000
1!
b0 %
1'
b0 +
#838280000000
1"
1(
#838290000000
0!
0"
b100 &
0'
0(
b100 ,
#838300000000
1!
1$
b1 %
1'
1*
b1 +
#838310000000
0!
0'
#838320000000
1!
b10 %
1'
b10 +
#838330000000
0!
0'
#838340000000
1!
b11 %
1'
b11 +
#838350000000
0!
0'
#838360000000
1!
b100 %
1'
b100 +
#838370000000
0!
0'
#838380000000
1!
b101 %
1'
b101 +
#838390000000
0!
0'
#838400000000
1!
b110 %
1'
b110 +
#838410000000
0!
0'
#838420000000
1!
b111 %
1'
b111 +
#838430000000
0!
0'
#838440000000
1!
0$
b1000 %
1'
0*
b1000 +
#838450000000
0!
0'
#838460000000
1!
b1001 %
1'
b1001 +
#838470000000
0!
0'
#838480000000
1!
b0 %
1'
b0 +
#838490000000
0!
0'
#838500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#838510000000
0!
0'
#838520000000
1!
b10 %
1'
b10 +
#838530000000
0!
0'
#838540000000
1!
b11 %
1'
b11 +
#838550000000
0!
0'
#838560000000
1!
b100 %
1'
b100 +
#838570000000
0!
0'
#838580000000
1!
b101 %
1'
b101 +
#838590000000
0!
0'
#838600000000
1!
0$
b110 %
1'
0*
b110 +
#838610000000
0!
0'
#838620000000
1!
b111 %
1'
b111 +
#838630000000
0!
0'
#838640000000
1!
b1000 %
1'
b1000 +
#838650000000
0!
0'
#838660000000
1!
b1001 %
1'
b1001 +
#838670000000
0!
0'
#838680000000
1!
b0 %
1'
b0 +
#838690000000
0!
0'
#838700000000
1!
1$
b1 %
1'
1*
b1 +
#838710000000
1"
1(
#838720000000
0!
0"
b100 &
0'
0(
b100 ,
#838730000000
1!
b10 %
1'
b10 +
#838740000000
0!
0'
#838750000000
1!
b11 %
1'
b11 +
#838760000000
0!
0'
#838770000000
1!
b100 %
1'
b100 +
#838780000000
0!
0'
#838790000000
1!
b101 %
1'
b101 +
#838800000000
0!
0'
#838810000000
1!
b110 %
1'
b110 +
#838820000000
0!
0'
#838830000000
1!
b111 %
1'
b111 +
#838840000000
0!
0'
#838850000000
1!
0$
b1000 %
1'
0*
b1000 +
#838860000000
0!
0'
#838870000000
1!
b1001 %
1'
b1001 +
#838880000000
0!
0'
#838890000000
1!
b0 %
1'
b0 +
#838900000000
0!
0'
#838910000000
1!
1$
b1 %
1'
1*
b1 +
#838920000000
0!
0'
#838930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#838940000000
0!
0'
#838950000000
1!
b11 %
1'
b11 +
#838960000000
0!
0'
#838970000000
1!
b100 %
1'
b100 +
#838980000000
0!
0'
#838990000000
1!
b101 %
1'
b101 +
#839000000000
0!
0'
#839010000000
1!
0$
b110 %
1'
0*
b110 +
#839020000000
0!
0'
#839030000000
1!
b111 %
1'
b111 +
#839040000000
0!
0'
#839050000000
1!
b1000 %
1'
b1000 +
#839060000000
0!
0'
#839070000000
1!
b1001 %
1'
b1001 +
#839080000000
0!
0'
#839090000000
1!
b0 %
1'
b0 +
#839100000000
0!
0'
#839110000000
1!
1$
b1 %
1'
1*
b1 +
#839120000000
0!
0'
#839130000000
1!
b10 %
1'
b10 +
#839140000000
1"
1(
#839150000000
0!
0"
b100 &
0'
0(
b100 ,
#839160000000
1!
b11 %
1'
b11 +
#839170000000
0!
0'
#839180000000
1!
b100 %
1'
b100 +
#839190000000
0!
0'
#839200000000
1!
b101 %
1'
b101 +
#839210000000
0!
0'
#839220000000
1!
b110 %
1'
b110 +
#839230000000
0!
0'
#839240000000
1!
b111 %
1'
b111 +
#839250000000
0!
0'
#839260000000
1!
0$
b1000 %
1'
0*
b1000 +
#839270000000
0!
0'
#839280000000
1!
b1001 %
1'
b1001 +
#839290000000
0!
0'
#839300000000
1!
b0 %
1'
b0 +
#839310000000
0!
0'
#839320000000
1!
1$
b1 %
1'
1*
b1 +
#839330000000
0!
0'
#839340000000
1!
b10 %
1'
b10 +
#839350000000
0!
0'
#839360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#839370000000
0!
0'
#839380000000
1!
b100 %
1'
b100 +
#839390000000
0!
0'
#839400000000
1!
b101 %
1'
b101 +
#839410000000
0!
0'
#839420000000
1!
0$
b110 %
1'
0*
b110 +
#839430000000
0!
0'
#839440000000
1!
b111 %
1'
b111 +
#839450000000
0!
0'
#839460000000
1!
b1000 %
1'
b1000 +
#839470000000
0!
0'
#839480000000
1!
b1001 %
1'
b1001 +
#839490000000
0!
0'
#839500000000
1!
b0 %
1'
b0 +
#839510000000
0!
0'
#839520000000
1!
1$
b1 %
1'
1*
b1 +
#839530000000
0!
0'
#839540000000
1!
b10 %
1'
b10 +
#839550000000
0!
0'
#839560000000
1!
b11 %
1'
b11 +
#839570000000
1"
1(
#839580000000
0!
0"
b100 &
0'
0(
b100 ,
#839590000000
1!
b100 %
1'
b100 +
#839600000000
0!
0'
#839610000000
1!
b101 %
1'
b101 +
#839620000000
0!
0'
#839630000000
1!
b110 %
1'
b110 +
#839640000000
0!
0'
#839650000000
1!
b111 %
1'
b111 +
#839660000000
0!
0'
#839670000000
1!
0$
b1000 %
1'
0*
b1000 +
#839680000000
0!
0'
#839690000000
1!
b1001 %
1'
b1001 +
#839700000000
0!
0'
#839710000000
1!
b0 %
1'
b0 +
#839720000000
0!
0'
#839730000000
1!
1$
b1 %
1'
1*
b1 +
#839740000000
0!
0'
#839750000000
1!
b10 %
1'
b10 +
#839760000000
0!
0'
#839770000000
1!
b11 %
1'
b11 +
#839780000000
0!
0'
#839790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#839800000000
0!
0'
#839810000000
1!
b101 %
1'
b101 +
#839820000000
0!
0'
#839830000000
1!
0$
b110 %
1'
0*
b110 +
#839840000000
0!
0'
#839850000000
1!
b111 %
1'
b111 +
#839860000000
0!
0'
#839870000000
1!
b1000 %
1'
b1000 +
#839880000000
0!
0'
#839890000000
1!
b1001 %
1'
b1001 +
#839900000000
0!
0'
#839910000000
1!
b0 %
1'
b0 +
#839920000000
0!
0'
#839930000000
1!
1$
b1 %
1'
1*
b1 +
#839940000000
0!
0'
#839950000000
1!
b10 %
1'
b10 +
#839960000000
0!
0'
#839970000000
1!
b11 %
1'
b11 +
#839980000000
0!
0'
#839990000000
1!
b100 %
1'
b100 +
#840000000000
1"
1(
#840010000000
0!
0"
b100 &
0'
0(
b100 ,
#840020000000
1!
b101 %
1'
b101 +
#840030000000
0!
0'
#840040000000
1!
b110 %
1'
b110 +
#840050000000
0!
0'
#840060000000
1!
b111 %
1'
b111 +
#840070000000
0!
0'
#840080000000
1!
0$
b1000 %
1'
0*
b1000 +
#840090000000
0!
0'
#840100000000
1!
b1001 %
1'
b1001 +
#840110000000
0!
0'
#840120000000
1!
b0 %
1'
b0 +
#840130000000
0!
0'
#840140000000
1!
1$
b1 %
1'
1*
b1 +
#840150000000
0!
0'
#840160000000
1!
b10 %
1'
b10 +
#840170000000
0!
0'
#840180000000
1!
b11 %
1'
b11 +
#840190000000
0!
0'
#840200000000
1!
b100 %
1'
b100 +
#840210000000
0!
0'
#840220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#840230000000
0!
0'
#840240000000
1!
0$
b110 %
1'
0*
b110 +
#840250000000
0!
0'
#840260000000
1!
b111 %
1'
b111 +
#840270000000
0!
0'
#840280000000
1!
b1000 %
1'
b1000 +
#840290000000
0!
0'
#840300000000
1!
b1001 %
1'
b1001 +
#840310000000
0!
0'
#840320000000
1!
b0 %
1'
b0 +
#840330000000
0!
0'
#840340000000
1!
1$
b1 %
1'
1*
b1 +
#840350000000
0!
0'
#840360000000
1!
b10 %
1'
b10 +
#840370000000
0!
0'
#840380000000
1!
b11 %
1'
b11 +
#840390000000
0!
0'
#840400000000
1!
b100 %
1'
b100 +
#840410000000
0!
0'
#840420000000
1!
b101 %
1'
b101 +
#840430000000
1"
1(
#840440000000
0!
0"
b100 &
0'
0(
b100 ,
#840450000000
1!
b110 %
1'
b110 +
#840460000000
0!
0'
#840470000000
1!
b111 %
1'
b111 +
#840480000000
0!
0'
#840490000000
1!
0$
b1000 %
1'
0*
b1000 +
#840500000000
0!
0'
#840510000000
1!
b1001 %
1'
b1001 +
#840520000000
0!
0'
#840530000000
1!
b0 %
1'
b0 +
#840540000000
0!
0'
#840550000000
1!
1$
b1 %
1'
1*
b1 +
#840560000000
0!
0'
#840570000000
1!
b10 %
1'
b10 +
#840580000000
0!
0'
#840590000000
1!
b11 %
1'
b11 +
#840600000000
0!
0'
#840610000000
1!
b100 %
1'
b100 +
#840620000000
0!
0'
#840630000000
1!
b101 %
1'
b101 +
#840640000000
0!
0'
#840650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#840660000000
0!
0'
#840670000000
1!
b111 %
1'
b111 +
#840680000000
0!
0'
#840690000000
1!
b1000 %
1'
b1000 +
#840700000000
0!
0'
#840710000000
1!
b1001 %
1'
b1001 +
#840720000000
0!
0'
#840730000000
1!
b0 %
1'
b0 +
#840740000000
0!
0'
#840750000000
1!
1$
b1 %
1'
1*
b1 +
#840760000000
0!
0'
#840770000000
1!
b10 %
1'
b10 +
#840780000000
0!
0'
#840790000000
1!
b11 %
1'
b11 +
#840800000000
0!
0'
#840810000000
1!
b100 %
1'
b100 +
#840820000000
0!
0'
#840830000000
1!
b101 %
1'
b101 +
#840840000000
0!
0'
#840850000000
1!
0$
b110 %
1'
0*
b110 +
#840860000000
1"
1(
#840870000000
0!
0"
b100 &
0'
0(
b100 ,
#840880000000
1!
1$
b111 %
1'
1*
b111 +
#840890000000
0!
0'
#840900000000
1!
0$
b1000 %
1'
0*
b1000 +
#840910000000
0!
0'
#840920000000
1!
b1001 %
1'
b1001 +
#840930000000
0!
0'
#840940000000
1!
b0 %
1'
b0 +
#840950000000
0!
0'
#840960000000
1!
1$
b1 %
1'
1*
b1 +
#840970000000
0!
0'
#840980000000
1!
b10 %
1'
b10 +
#840990000000
0!
0'
#841000000000
1!
b11 %
1'
b11 +
#841010000000
0!
0'
#841020000000
1!
b100 %
1'
b100 +
#841030000000
0!
0'
#841040000000
1!
b101 %
1'
b101 +
#841050000000
0!
0'
#841060000000
1!
b110 %
1'
b110 +
#841070000000
0!
0'
#841080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#841090000000
0!
0'
#841100000000
1!
b1000 %
1'
b1000 +
#841110000000
0!
0'
#841120000000
1!
b1001 %
1'
b1001 +
#841130000000
0!
0'
#841140000000
1!
b0 %
1'
b0 +
#841150000000
0!
0'
#841160000000
1!
1$
b1 %
1'
1*
b1 +
#841170000000
0!
0'
#841180000000
1!
b10 %
1'
b10 +
#841190000000
0!
0'
#841200000000
1!
b11 %
1'
b11 +
#841210000000
0!
0'
#841220000000
1!
b100 %
1'
b100 +
#841230000000
0!
0'
#841240000000
1!
b101 %
1'
b101 +
#841250000000
0!
0'
#841260000000
1!
0$
b110 %
1'
0*
b110 +
#841270000000
0!
0'
#841280000000
1!
b111 %
1'
b111 +
#841290000000
1"
1(
#841300000000
0!
0"
b100 &
0'
0(
b100 ,
#841310000000
1!
b1000 %
1'
b1000 +
#841320000000
0!
0'
#841330000000
1!
b1001 %
1'
b1001 +
#841340000000
0!
0'
#841350000000
1!
b0 %
1'
b0 +
#841360000000
0!
0'
#841370000000
1!
1$
b1 %
1'
1*
b1 +
#841380000000
0!
0'
#841390000000
1!
b10 %
1'
b10 +
#841400000000
0!
0'
#841410000000
1!
b11 %
1'
b11 +
#841420000000
0!
0'
#841430000000
1!
b100 %
1'
b100 +
#841440000000
0!
0'
#841450000000
1!
b101 %
1'
b101 +
#841460000000
0!
0'
#841470000000
1!
b110 %
1'
b110 +
#841480000000
0!
0'
#841490000000
1!
b111 %
1'
b111 +
#841500000000
0!
0'
#841510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#841520000000
0!
0'
#841530000000
1!
b1001 %
1'
b1001 +
#841540000000
0!
0'
#841550000000
1!
b0 %
1'
b0 +
#841560000000
0!
0'
#841570000000
1!
1$
b1 %
1'
1*
b1 +
#841580000000
0!
0'
#841590000000
1!
b10 %
1'
b10 +
#841600000000
0!
0'
#841610000000
1!
b11 %
1'
b11 +
#841620000000
0!
0'
#841630000000
1!
b100 %
1'
b100 +
#841640000000
0!
0'
#841650000000
1!
b101 %
1'
b101 +
#841660000000
0!
0'
#841670000000
1!
0$
b110 %
1'
0*
b110 +
#841680000000
0!
0'
#841690000000
1!
b111 %
1'
b111 +
#841700000000
0!
0'
#841710000000
1!
b1000 %
1'
b1000 +
#841720000000
1"
1(
#841730000000
0!
0"
b100 &
0'
0(
b100 ,
#841740000000
1!
b1001 %
1'
b1001 +
#841750000000
0!
0'
#841760000000
1!
b0 %
1'
b0 +
#841770000000
0!
0'
#841780000000
1!
1$
b1 %
1'
1*
b1 +
#841790000000
0!
0'
#841800000000
1!
b10 %
1'
b10 +
#841810000000
0!
0'
#841820000000
1!
b11 %
1'
b11 +
#841830000000
0!
0'
#841840000000
1!
b100 %
1'
b100 +
#841850000000
0!
0'
#841860000000
1!
b101 %
1'
b101 +
#841870000000
0!
0'
#841880000000
1!
b110 %
1'
b110 +
#841890000000
0!
0'
#841900000000
1!
b111 %
1'
b111 +
#841910000000
0!
0'
#841920000000
1!
0$
b1000 %
1'
0*
b1000 +
#841930000000
0!
0'
#841940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#841950000000
0!
0'
#841960000000
1!
b0 %
1'
b0 +
#841970000000
0!
0'
#841980000000
1!
1$
b1 %
1'
1*
b1 +
#841990000000
0!
0'
#842000000000
1!
b10 %
1'
b10 +
#842010000000
0!
0'
#842020000000
1!
b11 %
1'
b11 +
#842030000000
0!
0'
#842040000000
1!
b100 %
1'
b100 +
#842050000000
0!
0'
#842060000000
1!
b101 %
1'
b101 +
#842070000000
0!
0'
#842080000000
1!
0$
b110 %
1'
0*
b110 +
#842090000000
0!
0'
#842100000000
1!
b111 %
1'
b111 +
#842110000000
0!
0'
#842120000000
1!
b1000 %
1'
b1000 +
#842130000000
0!
0'
#842140000000
1!
b1001 %
1'
b1001 +
#842150000000
1"
1(
#842160000000
0!
0"
b100 &
0'
0(
b100 ,
#842170000000
1!
b0 %
1'
b0 +
#842180000000
0!
0'
#842190000000
1!
1$
b1 %
1'
1*
b1 +
#842200000000
0!
0'
#842210000000
1!
b10 %
1'
b10 +
#842220000000
0!
0'
#842230000000
1!
b11 %
1'
b11 +
#842240000000
0!
0'
#842250000000
1!
b100 %
1'
b100 +
#842260000000
0!
0'
#842270000000
1!
b101 %
1'
b101 +
#842280000000
0!
0'
#842290000000
1!
b110 %
1'
b110 +
#842300000000
0!
0'
#842310000000
1!
b111 %
1'
b111 +
#842320000000
0!
0'
#842330000000
1!
0$
b1000 %
1'
0*
b1000 +
#842340000000
0!
0'
#842350000000
1!
b1001 %
1'
b1001 +
#842360000000
0!
0'
#842370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#842380000000
0!
0'
#842390000000
1!
1$
b1 %
1'
1*
b1 +
#842400000000
0!
0'
#842410000000
1!
b10 %
1'
b10 +
#842420000000
0!
0'
#842430000000
1!
b11 %
1'
b11 +
#842440000000
0!
0'
#842450000000
1!
b100 %
1'
b100 +
#842460000000
0!
0'
#842470000000
1!
b101 %
1'
b101 +
#842480000000
0!
0'
#842490000000
1!
0$
b110 %
1'
0*
b110 +
#842500000000
0!
0'
#842510000000
1!
b111 %
1'
b111 +
#842520000000
0!
0'
#842530000000
1!
b1000 %
1'
b1000 +
#842540000000
0!
0'
#842550000000
1!
b1001 %
1'
b1001 +
#842560000000
0!
0'
#842570000000
1!
b0 %
1'
b0 +
#842580000000
1"
1(
#842590000000
0!
0"
b100 &
0'
0(
b100 ,
#842600000000
1!
1$
b1 %
1'
1*
b1 +
#842610000000
0!
0'
#842620000000
1!
b10 %
1'
b10 +
#842630000000
0!
0'
#842640000000
1!
b11 %
1'
b11 +
#842650000000
0!
0'
#842660000000
1!
b100 %
1'
b100 +
#842670000000
0!
0'
#842680000000
1!
b101 %
1'
b101 +
#842690000000
0!
0'
#842700000000
1!
b110 %
1'
b110 +
#842710000000
0!
0'
#842720000000
1!
b111 %
1'
b111 +
#842730000000
0!
0'
#842740000000
1!
0$
b1000 %
1'
0*
b1000 +
#842750000000
0!
0'
#842760000000
1!
b1001 %
1'
b1001 +
#842770000000
0!
0'
#842780000000
1!
b0 %
1'
b0 +
#842790000000
0!
0'
#842800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#842810000000
0!
0'
#842820000000
1!
b10 %
1'
b10 +
#842830000000
0!
0'
#842840000000
1!
b11 %
1'
b11 +
#842850000000
0!
0'
#842860000000
1!
b100 %
1'
b100 +
#842870000000
0!
0'
#842880000000
1!
b101 %
1'
b101 +
#842890000000
0!
0'
#842900000000
1!
0$
b110 %
1'
0*
b110 +
#842910000000
0!
0'
#842920000000
1!
b111 %
1'
b111 +
#842930000000
0!
0'
#842940000000
1!
b1000 %
1'
b1000 +
#842950000000
0!
0'
#842960000000
1!
b1001 %
1'
b1001 +
#842970000000
0!
0'
#842980000000
1!
b0 %
1'
b0 +
#842990000000
0!
0'
#843000000000
1!
1$
b1 %
1'
1*
b1 +
#843010000000
1"
1(
#843020000000
0!
0"
b100 &
0'
0(
b100 ,
#843030000000
1!
b10 %
1'
b10 +
#843040000000
0!
0'
#843050000000
1!
b11 %
1'
b11 +
#843060000000
0!
0'
#843070000000
1!
b100 %
1'
b100 +
#843080000000
0!
0'
#843090000000
1!
b101 %
1'
b101 +
#843100000000
0!
0'
#843110000000
1!
b110 %
1'
b110 +
#843120000000
0!
0'
#843130000000
1!
b111 %
1'
b111 +
#843140000000
0!
0'
#843150000000
1!
0$
b1000 %
1'
0*
b1000 +
#843160000000
0!
0'
#843170000000
1!
b1001 %
1'
b1001 +
#843180000000
0!
0'
#843190000000
1!
b0 %
1'
b0 +
#843200000000
0!
0'
#843210000000
1!
1$
b1 %
1'
1*
b1 +
#843220000000
0!
0'
#843230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#843240000000
0!
0'
#843250000000
1!
b11 %
1'
b11 +
#843260000000
0!
0'
#843270000000
1!
b100 %
1'
b100 +
#843280000000
0!
0'
#843290000000
1!
b101 %
1'
b101 +
#843300000000
0!
0'
#843310000000
1!
0$
b110 %
1'
0*
b110 +
#843320000000
0!
0'
#843330000000
1!
b111 %
1'
b111 +
#843340000000
0!
0'
#843350000000
1!
b1000 %
1'
b1000 +
#843360000000
0!
0'
#843370000000
1!
b1001 %
1'
b1001 +
#843380000000
0!
0'
#843390000000
1!
b0 %
1'
b0 +
#843400000000
0!
0'
#843410000000
1!
1$
b1 %
1'
1*
b1 +
#843420000000
0!
0'
#843430000000
1!
b10 %
1'
b10 +
#843440000000
1"
1(
#843450000000
0!
0"
b100 &
0'
0(
b100 ,
#843460000000
1!
b11 %
1'
b11 +
#843470000000
0!
0'
#843480000000
1!
b100 %
1'
b100 +
#843490000000
0!
0'
#843500000000
1!
b101 %
1'
b101 +
#843510000000
0!
0'
#843520000000
1!
b110 %
1'
b110 +
#843530000000
0!
0'
#843540000000
1!
b111 %
1'
b111 +
#843550000000
0!
0'
#843560000000
1!
0$
b1000 %
1'
0*
b1000 +
#843570000000
0!
0'
#843580000000
1!
b1001 %
1'
b1001 +
#843590000000
0!
0'
#843600000000
1!
b0 %
1'
b0 +
#843610000000
0!
0'
#843620000000
1!
1$
b1 %
1'
1*
b1 +
#843630000000
0!
0'
#843640000000
1!
b10 %
1'
b10 +
#843650000000
0!
0'
#843660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#843670000000
0!
0'
#843680000000
1!
b100 %
1'
b100 +
#843690000000
0!
0'
#843700000000
1!
b101 %
1'
b101 +
#843710000000
0!
0'
#843720000000
1!
0$
b110 %
1'
0*
b110 +
#843730000000
0!
0'
#843740000000
1!
b111 %
1'
b111 +
#843750000000
0!
0'
#843760000000
1!
b1000 %
1'
b1000 +
#843770000000
0!
0'
#843780000000
1!
b1001 %
1'
b1001 +
#843790000000
0!
0'
#843800000000
1!
b0 %
1'
b0 +
#843810000000
0!
0'
#843820000000
1!
1$
b1 %
1'
1*
b1 +
#843830000000
0!
0'
#843840000000
1!
b10 %
1'
b10 +
#843850000000
0!
0'
#843860000000
1!
b11 %
1'
b11 +
#843870000000
1"
1(
#843880000000
0!
0"
b100 &
0'
0(
b100 ,
#843890000000
1!
b100 %
1'
b100 +
#843900000000
0!
0'
#843910000000
1!
b101 %
1'
b101 +
#843920000000
0!
0'
#843930000000
1!
b110 %
1'
b110 +
#843940000000
0!
0'
#843950000000
1!
b111 %
1'
b111 +
#843960000000
0!
0'
#843970000000
1!
0$
b1000 %
1'
0*
b1000 +
#843980000000
0!
0'
#843990000000
1!
b1001 %
1'
b1001 +
#844000000000
0!
0'
#844010000000
1!
b0 %
1'
b0 +
#844020000000
0!
0'
#844030000000
1!
1$
b1 %
1'
1*
b1 +
#844040000000
0!
0'
#844050000000
1!
b10 %
1'
b10 +
#844060000000
0!
0'
#844070000000
1!
b11 %
1'
b11 +
#844080000000
0!
0'
#844090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#844100000000
0!
0'
#844110000000
1!
b101 %
1'
b101 +
#844120000000
0!
0'
#844130000000
1!
0$
b110 %
1'
0*
b110 +
#844140000000
0!
0'
#844150000000
1!
b111 %
1'
b111 +
#844160000000
0!
0'
#844170000000
1!
b1000 %
1'
b1000 +
#844180000000
0!
0'
#844190000000
1!
b1001 %
1'
b1001 +
#844200000000
0!
0'
#844210000000
1!
b0 %
1'
b0 +
#844220000000
0!
0'
#844230000000
1!
1$
b1 %
1'
1*
b1 +
#844240000000
0!
0'
#844250000000
1!
b10 %
1'
b10 +
#844260000000
0!
0'
#844270000000
1!
b11 %
1'
b11 +
#844280000000
0!
0'
#844290000000
1!
b100 %
1'
b100 +
#844300000000
1"
1(
#844310000000
0!
0"
b100 &
0'
0(
b100 ,
#844320000000
1!
b101 %
1'
b101 +
#844330000000
0!
0'
#844340000000
1!
b110 %
1'
b110 +
#844350000000
0!
0'
#844360000000
1!
b111 %
1'
b111 +
#844370000000
0!
0'
#844380000000
1!
0$
b1000 %
1'
0*
b1000 +
#844390000000
0!
0'
#844400000000
1!
b1001 %
1'
b1001 +
#844410000000
0!
0'
#844420000000
1!
b0 %
1'
b0 +
#844430000000
0!
0'
#844440000000
1!
1$
b1 %
1'
1*
b1 +
#844450000000
0!
0'
#844460000000
1!
b10 %
1'
b10 +
#844470000000
0!
0'
#844480000000
1!
b11 %
1'
b11 +
#844490000000
0!
0'
#844500000000
1!
b100 %
1'
b100 +
#844510000000
0!
0'
#844520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#844530000000
0!
0'
#844540000000
1!
0$
b110 %
1'
0*
b110 +
#844550000000
0!
0'
#844560000000
1!
b111 %
1'
b111 +
#844570000000
0!
0'
#844580000000
1!
b1000 %
1'
b1000 +
#844590000000
0!
0'
#844600000000
1!
b1001 %
1'
b1001 +
#844610000000
0!
0'
#844620000000
1!
b0 %
1'
b0 +
#844630000000
0!
0'
#844640000000
1!
1$
b1 %
1'
1*
b1 +
#844650000000
0!
0'
#844660000000
1!
b10 %
1'
b10 +
#844670000000
0!
0'
#844680000000
1!
b11 %
1'
b11 +
#844690000000
0!
0'
#844700000000
1!
b100 %
1'
b100 +
#844710000000
0!
0'
#844720000000
1!
b101 %
1'
b101 +
#844730000000
1"
1(
#844740000000
0!
0"
b100 &
0'
0(
b100 ,
#844750000000
1!
b110 %
1'
b110 +
#844760000000
0!
0'
#844770000000
1!
b111 %
1'
b111 +
#844780000000
0!
0'
#844790000000
1!
0$
b1000 %
1'
0*
b1000 +
#844800000000
0!
0'
#844810000000
1!
b1001 %
1'
b1001 +
#844820000000
0!
0'
#844830000000
1!
b0 %
1'
b0 +
#844840000000
0!
0'
#844850000000
1!
1$
b1 %
1'
1*
b1 +
#844860000000
0!
0'
#844870000000
1!
b10 %
1'
b10 +
#844880000000
0!
0'
#844890000000
1!
b11 %
1'
b11 +
#844900000000
0!
0'
#844910000000
1!
b100 %
1'
b100 +
#844920000000
0!
0'
#844930000000
1!
b101 %
1'
b101 +
#844940000000
0!
0'
#844950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#844960000000
0!
0'
#844970000000
1!
b111 %
1'
b111 +
#844980000000
0!
0'
#844990000000
1!
b1000 %
1'
b1000 +
#845000000000
0!
0'
#845010000000
1!
b1001 %
1'
b1001 +
#845020000000
0!
0'
#845030000000
1!
b0 %
1'
b0 +
#845040000000
0!
0'
#845050000000
1!
1$
b1 %
1'
1*
b1 +
#845060000000
0!
0'
#845070000000
1!
b10 %
1'
b10 +
#845080000000
0!
0'
#845090000000
1!
b11 %
1'
b11 +
#845100000000
0!
0'
#845110000000
1!
b100 %
1'
b100 +
#845120000000
0!
0'
#845130000000
1!
b101 %
1'
b101 +
#845140000000
0!
0'
#845150000000
1!
0$
b110 %
1'
0*
b110 +
#845160000000
1"
1(
#845170000000
0!
0"
b100 &
0'
0(
b100 ,
#845180000000
1!
1$
b111 %
1'
1*
b111 +
#845190000000
0!
0'
#845200000000
1!
0$
b1000 %
1'
0*
b1000 +
#845210000000
0!
0'
#845220000000
1!
b1001 %
1'
b1001 +
#845230000000
0!
0'
#845240000000
1!
b0 %
1'
b0 +
#845250000000
0!
0'
#845260000000
1!
1$
b1 %
1'
1*
b1 +
#845270000000
0!
0'
#845280000000
1!
b10 %
1'
b10 +
#845290000000
0!
0'
#845300000000
1!
b11 %
1'
b11 +
#845310000000
0!
0'
#845320000000
1!
b100 %
1'
b100 +
#845330000000
0!
0'
#845340000000
1!
b101 %
1'
b101 +
#845350000000
0!
0'
#845360000000
1!
b110 %
1'
b110 +
#845370000000
0!
0'
#845380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#845390000000
0!
0'
#845400000000
1!
b1000 %
1'
b1000 +
#845410000000
0!
0'
#845420000000
1!
b1001 %
1'
b1001 +
#845430000000
0!
0'
#845440000000
1!
b0 %
1'
b0 +
#845450000000
0!
0'
#845460000000
1!
1$
b1 %
1'
1*
b1 +
#845470000000
0!
0'
#845480000000
1!
b10 %
1'
b10 +
#845490000000
0!
0'
#845500000000
1!
b11 %
1'
b11 +
#845510000000
0!
0'
#845520000000
1!
b100 %
1'
b100 +
#845530000000
0!
0'
#845540000000
1!
b101 %
1'
b101 +
#845550000000
0!
0'
#845560000000
1!
0$
b110 %
1'
0*
b110 +
#845570000000
0!
0'
#845580000000
1!
b111 %
1'
b111 +
#845590000000
1"
1(
#845600000000
0!
0"
b100 &
0'
0(
b100 ,
#845610000000
1!
b1000 %
1'
b1000 +
#845620000000
0!
0'
#845630000000
1!
b1001 %
1'
b1001 +
#845640000000
0!
0'
#845650000000
1!
b0 %
1'
b0 +
#845660000000
0!
0'
#845670000000
1!
1$
b1 %
1'
1*
b1 +
#845680000000
0!
0'
#845690000000
1!
b10 %
1'
b10 +
#845700000000
0!
0'
#845710000000
1!
b11 %
1'
b11 +
#845720000000
0!
0'
#845730000000
1!
b100 %
1'
b100 +
#845740000000
0!
0'
#845750000000
1!
b101 %
1'
b101 +
#845760000000
0!
0'
#845770000000
1!
b110 %
1'
b110 +
#845780000000
0!
0'
#845790000000
1!
b111 %
1'
b111 +
#845800000000
0!
0'
#845810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#845820000000
0!
0'
#845830000000
1!
b1001 %
1'
b1001 +
#845840000000
0!
0'
#845850000000
1!
b0 %
1'
b0 +
#845860000000
0!
0'
#845870000000
1!
1$
b1 %
1'
1*
b1 +
#845880000000
0!
0'
#845890000000
1!
b10 %
1'
b10 +
#845900000000
0!
0'
#845910000000
1!
b11 %
1'
b11 +
#845920000000
0!
0'
#845930000000
1!
b100 %
1'
b100 +
#845940000000
0!
0'
#845950000000
1!
b101 %
1'
b101 +
#845960000000
0!
0'
#845970000000
1!
0$
b110 %
1'
0*
b110 +
#845980000000
0!
0'
#845990000000
1!
b111 %
1'
b111 +
#846000000000
0!
0'
#846010000000
1!
b1000 %
1'
b1000 +
#846020000000
1"
1(
#846030000000
0!
0"
b100 &
0'
0(
b100 ,
#846040000000
1!
b1001 %
1'
b1001 +
#846050000000
0!
0'
#846060000000
1!
b0 %
1'
b0 +
#846070000000
0!
0'
#846080000000
1!
1$
b1 %
1'
1*
b1 +
#846090000000
0!
0'
#846100000000
1!
b10 %
1'
b10 +
#846110000000
0!
0'
#846120000000
1!
b11 %
1'
b11 +
#846130000000
0!
0'
#846140000000
1!
b100 %
1'
b100 +
#846150000000
0!
0'
#846160000000
1!
b101 %
1'
b101 +
#846170000000
0!
0'
#846180000000
1!
b110 %
1'
b110 +
#846190000000
0!
0'
#846200000000
1!
b111 %
1'
b111 +
#846210000000
0!
0'
#846220000000
1!
0$
b1000 %
1'
0*
b1000 +
#846230000000
0!
0'
#846240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#846250000000
0!
0'
#846260000000
1!
b0 %
1'
b0 +
#846270000000
0!
0'
#846280000000
1!
1$
b1 %
1'
1*
b1 +
#846290000000
0!
0'
#846300000000
1!
b10 %
1'
b10 +
#846310000000
0!
0'
#846320000000
1!
b11 %
1'
b11 +
#846330000000
0!
0'
#846340000000
1!
b100 %
1'
b100 +
#846350000000
0!
0'
#846360000000
1!
b101 %
1'
b101 +
#846370000000
0!
0'
#846380000000
1!
0$
b110 %
1'
0*
b110 +
#846390000000
0!
0'
#846400000000
1!
b111 %
1'
b111 +
#846410000000
0!
0'
#846420000000
1!
b1000 %
1'
b1000 +
#846430000000
0!
0'
#846440000000
1!
b1001 %
1'
b1001 +
#846450000000
1"
1(
#846460000000
0!
0"
b100 &
0'
0(
b100 ,
#846470000000
1!
b0 %
1'
b0 +
#846480000000
0!
0'
#846490000000
1!
1$
b1 %
1'
1*
b1 +
#846500000000
0!
0'
#846510000000
1!
b10 %
1'
b10 +
#846520000000
0!
0'
#846530000000
1!
b11 %
1'
b11 +
#846540000000
0!
0'
#846550000000
1!
b100 %
1'
b100 +
#846560000000
0!
0'
#846570000000
1!
b101 %
1'
b101 +
#846580000000
0!
0'
#846590000000
1!
b110 %
1'
b110 +
#846600000000
0!
0'
#846610000000
1!
b111 %
1'
b111 +
#846620000000
0!
0'
#846630000000
1!
0$
b1000 %
1'
0*
b1000 +
#846640000000
0!
0'
#846650000000
1!
b1001 %
1'
b1001 +
#846660000000
0!
0'
#846670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#846680000000
0!
0'
#846690000000
1!
1$
b1 %
1'
1*
b1 +
#846700000000
0!
0'
#846710000000
1!
b10 %
1'
b10 +
#846720000000
0!
0'
#846730000000
1!
b11 %
1'
b11 +
#846740000000
0!
0'
#846750000000
1!
b100 %
1'
b100 +
#846760000000
0!
0'
#846770000000
1!
b101 %
1'
b101 +
#846780000000
0!
0'
#846790000000
1!
0$
b110 %
1'
0*
b110 +
#846800000000
0!
0'
#846810000000
1!
b111 %
1'
b111 +
#846820000000
0!
0'
#846830000000
1!
b1000 %
1'
b1000 +
#846840000000
0!
0'
#846850000000
1!
b1001 %
1'
b1001 +
#846860000000
0!
0'
#846870000000
1!
b0 %
1'
b0 +
#846880000000
1"
1(
#846890000000
0!
0"
b100 &
0'
0(
b100 ,
#846900000000
1!
1$
b1 %
1'
1*
b1 +
#846910000000
0!
0'
#846920000000
1!
b10 %
1'
b10 +
#846930000000
0!
0'
#846940000000
1!
b11 %
1'
b11 +
#846950000000
0!
0'
#846960000000
1!
b100 %
1'
b100 +
#846970000000
0!
0'
#846980000000
1!
b101 %
1'
b101 +
#846990000000
0!
0'
#847000000000
1!
b110 %
1'
b110 +
#847010000000
0!
0'
#847020000000
1!
b111 %
1'
b111 +
#847030000000
0!
0'
#847040000000
1!
0$
b1000 %
1'
0*
b1000 +
#847050000000
0!
0'
#847060000000
1!
b1001 %
1'
b1001 +
#847070000000
0!
0'
#847080000000
1!
b0 %
1'
b0 +
#847090000000
0!
0'
#847100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#847110000000
0!
0'
#847120000000
1!
b10 %
1'
b10 +
#847130000000
0!
0'
#847140000000
1!
b11 %
1'
b11 +
#847150000000
0!
0'
#847160000000
1!
b100 %
1'
b100 +
#847170000000
0!
0'
#847180000000
1!
b101 %
1'
b101 +
#847190000000
0!
0'
#847200000000
1!
0$
b110 %
1'
0*
b110 +
#847210000000
0!
0'
#847220000000
1!
b111 %
1'
b111 +
#847230000000
0!
0'
#847240000000
1!
b1000 %
1'
b1000 +
#847250000000
0!
0'
#847260000000
1!
b1001 %
1'
b1001 +
#847270000000
0!
0'
#847280000000
1!
b0 %
1'
b0 +
#847290000000
0!
0'
#847300000000
1!
1$
b1 %
1'
1*
b1 +
#847310000000
1"
1(
#847320000000
0!
0"
b100 &
0'
0(
b100 ,
#847330000000
1!
b10 %
1'
b10 +
#847340000000
0!
0'
#847350000000
1!
b11 %
1'
b11 +
#847360000000
0!
0'
#847370000000
1!
b100 %
1'
b100 +
#847380000000
0!
0'
#847390000000
1!
b101 %
1'
b101 +
#847400000000
0!
0'
#847410000000
1!
b110 %
1'
b110 +
#847420000000
0!
0'
#847430000000
1!
b111 %
1'
b111 +
#847440000000
0!
0'
#847450000000
1!
0$
b1000 %
1'
0*
b1000 +
#847460000000
0!
0'
#847470000000
1!
b1001 %
1'
b1001 +
#847480000000
0!
0'
#847490000000
1!
b0 %
1'
b0 +
#847500000000
0!
0'
#847510000000
1!
1$
b1 %
1'
1*
b1 +
#847520000000
0!
0'
#847530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#847540000000
0!
0'
#847550000000
1!
b11 %
1'
b11 +
#847560000000
0!
0'
#847570000000
1!
b100 %
1'
b100 +
#847580000000
0!
0'
#847590000000
1!
b101 %
1'
b101 +
#847600000000
0!
0'
#847610000000
1!
0$
b110 %
1'
0*
b110 +
#847620000000
0!
0'
#847630000000
1!
b111 %
1'
b111 +
#847640000000
0!
0'
#847650000000
1!
b1000 %
1'
b1000 +
#847660000000
0!
0'
#847670000000
1!
b1001 %
1'
b1001 +
#847680000000
0!
0'
#847690000000
1!
b0 %
1'
b0 +
#847700000000
0!
0'
#847710000000
1!
1$
b1 %
1'
1*
b1 +
#847720000000
0!
0'
#847730000000
1!
b10 %
1'
b10 +
#847740000000
1"
1(
#847750000000
0!
0"
b100 &
0'
0(
b100 ,
#847760000000
1!
b11 %
1'
b11 +
#847770000000
0!
0'
#847780000000
1!
b100 %
1'
b100 +
#847790000000
0!
0'
#847800000000
1!
b101 %
1'
b101 +
#847810000000
0!
0'
#847820000000
1!
b110 %
1'
b110 +
#847830000000
0!
0'
#847840000000
1!
b111 %
1'
b111 +
#847850000000
0!
0'
#847860000000
1!
0$
b1000 %
1'
0*
b1000 +
#847870000000
0!
0'
#847880000000
1!
b1001 %
1'
b1001 +
#847890000000
0!
0'
#847900000000
1!
b0 %
1'
b0 +
#847910000000
0!
0'
#847920000000
1!
1$
b1 %
1'
1*
b1 +
#847930000000
0!
0'
#847940000000
1!
b10 %
1'
b10 +
#847950000000
0!
0'
#847960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#847970000000
0!
0'
#847980000000
1!
b100 %
1'
b100 +
#847990000000
0!
0'
#848000000000
1!
b101 %
1'
b101 +
#848010000000
0!
0'
#848020000000
1!
0$
b110 %
1'
0*
b110 +
#848030000000
0!
0'
#848040000000
1!
b111 %
1'
b111 +
#848050000000
0!
0'
#848060000000
1!
b1000 %
1'
b1000 +
#848070000000
0!
0'
#848080000000
1!
b1001 %
1'
b1001 +
#848090000000
0!
0'
#848100000000
1!
b0 %
1'
b0 +
#848110000000
0!
0'
#848120000000
1!
1$
b1 %
1'
1*
b1 +
#848130000000
0!
0'
#848140000000
1!
b10 %
1'
b10 +
#848150000000
0!
0'
#848160000000
1!
b11 %
1'
b11 +
#848170000000
1"
1(
#848180000000
0!
0"
b100 &
0'
0(
b100 ,
#848190000000
1!
b100 %
1'
b100 +
#848200000000
0!
0'
#848210000000
1!
b101 %
1'
b101 +
#848220000000
0!
0'
#848230000000
1!
b110 %
1'
b110 +
#848240000000
0!
0'
#848250000000
1!
b111 %
1'
b111 +
#848260000000
0!
0'
#848270000000
1!
0$
b1000 %
1'
0*
b1000 +
#848280000000
0!
0'
#848290000000
1!
b1001 %
1'
b1001 +
#848300000000
0!
0'
#848310000000
1!
b0 %
1'
b0 +
#848320000000
0!
0'
#848330000000
1!
1$
b1 %
1'
1*
b1 +
#848340000000
0!
0'
#848350000000
1!
b10 %
1'
b10 +
#848360000000
0!
0'
#848370000000
1!
b11 %
1'
b11 +
#848380000000
0!
0'
#848390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#848400000000
0!
0'
#848410000000
1!
b101 %
1'
b101 +
#848420000000
0!
0'
#848430000000
1!
0$
b110 %
1'
0*
b110 +
#848440000000
0!
0'
#848450000000
1!
b111 %
1'
b111 +
#848460000000
0!
0'
#848470000000
1!
b1000 %
1'
b1000 +
#848480000000
0!
0'
#848490000000
1!
b1001 %
1'
b1001 +
#848500000000
0!
0'
#848510000000
1!
b0 %
1'
b0 +
#848520000000
0!
0'
#848530000000
1!
1$
b1 %
1'
1*
b1 +
#848540000000
0!
0'
#848550000000
1!
b10 %
1'
b10 +
#848560000000
0!
0'
#848570000000
1!
b11 %
1'
b11 +
#848580000000
0!
0'
#848590000000
1!
b100 %
1'
b100 +
#848600000000
1"
1(
#848610000000
0!
0"
b100 &
0'
0(
b100 ,
#848620000000
1!
b101 %
1'
b101 +
#848630000000
0!
0'
#848640000000
1!
b110 %
1'
b110 +
#848650000000
0!
0'
#848660000000
1!
b111 %
1'
b111 +
#848670000000
0!
0'
#848680000000
1!
0$
b1000 %
1'
0*
b1000 +
#848690000000
0!
0'
#848700000000
1!
b1001 %
1'
b1001 +
#848710000000
0!
0'
#848720000000
1!
b0 %
1'
b0 +
#848730000000
0!
0'
#848740000000
1!
1$
b1 %
1'
1*
b1 +
#848750000000
0!
0'
#848760000000
1!
b10 %
1'
b10 +
#848770000000
0!
0'
#848780000000
1!
b11 %
1'
b11 +
#848790000000
0!
0'
#848800000000
1!
b100 %
1'
b100 +
#848810000000
0!
0'
#848820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#848830000000
0!
0'
#848840000000
1!
0$
b110 %
1'
0*
b110 +
#848850000000
0!
0'
#848860000000
1!
b111 %
1'
b111 +
#848870000000
0!
0'
#848880000000
1!
b1000 %
1'
b1000 +
#848890000000
0!
0'
#848900000000
1!
b1001 %
1'
b1001 +
#848910000000
0!
0'
#848920000000
1!
b0 %
1'
b0 +
#848930000000
0!
0'
#848940000000
1!
1$
b1 %
1'
1*
b1 +
#848950000000
0!
0'
#848960000000
1!
b10 %
1'
b10 +
#848970000000
0!
0'
#848980000000
1!
b11 %
1'
b11 +
#848990000000
0!
0'
#849000000000
1!
b100 %
1'
b100 +
#849010000000
0!
0'
#849020000000
1!
b101 %
1'
b101 +
#849030000000
1"
1(
#849040000000
0!
0"
b100 &
0'
0(
b100 ,
#849050000000
1!
b110 %
1'
b110 +
#849060000000
0!
0'
#849070000000
1!
b111 %
1'
b111 +
#849080000000
0!
0'
#849090000000
1!
0$
b1000 %
1'
0*
b1000 +
#849100000000
0!
0'
#849110000000
1!
b1001 %
1'
b1001 +
#849120000000
0!
0'
#849130000000
1!
b0 %
1'
b0 +
#849140000000
0!
0'
#849150000000
1!
1$
b1 %
1'
1*
b1 +
#849160000000
0!
0'
#849170000000
1!
b10 %
1'
b10 +
#849180000000
0!
0'
#849190000000
1!
b11 %
1'
b11 +
#849200000000
0!
0'
#849210000000
1!
b100 %
1'
b100 +
#849220000000
0!
0'
#849230000000
1!
b101 %
1'
b101 +
#849240000000
0!
0'
#849250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#849260000000
0!
0'
#849270000000
1!
b111 %
1'
b111 +
#849280000000
0!
0'
#849290000000
1!
b1000 %
1'
b1000 +
#849300000000
0!
0'
#849310000000
1!
b1001 %
1'
b1001 +
#849320000000
0!
0'
#849330000000
1!
b0 %
1'
b0 +
#849340000000
0!
0'
#849350000000
1!
1$
b1 %
1'
1*
b1 +
#849360000000
0!
0'
#849370000000
1!
b10 %
1'
b10 +
#849380000000
0!
0'
#849390000000
1!
b11 %
1'
b11 +
#849400000000
0!
0'
#849410000000
1!
b100 %
1'
b100 +
#849420000000
0!
0'
#849430000000
1!
b101 %
1'
b101 +
#849440000000
0!
0'
#849450000000
1!
0$
b110 %
1'
0*
b110 +
#849460000000
1"
1(
#849470000000
0!
0"
b100 &
0'
0(
b100 ,
#849480000000
1!
1$
b111 %
1'
1*
b111 +
#849490000000
0!
0'
#849500000000
1!
0$
b1000 %
1'
0*
b1000 +
#849510000000
0!
0'
#849520000000
1!
b1001 %
1'
b1001 +
#849530000000
0!
0'
#849540000000
1!
b0 %
1'
b0 +
#849550000000
0!
0'
#849560000000
1!
1$
b1 %
1'
1*
b1 +
#849570000000
0!
0'
#849580000000
1!
b10 %
1'
b10 +
#849590000000
0!
0'
#849600000000
1!
b11 %
1'
b11 +
#849610000000
0!
0'
#849620000000
1!
b100 %
1'
b100 +
#849630000000
0!
0'
#849640000000
1!
b101 %
1'
b101 +
#849650000000
0!
0'
#849660000000
1!
b110 %
1'
b110 +
#849670000000
0!
0'
#849680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#849690000000
0!
0'
#849700000000
1!
b1000 %
1'
b1000 +
#849710000000
0!
0'
#849720000000
1!
b1001 %
1'
b1001 +
#849730000000
0!
0'
#849740000000
1!
b0 %
1'
b0 +
#849750000000
0!
0'
#849760000000
1!
1$
b1 %
1'
1*
b1 +
#849770000000
0!
0'
#849780000000
1!
b10 %
1'
b10 +
#849790000000
0!
0'
#849800000000
1!
b11 %
1'
b11 +
#849810000000
0!
0'
#849820000000
1!
b100 %
1'
b100 +
#849830000000
0!
0'
#849840000000
1!
b101 %
1'
b101 +
#849850000000
0!
0'
#849860000000
1!
0$
b110 %
1'
0*
b110 +
#849870000000
0!
0'
#849880000000
1!
b111 %
1'
b111 +
#849890000000
1"
1(
#849900000000
0!
0"
b100 &
0'
0(
b100 ,
#849910000000
1!
b1000 %
1'
b1000 +
#849920000000
0!
0'
#849930000000
1!
b1001 %
1'
b1001 +
#849940000000
0!
0'
#849950000000
1!
b0 %
1'
b0 +
#849960000000
0!
0'
#849970000000
1!
1$
b1 %
1'
1*
b1 +
#849980000000
0!
0'
#849990000000
1!
b10 %
1'
b10 +
#850000000000
0!
0'
#850010000000
1!
b11 %
1'
b11 +
#850020000000
0!
0'
#850030000000
1!
b100 %
1'
b100 +
#850040000000
0!
0'
#850050000000
1!
b101 %
1'
b101 +
#850060000000
0!
0'
#850070000000
1!
b110 %
1'
b110 +
#850080000000
0!
0'
#850090000000
1!
b111 %
1'
b111 +
#850100000000
0!
0'
#850110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#850120000000
0!
0'
#850130000000
1!
b1001 %
1'
b1001 +
#850140000000
0!
0'
#850150000000
1!
b0 %
1'
b0 +
#850160000000
0!
0'
#850170000000
1!
1$
b1 %
1'
1*
b1 +
#850180000000
0!
0'
#850190000000
1!
b10 %
1'
b10 +
#850200000000
0!
0'
#850210000000
1!
b11 %
1'
b11 +
#850220000000
0!
0'
#850230000000
1!
b100 %
1'
b100 +
#850240000000
0!
0'
#850250000000
1!
b101 %
1'
b101 +
#850260000000
0!
0'
#850270000000
1!
0$
b110 %
1'
0*
b110 +
#850280000000
0!
0'
#850290000000
1!
b111 %
1'
b111 +
#850300000000
0!
0'
#850310000000
1!
b1000 %
1'
b1000 +
#850320000000
1"
1(
#850330000000
0!
0"
b100 &
0'
0(
b100 ,
#850340000000
1!
b1001 %
1'
b1001 +
#850350000000
0!
0'
#850360000000
1!
b0 %
1'
b0 +
#850370000000
0!
0'
#850380000000
1!
1$
b1 %
1'
1*
b1 +
#850390000000
0!
0'
#850400000000
1!
b10 %
1'
b10 +
#850410000000
0!
0'
#850420000000
1!
b11 %
1'
b11 +
#850430000000
0!
0'
#850440000000
1!
b100 %
1'
b100 +
#850450000000
0!
0'
#850460000000
1!
b101 %
1'
b101 +
#850470000000
0!
0'
#850480000000
1!
b110 %
1'
b110 +
#850490000000
0!
0'
#850500000000
1!
b111 %
1'
b111 +
#850510000000
0!
0'
#850520000000
1!
0$
b1000 %
1'
0*
b1000 +
#850530000000
0!
0'
#850540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#850550000000
0!
0'
#850560000000
1!
b0 %
1'
b0 +
#850570000000
0!
0'
#850580000000
1!
1$
b1 %
1'
1*
b1 +
#850590000000
0!
0'
#850600000000
1!
b10 %
1'
b10 +
#850610000000
0!
0'
#850620000000
1!
b11 %
1'
b11 +
#850630000000
0!
0'
#850640000000
1!
b100 %
1'
b100 +
#850650000000
0!
0'
#850660000000
1!
b101 %
1'
b101 +
#850670000000
0!
0'
#850680000000
1!
0$
b110 %
1'
0*
b110 +
#850690000000
0!
0'
#850700000000
1!
b111 %
1'
b111 +
#850710000000
0!
0'
#850720000000
1!
b1000 %
1'
b1000 +
#850730000000
0!
0'
#850740000000
1!
b1001 %
1'
b1001 +
#850750000000
1"
1(
#850760000000
0!
0"
b100 &
0'
0(
b100 ,
#850770000000
1!
b0 %
1'
b0 +
#850780000000
0!
0'
#850790000000
1!
1$
b1 %
1'
1*
b1 +
#850800000000
0!
0'
#850810000000
1!
b10 %
1'
b10 +
#850820000000
0!
0'
#850830000000
1!
b11 %
1'
b11 +
#850840000000
0!
0'
#850850000000
1!
b100 %
1'
b100 +
#850860000000
0!
0'
#850870000000
1!
b101 %
1'
b101 +
#850880000000
0!
0'
#850890000000
1!
b110 %
1'
b110 +
#850900000000
0!
0'
#850910000000
1!
b111 %
1'
b111 +
#850920000000
0!
0'
#850930000000
1!
0$
b1000 %
1'
0*
b1000 +
#850940000000
0!
0'
#850950000000
1!
b1001 %
1'
b1001 +
#850960000000
0!
0'
#850970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#850980000000
0!
0'
#850990000000
1!
1$
b1 %
1'
1*
b1 +
#851000000000
0!
0'
#851010000000
1!
b10 %
1'
b10 +
#851020000000
0!
0'
#851030000000
1!
b11 %
1'
b11 +
#851040000000
0!
0'
#851050000000
1!
b100 %
1'
b100 +
#851060000000
0!
0'
#851070000000
1!
b101 %
1'
b101 +
#851080000000
0!
0'
#851090000000
1!
0$
b110 %
1'
0*
b110 +
#851100000000
0!
0'
#851110000000
1!
b111 %
1'
b111 +
#851120000000
0!
0'
#851130000000
1!
b1000 %
1'
b1000 +
#851140000000
0!
0'
#851150000000
1!
b1001 %
1'
b1001 +
#851160000000
0!
0'
#851170000000
1!
b0 %
1'
b0 +
#851180000000
1"
1(
#851190000000
0!
0"
b100 &
0'
0(
b100 ,
#851200000000
1!
1$
b1 %
1'
1*
b1 +
#851210000000
0!
0'
#851220000000
1!
b10 %
1'
b10 +
#851230000000
0!
0'
#851240000000
1!
b11 %
1'
b11 +
#851250000000
0!
0'
#851260000000
1!
b100 %
1'
b100 +
#851270000000
0!
0'
#851280000000
1!
b101 %
1'
b101 +
#851290000000
0!
0'
#851300000000
1!
b110 %
1'
b110 +
#851310000000
0!
0'
#851320000000
1!
b111 %
1'
b111 +
#851330000000
0!
0'
#851340000000
1!
0$
b1000 %
1'
0*
b1000 +
#851350000000
0!
0'
#851360000000
1!
b1001 %
1'
b1001 +
#851370000000
0!
0'
#851380000000
1!
b0 %
1'
b0 +
#851390000000
0!
0'
#851400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#851410000000
0!
0'
#851420000000
1!
b10 %
1'
b10 +
#851430000000
0!
0'
#851440000000
1!
b11 %
1'
b11 +
#851450000000
0!
0'
#851460000000
1!
b100 %
1'
b100 +
#851470000000
0!
0'
#851480000000
1!
b101 %
1'
b101 +
#851490000000
0!
0'
#851500000000
1!
0$
b110 %
1'
0*
b110 +
#851510000000
0!
0'
#851520000000
1!
b111 %
1'
b111 +
#851530000000
0!
0'
#851540000000
1!
b1000 %
1'
b1000 +
#851550000000
0!
0'
#851560000000
1!
b1001 %
1'
b1001 +
#851570000000
0!
0'
#851580000000
1!
b0 %
1'
b0 +
#851590000000
0!
0'
#851600000000
1!
1$
b1 %
1'
1*
b1 +
#851610000000
1"
1(
#851620000000
0!
0"
b100 &
0'
0(
b100 ,
#851630000000
1!
b10 %
1'
b10 +
#851640000000
0!
0'
#851650000000
1!
b11 %
1'
b11 +
#851660000000
0!
0'
#851670000000
1!
b100 %
1'
b100 +
#851680000000
0!
0'
#851690000000
1!
b101 %
1'
b101 +
#851700000000
0!
0'
#851710000000
1!
b110 %
1'
b110 +
#851720000000
0!
0'
#851730000000
1!
b111 %
1'
b111 +
#851740000000
0!
0'
#851750000000
1!
0$
b1000 %
1'
0*
b1000 +
#851760000000
0!
0'
#851770000000
1!
b1001 %
1'
b1001 +
#851780000000
0!
0'
#851790000000
1!
b0 %
1'
b0 +
#851800000000
0!
0'
#851810000000
1!
1$
b1 %
1'
1*
b1 +
#851820000000
0!
0'
#851830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#851840000000
0!
0'
#851850000000
1!
b11 %
1'
b11 +
#851860000000
0!
0'
#851870000000
1!
b100 %
1'
b100 +
#851880000000
0!
0'
#851890000000
1!
b101 %
1'
b101 +
#851900000000
0!
0'
#851910000000
1!
0$
b110 %
1'
0*
b110 +
#851920000000
0!
0'
#851930000000
1!
b111 %
1'
b111 +
#851940000000
0!
0'
#851950000000
1!
b1000 %
1'
b1000 +
#851960000000
0!
0'
#851970000000
1!
b1001 %
1'
b1001 +
#851980000000
0!
0'
#851990000000
1!
b0 %
1'
b0 +
#852000000000
0!
0'
#852010000000
1!
1$
b1 %
1'
1*
b1 +
#852020000000
0!
0'
#852030000000
1!
b10 %
1'
b10 +
#852040000000
1"
1(
#852050000000
0!
0"
b100 &
0'
0(
b100 ,
#852060000000
1!
b11 %
1'
b11 +
#852070000000
0!
0'
#852080000000
1!
b100 %
1'
b100 +
#852090000000
0!
0'
#852100000000
1!
b101 %
1'
b101 +
#852110000000
0!
0'
#852120000000
1!
b110 %
1'
b110 +
#852130000000
0!
0'
#852140000000
1!
b111 %
1'
b111 +
#852150000000
0!
0'
#852160000000
1!
0$
b1000 %
1'
0*
b1000 +
#852170000000
0!
0'
#852180000000
1!
b1001 %
1'
b1001 +
#852190000000
0!
0'
#852200000000
1!
b0 %
1'
b0 +
#852210000000
0!
0'
#852220000000
1!
1$
b1 %
1'
1*
b1 +
#852230000000
0!
0'
#852240000000
1!
b10 %
1'
b10 +
#852250000000
0!
0'
#852260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#852270000000
0!
0'
#852280000000
1!
b100 %
1'
b100 +
#852290000000
0!
0'
#852300000000
1!
b101 %
1'
b101 +
#852310000000
0!
0'
#852320000000
1!
0$
b110 %
1'
0*
b110 +
#852330000000
0!
0'
#852340000000
1!
b111 %
1'
b111 +
#852350000000
0!
0'
#852360000000
1!
b1000 %
1'
b1000 +
#852370000000
0!
0'
#852380000000
1!
b1001 %
1'
b1001 +
#852390000000
0!
0'
#852400000000
1!
b0 %
1'
b0 +
#852410000000
0!
0'
#852420000000
1!
1$
b1 %
1'
1*
b1 +
#852430000000
0!
0'
#852440000000
1!
b10 %
1'
b10 +
#852450000000
0!
0'
#852460000000
1!
b11 %
1'
b11 +
#852470000000
1"
1(
#852480000000
0!
0"
b100 &
0'
0(
b100 ,
#852490000000
1!
b100 %
1'
b100 +
#852500000000
0!
0'
#852510000000
1!
b101 %
1'
b101 +
#852520000000
0!
0'
#852530000000
1!
b110 %
1'
b110 +
#852540000000
0!
0'
#852550000000
1!
b111 %
1'
b111 +
#852560000000
0!
0'
#852570000000
1!
0$
b1000 %
1'
0*
b1000 +
#852580000000
0!
0'
#852590000000
1!
b1001 %
1'
b1001 +
#852600000000
0!
0'
#852610000000
1!
b0 %
1'
b0 +
#852620000000
0!
0'
#852630000000
1!
1$
b1 %
1'
1*
b1 +
#852640000000
0!
0'
#852650000000
1!
b10 %
1'
b10 +
#852660000000
0!
0'
#852670000000
1!
b11 %
1'
b11 +
#852680000000
0!
0'
#852690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#852700000000
0!
0'
#852710000000
1!
b101 %
1'
b101 +
#852720000000
0!
0'
#852730000000
1!
0$
b110 %
1'
0*
b110 +
#852740000000
0!
0'
#852750000000
1!
b111 %
1'
b111 +
#852760000000
0!
0'
#852770000000
1!
b1000 %
1'
b1000 +
#852780000000
0!
0'
#852790000000
1!
b1001 %
1'
b1001 +
#852800000000
0!
0'
#852810000000
1!
b0 %
1'
b0 +
#852820000000
0!
0'
#852830000000
1!
1$
b1 %
1'
1*
b1 +
#852840000000
0!
0'
#852850000000
1!
b10 %
1'
b10 +
#852860000000
0!
0'
#852870000000
1!
b11 %
1'
b11 +
#852880000000
0!
0'
#852890000000
1!
b100 %
1'
b100 +
#852900000000
1"
1(
#852910000000
0!
0"
b100 &
0'
0(
b100 ,
#852920000000
1!
b101 %
1'
b101 +
#852930000000
0!
0'
#852940000000
1!
b110 %
1'
b110 +
#852950000000
0!
0'
#852960000000
1!
b111 %
1'
b111 +
#852970000000
0!
0'
#852980000000
1!
0$
b1000 %
1'
0*
b1000 +
#852990000000
0!
0'
#853000000000
1!
b1001 %
1'
b1001 +
#853010000000
0!
0'
#853020000000
1!
b0 %
1'
b0 +
#853030000000
0!
0'
#853040000000
1!
1$
b1 %
1'
1*
b1 +
#853050000000
0!
0'
#853060000000
1!
b10 %
1'
b10 +
#853070000000
0!
0'
#853080000000
1!
b11 %
1'
b11 +
#853090000000
0!
0'
#853100000000
1!
b100 %
1'
b100 +
#853110000000
0!
0'
#853120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#853130000000
0!
0'
#853140000000
1!
0$
b110 %
1'
0*
b110 +
#853150000000
0!
0'
#853160000000
1!
b111 %
1'
b111 +
#853170000000
0!
0'
#853180000000
1!
b1000 %
1'
b1000 +
#853190000000
0!
0'
#853200000000
1!
b1001 %
1'
b1001 +
#853210000000
0!
0'
#853220000000
1!
b0 %
1'
b0 +
#853230000000
0!
0'
#853240000000
1!
1$
b1 %
1'
1*
b1 +
#853250000000
0!
0'
#853260000000
1!
b10 %
1'
b10 +
#853270000000
0!
0'
#853280000000
1!
b11 %
1'
b11 +
#853290000000
0!
0'
#853300000000
1!
b100 %
1'
b100 +
#853310000000
0!
0'
#853320000000
1!
b101 %
1'
b101 +
#853330000000
1"
1(
#853340000000
0!
0"
b100 &
0'
0(
b100 ,
#853350000000
1!
b110 %
1'
b110 +
#853360000000
0!
0'
#853370000000
1!
b111 %
1'
b111 +
#853380000000
0!
0'
#853390000000
1!
0$
b1000 %
1'
0*
b1000 +
#853400000000
0!
0'
#853410000000
1!
b1001 %
1'
b1001 +
#853420000000
0!
0'
#853430000000
1!
b0 %
1'
b0 +
#853440000000
0!
0'
#853450000000
1!
1$
b1 %
1'
1*
b1 +
#853460000000
0!
0'
#853470000000
1!
b10 %
1'
b10 +
#853480000000
0!
0'
#853490000000
1!
b11 %
1'
b11 +
#853500000000
0!
0'
#853510000000
1!
b100 %
1'
b100 +
#853520000000
0!
0'
#853530000000
1!
b101 %
1'
b101 +
#853540000000
0!
0'
#853550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#853560000000
0!
0'
#853570000000
1!
b111 %
1'
b111 +
#853580000000
0!
0'
#853590000000
1!
b1000 %
1'
b1000 +
#853600000000
0!
0'
#853610000000
1!
b1001 %
1'
b1001 +
#853620000000
0!
0'
#853630000000
1!
b0 %
1'
b0 +
#853640000000
0!
0'
#853650000000
1!
1$
b1 %
1'
1*
b1 +
#853660000000
0!
0'
#853670000000
1!
b10 %
1'
b10 +
#853680000000
0!
0'
#853690000000
1!
b11 %
1'
b11 +
#853700000000
0!
0'
#853710000000
1!
b100 %
1'
b100 +
#853720000000
0!
0'
#853730000000
1!
b101 %
1'
b101 +
#853740000000
0!
0'
#853750000000
1!
0$
b110 %
1'
0*
b110 +
#853760000000
1"
1(
#853770000000
0!
0"
b100 &
0'
0(
b100 ,
#853780000000
1!
1$
b111 %
1'
1*
b111 +
#853790000000
0!
0'
#853800000000
1!
0$
b1000 %
1'
0*
b1000 +
#853810000000
0!
0'
#853820000000
1!
b1001 %
1'
b1001 +
#853830000000
0!
0'
#853840000000
1!
b0 %
1'
b0 +
#853850000000
0!
0'
#853860000000
1!
1$
b1 %
1'
1*
b1 +
#853870000000
0!
0'
#853880000000
1!
b10 %
1'
b10 +
#853890000000
0!
0'
#853900000000
1!
b11 %
1'
b11 +
#853910000000
0!
0'
#853920000000
1!
b100 %
1'
b100 +
#853930000000
0!
0'
#853940000000
1!
b101 %
1'
b101 +
#853950000000
0!
0'
#853960000000
1!
b110 %
1'
b110 +
#853970000000
0!
0'
#853980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#853990000000
0!
0'
#854000000000
1!
b1000 %
1'
b1000 +
#854010000000
0!
0'
#854020000000
1!
b1001 %
1'
b1001 +
#854030000000
0!
0'
#854040000000
1!
b0 %
1'
b0 +
#854050000000
0!
0'
#854060000000
1!
1$
b1 %
1'
1*
b1 +
#854070000000
0!
0'
#854080000000
1!
b10 %
1'
b10 +
#854090000000
0!
0'
#854100000000
1!
b11 %
1'
b11 +
#854110000000
0!
0'
#854120000000
1!
b100 %
1'
b100 +
#854130000000
0!
0'
#854140000000
1!
b101 %
1'
b101 +
#854150000000
0!
0'
#854160000000
1!
0$
b110 %
1'
0*
b110 +
#854170000000
0!
0'
#854180000000
1!
b111 %
1'
b111 +
#854190000000
1"
1(
#854200000000
0!
0"
b100 &
0'
0(
b100 ,
#854210000000
1!
b1000 %
1'
b1000 +
#854220000000
0!
0'
#854230000000
1!
b1001 %
1'
b1001 +
#854240000000
0!
0'
#854250000000
1!
b0 %
1'
b0 +
#854260000000
0!
0'
#854270000000
1!
1$
b1 %
1'
1*
b1 +
#854280000000
0!
0'
#854290000000
1!
b10 %
1'
b10 +
#854300000000
0!
0'
#854310000000
1!
b11 %
1'
b11 +
#854320000000
0!
0'
#854330000000
1!
b100 %
1'
b100 +
#854340000000
0!
0'
#854350000000
1!
b101 %
1'
b101 +
#854360000000
0!
0'
#854370000000
1!
b110 %
1'
b110 +
#854380000000
0!
0'
#854390000000
1!
b111 %
1'
b111 +
#854400000000
0!
0'
#854410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#854420000000
0!
0'
#854430000000
1!
b1001 %
1'
b1001 +
#854440000000
0!
0'
#854450000000
1!
b0 %
1'
b0 +
#854460000000
0!
0'
#854470000000
1!
1$
b1 %
1'
1*
b1 +
#854480000000
0!
0'
#854490000000
1!
b10 %
1'
b10 +
#854500000000
0!
0'
#854510000000
1!
b11 %
1'
b11 +
#854520000000
0!
0'
#854530000000
1!
b100 %
1'
b100 +
#854540000000
0!
0'
#854550000000
1!
b101 %
1'
b101 +
#854560000000
0!
0'
#854570000000
1!
0$
b110 %
1'
0*
b110 +
#854580000000
0!
0'
#854590000000
1!
b111 %
1'
b111 +
#854600000000
0!
0'
#854610000000
1!
b1000 %
1'
b1000 +
#854620000000
1"
1(
#854630000000
0!
0"
b100 &
0'
0(
b100 ,
#854640000000
1!
b1001 %
1'
b1001 +
#854650000000
0!
0'
#854660000000
1!
b0 %
1'
b0 +
#854670000000
0!
0'
#854680000000
1!
1$
b1 %
1'
1*
b1 +
#854690000000
0!
0'
#854700000000
1!
b10 %
1'
b10 +
#854710000000
0!
0'
#854720000000
1!
b11 %
1'
b11 +
#854730000000
0!
0'
#854740000000
1!
b100 %
1'
b100 +
#854750000000
0!
0'
#854760000000
1!
b101 %
1'
b101 +
#854770000000
0!
0'
#854780000000
1!
b110 %
1'
b110 +
#854790000000
0!
0'
#854800000000
1!
b111 %
1'
b111 +
#854810000000
0!
0'
#854820000000
1!
0$
b1000 %
1'
0*
b1000 +
#854830000000
0!
0'
#854840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#854850000000
0!
0'
#854860000000
1!
b0 %
1'
b0 +
#854870000000
0!
0'
#854880000000
1!
1$
b1 %
1'
1*
b1 +
#854890000000
0!
0'
#854900000000
1!
b10 %
1'
b10 +
#854910000000
0!
0'
#854920000000
1!
b11 %
1'
b11 +
#854930000000
0!
0'
#854940000000
1!
b100 %
1'
b100 +
#854950000000
0!
0'
#854960000000
1!
b101 %
1'
b101 +
#854970000000
0!
0'
#854980000000
1!
0$
b110 %
1'
0*
b110 +
#854990000000
0!
0'
#855000000000
1!
b111 %
1'
b111 +
#855010000000
0!
0'
#855020000000
1!
b1000 %
1'
b1000 +
#855030000000
0!
0'
#855040000000
1!
b1001 %
1'
b1001 +
#855050000000
1"
1(
#855060000000
0!
0"
b100 &
0'
0(
b100 ,
#855070000000
1!
b0 %
1'
b0 +
#855080000000
0!
0'
#855090000000
1!
1$
b1 %
1'
1*
b1 +
#855100000000
0!
0'
#855110000000
1!
b10 %
1'
b10 +
#855120000000
0!
0'
#855130000000
1!
b11 %
1'
b11 +
#855140000000
0!
0'
#855150000000
1!
b100 %
1'
b100 +
#855160000000
0!
0'
#855170000000
1!
b101 %
1'
b101 +
#855180000000
0!
0'
#855190000000
1!
b110 %
1'
b110 +
#855200000000
0!
0'
#855210000000
1!
b111 %
1'
b111 +
#855220000000
0!
0'
#855230000000
1!
0$
b1000 %
1'
0*
b1000 +
#855240000000
0!
0'
#855250000000
1!
b1001 %
1'
b1001 +
#855260000000
0!
0'
#855270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#855280000000
0!
0'
#855290000000
1!
1$
b1 %
1'
1*
b1 +
#855300000000
0!
0'
#855310000000
1!
b10 %
1'
b10 +
#855320000000
0!
0'
#855330000000
1!
b11 %
1'
b11 +
#855340000000
0!
0'
#855350000000
1!
b100 %
1'
b100 +
#855360000000
0!
0'
#855370000000
1!
b101 %
1'
b101 +
#855380000000
0!
0'
#855390000000
1!
0$
b110 %
1'
0*
b110 +
#855400000000
0!
0'
#855410000000
1!
b111 %
1'
b111 +
#855420000000
0!
0'
#855430000000
1!
b1000 %
1'
b1000 +
#855440000000
0!
0'
#855450000000
1!
b1001 %
1'
b1001 +
#855460000000
0!
0'
#855470000000
1!
b0 %
1'
b0 +
#855480000000
1"
1(
#855490000000
0!
0"
b100 &
0'
0(
b100 ,
#855500000000
1!
1$
b1 %
1'
1*
b1 +
#855510000000
0!
0'
#855520000000
1!
b10 %
1'
b10 +
#855530000000
0!
0'
#855540000000
1!
b11 %
1'
b11 +
#855550000000
0!
0'
#855560000000
1!
b100 %
1'
b100 +
#855570000000
0!
0'
#855580000000
1!
b101 %
1'
b101 +
#855590000000
0!
0'
#855600000000
1!
b110 %
1'
b110 +
#855610000000
0!
0'
#855620000000
1!
b111 %
1'
b111 +
#855630000000
0!
0'
#855640000000
1!
0$
b1000 %
1'
0*
b1000 +
#855650000000
0!
0'
#855660000000
1!
b1001 %
1'
b1001 +
#855670000000
0!
0'
#855680000000
1!
b0 %
1'
b0 +
#855690000000
0!
0'
#855700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#855710000000
0!
0'
#855720000000
1!
b10 %
1'
b10 +
#855730000000
0!
0'
#855740000000
1!
b11 %
1'
b11 +
#855750000000
0!
0'
#855760000000
1!
b100 %
1'
b100 +
#855770000000
0!
0'
#855780000000
1!
b101 %
1'
b101 +
#855790000000
0!
0'
#855800000000
1!
0$
b110 %
1'
0*
b110 +
#855810000000
0!
0'
#855820000000
1!
b111 %
1'
b111 +
#855830000000
0!
0'
#855840000000
1!
b1000 %
1'
b1000 +
#855850000000
0!
0'
#855860000000
1!
b1001 %
1'
b1001 +
#855870000000
0!
0'
#855880000000
1!
b0 %
1'
b0 +
#855890000000
0!
0'
#855900000000
1!
1$
b1 %
1'
1*
b1 +
#855910000000
1"
1(
#855920000000
0!
0"
b100 &
0'
0(
b100 ,
#855930000000
1!
b10 %
1'
b10 +
#855940000000
0!
0'
#855950000000
1!
b11 %
1'
b11 +
#855960000000
0!
0'
#855970000000
1!
b100 %
1'
b100 +
#855980000000
0!
0'
#855990000000
1!
b101 %
1'
b101 +
#856000000000
0!
0'
#856010000000
1!
b110 %
1'
b110 +
#856020000000
0!
0'
#856030000000
1!
b111 %
1'
b111 +
#856040000000
0!
0'
#856050000000
1!
0$
b1000 %
1'
0*
b1000 +
#856060000000
0!
0'
#856070000000
1!
b1001 %
1'
b1001 +
#856080000000
0!
0'
#856090000000
1!
b0 %
1'
b0 +
#856100000000
0!
0'
#856110000000
1!
1$
b1 %
1'
1*
b1 +
#856120000000
0!
0'
#856130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#856140000000
0!
0'
#856150000000
1!
b11 %
1'
b11 +
#856160000000
0!
0'
#856170000000
1!
b100 %
1'
b100 +
#856180000000
0!
0'
#856190000000
1!
b101 %
1'
b101 +
#856200000000
0!
0'
#856210000000
1!
0$
b110 %
1'
0*
b110 +
#856220000000
0!
0'
#856230000000
1!
b111 %
1'
b111 +
#856240000000
0!
0'
#856250000000
1!
b1000 %
1'
b1000 +
#856260000000
0!
0'
#856270000000
1!
b1001 %
1'
b1001 +
#856280000000
0!
0'
#856290000000
1!
b0 %
1'
b0 +
#856300000000
0!
0'
#856310000000
1!
1$
b1 %
1'
1*
b1 +
#856320000000
0!
0'
#856330000000
1!
b10 %
1'
b10 +
#856340000000
1"
1(
#856350000000
0!
0"
b100 &
0'
0(
b100 ,
#856360000000
1!
b11 %
1'
b11 +
#856370000000
0!
0'
#856380000000
1!
b100 %
1'
b100 +
#856390000000
0!
0'
#856400000000
1!
b101 %
1'
b101 +
#856410000000
0!
0'
#856420000000
1!
b110 %
1'
b110 +
#856430000000
0!
0'
#856440000000
1!
b111 %
1'
b111 +
#856450000000
0!
0'
#856460000000
1!
0$
b1000 %
1'
0*
b1000 +
#856470000000
0!
0'
#856480000000
1!
b1001 %
1'
b1001 +
#856490000000
0!
0'
#856500000000
1!
b0 %
1'
b0 +
#856510000000
0!
0'
#856520000000
1!
1$
b1 %
1'
1*
b1 +
#856530000000
0!
0'
#856540000000
1!
b10 %
1'
b10 +
#856550000000
0!
0'
#856560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#856570000000
0!
0'
#856580000000
1!
b100 %
1'
b100 +
#856590000000
0!
0'
#856600000000
1!
b101 %
1'
b101 +
#856610000000
0!
0'
#856620000000
1!
0$
b110 %
1'
0*
b110 +
#856630000000
0!
0'
#856640000000
1!
b111 %
1'
b111 +
#856650000000
0!
0'
#856660000000
1!
b1000 %
1'
b1000 +
#856670000000
0!
0'
#856680000000
1!
b1001 %
1'
b1001 +
#856690000000
0!
0'
#856700000000
1!
b0 %
1'
b0 +
#856710000000
0!
0'
#856720000000
1!
1$
b1 %
1'
1*
b1 +
#856730000000
0!
0'
#856740000000
1!
b10 %
1'
b10 +
#856750000000
0!
0'
#856760000000
1!
b11 %
1'
b11 +
#856770000000
1"
1(
#856780000000
0!
0"
b100 &
0'
0(
b100 ,
#856790000000
1!
b100 %
1'
b100 +
#856800000000
0!
0'
#856810000000
1!
b101 %
1'
b101 +
#856820000000
0!
0'
#856830000000
1!
b110 %
1'
b110 +
#856840000000
0!
0'
#856850000000
1!
b111 %
1'
b111 +
#856860000000
0!
0'
#856870000000
1!
0$
b1000 %
1'
0*
b1000 +
#856880000000
0!
0'
#856890000000
1!
b1001 %
1'
b1001 +
#856900000000
0!
0'
#856910000000
1!
b0 %
1'
b0 +
#856920000000
0!
0'
#856930000000
1!
1$
b1 %
1'
1*
b1 +
#856940000000
0!
0'
#856950000000
1!
b10 %
1'
b10 +
#856960000000
0!
0'
#856970000000
1!
b11 %
1'
b11 +
#856980000000
0!
0'
#856990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#857000000000
0!
0'
#857010000000
1!
b101 %
1'
b101 +
#857020000000
0!
0'
#857030000000
1!
0$
b110 %
1'
0*
b110 +
#857040000000
0!
0'
#857050000000
1!
b111 %
1'
b111 +
#857060000000
0!
0'
#857070000000
1!
b1000 %
1'
b1000 +
#857080000000
0!
0'
#857090000000
1!
b1001 %
1'
b1001 +
#857100000000
0!
0'
#857110000000
1!
b0 %
1'
b0 +
#857120000000
0!
0'
#857130000000
1!
1$
b1 %
1'
1*
b1 +
#857140000000
0!
0'
#857150000000
1!
b10 %
1'
b10 +
#857160000000
0!
0'
#857170000000
1!
b11 %
1'
b11 +
#857180000000
0!
0'
#857190000000
1!
b100 %
1'
b100 +
#857200000000
1"
1(
#857210000000
0!
0"
b100 &
0'
0(
b100 ,
#857220000000
1!
b101 %
1'
b101 +
#857230000000
0!
0'
#857240000000
1!
b110 %
1'
b110 +
#857250000000
0!
0'
#857260000000
1!
b111 %
1'
b111 +
#857270000000
0!
0'
#857280000000
1!
0$
b1000 %
1'
0*
b1000 +
#857290000000
0!
0'
#857300000000
1!
b1001 %
1'
b1001 +
#857310000000
0!
0'
#857320000000
1!
b0 %
1'
b0 +
#857330000000
0!
0'
#857340000000
1!
1$
b1 %
1'
1*
b1 +
#857350000000
0!
0'
#857360000000
1!
b10 %
1'
b10 +
#857370000000
0!
0'
#857380000000
1!
b11 %
1'
b11 +
#857390000000
0!
0'
#857400000000
1!
b100 %
1'
b100 +
#857410000000
0!
0'
#857420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#857430000000
0!
0'
#857440000000
1!
0$
b110 %
1'
0*
b110 +
#857450000000
0!
0'
#857460000000
1!
b111 %
1'
b111 +
#857470000000
0!
0'
#857480000000
1!
b1000 %
1'
b1000 +
#857490000000
0!
0'
#857500000000
1!
b1001 %
1'
b1001 +
#857510000000
0!
0'
#857520000000
1!
b0 %
1'
b0 +
#857530000000
0!
0'
#857540000000
1!
1$
b1 %
1'
1*
b1 +
#857550000000
0!
0'
#857560000000
1!
b10 %
1'
b10 +
#857570000000
0!
0'
#857580000000
1!
b11 %
1'
b11 +
#857590000000
0!
0'
#857600000000
1!
b100 %
1'
b100 +
#857610000000
0!
0'
#857620000000
1!
b101 %
1'
b101 +
#857630000000
1"
1(
#857640000000
0!
0"
b100 &
0'
0(
b100 ,
#857650000000
1!
b110 %
1'
b110 +
#857660000000
0!
0'
#857670000000
1!
b111 %
1'
b111 +
#857680000000
0!
0'
#857690000000
1!
0$
b1000 %
1'
0*
b1000 +
#857700000000
0!
0'
#857710000000
1!
b1001 %
1'
b1001 +
#857720000000
0!
0'
#857730000000
1!
b0 %
1'
b0 +
#857740000000
0!
0'
#857750000000
1!
1$
b1 %
1'
1*
b1 +
#857760000000
0!
0'
#857770000000
1!
b10 %
1'
b10 +
#857780000000
0!
0'
#857790000000
1!
b11 %
1'
b11 +
#857800000000
0!
0'
#857810000000
1!
b100 %
1'
b100 +
#857820000000
0!
0'
#857830000000
1!
b101 %
1'
b101 +
#857840000000
0!
0'
#857850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#857860000000
0!
0'
#857870000000
1!
b111 %
1'
b111 +
#857880000000
0!
0'
#857890000000
1!
b1000 %
1'
b1000 +
#857900000000
0!
0'
#857910000000
1!
b1001 %
1'
b1001 +
#857920000000
0!
0'
#857930000000
1!
b0 %
1'
b0 +
#857940000000
0!
0'
#857950000000
1!
1$
b1 %
1'
1*
b1 +
#857960000000
0!
0'
#857970000000
1!
b10 %
1'
b10 +
#857980000000
0!
0'
#857990000000
1!
b11 %
1'
b11 +
#858000000000
0!
0'
#858010000000
1!
b100 %
1'
b100 +
#858020000000
0!
0'
#858030000000
1!
b101 %
1'
b101 +
#858040000000
0!
0'
#858050000000
1!
0$
b110 %
1'
0*
b110 +
#858060000000
1"
1(
#858070000000
0!
0"
b100 &
0'
0(
b100 ,
#858080000000
1!
1$
b111 %
1'
1*
b111 +
#858090000000
0!
0'
#858100000000
1!
0$
b1000 %
1'
0*
b1000 +
#858110000000
0!
0'
#858120000000
1!
b1001 %
1'
b1001 +
#858130000000
0!
0'
#858140000000
1!
b0 %
1'
b0 +
#858150000000
0!
0'
#858160000000
1!
1$
b1 %
1'
1*
b1 +
#858170000000
0!
0'
#858180000000
1!
b10 %
1'
b10 +
#858190000000
0!
0'
#858200000000
1!
b11 %
1'
b11 +
#858210000000
0!
0'
#858220000000
1!
b100 %
1'
b100 +
#858230000000
0!
0'
#858240000000
1!
b101 %
1'
b101 +
#858250000000
0!
0'
#858260000000
1!
b110 %
1'
b110 +
#858270000000
0!
0'
#858280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#858290000000
0!
0'
#858300000000
1!
b1000 %
1'
b1000 +
#858310000000
0!
0'
#858320000000
1!
b1001 %
1'
b1001 +
#858330000000
0!
0'
#858340000000
1!
b0 %
1'
b0 +
#858350000000
0!
0'
#858360000000
1!
1$
b1 %
1'
1*
b1 +
#858370000000
0!
0'
#858380000000
1!
b10 %
1'
b10 +
#858390000000
0!
0'
#858400000000
1!
b11 %
1'
b11 +
#858410000000
0!
0'
#858420000000
1!
b100 %
1'
b100 +
#858430000000
0!
0'
#858440000000
1!
b101 %
1'
b101 +
#858450000000
0!
0'
#858460000000
1!
0$
b110 %
1'
0*
b110 +
#858470000000
0!
0'
#858480000000
1!
b111 %
1'
b111 +
#858490000000
1"
1(
#858500000000
0!
0"
b100 &
0'
0(
b100 ,
#858510000000
1!
b1000 %
1'
b1000 +
#858520000000
0!
0'
#858530000000
1!
b1001 %
1'
b1001 +
#858540000000
0!
0'
#858550000000
1!
b0 %
1'
b0 +
#858560000000
0!
0'
#858570000000
1!
1$
b1 %
1'
1*
b1 +
#858580000000
0!
0'
#858590000000
1!
b10 %
1'
b10 +
#858600000000
0!
0'
#858610000000
1!
b11 %
1'
b11 +
#858620000000
0!
0'
#858630000000
1!
b100 %
1'
b100 +
#858640000000
0!
0'
#858650000000
1!
b101 %
1'
b101 +
#858660000000
0!
0'
#858670000000
1!
b110 %
1'
b110 +
#858680000000
0!
0'
#858690000000
1!
b111 %
1'
b111 +
#858700000000
0!
0'
#858710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#858720000000
0!
0'
#858730000000
1!
b1001 %
1'
b1001 +
#858740000000
0!
0'
#858750000000
1!
b0 %
1'
b0 +
#858760000000
0!
0'
#858770000000
1!
1$
b1 %
1'
1*
b1 +
#858780000000
0!
0'
#858790000000
1!
b10 %
1'
b10 +
#858800000000
0!
0'
#858810000000
1!
b11 %
1'
b11 +
#858820000000
0!
0'
#858830000000
1!
b100 %
1'
b100 +
#858840000000
0!
0'
#858850000000
1!
b101 %
1'
b101 +
#858860000000
0!
0'
#858870000000
1!
0$
b110 %
1'
0*
b110 +
#858880000000
0!
0'
#858890000000
1!
b111 %
1'
b111 +
#858900000000
0!
0'
#858910000000
1!
b1000 %
1'
b1000 +
#858920000000
1"
1(
#858930000000
0!
0"
b100 &
0'
0(
b100 ,
#858940000000
1!
b1001 %
1'
b1001 +
#858950000000
0!
0'
#858960000000
1!
b0 %
1'
b0 +
#858970000000
0!
0'
#858980000000
1!
1$
b1 %
1'
1*
b1 +
#858990000000
0!
0'
#859000000000
1!
b10 %
1'
b10 +
#859010000000
0!
0'
#859020000000
1!
b11 %
1'
b11 +
#859030000000
0!
0'
#859040000000
1!
b100 %
1'
b100 +
#859050000000
0!
0'
#859060000000
1!
b101 %
1'
b101 +
#859070000000
0!
0'
#859080000000
1!
b110 %
1'
b110 +
#859090000000
0!
0'
#859100000000
1!
b111 %
1'
b111 +
#859110000000
0!
0'
#859120000000
1!
0$
b1000 %
1'
0*
b1000 +
#859130000000
0!
0'
#859140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#859150000000
0!
0'
#859160000000
1!
b0 %
1'
b0 +
#859170000000
0!
0'
#859180000000
1!
1$
b1 %
1'
1*
b1 +
#859190000000
0!
0'
#859200000000
1!
b10 %
1'
b10 +
#859210000000
0!
0'
#859220000000
1!
b11 %
1'
b11 +
#859230000000
0!
0'
#859240000000
1!
b100 %
1'
b100 +
#859250000000
0!
0'
#859260000000
1!
b101 %
1'
b101 +
#859270000000
0!
0'
#859280000000
1!
0$
b110 %
1'
0*
b110 +
#859290000000
0!
0'
#859300000000
1!
b111 %
1'
b111 +
#859310000000
0!
0'
#859320000000
1!
b1000 %
1'
b1000 +
#859330000000
0!
0'
#859340000000
1!
b1001 %
1'
b1001 +
#859350000000
1"
1(
#859360000000
0!
0"
b100 &
0'
0(
b100 ,
#859370000000
1!
b0 %
1'
b0 +
#859380000000
0!
0'
#859390000000
1!
1$
b1 %
1'
1*
b1 +
#859400000000
0!
0'
#859410000000
1!
b10 %
1'
b10 +
#859420000000
0!
0'
#859430000000
1!
b11 %
1'
b11 +
#859440000000
0!
0'
#859450000000
1!
b100 %
1'
b100 +
#859460000000
0!
0'
#859470000000
1!
b101 %
1'
b101 +
#859480000000
0!
0'
#859490000000
1!
b110 %
1'
b110 +
#859500000000
0!
0'
#859510000000
1!
b111 %
1'
b111 +
#859520000000
0!
0'
#859530000000
1!
0$
b1000 %
1'
0*
b1000 +
#859540000000
0!
0'
#859550000000
1!
b1001 %
1'
b1001 +
#859560000000
0!
0'
#859570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#859580000000
0!
0'
#859590000000
1!
1$
b1 %
1'
1*
b1 +
#859600000000
0!
0'
#859610000000
1!
b10 %
1'
b10 +
#859620000000
0!
0'
#859630000000
1!
b11 %
1'
b11 +
#859640000000
0!
0'
#859650000000
1!
b100 %
1'
b100 +
#859660000000
0!
0'
#859670000000
1!
b101 %
1'
b101 +
#859680000000
0!
0'
#859690000000
1!
0$
b110 %
1'
0*
b110 +
#859700000000
0!
0'
#859710000000
1!
b111 %
1'
b111 +
#859720000000
0!
0'
#859730000000
1!
b1000 %
1'
b1000 +
#859740000000
0!
0'
#859750000000
1!
b1001 %
1'
b1001 +
#859760000000
0!
0'
#859770000000
1!
b0 %
1'
b0 +
#859780000000
1"
1(
#859790000000
0!
0"
b100 &
0'
0(
b100 ,
#859800000000
1!
1$
b1 %
1'
1*
b1 +
#859810000000
0!
0'
#859820000000
1!
b10 %
1'
b10 +
#859830000000
0!
0'
#859840000000
1!
b11 %
1'
b11 +
#859850000000
0!
0'
#859860000000
1!
b100 %
1'
b100 +
#859870000000
0!
0'
#859880000000
1!
b101 %
1'
b101 +
#859890000000
0!
0'
#859900000000
1!
b110 %
1'
b110 +
#859910000000
0!
0'
#859920000000
1!
b111 %
1'
b111 +
#859930000000
0!
0'
#859940000000
1!
0$
b1000 %
1'
0*
b1000 +
#859950000000
0!
0'
#859960000000
1!
b1001 %
1'
b1001 +
#859970000000
0!
0'
#859980000000
1!
b0 %
1'
b0 +
#859990000000
0!
0'
#860000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#860010000000
0!
0'
#860020000000
1!
b10 %
1'
b10 +
#860030000000
0!
0'
#860040000000
1!
b11 %
1'
b11 +
#860050000000
0!
0'
#860060000000
1!
b100 %
1'
b100 +
#860070000000
0!
0'
#860080000000
1!
b101 %
1'
b101 +
#860090000000
0!
0'
#860100000000
1!
0$
b110 %
1'
0*
b110 +
#860110000000
0!
0'
#860120000000
1!
b111 %
1'
b111 +
#860130000000
0!
0'
#860140000000
1!
b1000 %
1'
b1000 +
#860150000000
0!
0'
#860160000000
1!
b1001 %
1'
b1001 +
#860170000000
0!
0'
#860180000000
1!
b0 %
1'
b0 +
#860190000000
0!
0'
#860200000000
1!
1$
b1 %
1'
1*
b1 +
#860210000000
1"
1(
#860220000000
0!
0"
b100 &
0'
0(
b100 ,
#860230000000
1!
b10 %
1'
b10 +
#860240000000
0!
0'
#860250000000
1!
b11 %
1'
b11 +
#860260000000
0!
0'
#860270000000
1!
b100 %
1'
b100 +
#860280000000
0!
0'
#860290000000
1!
b101 %
1'
b101 +
#860300000000
0!
0'
#860310000000
1!
b110 %
1'
b110 +
#860320000000
0!
0'
#860330000000
1!
b111 %
1'
b111 +
#860340000000
0!
0'
#860350000000
1!
0$
b1000 %
1'
0*
b1000 +
#860360000000
0!
0'
#860370000000
1!
b1001 %
1'
b1001 +
#860380000000
0!
0'
#860390000000
1!
b0 %
1'
b0 +
#860400000000
0!
0'
#860410000000
1!
1$
b1 %
1'
1*
b1 +
#860420000000
0!
0'
#860430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#860440000000
0!
0'
#860450000000
1!
b11 %
1'
b11 +
#860460000000
0!
0'
#860470000000
1!
b100 %
1'
b100 +
#860480000000
0!
0'
#860490000000
1!
b101 %
1'
b101 +
#860500000000
0!
0'
#860510000000
1!
0$
b110 %
1'
0*
b110 +
#860520000000
0!
0'
#860530000000
1!
b111 %
1'
b111 +
#860540000000
0!
0'
#860550000000
1!
b1000 %
1'
b1000 +
#860560000000
0!
0'
#860570000000
1!
b1001 %
1'
b1001 +
#860580000000
0!
0'
#860590000000
1!
b0 %
1'
b0 +
#860600000000
0!
0'
#860610000000
1!
1$
b1 %
1'
1*
b1 +
#860620000000
0!
0'
#860630000000
1!
b10 %
1'
b10 +
#860640000000
1"
1(
#860650000000
0!
0"
b100 &
0'
0(
b100 ,
#860660000000
1!
b11 %
1'
b11 +
#860670000000
0!
0'
#860680000000
1!
b100 %
1'
b100 +
#860690000000
0!
0'
#860700000000
1!
b101 %
1'
b101 +
#860710000000
0!
0'
#860720000000
1!
b110 %
1'
b110 +
#860730000000
0!
0'
#860740000000
1!
b111 %
1'
b111 +
#860750000000
0!
0'
#860760000000
1!
0$
b1000 %
1'
0*
b1000 +
#860770000000
0!
0'
#860780000000
1!
b1001 %
1'
b1001 +
#860790000000
0!
0'
#860800000000
1!
b0 %
1'
b0 +
#860810000000
0!
0'
#860820000000
1!
1$
b1 %
1'
1*
b1 +
#860830000000
0!
0'
#860840000000
1!
b10 %
1'
b10 +
#860850000000
0!
0'
#860860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#860870000000
0!
0'
#860880000000
1!
b100 %
1'
b100 +
#860890000000
0!
0'
#860900000000
1!
b101 %
1'
b101 +
#860910000000
0!
0'
#860920000000
1!
0$
b110 %
1'
0*
b110 +
#860930000000
0!
0'
#860940000000
1!
b111 %
1'
b111 +
#860950000000
0!
0'
#860960000000
1!
b1000 %
1'
b1000 +
#860970000000
0!
0'
#860980000000
1!
b1001 %
1'
b1001 +
#860990000000
0!
0'
#861000000000
1!
b0 %
1'
b0 +
#861010000000
0!
0'
#861020000000
1!
1$
b1 %
1'
1*
b1 +
#861030000000
0!
0'
#861040000000
1!
b10 %
1'
b10 +
#861050000000
0!
0'
#861060000000
1!
b11 %
1'
b11 +
#861070000000
1"
1(
#861080000000
0!
0"
b100 &
0'
0(
b100 ,
#861090000000
1!
b100 %
1'
b100 +
#861100000000
0!
0'
#861110000000
1!
b101 %
1'
b101 +
#861120000000
0!
0'
#861130000000
1!
b110 %
1'
b110 +
#861140000000
0!
0'
#861150000000
1!
b111 %
1'
b111 +
#861160000000
0!
0'
#861170000000
1!
0$
b1000 %
1'
0*
b1000 +
#861180000000
0!
0'
#861190000000
1!
b1001 %
1'
b1001 +
#861200000000
0!
0'
#861210000000
1!
b0 %
1'
b0 +
#861220000000
0!
0'
#861230000000
1!
1$
b1 %
1'
1*
b1 +
#861240000000
0!
0'
#861250000000
1!
b10 %
1'
b10 +
#861260000000
0!
0'
#861270000000
1!
b11 %
1'
b11 +
#861280000000
0!
0'
#861290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#861300000000
0!
0'
#861310000000
1!
b101 %
1'
b101 +
#861320000000
0!
0'
#861330000000
1!
0$
b110 %
1'
0*
b110 +
#861340000000
0!
0'
#861350000000
1!
b111 %
1'
b111 +
#861360000000
0!
0'
#861370000000
1!
b1000 %
1'
b1000 +
#861380000000
0!
0'
#861390000000
1!
b1001 %
1'
b1001 +
#861400000000
0!
0'
#861410000000
1!
b0 %
1'
b0 +
#861420000000
0!
0'
#861430000000
1!
1$
b1 %
1'
1*
b1 +
#861440000000
0!
0'
#861450000000
1!
b10 %
1'
b10 +
#861460000000
0!
0'
#861470000000
1!
b11 %
1'
b11 +
#861480000000
0!
0'
#861490000000
1!
b100 %
1'
b100 +
#861500000000
1"
1(
#861510000000
0!
0"
b100 &
0'
0(
b100 ,
#861520000000
1!
b101 %
1'
b101 +
#861530000000
0!
0'
#861540000000
1!
b110 %
1'
b110 +
#861550000000
0!
0'
#861560000000
1!
b111 %
1'
b111 +
#861570000000
0!
0'
#861580000000
1!
0$
b1000 %
1'
0*
b1000 +
#861590000000
0!
0'
#861600000000
1!
b1001 %
1'
b1001 +
#861610000000
0!
0'
#861620000000
1!
b0 %
1'
b0 +
#861630000000
0!
0'
#861640000000
1!
1$
b1 %
1'
1*
b1 +
#861650000000
0!
0'
#861660000000
1!
b10 %
1'
b10 +
#861670000000
0!
0'
#861680000000
1!
b11 %
1'
b11 +
#861690000000
0!
0'
#861700000000
1!
b100 %
1'
b100 +
#861710000000
0!
0'
#861720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#861730000000
0!
0'
#861740000000
1!
0$
b110 %
1'
0*
b110 +
#861750000000
0!
0'
#861760000000
1!
b111 %
1'
b111 +
#861770000000
0!
0'
#861780000000
1!
b1000 %
1'
b1000 +
#861790000000
0!
0'
#861800000000
1!
b1001 %
1'
b1001 +
#861810000000
0!
0'
#861820000000
1!
b0 %
1'
b0 +
#861830000000
0!
0'
#861840000000
1!
1$
b1 %
1'
1*
b1 +
#861850000000
0!
0'
#861860000000
1!
b10 %
1'
b10 +
#861870000000
0!
0'
#861880000000
1!
b11 %
1'
b11 +
#861890000000
0!
0'
#861900000000
1!
b100 %
1'
b100 +
#861910000000
0!
0'
#861920000000
1!
b101 %
1'
b101 +
#861930000000
1"
1(
#861940000000
0!
0"
b100 &
0'
0(
b100 ,
#861950000000
1!
b110 %
1'
b110 +
#861960000000
0!
0'
#861970000000
1!
b111 %
1'
b111 +
#861980000000
0!
0'
#861990000000
1!
0$
b1000 %
1'
0*
b1000 +
#862000000000
0!
0'
#862010000000
1!
b1001 %
1'
b1001 +
#862020000000
0!
0'
#862030000000
1!
b0 %
1'
b0 +
#862040000000
0!
0'
#862050000000
1!
1$
b1 %
1'
1*
b1 +
#862060000000
0!
0'
#862070000000
1!
b10 %
1'
b10 +
#862080000000
0!
0'
#862090000000
1!
b11 %
1'
b11 +
#862100000000
0!
0'
#862110000000
1!
b100 %
1'
b100 +
#862120000000
0!
0'
#862130000000
1!
b101 %
1'
b101 +
#862140000000
0!
0'
#862150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#862160000000
0!
0'
#862170000000
1!
b111 %
1'
b111 +
#862180000000
0!
0'
#862190000000
1!
b1000 %
1'
b1000 +
#862200000000
0!
0'
#862210000000
1!
b1001 %
1'
b1001 +
#862220000000
0!
0'
#862230000000
1!
b0 %
1'
b0 +
#862240000000
0!
0'
#862250000000
1!
1$
b1 %
1'
1*
b1 +
#862260000000
0!
0'
#862270000000
1!
b10 %
1'
b10 +
#862280000000
0!
0'
#862290000000
1!
b11 %
1'
b11 +
#862300000000
0!
0'
#862310000000
1!
b100 %
1'
b100 +
#862320000000
0!
0'
#862330000000
1!
b101 %
1'
b101 +
#862340000000
0!
0'
#862350000000
1!
0$
b110 %
1'
0*
b110 +
#862360000000
1"
1(
#862370000000
0!
0"
b100 &
0'
0(
b100 ,
#862380000000
1!
1$
b111 %
1'
1*
b111 +
#862390000000
0!
0'
#862400000000
1!
0$
b1000 %
1'
0*
b1000 +
#862410000000
0!
0'
#862420000000
1!
b1001 %
1'
b1001 +
#862430000000
0!
0'
#862440000000
1!
b0 %
1'
b0 +
#862450000000
0!
0'
#862460000000
1!
1$
b1 %
1'
1*
b1 +
#862470000000
0!
0'
#862480000000
1!
b10 %
1'
b10 +
#862490000000
0!
0'
#862500000000
1!
b11 %
1'
b11 +
#862510000000
0!
0'
#862520000000
1!
b100 %
1'
b100 +
#862530000000
0!
0'
#862540000000
1!
b101 %
1'
b101 +
#862550000000
0!
0'
#862560000000
1!
b110 %
1'
b110 +
#862570000000
0!
0'
#862580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#862590000000
0!
0'
#862600000000
1!
b1000 %
1'
b1000 +
#862610000000
0!
0'
#862620000000
1!
b1001 %
1'
b1001 +
#862630000000
0!
0'
#862640000000
1!
b0 %
1'
b0 +
#862650000000
0!
0'
#862660000000
1!
1$
b1 %
1'
1*
b1 +
#862670000000
0!
0'
#862680000000
1!
b10 %
1'
b10 +
#862690000000
0!
0'
#862700000000
1!
b11 %
1'
b11 +
#862710000000
0!
0'
#862720000000
1!
b100 %
1'
b100 +
#862730000000
0!
0'
#862740000000
1!
b101 %
1'
b101 +
#862750000000
0!
0'
#862760000000
1!
0$
b110 %
1'
0*
b110 +
#862770000000
0!
0'
#862780000000
1!
b111 %
1'
b111 +
#862790000000
1"
1(
#862800000000
0!
0"
b100 &
0'
0(
b100 ,
#862810000000
1!
b1000 %
1'
b1000 +
#862820000000
0!
0'
#862830000000
1!
b1001 %
1'
b1001 +
#862840000000
0!
0'
#862850000000
1!
b0 %
1'
b0 +
#862860000000
0!
0'
#862870000000
1!
1$
b1 %
1'
1*
b1 +
#862880000000
0!
0'
#862890000000
1!
b10 %
1'
b10 +
#862900000000
0!
0'
#862910000000
1!
b11 %
1'
b11 +
#862920000000
0!
0'
#862930000000
1!
b100 %
1'
b100 +
#862940000000
0!
0'
#862950000000
1!
b101 %
1'
b101 +
#862960000000
0!
0'
#862970000000
1!
b110 %
1'
b110 +
#862980000000
0!
0'
#862990000000
1!
b111 %
1'
b111 +
#863000000000
0!
0'
#863010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#863020000000
0!
0'
#863030000000
1!
b1001 %
1'
b1001 +
#863040000000
0!
0'
#863050000000
1!
b0 %
1'
b0 +
#863060000000
0!
0'
#863070000000
1!
1$
b1 %
1'
1*
b1 +
#863080000000
0!
0'
#863090000000
1!
b10 %
1'
b10 +
#863100000000
0!
0'
#863110000000
1!
b11 %
1'
b11 +
#863120000000
0!
0'
#863130000000
1!
b100 %
1'
b100 +
#863140000000
0!
0'
#863150000000
1!
b101 %
1'
b101 +
#863160000000
0!
0'
#863170000000
1!
0$
b110 %
1'
0*
b110 +
#863180000000
0!
0'
#863190000000
1!
b111 %
1'
b111 +
#863200000000
0!
0'
#863210000000
1!
b1000 %
1'
b1000 +
#863220000000
1"
1(
#863230000000
0!
0"
b100 &
0'
0(
b100 ,
#863240000000
1!
b1001 %
1'
b1001 +
#863250000000
0!
0'
#863260000000
1!
b0 %
1'
b0 +
#863270000000
0!
0'
#863280000000
1!
1$
b1 %
1'
1*
b1 +
#863290000000
0!
0'
#863300000000
1!
b10 %
1'
b10 +
#863310000000
0!
0'
#863320000000
1!
b11 %
1'
b11 +
#863330000000
0!
0'
#863340000000
1!
b100 %
1'
b100 +
#863350000000
0!
0'
#863360000000
1!
b101 %
1'
b101 +
#863370000000
0!
0'
#863380000000
1!
b110 %
1'
b110 +
#863390000000
0!
0'
#863400000000
1!
b111 %
1'
b111 +
#863410000000
0!
0'
#863420000000
1!
0$
b1000 %
1'
0*
b1000 +
#863430000000
0!
0'
#863440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#863450000000
0!
0'
#863460000000
1!
b0 %
1'
b0 +
#863470000000
0!
0'
#863480000000
1!
1$
b1 %
1'
1*
b1 +
#863490000000
0!
0'
#863500000000
1!
b10 %
1'
b10 +
#863510000000
0!
0'
#863520000000
1!
b11 %
1'
b11 +
#863530000000
0!
0'
#863540000000
1!
b100 %
1'
b100 +
#863550000000
0!
0'
#863560000000
1!
b101 %
1'
b101 +
#863570000000
0!
0'
#863580000000
1!
0$
b110 %
1'
0*
b110 +
#863590000000
0!
0'
#863600000000
1!
b111 %
1'
b111 +
#863610000000
0!
0'
#863620000000
1!
b1000 %
1'
b1000 +
#863630000000
0!
0'
#863640000000
1!
b1001 %
1'
b1001 +
#863650000000
1"
1(
#863660000000
0!
0"
b100 &
0'
0(
b100 ,
#863670000000
1!
b0 %
1'
b0 +
#863680000000
0!
0'
#863690000000
1!
1$
b1 %
1'
1*
b1 +
#863700000000
0!
0'
#863710000000
1!
b10 %
1'
b10 +
#863720000000
0!
0'
#863730000000
1!
b11 %
1'
b11 +
#863740000000
0!
0'
#863750000000
1!
b100 %
1'
b100 +
#863760000000
0!
0'
#863770000000
1!
b101 %
1'
b101 +
#863780000000
0!
0'
#863790000000
1!
b110 %
1'
b110 +
#863800000000
0!
0'
#863810000000
1!
b111 %
1'
b111 +
#863820000000
0!
0'
#863830000000
1!
0$
b1000 %
1'
0*
b1000 +
#863840000000
0!
0'
#863850000000
1!
b1001 %
1'
b1001 +
#863860000000
0!
0'
#863870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#863880000000
0!
0'
#863890000000
1!
1$
b1 %
1'
1*
b1 +
#863900000000
0!
0'
#863910000000
1!
b10 %
1'
b10 +
#863920000000
0!
0'
#863930000000
1!
b11 %
1'
b11 +
#863940000000
0!
0'
#863950000000
1!
b100 %
1'
b100 +
#863960000000
0!
0'
#863970000000
1!
b101 %
1'
b101 +
#863980000000
0!
0'
#863990000000
1!
0$
b110 %
1'
0*
b110 +
#864000000000
0!
0'
#864010000000
1!
b111 %
1'
b111 +
#864020000000
0!
0'
#864030000000
1!
b1000 %
1'
b1000 +
#864040000000
0!
0'
#864050000000
1!
b1001 %
1'
b1001 +
#864060000000
0!
0'
#864070000000
1!
b0 %
1'
b0 +
#864080000000
1"
1(
#864090000000
0!
0"
b100 &
0'
0(
b100 ,
#864100000000
1!
1$
b1 %
1'
1*
b1 +
#864110000000
0!
0'
#864120000000
1!
b10 %
1'
b10 +
#864130000000
0!
0'
#864140000000
1!
b11 %
1'
b11 +
#864150000000
0!
0'
#864160000000
1!
b100 %
1'
b100 +
#864170000000
0!
0'
#864180000000
1!
b101 %
1'
b101 +
#864190000000
0!
0'
#864200000000
1!
b110 %
1'
b110 +
#864210000000
0!
0'
#864220000000
1!
b111 %
1'
b111 +
#864230000000
0!
0'
#864240000000
1!
0$
b1000 %
1'
0*
b1000 +
#864250000000
0!
0'
#864260000000
1!
b1001 %
1'
b1001 +
#864270000000
0!
0'
#864280000000
1!
b0 %
1'
b0 +
#864290000000
0!
0'
#864300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#864310000000
0!
0'
#864320000000
1!
b10 %
1'
b10 +
#864330000000
0!
0'
#864340000000
1!
b11 %
1'
b11 +
#864350000000
0!
0'
#864360000000
1!
b100 %
1'
b100 +
#864370000000
0!
0'
#864380000000
1!
b101 %
1'
b101 +
#864390000000
0!
0'
#864400000000
1!
0$
b110 %
1'
0*
b110 +
#864410000000
0!
0'
#864420000000
1!
b111 %
1'
b111 +
#864430000000
0!
0'
#864440000000
1!
b1000 %
1'
b1000 +
#864450000000
0!
0'
#864460000000
1!
b1001 %
1'
b1001 +
#864470000000
0!
0'
#864480000000
1!
b0 %
1'
b0 +
#864490000000
0!
0'
#864500000000
1!
1$
b1 %
1'
1*
b1 +
#864510000000
1"
1(
#864520000000
0!
0"
b100 &
0'
0(
b100 ,
#864530000000
1!
b10 %
1'
b10 +
#864540000000
0!
0'
#864550000000
1!
b11 %
1'
b11 +
#864560000000
0!
0'
#864570000000
1!
b100 %
1'
b100 +
#864580000000
0!
0'
#864590000000
1!
b101 %
1'
b101 +
#864600000000
0!
0'
#864610000000
1!
b110 %
1'
b110 +
#864620000000
0!
0'
#864630000000
1!
b111 %
1'
b111 +
#864640000000
0!
0'
#864650000000
1!
0$
b1000 %
1'
0*
b1000 +
#864660000000
0!
0'
#864670000000
1!
b1001 %
1'
b1001 +
#864680000000
0!
0'
#864690000000
1!
b0 %
1'
b0 +
#864700000000
0!
0'
#864710000000
1!
1$
b1 %
1'
1*
b1 +
#864720000000
0!
0'
#864730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#864740000000
0!
0'
#864750000000
1!
b11 %
1'
b11 +
#864760000000
0!
0'
#864770000000
1!
b100 %
1'
b100 +
#864780000000
0!
0'
#864790000000
1!
b101 %
1'
b101 +
#864800000000
0!
0'
#864810000000
1!
0$
b110 %
1'
0*
b110 +
#864820000000
0!
0'
#864830000000
1!
b111 %
1'
b111 +
#864840000000
0!
0'
#864850000000
1!
b1000 %
1'
b1000 +
#864860000000
0!
0'
#864870000000
1!
b1001 %
1'
b1001 +
#864880000000
0!
0'
#864890000000
1!
b0 %
1'
b0 +
#864900000000
0!
0'
#864910000000
1!
1$
b1 %
1'
1*
b1 +
#864920000000
0!
0'
#864930000000
1!
b10 %
1'
b10 +
#864940000000
1"
1(
#864950000000
0!
0"
b100 &
0'
0(
b100 ,
#864960000000
1!
b11 %
1'
b11 +
#864970000000
0!
0'
#864980000000
1!
b100 %
1'
b100 +
#864990000000
0!
0'
#865000000000
1!
b101 %
1'
b101 +
#865010000000
0!
0'
#865020000000
1!
b110 %
1'
b110 +
#865030000000
0!
0'
#865040000000
1!
b111 %
1'
b111 +
#865050000000
0!
0'
#865060000000
1!
0$
b1000 %
1'
0*
b1000 +
#865070000000
0!
0'
#865080000000
1!
b1001 %
1'
b1001 +
#865090000000
0!
0'
#865100000000
1!
b0 %
1'
b0 +
#865110000000
0!
0'
#865120000000
1!
1$
b1 %
1'
1*
b1 +
#865130000000
0!
0'
#865140000000
1!
b10 %
1'
b10 +
#865150000000
0!
0'
#865160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#865170000000
0!
0'
#865180000000
1!
b100 %
1'
b100 +
#865190000000
0!
0'
#865200000000
1!
b101 %
1'
b101 +
#865210000000
0!
0'
#865220000000
1!
0$
b110 %
1'
0*
b110 +
#865230000000
0!
0'
#865240000000
1!
b111 %
1'
b111 +
#865250000000
0!
0'
#865260000000
1!
b1000 %
1'
b1000 +
#865270000000
0!
0'
#865280000000
1!
b1001 %
1'
b1001 +
#865290000000
0!
0'
#865300000000
1!
b0 %
1'
b0 +
#865310000000
0!
0'
#865320000000
1!
1$
b1 %
1'
1*
b1 +
#865330000000
0!
0'
#865340000000
1!
b10 %
1'
b10 +
#865350000000
0!
0'
#865360000000
1!
b11 %
1'
b11 +
#865370000000
1"
1(
#865380000000
0!
0"
b100 &
0'
0(
b100 ,
#865390000000
1!
b100 %
1'
b100 +
#865400000000
0!
0'
#865410000000
1!
b101 %
1'
b101 +
#865420000000
0!
0'
#865430000000
1!
b110 %
1'
b110 +
#865440000000
0!
0'
#865450000000
1!
b111 %
1'
b111 +
#865460000000
0!
0'
#865470000000
1!
0$
b1000 %
1'
0*
b1000 +
#865480000000
0!
0'
#865490000000
1!
b1001 %
1'
b1001 +
#865500000000
0!
0'
#865510000000
1!
b0 %
1'
b0 +
#865520000000
0!
0'
#865530000000
1!
1$
b1 %
1'
1*
b1 +
#865540000000
0!
0'
#865550000000
1!
b10 %
1'
b10 +
#865560000000
0!
0'
#865570000000
1!
b11 %
1'
b11 +
#865580000000
0!
0'
#865590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#865600000000
0!
0'
#865610000000
1!
b101 %
1'
b101 +
#865620000000
0!
0'
#865630000000
1!
0$
b110 %
1'
0*
b110 +
#865640000000
0!
0'
#865650000000
1!
b111 %
1'
b111 +
#865660000000
0!
0'
#865670000000
1!
b1000 %
1'
b1000 +
#865680000000
0!
0'
#865690000000
1!
b1001 %
1'
b1001 +
#865700000000
0!
0'
#865710000000
1!
b0 %
1'
b0 +
#865720000000
0!
0'
#865730000000
1!
1$
b1 %
1'
1*
b1 +
#865740000000
0!
0'
#865750000000
1!
b10 %
1'
b10 +
#865760000000
0!
0'
#865770000000
1!
b11 %
1'
b11 +
#865780000000
0!
0'
#865790000000
1!
b100 %
1'
b100 +
#865800000000
1"
1(
#865810000000
0!
0"
b100 &
0'
0(
b100 ,
#865820000000
1!
b101 %
1'
b101 +
#865830000000
0!
0'
#865840000000
1!
b110 %
1'
b110 +
#865850000000
0!
0'
#865860000000
1!
b111 %
1'
b111 +
#865870000000
0!
0'
#865880000000
1!
0$
b1000 %
1'
0*
b1000 +
#865890000000
0!
0'
#865900000000
1!
b1001 %
1'
b1001 +
#865910000000
0!
0'
#865920000000
1!
b0 %
1'
b0 +
#865930000000
0!
0'
#865940000000
1!
1$
b1 %
1'
1*
b1 +
#865950000000
0!
0'
#865960000000
1!
b10 %
1'
b10 +
#865970000000
0!
0'
#865980000000
1!
b11 %
1'
b11 +
#865990000000
0!
0'
#866000000000
1!
b100 %
1'
b100 +
#866010000000
0!
0'
#866020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#866030000000
0!
0'
#866040000000
1!
0$
b110 %
1'
0*
b110 +
#866050000000
0!
0'
#866060000000
1!
b111 %
1'
b111 +
#866070000000
0!
0'
#866080000000
1!
b1000 %
1'
b1000 +
#866090000000
0!
0'
#866100000000
1!
b1001 %
1'
b1001 +
#866110000000
0!
0'
#866120000000
1!
b0 %
1'
b0 +
#866130000000
0!
0'
#866140000000
1!
1$
b1 %
1'
1*
b1 +
#866150000000
0!
0'
#866160000000
1!
b10 %
1'
b10 +
#866170000000
0!
0'
#866180000000
1!
b11 %
1'
b11 +
#866190000000
0!
0'
#866200000000
1!
b100 %
1'
b100 +
#866210000000
0!
0'
#866220000000
1!
b101 %
1'
b101 +
#866230000000
1"
1(
#866240000000
0!
0"
b100 &
0'
0(
b100 ,
#866250000000
1!
b110 %
1'
b110 +
#866260000000
0!
0'
#866270000000
1!
b111 %
1'
b111 +
#866280000000
0!
0'
#866290000000
1!
0$
b1000 %
1'
0*
b1000 +
#866300000000
0!
0'
#866310000000
1!
b1001 %
1'
b1001 +
#866320000000
0!
0'
#866330000000
1!
b0 %
1'
b0 +
#866340000000
0!
0'
#866350000000
1!
1$
b1 %
1'
1*
b1 +
#866360000000
0!
0'
#866370000000
1!
b10 %
1'
b10 +
#866380000000
0!
0'
#866390000000
1!
b11 %
1'
b11 +
#866400000000
0!
0'
#866410000000
1!
b100 %
1'
b100 +
#866420000000
0!
0'
#866430000000
1!
b101 %
1'
b101 +
#866440000000
0!
0'
#866450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#866460000000
0!
0'
#866470000000
1!
b111 %
1'
b111 +
#866480000000
0!
0'
#866490000000
1!
b1000 %
1'
b1000 +
#866500000000
0!
0'
#866510000000
1!
b1001 %
1'
b1001 +
#866520000000
0!
0'
#866530000000
1!
b0 %
1'
b0 +
#866540000000
0!
0'
#866550000000
1!
1$
b1 %
1'
1*
b1 +
#866560000000
0!
0'
#866570000000
1!
b10 %
1'
b10 +
#866580000000
0!
0'
#866590000000
1!
b11 %
1'
b11 +
#866600000000
0!
0'
#866610000000
1!
b100 %
1'
b100 +
#866620000000
0!
0'
#866630000000
1!
b101 %
1'
b101 +
#866640000000
0!
0'
#866650000000
1!
0$
b110 %
1'
0*
b110 +
#866660000000
1"
1(
#866670000000
0!
0"
b100 &
0'
0(
b100 ,
#866680000000
1!
1$
b111 %
1'
1*
b111 +
#866690000000
0!
0'
#866700000000
1!
0$
b1000 %
1'
0*
b1000 +
#866710000000
0!
0'
#866720000000
1!
b1001 %
1'
b1001 +
#866730000000
0!
0'
#866740000000
1!
b0 %
1'
b0 +
#866750000000
0!
0'
#866760000000
1!
1$
b1 %
1'
1*
b1 +
#866770000000
0!
0'
#866780000000
1!
b10 %
1'
b10 +
#866790000000
0!
0'
#866800000000
1!
b11 %
1'
b11 +
#866810000000
0!
0'
#866820000000
1!
b100 %
1'
b100 +
#866830000000
0!
0'
#866840000000
1!
b101 %
1'
b101 +
#866850000000
0!
0'
#866860000000
1!
b110 %
1'
b110 +
#866870000000
0!
0'
#866880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#866890000000
0!
0'
#866900000000
1!
b1000 %
1'
b1000 +
#866910000000
0!
0'
#866920000000
1!
b1001 %
1'
b1001 +
#866930000000
0!
0'
#866940000000
1!
b0 %
1'
b0 +
#866950000000
0!
0'
#866960000000
1!
1$
b1 %
1'
1*
b1 +
#866970000000
0!
0'
#866980000000
1!
b10 %
1'
b10 +
#866990000000
0!
0'
#867000000000
1!
b11 %
1'
b11 +
#867010000000
0!
0'
#867020000000
1!
b100 %
1'
b100 +
#867030000000
0!
0'
#867040000000
1!
b101 %
1'
b101 +
#867050000000
0!
0'
#867060000000
1!
0$
b110 %
1'
0*
b110 +
#867070000000
0!
0'
#867080000000
1!
b111 %
1'
b111 +
#867090000000
1"
1(
#867100000000
0!
0"
b100 &
0'
0(
b100 ,
#867110000000
1!
b1000 %
1'
b1000 +
#867120000000
0!
0'
#867130000000
1!
b1001 %
1'
b1001 +
#867140000000
0!
0'
#867150000000
1!
b0 %
1'
b0 +
#867160000000
0!
0'
#867170000000
1!
1$
b1 %
1'
1*
b1 +
#867180000000
0!
0'
#867190000000
1!
b10 %
1'
b10 +
#867200000000
0!
0'
#867210000000
1!
b11 %
1'
b11 +
#867220000000
0!
0'
#867230000000
1!
b100 %
1'
b100 +
#867240000000
0!
0'
#867250000000
1!
b101 %
1'
b101 +
#867260000000
0!
0'
#867270000000
1!
b110 %
1'
b110 +
#867280000000
0!
0'
#867290000000
1!
b111 %
1'
b111 +
#867300000000
0!
0'
#867310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#867320000000
0!
0'
#867330000000
1!
b1001 %
1'
b1001 +
#867340000000
0!
0'
#867350000000
1!
b0 %
1'
b0 +
#867360000000
0!
0'
#867370000000
1!
1$
b1 %
1'
1*
b1 +
#867380000000
0!
0'
#867390000000
1!
b10 %
1'
b10 +
#867400000000
0!
0'
#867410000000
1!
b11 %
1'
b11 +
#867420000000
0!
0'
#867430000000
1!
b100 %
1'
b100 +
#867440000000
0!
0'
#867450000000
1!
b101 %
1'
b101 +
#867460000000
0!
0'
#867470000000
1!
0$
b110 %
1'
0*
b110 +
#867480000000
0!
0'
#867490000000
1!
b111 %
1'
b111 +
#867500000000
0!
0'
#867510000000
1!
b1000 %
1'
b1000 +
#867520000000
1"
1(
#867530000000
0!
0"
b100 &
0'
0(
b100 ,
#867540000000
1!
b1001 %
1'
b1001 +
#867550000000
0!
0'
#867560000000
1!
b0 %
1'
b0 +
#867570000000
0!
0'
#867580000000
1!
1$
b1 %
1'
1*
b1 +
#867590000000
0!
0'
#867600000000
1!
b10 %
1'
b10 +
#867610000000
0!
0'
#867620000000
1!
b11 %
1'
b11 +
#867630000000
0!
0'
#867640000000
1!
b100 %
1'
b100 +
#867650000000
0!
0'
#867660000000
1!
b101 %
1'
b101 +
#867670000000
0!
0'
#867680000000
1!
b110 %
1'
b110 +
#867690000000
0!
0'
#867700000000
1!
b111 %
1'
b111 +
#867710000000
0!
0'
#867720000000
1!
0$
b1000 %
1'
0*
b1000 +
#867730000000
0!
0'
#867740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#867750000000
0!
0'
#867760000000
1!
b0 %
1'
b0 +
#867770000000
0!
0'
#867780000000
1!
1$
b1 %
1'
1*
b1 +
#867790000000
0!
0'
#867800000000
1!
b10 %
1'
b10 +
#867810000000
0!
0'
#867820000000
1!
b11 %
1'
b11 +
#867830000000
0!
0'
#867840000000
1!
b100 %
1'
b100 +
#867850000000
0!
0'
#867860000000
1!
b101 %
1'
b101 +
#867870000000
0!
0'
#867880000000
1!
0$
b110 %
1'
0*
b110 +
#867890000000
0!
0'
#867900000000
1!
b111 %
1'
b111 +
#867910000000
0!
0'
#867920000000
1!
b1000 %
1'
b1000 +
#867930000000
0!
0'
#867940000000
1!
b1001 %
1'
b1001 +
#867950000000
1"
1(
#867960000000
0!
0"
b100 &
0'
0(
b100 ,
#867970000000
1!
b0 %
1'
b0 +
#867980000000
0!
0'
#867990000000
1!
1$
b1 %
1'
1*
b1 +
#868000000000
0!
0'
#868010000000
1!
b10 %
1'
b10 +
#868020000000
0!
0'
#868030000000
1!
b11 %
1'
b11 +
#868040000000
0!
0'
#868050000000
1!
b100 %
1'
b100 +
#868060000000
0!
0'
#868070000000
1!
b101 %
1'
b101 +
#868080000000
0!
0'
#868090000000
1!
b110 %
1'
b110 +
#868100000000
0!
0'
#868110000000
1!
b111 %
1'
b111 +
#868120000000
0!
0'
#868130000000
1!
0$
b1000 %
1'
0*
b1000 +
#868140000000
0!
0'
#868150000000
1!
b1001 %
1'
b1001 +
#868160000000
0!
0'
#868170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#868180000000
0!
0'
#868190000000
1!
1$
b1 %
1'
1*
b1 +
#868200000000
0!
0'
#868210000000
1!
b10 %
1'
b10 +
#868220000000
0!
0'
#868230000000
1!
b11 %
1'
b11 +
#868240000000
0!
0'
#868250000000
1!
b100 %
1'
b100 +
#868260000000
0!
0'
#868270000000
1!
b101 %
1'
b101 +
#868280000000
0!
0'
#868290000000
1!
0$
b110 %
1'
0*
b110 +
#868300000000
0!
0'
#868310000000
1!
b111 %
1'
b111 +
#868320000000
0!
0'
#868330000000
1!
b1000 %
1'
b1000 +
#868340000000
0!
0'
#868350000000
1!
b1001 %
1'
b1001 +
#868360000000
0!
0'
#868370000000
1!
b0 %
1'
b0 +
#868380000000
1"
1(
#868390000000
0!
0"
b100 &
0'
0(
b100 ,
#868400000000
1!
1$
b1 %
1'
1*
b1 +
#868410000000
0!
0'
#868420000000
1!
b10 %
1'
b10 +
#868430000000
0!
0'
#868440000000
1!
b11 %
1'
b11 +
#868450000000
0!
0'
#868460000000
1!
b100 %
1'
b100 +
#868470000000
0!
0'
#868480000000
1!
b101 %
1'
b101 +
#868490000000
0!
0'
#868500000000
1!
b110 %
1'
b110 +
#868510000000
0!
0'
#868520000000
1!
b111 %
1'
b111 +
#868530000000
0!
0'
#868540000000
1!
0$
b1000 %
1'
0*
b1000 +
#868550000000
0!
0'
#868560000000
1!
b1001 %
1'
b1001 +
#868570000000
0!
0'
#868580000000
1!
b0 %
1'
b0 +
#868590000000
0!
0'
#868600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#868610000000
0!
0'
#868620000000
1!
b10 %
1'
b10 +
#868630000000
0!
0'
#868640000000
1!
b11 %
1'
b11 +
#868650000000
0!
0'
#868660000000
1!
b100 %
1'
b100 +
#868670000000
0!
0'
#868680000000
1!
b101 %
1'
b101 +
#868690000000
0!
0'
#868700000000
1!
0$
b110 %
1'
0*
b110 +
#868710000000
0!
0'
#868720000000
1!
b111 %
1'
b111 +
#868730000000
0!
0'
#868740000000
1!
b1000 %
1'
b1000 +
#868750000000
0!
0'
#868760000000
1!
b1001 %
1'
b1001 +
#868770000000
0!
0'
#868780000000
1!
b0 %
1'
b0 +
#868790000000
0!
0'
#868800000000
1!
1$
b1 %
1'
1*
b1 +
#868810000000
1"
1(
#868820000000
0!
0"
b100 &
0'
0(
b100 ,
#868830000000
1!
b10 %
1'
b10 +
#868840000000
0!
0'
#868850000000
1!
b11 %
1'
b11 +
#868860000000
0!
0'
#868870000000
1!
b100 %
1'
b100 +
#868880000000
0!
0'
#868890000000
1!
b101 %
1'
b101 +
#868900000000
0!
0'
#868910000000
1!
b110 %
1'
b110 +
#868920000000
0!
0'
#868930000000
1!
b111 %
1'
b111 +
#868940000000
0!
0'
#868950000000
1!
0$
b1000 %
1'
0*
b1000 +
#868960000000
0!
0'
#868970000000
1!
b1001 %
1'
b1001 +
#868980000000
0!
0'
#868990000000
1!
b0 %
1'
b0 +
#869000000000
0!
0'
#869010000000
1!
1$
b1 %
1'
1*
b1 +
#869020000000
0!
0'
#869030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#869040000000
0!
0'
#869050000000
1!
b11 %
1'
b11 +
#869060000000
0!
0'
#869070000000
1!
b100 %
1'
b100 +
#869080000000
0!
0'
#869090000000
1!
b101 %
1'
b101 +
#869100000000
0!
0'
#869110000000
1!
0$
b110 %
1'
0*
b110 +
#869120000000
0!
0'
#869130000000
1!
b111 %
1'
b111 +
#869140000000
0!
0'
#869150000000
1!
b1000 %
1'
b1000 +
#869160000000
0!
0'
#869170000000
1!
b1001 %
1'
b1001 +
#869180000000
0!
0'
#869190000000
1!
b0 %
1'
b0 +
#869200000000
0!
0'
#869210000000
1!
1$
b1 %
1'
1*
b1 +
#869220000000
0!
0'
#869230000000
1!
b10 %
1'
b10 +
#869240000000
1"
1(
#869250000000
0!
0"
b100 &
0'
0(
b100 ,
#869260000000
1!
b11 %
1'
b11 +
#869270000000
0!
0'
#869280000000
1!
b100 %
1'
b100 +
#869290000000
0!
0'
#869300000000
1!
b101 %
1'
b101 +
#869310000000
0!
0'
#869320000000
1!
b110 %
1'
b110 +
#869330000000
0!
0'
#869340000000
1!
b111 %
1'
b111 +
#869350000000
0!
0'
#869360000000
1!
0$
b1000 %
1'
0*
b1000 +
#869370000000
0!
0'
#869380000000
1!
b1001 %
1'
b1001 +
#869390000000
0!
0'
#869400000000
1!
b0 %
1'
b0 +
#869410000000
0!
0'
#869420000000
1!
1$
b1 %
1'
1*
b1 +
#869430000000
0!
0'
#869440000000
1!
b10 %
1'
b10 +
#869450000000
0!
0'
#869460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#869470000000
0!
0'
#869480000000
1!
b100 %
1'
b100 +
#869490000000
0!
0'
#869500000000
1!
b101 %
1'
b101 +
#869510000000
0!
0'
#869520000000
1!
0$
b110 %
1'
0*
b110 +
#869530000000
0!
0'
#869540000000
1!
b111 %
1'
b111 +
#869550000000
0!
0'
#869560000000
1!
b1000 %
1'
b1000 +
#869570000000
0!
0'
#869580000000
1!
b1001 %
1'
b1001 +
#869590000000
0!
0'
#869600000000
1!
b0 %
1'
b0 +
#869610000000
0!
0'
#869620000000
1!
1$
b1 %
1'
1*
b1 +
#869630000000
0!
0'
#869640000000
1!
b10 %
1'
b10 +
#869650000000
0!
0'
#869660000000
1!
b11 %
1'
b11 +
#869670000000
1"
1(
#869680000000
0!
0"
b100 &
0'
0(
b100 ,
#869690000000
1!
b100 %
1'
b100 +
#869700000000
0!
0'
#869710000000
1!
b101 %
1'
b101 +
#869720000000
0!
0'
#869730000000
1!
b110 %
1'
b110 +
#869740000000
0!
0'
#869750000000
1!
b111 %
1'
b111 +
#869760000000
0!
0'
#869770000000
1!
0$
b1000 %
1'
0*
b1000 +
#869780000000
0!
0'
#869790000000
1!
b1001 %
1'
b1001 +
#869800000000
0!
0'
#869810000000
1!
b0 %
1'
b0 +
#869820000000
0!
0'
#869830000000
1!
1$
b1 %
1'
1*
b1 +
#869840000000
0!
0'
#869850000000
1!
b10 %
1'
b10 +
#869860000000
0!
0'
#869870000000
1!
b11 %
1'
b11 +
#869880000000
0!
0'
#869890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#869900000000
0!
0'
#869910000000
1!
b101 %
1'
b101 +
#869920000000
0!
0'
#869930000000
1!
0$
b110 %
1'
0*
b110 +
#869940000000
0!
0'
#869950000000
1!
b111 %
1'
b111 +
#869960000000
0!
0'
#869970000000
1!
b1000 %
1'
b1000 +
#869980000000
0!
0'
#869990000000
1!
b1001 %
1'
b1001 +
#870000000000
0!
0'
#870010000000
1!
b0 %
1'
b0 +
#870020000000
0!
0'
#870030000000
1!
1$
b1 %
1'
1*
b1 +
#870040000000
0!
0'
#870050000000
1!
b10 %
1'
b10 +
#870060000000
0!
0'
#870070000000
1!
b11 %
1'
b11 +
#870080000000
0!
0'
#870090000000
1!
b100 %
1'
b100 +
#870100000000
1"
1(
#870110000000
0!
0"
b100 &
0'
0(
b100 ,
#870120000000
1!
b101 %
1'
b101 +
#870130000000
0!
0'
#870140000000
1!
b110 %
1'
b110 +
#870150000000
0!
0'
#870160000000
1!
b111 %
1'
b111 +
#870170000000
0!
0'
#870180000000
1!
0$
b1000 %
1'
0*
b1000 +
#870190000000
0!
0'
#870200000000
1!
b1001 %
1'
b1001 +
#870210000000
0!
0'
#870220000000
1!
b0 %
1'
b0 +
#870230000000
0!
0'
#870240000000
1!
1$
b1 %
1'
1*
b1 +
#870250000000
0!
0'
#870260000000
1!
b10 %
1'
b10 +
#870270000000
0!
0'
#870280000000
1!
b11 %
1'
b11 +
#870290000000
0!
0'
#870300000000
1!
b100 %
1'
b100 +
#870310000000
0!
0'
#870320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#870330000000
0!
0'
#870340000000
1!
0$
b110 %
1'
0*
b110 +
#870350000000
0!
0'
#870360000000
1!
b111 %
1'
b111 +
#870370000000
0!
0'
#870380000000
1!
b1000 %
1'
b1000 +
#870390000000
0!
0'
#870400000000
1!
b1001 %
1'
b1001 +
#870410000000
0!
0'
#870420000000
1!
b0 %
1'
b0 +
#870430000000
0!
0'
#870440000000
1!
1$
b1 %
1'
1*
b1 +
#870450000000
0!
0'
#870460000000
1!
b10 %
1'
b10 +
#870470000000
0!
0'
#870480000000
1!
b11 %
1'
b11 +
#870490000000
0!
0'
#870500000000
1!
b100 %
1'
b100 +
#870510000000
0!
0'
#870520000000
1!
b101 %
1'
b101 +
#870530000000
1"
1(
#870540000000
0!
0"
b100 &
0'
0(
b100 ,
#870550000000
1!
b110 %
1'
b110 +
#870560000000
0!
0'
#870570000000
1!
b111 %
1'
b111 +
#870580000000
0!
0'
#870590000000
1!
0$
b1000 %
1'
0*
b1000 +
#870600000000
0!
0'
#870610000000
1!
b1001 %
1'
b1001 +
#870620000000
0!
0'
#870630000000
1!
b0 %
1'
b0 +
#870640000000
0!
0'
#870650000000
1!
1$
b1 %
1'
1*
b1 +
#870660000000
0!
0'
#870670000000
1!
b10 %
1'
b10 +
#870680000000
0!
0'
#870690000000
1!
b11 %
1'
b11 +
#870700000000
0!
0'
#870710000000
1!
b100 %
1'
b100 +
#870720000000
0!
0'
#870730000000
1!
b101 %
1'
b101 +
#870740000000
0!
0'
#870750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#870760000000
0!
0'
#870770000000
1!
b111 %
1'
b111 +
#870780000000
0!
0'
#870790000000
1!
b1000 %
1'
b1000 +
#870800000000
0!
0'
#870810000000
1!
b1001 %
1'
b1001 +
#870820000000
0!
0'
#870830000000
1!
b0 %
1'
b0 +
#870840000000
0!
0'
#870850000000
1!
1$
b1 %
1'
1*
b1 +
#870860000000
0!
0'
#870870000000
1!
b10 %
1'
b10 +
#870880000000
0!
0'
#870890000000
1!
b11 %
1'
b11 +
#870900000000
0!
0'
#870910000000
1!
b100 %
1'
b100 +
#870920000000
0!
0'
#870930000000
1!
b101 %
1'
b101 +
#870940000000
0!
0'
#870950000000
1!
0$
b110 %
1'
0*
b110 +
#870960000000
1"
1(
#870970000000
0!
0"
b100 &
0'
0(
b100 ,
#870980000000
1!
1$
b111 %
1'
1*
b111 +
#870990000000
0!
0'
#871000000000
1!
0$
b1000 %
1'
0*
b1000 +
#871010000000
0!
0'
#871020000000
1!
b1001 %
1'
b1001 +
#871030000000
0!
0'
#871040000000
1!
b0 %
1'
b0 +
#871050000000
0!
0'
#871060000000
1!
1$
b1 %
1'
1*
b1 +
#871070000000
0!
0'
#871080000000
1!
b10 %
1'
b10 +
#871090000000
0!
0'
#871100000000
1!
b11 %
1'
b11 +
#871110000000
0!
0'
#871120000000
1!
b100 %
1'
b100 +
#871130000000
0!
0'
#871140000000
1!
b101 %
1'
b101 +
#871150000000
0!
0'
#871160000000
1!
b110 %
1'
b110 +
#871170000000
0!
0'
#871180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#871190000000
0!
0'
#871200000000
1!
b1000 %
1'
b1000 +
#871210000000
0!
0'
#871220000000
1!
b1001 %
1'
b1001 +
#871230000000
0!
0'
#871240000000
1!
b0 %
1'
b0 +
#871250000000
0!
0'
#871260000000
1!
1$
b1 %
1'
1*
b1 +
#871270000000
0!
0'
#871280000000
1!
b10 %
1'
b10 +
#871290000000
0!
0'
#871300000000
1!
b11 %
1'
b11 +
#871310000000
0!
0'
#871320000000
1!
b100 %
1'
b100 +
#871330000000
0!
0'
#871340000000
1!
b101 %
1'
b101 +
#871350000000
0!
0'
#871360000000
1!
0$
b110 %
1'
0*
b110 +
#871370000000
0!
0'
#871380000000
1!
b111 %
1'
b111 +
#871390000000
1"
1(
#871400000000
0!
0"
b100 &
0'
0(
b100 ,
#871410000000
1!
b1000 %
1'
b1000 +
#871420000000
0!
0'
#871430000000
1!
b1001 %
1'
b1001 +
#871440000000
0!
0'
#871450000000
1!
b0 %
1'
b0 +
#871460000000
0!
0'
#871470000000
1!
1$
b1 %
1'
1*
b1 +
#871480000000
0!
0'
#871490000000
1!
b10 %
1'
b10 +
#871500000000
0!
0'
#871510000000
1!
b11 %
1'
b11 +
#871520000000
0!
0'
#871530000000
1!
b100 %
1'
b100 +
#871540000000
0!
0'
#871550000000
1!
b101 %
1'
b101 +
#871560000000
0!
0'
#871570000000
1!
b110 %
1'
b110 +
#871580000000
0!
0'
#871590000000
1!
b111 %
1'
b111 +
#871600000000
0!
0'
#871610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#871620000000
0!
0'
#871630000000
1!
b1001 %
1'
b1001 +
#871640000000
0!
0'
#871650000000
1!
b0 %
1'
b0 +
#871660000000
0!
0'
#871670000000
1!
1$
b1 %
1'
1*
b1 +
#871680000000
0!
0'
#871690000000
1!
b10 %
1'
b10 +
#871700000000
0!
0'
#871710000000
1!
b11 %
1'
b11 +
#871720000000
0!
0'
#871730000000
1!
b100 %
1'
b100 +
#871740000000
0!
0'
#871750000000
1!
b101 %
1'
b101 +
#871760000000
0!
0'
#871770000000
1!
0$
b110 %
1'
0*
b110 +
#871780000000
0!
0'
#871790000000
1!
b111 %
1'
b111 +
#871800000000
0!
0'
#871810000000
1!
b1000 %
1'
b1000 +
#871820000000
1"
1(
#871830000000
0!
0"
b100 &
0'
0(
b100 ,
#871840000000
1!
b1001 %
1'
b1001 +
#871850000000
0!
0'
#871860000000
1!
b0 %
1'
b0 +
#871870000000
0!
0'
#871880000000
1!
1$
b1 %
1'
1*
b1 +
#871890000000
0!
0'
#871900000000
1!
b10 %
1'
b10 +
#871910000000
0!
0'
#871920000000
1!
b11 %
1'
b11 +
#871930000000
0!
0'
#871940000000
1!
b100 %
1'
b100 +
#871950000000
0!
0'
#871960000000
1!
b101 %
1'
b101 +
#871970000000
0!
0'
#871980000000
1!
b110 %
1'
b110 +
#871990000000
0!
0'
#872000000000
1!
b111 %
1'
b111 +
#872010000000
0!
0'
#872020000000
1!
0$
b1000 %
1'
0*
b1000 +
#872030000000
0!
0'
#872040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#872050000000
0!
0'
#872060000000
1!
b0 %
1'
b0 +
#872070000000
0!
0'
#872080000000
1!
1$
b1 %
1'
1*
b1 +
#872090000000
0!
0'
#872100000000
1!
b10 %
1'
b10 +
#872110000000
0!
0'
#872120000000
1!
b11 %
1'
b11 +
#872130000000
0!
0'
#872140000000
1!
b100 %
1'
b100 +
#872150000000
0!
0'
#872160000000
1!
b101 %
1'
b101 +
#872170000000
0!
0'
#872180000000
1!
0$
b110 %
1'
0*
b110 +
#872190000000
0!
0'
#872200000000
1!
b111 %
1'
b111 +
#872210000000
0!
0'
#872220000000
1!
b1000 %
1'
b1000 +
#872230000000
0!
0'
#872240000000
1!
b1001 %
1'
b1001 +
#872250000000
1"
1(
#872260000000
0!
0"
b100 &
0'
0(
b100 ,
#872270000000
1!
b0 %
1'
b0 +
#872280000000
0!
0'
#872290000000
1!
1$
b1 %
1'
1*
b1 +
#872300000000
0!
0'
#872310000000
1!
b10 %
1'
b10 +
#872320000000
0!
0'
#872330000000
1!
b11 %
1'
b11 +
#872340000000
0!
0'
#872350000000
1!
b100 %
1'
b100 +
#872360000000
0!
0'
#872370000000
1!
b101 %
1'
b101 +
#872380000000
0!
0'
#872390000000
1!
b110 %
1'
b110 +
#872400000000
0!
0'
#872410000000
1!
b111 %
1'
b111 +
#872420000000
0!
0'
#872430000000
1!
0$
b1000 %
1'
0*
b1000 +
#872440000000
0!
0'
#872450000000
1!
b1001 %
1'
b1001 +
#872460000000
0!
0'
#872470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#872480000000
0!
0'
#872490000000
1!
1$
b1 %
1'
1*
b1 +
#872500000000
0!
0'
#872510000000
1!
b10 %
1'
b10 +
#872520000000
0!
0'
#872530000000
1!
b11 %
1'
b11 +
#872540000000
0!
0'
#872550000000
1!
b100 %
1'
b100 +
#872560000000
0!
0'
#872570000000
1!
b101 %
1'
b101 +
#872580000000
0!
0'
#872590000000
1!
0$
b110 %
1'
0*
b110 +
#872600000000
0!
0'
#872610000000
1!
b111 %
1'
b111 +
#872620000000
0!
0'
#872630000000
1!
b1000 %
1'
b1000 +
#872640000000
0!
0'
#872650000000
1!
b1001 %
1'
b1001 +
#872660000000
0!
0'
#872670000000
1!
b0 %
1'
b0 +
#872680000000
1"
1(
#872690000000
0!
0"
b100 &
0'
0(
b100 ,
#872700000000
1!
1$
b1 %
1'
1*
b1 +
#872710000000
0!
0'
#872720000000
1!
b10 %
1'
b10 +
#872730000000
0!
0'
#872740000000
1!
b11 %
1'
b11 +
#872750000000
0!
0'
#872760000000
1!
b100 %
1'
b100 +
#872770000000
0!
0'
#872780000000
1!
b101 %
1'
b101 +
#872790000000
0!
0'
#872800000000
1!
b110 %
1'
b110 +
#872810000000
0!
0'
#872820000000
1!
b111 %
1'
b111 +
#872830000000
0!
0'
#872840000000
1!
0$
b1000 %
1'
0*
b1000 +
#872850000000
0!
0'
#872860000000
1!
b1001 %
1'
b1001 +
#872870000000
0!
0'
#872880000000
1!
b0 %
1'
b0 +
#872890000000
0!
0'
#872900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#872910000000
0!
0'
#872920000000
1!
b10 %
1'
b10 +
#872930000000
0!
0'
#872940000000
1!
b11 %
1'
b11 +
#872950000000
0!
0'
#872960000000
1!
b100 %
1'
b100 +
#872970000000
0!
0'
#872980000000
1!
b101 %
1'
b101 +
#872990000000
0!
0'
#873000000000
1!
0$
b110 %
1'
0*
b110 +
#873010000000
0!
0'
#873020000000
1!
b111 %
1'
b111 +
#873030000000
0!
0'
#873040000000
1!
b1000 %
1'
b1000 +
#873050000000
0!
0'
#873060000000
1!
b1001 %
1'
b1001 +
#873070000000
0!
0'
#873080000000
1!
b0 %
1'
b0 +
#873090000000
0!
0'
#873100000000
1!
1$
b1 %
1'
1*
b1 +
#873110000000
1"
1(
#873120000000
0!
0"
b100 &
0'
0(
b100 ,
#873130000000
1!
b10 %
1'
b10 +
#873140000000
0!
0'
#873150000000
1!
b11 %
1'
b11 +
#873160000000
0!
0'
#873170000000
1!
b100 %
1'
b100 +
#873180000000
0!
0'
#873190000000
1!
b101 %
1'
b101 +
#873200000000
0!
0'
#873210000000
1!
b110 %
1'
b110 +
#873220000000
0!
0'
#873230000000
1!
b111 %
1'
b111 +
#873240000000
0!
0'
#873250000000
1!
0$
b1000 %
1'
0*
b1000 +
#873260000000
0!
0'
#873270000000
1!
b1001 %
1'
b1001 +
#873280000000
0!
0'
#873290000000
1!
b0 %
1'
b0 +
#873300000000
0!
0'
#873310000000
1!
1$
b1 %
1'
1*
b1 +
#873320000000
0!
0'
#873330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#873340000000
0!
0'
#873350000000
1!
b11 %
1'
b11 +
#873360000000
0!
0'
#873370000000
1!
b100 %
1'
b100 +
#873380000000
0!
0'
#873390000000
1!
b101 %
1'
b101 +
#873400000000
0!
0'
#873410000000
1!
0$
b110 %
1'
0*
b110 +
#873420000000
0!
0'
#873430000000
1!
b111 %
1'
b111 +
#873440000000
0!
0'
#873450000000
1!
b1000 %
1'
b1000 +
#873460000000
0!
0'
#873470000000
1!
b1001 %
1'
b1001 +
#873480000000
0!
0'
#873490000000
1!
b0 %
1'
b0 +
#873500000000
0!
0'
#873510000000
1!
1$
b1 %
1'
1*
b1 +
#873520000000
0!
0'
#873530000000
1!
b10 %
1'
b10 +
#873540000000
1"
1(
#873550000000
0!
0"
b100 &
0'
0(
b100 ,
#873560000000
1!
b11 %
1'
b11 +
#873570000000
0!
0'
#873580000000
1!
b100 %
1'
b100 +
#873590000000
0!
0'
#873600000000
1!
b101 %
1'
b101 +
#873610000000
0!
0'
#873620000000
1!
b110 %
1'
b110 +
#873630000000
0!
0'
#873640000000
1!
b111 %
1'
b111 +
#873650000000
0!
0'
#873660000000
1!
0$
b1000 %
1'
0*
b1000 +
#873670000000
0!
0'
#873680000000
1!
b1001 %
1'
b1001 +
#873690000000
0!
0'
#873700000000
1!
b0 %
1'
b0 +
#873710000000
0!
0'
#873720000000
1!
1$
b1 %
1'
1*
b1 +
#873730000000
0!
0'
#873740000000
1!
b10 %
1'
b10 +
#873750000000
0!
0'
#873760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#873770000000
0!
0'
#873780000000
1!
b100 %
1'
b100 +
#873790000000
0!
0'
#873800000000
1!
b101 %
1'
b101 +
#873810000000
0!
0'
#873820000000
1!
0$
b110 %
1'
0*
b110 +
#873830000000
0!
0'
#873840000000
1!
b111 %
1'
b111 +
#873850000000
0!
0'
#873860000000
1!
b1000 %
1'
b1000 +
#873870000000
0!
0'
#873880000000
1!
b1001 %
1'
b1001 +
#873890000000
0!
0'
#873900000000
1!
b0 %
1'
b0 +
#873910000000
0!
0'
#873920000000
1!
1$
b1 %
1'
1*
b1 +
#873930000000
0!
0'
#873940000000
1!
b10 %
1'
b10 +
#873950000000
0!
0'
#873960000000
1!
b11 %
1'
b11 +
#873970000000
1"
1(
#873980000000
0!
0"
b100 &
0'
0(
b100 ,
#873990000000
1!
b100 %
1'
b100 +
#874000000000
0!
0'
#874010000000
1!
b101 %
1'
b101 +
#874020000000
0!
0'
#874030000000
1!
b110 %
1'
b110 +
#874040000000
0!
0'
#874050000000
1!
b111 %
1'
b111 +
#874060000000
0!
0'
#874070000000
1!
0$
b1000 %
1'
0*
b1000 +
#874080000000
0!
0'
#874090000000
1!
b1001 %
1'
b1001 +
#874100000000
0!
0'
#874110000000
1!
b0 %
1'
b0 +
#874120000000
0!
0'
#874130000000
1!
1$
b1 %
1'
1*
b1 +
#874140000000
0!
0'
#874150000000
1!
b10 %
1'
b10 +
#874160000000
0!
0'
#874170000000
1!
b11 %
1'
b11 +
#874180000000
0!
0'
#874190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#874200000000
0!
0'
#874210000000
1!
b101 %
1'
b101 +
#874220000000
0!
0'
#874230000000
1!
0$
b110 %
1'
0*
b110 +
#874240000000
0!
0'
#874250000000
1!
b111 %
1'
b111 +
#874260000000
0!
0'
#874270000000
1!
b1000 %
1'
b1000 +
#874280000000
0!
0'
#874290000000
1!
b1001 %
1'
b1001 +
#874300000000
0!
0'
#874310000000
1!
b0 %
1'
b0 +
#874320000000
0!
0'
#874330000000
1!
1$
b1 %
1'
1*
b1 +
#874340000000
0!
0'
#874350000000
1!
b10 %
1'
b10 +
#874360000000
0!
0'
#874370000000
1!
b11 %
1'
b11 +
#874380000000
0!
0'
#874390000000
1!
b100 %
1'
b100 +
#874400000000
1"
1(
#874410000000
0!
0"
b100 &
0'
0(
b100 ,
#874420000000
1!
b101 %
1'
b101 +
#874430000000
0!
0'
#874440000000
1!
b110 %
1'
b110 +
#874450000000
0!
0'
#874460000000
1!
b111 %
1'
b111 +
#874470000000
0!
0'
#874480000000
1!
0$
b1000 %
1'
0*
b1000 +
#874490000000
0!
0'
#874500000000
1!
b1001 %
1'
b1001 +
#874510000000
0!
0'
#874520000000
1!
b0 %
1'
b0 +
#874530000000
0!
0'
#874540000000
1!
1$
b1 %
1'
1*
b1 +
#874550000000
0!
0'
#874560000000
1!
b10 %
1'
b10 +
#874570000000
0!
0'
#874580000000
1!
b11 %
1'
b11 +
#874590000000
0!
0'
#874600000000
1!
b100 %
1'
b100 +
#874610000000
0!
0'
#874620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#874630000000
0!
0'
#874640000000
1!
0$
b110 %
1'
0*
b110 +
#874650000000
0!
0'
#874660000000
1!
b111 %
1'
b111 +
#874670000000
0!
0'
#874680000000
1!
b1000 %
1'
b1000 +
#874690000000
0!
0'
#874700000000
1!
b1001 %
1'
b1001 +
#874710000000
0!
0'
#874720000000
1!
b0 %
1'
b0 +
#874730000000
0!
0'
#874740000000
1!
1$
b1 %
1'
1*
b1 +
#874750000000
0!
0'
#874760000000
1!
b10 %
1'
b10 +
#874770000000
0!
0'
#874780000000
1!
b11 %
1'
b11 +
#874790000000
0!
0'
#874800000000
1!
b100 %
1'
b100 +
#874810000000
0!
0'
#874820000000
1!
b101 %
1'
b101 +
#874830000000
1"
1(
#874840000000
0!
0"
b100 &
0'
0(
b100 ,
#874850000000
1!
b110 %
1'
b110 +
#874860000000
0!
0'
#874870000000
1!
b111 %
1'
b111 +
#874880000000
0!
0'
#874890000000
1!
0$
b1000 %
1'
0*
b1000 +
#874900000000
0!
0'
#874910000000
1!
b1001 %
1'
b1001 +
#874920000000
0!
0'
#874930000000
1!
b0 %
1'
b0 +
#874940000000
0!
0'
#874950000000
1!
1$
b1 %
1'
1*
b1 +
#874960000000
0!
0'
#874970000000
1!
b10 %
1'
b10 +
#874980000000
0!
0'
#874990000000
1!
b11 %
1'
b11 +
#875000000000
0!
0'
#875010000000
1!
b100 %
1'
b100 +
#875020000000
0!
0'
#875030000000
1!
b101 %
1'
b101 +
#875040000000
0!
0'
#875050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#875060000000
0!
0'
#875070000000
1!
b111 %
1'
b111 +
#875080000000
0!
0'
#875090000000
1!
b1000 %
1'
b1000 +
#875100000000
0!
0'
#875110000000
1!
b1001 %
1'
b1001 +
#875120000000
0!
0'
#875130000000
1!
b0 %
1'
b0 +
#875140000000
0!
0'
#875150000000
1!
1$
b1 %
1'
1*
b1 +
#875160000000
0!
0'
#875170000000
1!
b10 %
1'
b10 +
#875180000000
0!
0'
#875190000000
1!
b11 %
1'
b11 +
#875200000000
0!
0'
#875210000000
1!
b100 %
1'
b100 +
#875220000000
0!
0'
#875230000000
1!
b101 %
1'
b101 +
#875240000000
0!
0'
#875250000000
1!
0$
b110 %
1'
0*
b110 +
#875260000000
1"
1(
#875270000000
0!
0"
b100 &
0'
0(
b100 ,
#875280000000
1!
1$
b111 %
1'
1*
b111 +
#875290000000
0!
0'
#875300000000
1!
0$
b1000 %
1'
0*
b1000 +
#875310000000
0!
0'
#875320000000
1!
b1001 %
1'
b1001 +
#875330000000
0!
0'
#875340000000
1!
b0 %
1'
b0 +
#875350000000
0!
0'
#875360000000
1!
1$
b1 %
1'
1*
b1 +
#875370000000
0!
0'
#875380000000
1!
b10 %
1'
b10 +
#875390000000
0!
0'
#875400000000
1!
b11 %
1'
b11 +
#875410000000
0!
0'
#875420000000
1!
b100 %
1'
b100 +
#875430000000
0!
0'
#875440000000
1!
b101 %
1'
b101 +
#875450000000
0!
0'
#875460000000
1!
b110 %
1'
b110 +
#875470000000
0!
0'
#875480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#875490000000
0!
0'
#875500000000
1!
b1000 %
1'
b1000 +
#875510000000
0!
0'
#875520000000
1!
b1001 %
1'
b1001 +
#875530000000
0!
0'
#875540000000
1!
b0 %
1'
b0 +
#875550000000
0!
0'
#875560000000
1!
1$
b1 %
1'
1*
b1 +
#875570000000
0!
0'
#875580000000
1!
b10 %
1'
b10 +
#875590000000
0!
0'
#875600000000
1!
b11 %
1'
b11 +
#875610000000
0!
0'
#875620000000
1!
b100 %
1'
b100 +
#875630000000
0!
0'
#875640000000
1!
b101 %
1'
b101 +
#875650000000
0!
0'
#875660000000
1!
0$
b110 %
1'
0*
b110 +
#875670000000
0!
0'
#875680000000
1!
b111 %
1'
b111 +
#875690000000
1"
1(
#875700000000
0!
0"
b100 &
0'
0(
b100 ,
#875710000000
1!
b1000 %
1'
b1000 +
#875720000000
0!
0'
#875730000000
1!
b1001 %
1'
b1001 +
#875740000000
0!
0'
#875750000000
1!
b0 %
1'
b0 +
#875760000000
0!
0'
#875770000000
1!
1$
b1 %
1'
1*
b1 +
#875780000000
0!
0'
#875790000000
1!
b10 %
1'
b10 +
#875800000000
0!
0'
#875810000000
1!
b11 %
1'
b11 +
#875820000000
0!
0'
#875830000000
1!
b100 %
1'
b100 +
#875840000000
0!
0'
#875850000000
1!
b101 %
1'
b101 +
#875860000000
0!
0'
#875870000000
1!
b110 %
1'
b110 +
#875880000000
0!
0'
#875890000000
1!
b111 %
1'
b111 +
#875900000000
0!
0'
#875910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#875920000000
0!
0'
#875930000000
1!
b1001 %
1'
b1001 +
#875940000000
0!
0'
#875950000000
1!
b0 %
1'
b0 +
#875960000000
0!
0'
#875970000000
1!
1$
b1 %
1'
1*
b1 +
#875980000000
0!
0'
#875990000000
1!
b10 %
1'
b10 +
#876000000000
0!
0'
#876010000000
1!
b11 %
1'
b11 +
#876020000000
0!
0'
#876030000000
1!
b100 %
1'
b100 +
#876040000000
0!
0'
#876050000000
1!
b101 %
1'
b101 +
#876060000000
0!
0'
#876070000000
1!
0$
b110 %
1'
0*
b110 +
#876080000000
0!
0'
#876090000000
1!
b111 %
1'
b111 +
#876100000000
0!
0'
#876110000000
1!
b1000 %
1'
b1000 +
#876120000000
1"
1(
#876130000000
0!
0"
b100 &
0'
0(
b100 ,
#876140000000
1!
b1001 %
1'
b1001 +
#876150000000
0!
0'
#876160000000
1!
b0 %
1'
b0 +
#876170000000
0!
0'
#876180000000
1!
1$
b1 %
1'
1*
b1 +
#876190000000
0!
0'
#876200000000
1!
b10 %
1'
b10 +
#876210000000
0!
0'
#876220000000
1!
b11 %
1'
b11 +
#876230000000
0!
0'
#876240000000
1!
b100 %
1'
b100 +
#876250000000
0!
0'
#876260000000
1!
b101 %
1'
b101 +
#876270000000
0!
0'
#876280000000
1!
b110 %
1'
b110 +
#876290000000
0!
0'
#876300000000
1!
b111 %
1'
b111 +
#876310000000
0!
0'
#876320000000
1!
0$
b1000 %
1'
0*
b1000 +
#876330000000
0!
0'
#876340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#876350000000
0!
0'
#876360000000
1!
b0 %
1'
b0 +
#876370000000
0!
0'
#876380000000
1!
1$
b1 %
1'
1*
b1 +
#876390000000
0!
0'
#876400000000
1!
b10 %
1'
b10 +
#876410000000
0!
0'
#876420000000
1!
b11 %
1'
b11 +
#876430000000
0!
0'
#876440000000
1!
b100 %
1'
b100 +
#876450000000
0!
0'
#876460000000
1!
b101 %
1'
b101 +
#876470000000
0!
0'
#876480000000
1!
0$
b110 %
1'
0*
b110 +
#876490000000
0!
0'
#876500000000
1!
b111 %
1'
b111 +
#876510000000
0!
0'
#876520000000
1!
b1000 %
1'
b1000 +
#876530000000
0!
0'
#876540000000
1!
b1001 %
1'
b1001 +
#876550000000
1"
1(
#876560000000
0!
0"
b100 &
0'
0(
b100 ,
#876570000000
1!
b0 %
1'
b0 +
#876580000000
0!
0'
#876590000000
1!
1$
b1 %
1'
1*
b1 +
#876600000000
0!
0'
#876610000000
1!
b10 %
1'
b10 +
#876620000000
0!
0'
#876630000000
1!
b11 %
1'
b11 +
#876640000000
0!
0'
#876650000000
1!
b100 %
1'
b100 +
#876660000000
0!
0'
#876670000000
1!
b101 %
1'
b101 +
#876680000000
0!
0'
#876690000000
1!
b110 %
1'
b110 +
#876700000000
0!
0'
#876710000000
1!
b111 %
1'
b111 +
#876720000000
0!
0'
#876730000000
1!
0$
b1000 %
1'
0*
b1000 +
#876740000000
0!
0'
#876750000000
1!
b1001 %
1'
b1001 +
#876760000000
0!
0'
#876770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#876780000000
0!
0'
#876790000000
1!
1$
b1 %
1'
1*
b1 +
#876800000000
0!
0'
#876810000000
1!
b10 %
1'
b10 +
#876820000000
0!
0'
#876830000000
1!
b11 %
1'
b11 +
#876840000000
0!
0'
#876850000000
1!
b100 %
1'
b100 +
#876860000000
0!
0'
#876870000000
1!
b101 %
1'
b101 +
#876880000000
0!
0'
#876890000000
1!
0$
b110 %
1'
0*
b110 +
#876900000000
0!
0'
#876910000000
1!
b111 %
1'
b111 +
#876920000000
0!
0'
#876930000000
1!
b1000 %
1'
b1000 +
#876940000000
0!
0'
#876950000000
1!
b1001 %
1'
b1001 +
#876960000000
0!
0'
#876970000000
1!
b0 %
1'
b0 +
#876980000000
1"
1(
#876990000000
0!
0"
b100 &
0'
0(
b100 ,
#877000000000
1!
1$
b1 %
1'
1*
b1 +
#877010000000
0!
0'
#877020000000
1!
b10 %
1'
b10 +
#877030000000
0!
0'
#877040000000
1!
b11 %
1'
b11 +
#877050000000
0!
0'
#877060000000
1!
b100 %
1'
b100 +
#877070000000
0!
0'
#877080000000
1!
b101 %
1'
b101 +
#877090000000
0!
0'
#877100000000
1!
b110 %
1'
b110 +
#877110000000
0!
0'
#877120000000
1!
b111 %
1'
b111 +
#877130000000
0!
0'
#877140000000
1!
0$
b1000 %
1'
0*
b1000 +
#877150000000
0!
0'
#877160000000
1!
b1001 %
1'
b1001 +
#877170000000
0!
0'
#877180000000
1!
b0 %
1'
b0 +
#877190000000
0!
0'
#877200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#877210000000
0!
0'
#877220000000
1!
b10 %
1'
b10 +
#877230000000
0!
0'
#877240000000
1!
b11 %
1'
b11 +
#877250000000
0!
0'
#877260000000
1!
b100 %
1'
b100 +
#877270000000
0!
0'
#877280000000
1!
b101 %
1'
b101 +
#877290000000
0!
0'
#877300000000
1!
0$
b110 %
1'
0*
b110 +
#877310000000
0!
0'
#877320000000
1!
b111 %
1'
b111 +
#877330000000
0!
0'
#877340000000
1!
b1000 %
1'
b1000 +
#877350000000
0!
0'
#877360000000
1!
b1001 %
1'
b1001 +
#877370000000
0!
0'
#877380000000
1!
b0 %
1'
b0 +
#877390000000
0!
0'
#877400000000
1!
1$
b1 %
1'
1*
b1 +
#877410000000
1"
1(
#877420000000
0!
0"
b100 &
0'
0(
b100 ,
#877430000000
1!
b10 %
1'
b10 +
#877440000000
0!
0'
#877450000000
1!
b11 %
1'
b11 +
#877460000000
0!
0'
#877470000000
1!
b100 %
1'
b100 +
#877480000000
0!
0'
#877490000000
1!
b101 %
1'
b101 +
#877500000000
0!
0'
#877510000000
1!
b110 %
1'
b110 +
#877520000000
0!
0'
#877530000000
1!
b111 %
1'
b111 +
#877540000000
0!
0'
#877550000000
1!
0$
b1000 %
1'
0*
b1000 +
#877560000000
0!
0'
#877570000000
1!
b1001 %
1'
b1001 +
#877580000000
0!
0'
#877590000000
1!
b0 %
1'
b0 +
#877600000000
0!
0'
#877610000000
1!
1$
b1 %
1'
1*
b1 +
#877620000000
0!
0'
#877630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#877640000000
0!
0'
#877650000000
1!
b11 %
1'
b11 +
#877660000000
0!
0'
#877670000000
1!
b100 %
1'
b100 +
#877680000000
0!
0'
#877690000000
1!
b101 %
1'
b101 +
#877700000000
0!
0'
#877710000000
1!
0$
b110 %
1'
0*
b110 +
#877720000000
0!
0'
#877730000000
1!
b111 %
1'
b111 +
#877740000000
0!
0'
#877750000000
1!
b1000 %
1'
b1000 +
#877760000000
0!
0'
#877770000000
1!
b1001 %
1'
b1001 +
#877780000000
0!
0'
#877790000000
1!
b0 %
1'
b0 +
#877800000000
0!
0'
#877810000000
1!
1$
b1 %
1'
1*
b1 +
#877820000000
0!
0'
#877830000000
1!
b10 %
1'
b10 +
#877840000000
1"
1(
#877850000000
0!
0"
b100 &
0'
0(
b100 ,
#877860000000
1!
b11 %
1'
b11 +
#877870000000
0!
0'
#877880000000
1!
b100 %
1'
b100 +
#877890000000
0!
0'
#877900000000
1!
b101 %
1'
b101 +
#877910000000
0!
0'
#877920000000
1!
b110 %
1'
b110 +
#877930000000
0!
0'
#877940000000
1!
b111 %
1'
b111 +
#877950000000
0!
0'
#877960000000
1!
0$
b1000 %
1'
0*
b1000 +
#877970000000
0!
0'
#877980000000
1!
b1001 %
1'
b1001 +
#877990000000
0!
0'
#878000000000
1!
b0 %
1'
b0 +
#878010000000
0!
0'
#878020000000
1!
1$
b1 %
1'
1*
b1 +
#878030000000
0!
0'
#878040000000
1!
b10 %
1'
b10 +
#878050000000
0!
0'
#878060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#878070000000
0!
0'
#878080000000
1!
b100 %
1'
b100 +
#878090000000
0!
0'
#878100000000
1!
b101 %
1'
b101 +
#878110000000
0!
0'
#878120000000
1!
0$
b110 %
1'
0*
b110 +
#878130000000
0!
0'
#878140000000
1!
b111 %
1'
b111 +
#878150000000
0!
0'
#878160000000
1!
b1000 %
1'
b1000 +
#878170000000
0!
0'
#878180000000
1!
b1001 %
1'
b1001 +
#878190000000
0!
0'
#878200000000
1!
b0 %
1'
b0 +
#878210000000
0!
0'
#878220000000
1!
1$
b1 %
1'
1*
b1 +
#878230000000
0!
0'
#878240000000
1!
b10 %
1'
b10 +
#878250000000
0!
0'
#878260000000
1!
b11 %
1'
b11 +
#878270000000
1"
1(
#878280000000
0!
0"
b100 &
0'
0(
b100 ,
#878290000000
1!
b100 %
1'
b100 +
#878300000000
0!
0'
#878310000000
1!
b101 %
1'
b101 +
#878320000000
0!
0'
#878330000000
1!
b110 %
1'
b110 +
#878340000000
0!
0'
#878350000000
1!
b111 %
1'
b111 +
#878360000000
0!
0'
#878370000000
1!
0$
b1000 %
1'
0*
b1000 +
#878380000000
0!
0'
#878390000000
1!
b1001 %
1'
b1001 +
#878400000000
0!
0'
#878410000000
1!
b0 %
1'
b0 +
#878420000000
0!
0'
#878430000000
1!
1$
b1 %
1'
1*
b1 +
#878440000000
0!
0'
#878450000000
1!
b10 %
1'
b10 +
#878460000000
0!
0'
#878470000000
1!
b11 %
1'
b11 +
#878480000000
0!
0'
#878490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#878500000000
0!
0'
#878510000000
1!
b101 %
1'
b101 +
#878520000000
0!
0'
#878530000000
1!
0$
b110 %
1'
0*
b110 +
#878540000000
0!
0'
#878550000000
1!
b111 %
1'
b111 +
#878560000000
0!
0'
#878570000000
1!
b1000 %
1'
b1000 +
#878580000000
0!
0'
#878590000000
1!
b1001 %
1'
b1001 +
#878600000000
0!
0'
#878610000000
1!
b0 %
1'
b0 +
#878620000000
0!
0'
#878630000000
1!
1$
b1 %
1'
1*
b1 +
#878640000000
0!
0'
#878650000000
1!
b10 %
1'
b10 +
#878660000000
0!
0'
#878670000000
1!
b11 %
1'
b11 +
#878680000000
0!
0'
#878690000000
1!
b100 %
1'
b100 +
#878700000000
1"
1(
#878710000000
0!
0"
b100 &
0'
0(
b100 ,
#878720000000
1!
b101 %
1'
b101 +
#878730000000
0!
0'
#878740000000
1!
b110 %
1'
b110 +
#878750000000
0!
0'
#878760000000
1!
b111 %
1'
b111 +
#878770000000
0!
0'
#878780000000
1!
0$
b1000 %
1'
0*
b1000 +
#878790000000
0!
0'
#878800000000
1!
b1001 %
1'
b1001 +
#878810000000
0!
0'
#878820000000
1!
b0 %
1'
b0 +
#878830000000
0!
0'
#878840000000
1!
1$
b1 %
1'
1*
b1 +
#878850000000
0!
0'
#878860000000
1!
b10 %
1'
b10 +
#878870000000
0!
0'
#878880000000
1!
b11 %
1'
b11 +
#878890000000
0!
0'
#878900000000
1!
b100 %
1'
b100 +
#878910000000
0!
0'
#878920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#878930000000
0!
0'
#878940000000
1!
0$
b110 %
1'
0*
b110 +
#878950000000
0!
0'
#878960000000
1!
b111 %
1'
b111 +
#878970000000
0!
0'
#878980000000
1!
b1000 %
1'
b1000 +
#878990000000
0!
0'
#879000000000
1!
b1001 %
1'
b1001 +
#879010000000
0!
0'
#879020000000
1!
b0 %
1'
b0 +
#879030000000
0!
0'
#879040000000
1!
1$
b1 %
1'
1*
b1 +
#879050000000
0!
0'
#879060000000
1!
b10 %
1'
b10 +
#879070000000
0!
0'
#879080000000
1!
b11 %
1'
b11 +
#879090000000
0!
0'
#879100000000
1!
b100 %
1'
b100 +
#879110000000
0!
0'
#879120000000
1!
b101 %
1'
b101 +
#879130000000
1"
1(
#879140000000
0!
0"
b100 &
0'
0(
b100 ,
#879150000000
1!
b110 %
1'
b110 +
#879160000000
0!
0'
#879170000000
1!
b111 %
1'
b111 +
#879180000000
0!
0'
#879190000000
1!
0$
b1000 %
1'
0*
b1000 +
#879200000000
0!
0'
#879210000000
1!
b1001 %
1'
b1001 +
#879220000000
0!
0'
#879230000000
1!
b0 %
1'
b0 +
#879240000000
0!
0'
#879250000000
1!
1$
b1 %
1'
1*
b1 +
#879260000000
0!
0'
#879270000000
1!
b10 %
1'
b10 +
#879280000000
0!
0'
#879290000000
1!
b11 %
1'
b11 +
#879300000000
0!
0'
#879310000000
1!
b100 %
1'
b100 +
#879320000000
0!
0'
#879330000000
1!
b101 %
1'
b101 +
#879340000000
0!
0'
#879350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#879360000000
0!
0'
#879370000000
1!
b111 %
1'
b111 +
#879380000000
0!
0'
#879390000000
1!
b1000 %
1'
b1000 +
#879400000000
0!
0'
#879410000000
1!
b1001 %
1'
b1001 +
#879420000000
0!
0'
#879430000000
1!
b0 %
1'
b0 +
#879440000000
0!
0'
#879450000000
1!
1$
b1 %
1'
1*
b1 +
#879460000000
0!
0'
#879470000000
1!
b10 %
1'
b10 +
#879480000000
0!
0'
#879490000000
1!
b11 %
1'
b11 +
#879500000000
0!
0'
#879510000000
1!
b100 %
1'
b100 +
#879520000000
0!
0'
#879530000000
1!
b101 %
1'
b101 +
#879540000000
0!
0'
#879550000000
1!
0$
b110 %
1'
0*
b110 +
#879560000000
1"
1(
#879570000000
0!
0"
b100 &
0'
0(
b100 ,
#879580000000
1!
1$
b111 %
1'
1*
b111 +
#879590000000
0!
0'
#879600000000
1!
0$
b1000 %
1'
0*
b1000 +
#879610000000
0!
0'
#879620000000
1!
b1001 %
1'
b1001 +
#879630000000
0!
0'
#879640000000
1!
b0 %
1'
b0 +
#879650000000
0!
0'
#879660000000
1!
1$
b1 %
1'
1*
b1 +
#879670000000
0!
0'
#879680000000
1!
b10 %
1'
b10 +
#879690000000
0!
0'
#879700000000
1!
b11 %
1'
b11 +
#879710000000
0!
0'
#879720000000
1!
b100 %
1'
b100 +
#879730000000
0!
0'
#879740000000
1!
b101 %
1'
b101 +
#879750000000
0!
0'
#879760000000
1!
b110 %
1'
b110 +
#879770000000
0!
0'
#879780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#879790000000
0!
0'
#879800000000
1!
b1000 %
1'
b1000 +
#879810000000
0!
0'
#879820000000
1!
b1001 %
1'
b1001 +
#879830000000
0!
0'
#879840000000
1!
b0 %
1'
b0 +
#879850000000
0!
0'
#879860000000
1!
1$
b1 %
1'
1*
b1 +
#879870000000
0!
0'
#879880000000
1!
b10 %
1'
b10 +
#879890000000
0!
0'
#879900000000
1!
b11 %
1'
b11 +
#879910000000
0!
0'
#879920000000
1!
b100 %
1'
b100 +
#879930000000
0!
0'
#879940000000
1!
b101 %
1'
b101 +
#879950000000
0!
0'
#879960000000
1!
0$
b110 %
1'
0*
b110 +
#879970000000
0!
0'
#879980000000
1!
b111 %
1'
b111 +
#879990000000
1"
1(
#880000000000
0!
0"
b100 &
0'
0(
b100 ,
#880010000000
1!
b1000 %
1'
b1000 +
#880020000000
0!
0'
#880030000000
1!
b1001 %
1'
b1001 +
#880040000000
0!
0'
#880050000000
1!
b0 %
1'
b0 +
#880060000000
0!
0'
#880070000000
1!
1$
b1 %
1'
1*
b1 +
#880080000000
0!
0'
#880090000000
1!
b10 %
1'
b10 +
#880100000000
0!
0'
#880110000000
1!
b11 %
1'
b11 +
#880120000000
0!
0'
#880130000000
1!
b100 %
1'
b100 +
#880140000000
0!
0'
#880150000000
1!
b101 %
1'
b101 +
#880160000000
0!
0'
#880170000000
1!
b110 %
1'
b110 +
#880180000000
0!
0'
#880190000000
1!
b111 %
1'
b111 +
#880200000000
0!
0'
#880210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#880220000000
0!
0'
#880230000000
1!
b1001 %
1'
b1001 +
#880240000000
0!
0'
#880250000000
1!
b0 %
1'
b0 +
#880260000000
0!
0'
#880270000000
1!
1$
b1 %
1'
1*
b1 +
#880280000000
0!
0'
#880290000000
1!
b10 %
1'
b10 +
#880300000000
0!
0'
#880310000000
1!
b11 %
1'
b11 +
#880320000000
0!
0'
#880330000000
1!
b100 %
1'
b100 +
#880340000000
0!
0'
#880350000000
1!
b101 %
1'
b101 +
#880360000000
0!
0'
#880370000000
1!
0$
b110 %
1'
0*
b110 +
#880380000000
0!
0'
#880390000000
1!
b111 %
1'
b111 +
#880400000000
0!
0'
#880410000000
1!
b1000 %
1'
b1000 +
#880420000000
1"
1(
#880430000000
0!
0"
b100 &
0'
0(
b100 ,
#880440000000
1!
b1001 %
1'
b1001 +
#880450000000
0!
0'
#880460000000
1!
b0 %
1'
b0 +
#880470000000
0!
0'
#880480000000
1!
1$
b1 %
1'
1*
b1 +
#880490000000
0!
0'
#880500000000
1!
b10 %
1'
b10 +
#880510000000
0!
0'
#880520000000
1!
b11 %
1'
b11 +
#880530000000
0!
0'
#880540000000
1!
b100 %
1'
b100 +
#880550000000
0!
0'
#880560000000
1!
b101 %
1'
b101 +
#880570000000
0!
0'
#880580000000
1!
b110 %
1'
b110 +
#880590000000
0!
0'
#880600000000
1!
b111 %
1'
b111 +
#880610000000
0!
0'
#880620000000
1!
0$
b1000 %
1'
0*
b1000 +
#880630000000
0!
0'
#880640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#880650000000
0!
0'
#880660000000
1!
b0 %
1'
b0 +
#880670000000
0!
0'
#880680000000
1!
1$
b1 %
1'
1*
b1 +
#880690000000
0!
0'
#880700000000
1!
b10 %
1'
b10 +
#880710000000
0!
0'
#880720000000
1!
b11 %
1'
b11 +
#880730000000
0!
0'
#880740000000
1!
b100 %
1'
b100 +
#880750000000
0!
0'
#880760000000
1!
b101 %
1'
b101 +
#880770000000
0!
0'
#880780000000
1!
0$
b110 %
1'
0*
b110 +
#880790000000
0!
0'
#880800000000
1!
b111 %
1'
b111 +
#880810000000
0!
0'
#880820000000
1!
b1000 %
1'
b1000 +
#880830000000
0!
0'
#880840000000
1!
b1001 %
1'
b1001 +
#880850000000
1"
1(
#880860000000
0!
0"
b100 &
0'
0(
b100 ,
#880870000000
1!
b0 %
1'
b0 +
#880880000000
0!
0'
#880890000000
1!
1$
b1 %
1'
1*
b1 +
#880900000000
0!
0'
#880910000000
1!
b10 %
1'
b10 +
#880920000000
0!
0'
#880930000000
1!
b11 %
1'
b11 +
#880940000000
0!
0'
#880950000000
1!
b100 %
1'
b100 +
#880960000000
0!
0'
#880970000000
1!
b101 %
1'
b101 +
#880980000000
0!
0'
#880990000000
1!
b110 %
1'
b110 +
#881000000000
0!
0'
#881010000000
1!
b111 %
1'
b111 +
#881020000000
0!
0'
#881030000000
1!
0$
b1000 %
1'
0*
b1000 +
#881040000000
0!
0'
#881050000000
1!
b1001 %
1'
b1001 +
#881060000000
0!
0'
#881070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#881080000000
0!
0'
#881090000000
1!
1$
b1 %
1'
1*
b1 +
#881100000000
0!
0'
#881110000000
1!
b10 %
1'
b10 +
#881120000000
0!
0'
#881130000000
1!
b11 %
1'
b11 +
#881140000000
0!
0'
#881150000000
1!
b100 %
1'
b100 +
#881160000000
0!
0'
#881170000000
1!
b101 %
1'
b101 +
#881180000000
0!
0'
#881190000000
1!
0$
b110 %
1'
0*
b110 +
#881200000000
0!
0'
#881210000000
1!
b111 %
1'
b111 +
#881220000000
0!
0'
#881230000000
1!
b1000 %
1'
b1000 +
#881240000000
0!
0'
#881250000000
1!
b1001 %
1'
b1001 +
#881260000000
0!
0'
#881270000000
1!
b0 %
1'
b0 +
#881280000000
1"
1(
#881290000000
0!
0"
b100 &
0'
0(
b100 ,
#881300000000
1!
1$
b1 %
1'
1*
b1 +
#881310000000
0!
0'
#881320000000
1!
b10 %
1'
b10 +
#881330000000
0!
0'
#881340000000
1!
b11 %
1'
b11 +
#881350000000
0!
0'
#881360000000
1!
b100 %
1'
b100 +
#881370000000
0!
0'
#881380000000
1!
b101 %
1'
b101 +
#881390000000
0!
0'
#881400000000
1!
b110 %
1'
b110 +
#881410000000
0!
0'
#881420000000
1!
b111 %
1'
b111 +
#881430000000
0!
0'
#881440000000
1!
0$
b1000 %
1'
0*
b1000 +
#881450000000
0!
0'
#881460000000
1!
b1001 %
1'
b1001 +
#881470000000
0!
0'
#881480000000
1!
b0 %
1'
b0 +
#881490000000
0!
0'
#881500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#881510000000
0!
0'
#881520000000
1!
b10 %
1'
b10 +
#881530000000
0!
0'
#881540000000
1!
b11 %
1'
b11 +
#881550000000
0!
0'
#881560000000
1!
b100 %
1'
b100 +
#881570000000
0!
0'
#881580000000
1!
b101 %
1'
b101 +
#881590000000
0!
0'
#881600000000
1!
0$
b110 %
1'
0*
b110 +
#881610000000
0!
0'
#881620000000
1!
b111 %
1'
b111 +
#881630000000
0!
0'
#881640000000
1!
b1000 %
1'
b1000 +
#881650000000
0!
0'
#881660000000
1!
b1001 %
1'
b1001 +
#881670000000
0!
0'
#881680000000
1!
b0 %
1'
b0 +
#881690000000
0!
0'
#881700000000
1!
1$
b1 %
1'
1*
b1 +
#881710000000
1"
1(
#881720000000
0!
0"
b100 &
0'
0(
b100 ,
#881730000000
1!
b10 %
1'
b10 +
#881740000000
0!
0'
#881750000000
1!
b11 %
1'
b11 +
#881760000000
0!
0'
#881770000000
1!
b100 %
1'
b100 +
#881780000000
0!
0'
#881790000000
1!
b101 %
1'
b101 +
#881800000000
0!
0'
#881810000000
1!
b110 %
1'
b110 +
#881820000000
0!
0'
#881830000000
1!
b111 %
1'
b111 +
#881840000000
0!
0'
#881850000000
1!
0$
b1000 %
1'
0*
b1000 +
#881860000000
0!
0'
#881870000000
1!
b1001 %
1'
b1001 +
#881880000000
0!
0'
#881890000000
1!
b0 %
1'
b0 +
#881900000000
0!
0'
#881910000000
1!
1$
b1 %
1'
1*
b1 +
#881920000000
0!
0'
#881930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#881940000000
0!
0'
#881950000000
1!
b11 %
1'
b11 +
#881960000000
0!
0'
#881970000000
1!
b100 %
1'
b100 +
#881980000000
0!
0'
#881990000000
1!
b101 %
1'
b101 +
#882000000000
0!
0'
#882010000000
1!
0$
b110 %
1'
0*
b110 +
#882020000000
0!
0'
#882030000000
1!
b111 %
1'
b111 +
#882040000000
0!
0'
#882050000000
1!
b1000 %
1'
b1000 +
#882060000000
0!
0'
#882070000000
1!
b1001 %
1'
b1001 +
#882080000000
0!
0'
#882090000000
1!
b0 %
1'
b0 +
#882100000000
0!
0'
#882110000000
1!
1$
b1 %
1'
1*
b1 +
#882120000000
0!
0'
#882130000000
1!
b10 %
1'
b10 +
#882140000000
1"
1(
#882150000000
0!
0"
b100 &
0'
0(
b100 ,
#882160000000
1!
b11 %
1'
b11 +
#882170000000
0!
0'
#882180000000
1!
b100 %
1'
b100 +
#882190000000
0!
0'
#882200000000
1!
b101 %
1'
b101 +
#882210000000
0!
0'
#882220000000
1!
b110 %
1'
b110 +
#882230000000
0!
0'
#882240000000
1!
b111 %
1'
b111 +
#882250000000
0!
0'
#882260000000
1!
0$
b1000 %
1'
0*
b1000 +
#882270000000
0!
0'
#882280000000
1!
b1001 %
1'
b1001 +
#882290000000
0!
0'
#882300000000
1!
b0 %
1'
b0 +
#882310000000
0!
0'
#882320000000
1!
1$
b1 %
1'
1*
b1 +
#882330000000
0!
0'
#882340000000
1!
b10 %
1'
b10 +
#882350000000
0!
0'
#882360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#882370000000
0!
0'
#882380000000
1!
b100 %
1'
b100 +
#882390000000
0!
0'
#882400000000
1!
b101 %
1'
b101 +
#882410000000
0!
0'
#882420000000
1!
0$
b110 %
1'
0*
b110 +
#882430000000
0!
0'
#882440000000
1!
b111 %
1'
b111 +
#882450000000
0!
0'
#882460000000
1!
b1000 %
1'
b1000 +
#882470000000
0!
0'
#882480000000
1!
b1001 %
1'
b1001 +
#882490000000
0!
0'
#882500000000
1!
b0 %
1'
b0 +
#882510000000
0!
0'
#882520000000
1!
1$
b1 %
1'
1*
b1 +
#882530000000
0!
0'
#882540000000
1!
b10 %
1'
b10 +
#882550000000
0!
0'
#882560000000
1!
b11 %
1'
b11 +
#882570000000
1"
1(
#882580000000
0!
0"
b100 &
0'
0(
b100 ,
#882590000000
1!
b100 %
1'
b100 +
#882600000000
0!
0'
#882610000000
1!
b101 %
1'
b101 +
#882620000000
0!
0'
#882630000000
1!
b110 %
1'
b110 +
#882640000000
0!
0'
#882650000000
1!
b111 %
1'
b111 +
#882660000000
0!
0'
#882670000000
1!
0$
b1000 %
1'
0*
b1000 +
#882680000000
0!
0'
#882690000000
1!
b1001 %
1'
b1001 +
#882700000000
0!
0'
#882710000000
1!
b0 %
1'
b0 +
#882720000000
0!
0'
#882730000000
1!
1$
b1 %
1'
1*
b1 +
#882740000000
0!
0'
#882750000000
1!
b10 %
1'
b10 +
#882760000000
0!
0'
#882770000000
1!
b11 %
1'
b11 +
#882780000000
0!
0'
#882790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#882800000000
0!
0'
#882810000000
1!
b101 %
1'
b101 +
#882820000000
0!
0'
#882830000000
1!
0$
b110 %
1'
0*
b110 +
#882840000000
0!
0'
#882850000000
1!
b111 %
1'
b111 +
#882860000000
0!
0'
#882870000000
1!
b1000 %
1'
b1000 +
#882880000000
0!
0'
#882890000000
1!
b1001 %
1'
b1001 +
#882900000000
0!
0'
#882910000000
1!
b0 %
1'
b0 +
#882920000000
0!
0'
#882930000000
1!
1$
b1 %
1'
1*
b1 +
#882940000000
0!
0'
#882950000000
1!
b10 %
1'
b10 +
#882960000000
0!
0'
#882970000000
1!
b11 %
1'
b11 +
#882980000000
0!
0'
#882990000000
1!
b100 %
1'
b100 +
#883000000000
1"
1(
#883010000000
0!
0"
b100 &
0'
0(
b100 ,
#883020000000
1!
b101 %
1'
b101 +
#883030000000
0!
0'
#883040000000
1!
b110 %
1'
b110 +
#883050000000
0!
0'
#883060000000
1!
b111 %
1'
b111 +
#883070000000
0!
0'
#883080000000
1!
0$
b1000 %
1'
0*
b1000 +
#883090000000
0!
0'
#883100000000
1!
b1001 %
1'
b1001 +
#883110000000
0!
0'
#883120000000
1!
b0 %
1'
b0 +
#883130000000
0!
0'
#883140000000
1!
1$
b1 %
1'
1*
b1 +
#883150000000
0!
0'
#883160000000
1!
b10 %
1'
b10 +
#883170000000
0!
0'
#883180000000
1!
b11 %
1'
b11 +
#883190000000
0!
0'
#883200000000
1!
b100 %
1'
b100 +
#883210000000
0!
0'
#883220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#883230000000
0!
0'
#883240000000
1!
0$
b110 %
1'
0*
b110 +
#883250000000
0!
0'
#883260000000
1!
b111 %
1'
b111 +
#883270000000
0!
0'
#883280000000
1!
b1000 %
1'
b1000 +
#883290000000
0!
0'
#883300000000
1!
b1001 %
1'
b1001 +
#883310000000
0!
0'
#883320000000
1!
b0 %
1'
b0 +
#883330000000
0!
0'
#883340000000
1!
1$
b1 %
1'
1*
b1 +
#883350000000
0!
0'
#883360000000
1!
b10 %
1'
b10 +
#883370000000
0!
0'
#883380000000
1!
b11 %
1'
b11 +
#883390000000
0!
0'
#883400000000
1!
b100 %
1'
b100 +
#883410000000
0!
0'
#883420000000
1!
b101 %
1'
b101 +
#883430000000
1"
1(
#883440000000
0!
0"
b100 &
0'
0(
b100 ,
#883450000000
1!
b110 %
1'
b110 +
#883460000000
0!
0'
#883470000000
1!
b111 %
1'
b111 +
#883480000000
0!
0'
#883490000000
1!
0$
b1000 %
1'
0*
b1000 +
#883500000000
0!
0'
#883510000000
1!
b1001 %
1'
b1001 +
#883520000000
0!
0'
#883530000000
1!
b0 %
1'
b0 +
#883540000000
0!
0'
#883550000000
1!
1$
b1 %
1'
1*
b1 +
#883560000000
0!
0'
#883570000000
1!
b10 %
1'
b10 +
#883580000000
0!
0'
#883590000000
1!
b11 %
1'
b11 +
#883600000000
0!
0'
#883610000000
1!
b100 %
1'
b100 +
#883620000000
0!
0'
#883630000000
1!
b101 %
1'
b101 +
#883640000000
0!
0'
#883650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#883660000000
0!
0'
#883670000000
1!
b111 %
1'
b111 +
#883680000000
0!
0'
#883690000000
1!
b1000 %
1'
b1000 +
#883700000000
0!
0'
#883710000000
1!
b1001 %
1'
b1001 +
#883720000000
0!
0'
#883730000000
1!
b0 %
1'
b0 +
#883740000000
0!
0'
#883750000000
1!
1$
b1 %
1'
1*
b1 +
#883760000000
0!
0'
#883770000000
1!
b10 %
1'
b10 +
#883780000000
0!
0'
#883790000000
1!
b11 %
1'
b11 +
#883800000000
0!
0'
#883810000000
1!
b100 %
1'
b100 +
#883820000000
0!
0'
#883830000000
1!
b101 %
1'
b101 +
#883840000000
0!
0'
#883850000000
1!
0$
b110 %
1'
0*
b110 +
#883860000000
1"
1(
#883870000000
0!
0"
b100 &
0'
0(
b100 ,
#883880000000
1!
1$
b111 %
1'
1*
b111 +
#883890000000
0!
0'
#883900000000
1!
0$
b1000 %
1'
0*
b1000 +
#883910000000
0!
0'
#883920000000
1!
b1001 %
1'
b1001 +
#883930000000
0!
0'
#883940000000
1!
b0 %
1'
b0 +
#883950000000
0!
0'
#883960000000
1!
1$
b1 %
1'
1*
b1 +
#883970000000
0!
0'
#883980000000
1!
b10 %
1'
b10 +
#883990000000
0!
0'
#884000000000
1!
b11 %
1'
b11 +
#884010000000
0!
0'
#884020000000
1!
b100 %
1'
b100 +
#884030000000
0!
0'
#884040000000
1!
b101 %
1'
b101 +
#884050000000
0!
0'
#884060000000
1!
b110 %
1'
b110 +
#884070000000
0!
0'
#884080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#884090000000
0!
0'
#884100000000
1!
b1000 %
1'
b1000 +
#884110000000
0!
0'
#884120000000
1!
b1001 %
1'
b1001 +
#884130000000
0!
0'
#884140000000
1!
b0 %
1'
b0 +
#884150000000
0!
0'
#884160000000
1!
1$
b1 %
1'
1*
b1 +
#884170000000
0!
0'
#884180000000
1!
b10 %
1'
b10 +
#884190000000
0!
0'
#884200000000
1!
b11 %
1'
b11 +
#884210000000
0!
0'
#884220000000
1!
b100 %
1'
b100 +
#884230000000
0!
0'
#884240000000
1!
b101 %
1'
b101 +
#884250000000
0!
0'
#884260000000
1!
0$
b110 %
1'
0*
b110 +
#884270000000
0!
0'
#884280000000
1!
b111 %
1'
b111 +
#884290000000
1"
1(
#884300000000
0!
0"
b100 &
0'
0(
b100 ,
#884310000000
1!
b1000 %
1'
b1000 +
#884320000000
0!
0'
#884330000000
1!
b1001 %
1'
b1001 +
#884340000000
0!
0'
#884350000000
1!
b0 %
1'
b0 +
#884360000000
0!
0'
#884370000000
1!
1$
b1 %
1'
1*
b1 +
#884380000000
0!
0'
#884390000000
1!
b10 %
1'
b10 +
#884400000000
0!
0'
#884410000000
1!
b11 %
1'
b11 +
#884420000000
0!
0'
#884430000000
1!
b100 %
1'
b100 +
#884440000000
0!
0'
#884450000000
1!
b101 %
1'
b101 +
#884460000000
0!
0'
#884470000000
1!
b110 %
1'
b110 +
#884480000000
0!
0'
#884490000000
1!
b111 %
1'
b111 +
#884500000000
0!
0'
#884510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#884520000000
0!
0'
#884530000000
1!
b1001 %
1'
b1001 +
#884540000000
0!
0'
#884550000000
1!
b0 %
1'
b0 +
#884560000000
0!
0'
#884570000000
1!
1$
b1 %
1'
1*
b1 +
#884580000000
0!
0'
#884590000000
1!
b10 %
1'
b10 +
#884600000000
0!
0'
#884610000000
1!
b11 %
1'
b11 +
#884620000000
0!
0'
#884630000000
1!
b100 %
1'
b100 +
#884640000000
0!
0'
#884650000000
1!
b101 %
1'
b101 +
#884660000000
0!
0'
#884670000000
1!
0$
b110 %
1'
0*
b110 +
#884680000000
0!
0'
#884690000000
1!
b111 %
1'
b111 +
#884700000000
0!
0'
#884710000000
1!
b1000 %
1'
b1000 +
#884720000000
1"
1(
#884730000000
0!
0"
b100 &
0'
0(
b100 ,
#884740000000
1!
b1001 %
1'
b1001 +
#884750000000
0!
0'
#884760000000
1!
b0 %
1'
b0 +
#884770000000
0!
0'
#884780000000
1!
1$
b1 %
1'
1*
b1 +
#884790000000
0!
0'
#884800000000
1!
b10 %
1'
b10 +
#884810000000
0!
0'
#884820000000
1!
b11 %
1'
b11 +
#884830000000
0!
0'
#884840000000
1!
b100 %
1'
b100 +
#884850000000
0!
0'
#884860000000
1!
b101 %
1'
b101 +
#884870000000
0!
0'
#884880000000
1!
b110 %
1'
b110 +
#884890000000
0!
0'
#884900000000
1!
b111 %
1'
b111 +
#884910000000
0!
0'
#884920000000
1!
0$
b1000 %
1'
0*
b1000 +
#884930000000
0!
0'
#884940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#884950000000
0!
0'
#884960000000
1!
b0 %
1'
b0 +
#884970000000
0!
0'
#884980000000
1!
1$
b1 %
1'
1*
b1 +
#884990000000
0!
0'
#885000000000
1!
b10 %
1'
b10 +
#885010000000
0!
0'
#885020000000
1!
b11 %
1'
b11 +
#885030000000
0!
0'
#885040000000
1!
b100 %
1'
b100 +
#885050000000
0!
0'
#885060000000
1!
b101 %
1'
b101 +
#885070000000
0!
0'
#885080000000
1!
0$
b110 %
1'
0*
b110 +
#885090000000
0!
0'
#885100000000
1!
b111 %
1'
b111 +
#885110000000
0!
0'
#885120000000
1!
b1000 %
1'
b1000 +
#885130000000
0!
0'
#885140000000
1!
b1001 %
1'
b1001 +
#885150000000
1"
1(
#885160000000
0!
0"
b100 &
0'
0(
b100 ,
#885170000000
1!
b0 %
1'
b0 +
#885180000000
0!
0'
#885190000000
1!
1$
b1 %
1'
1*
b1 +
#885200000000
0!
0'
#885210000000
1!
b10 %
1'
b10 +
#885220000000
0!
0'
#885230000000
1!
b11 %
1'
b11 +
#885240000000
0!
0'
#885250000000
1!
b100 %
1'
b100 +
#885260000000
0!
0'
#885270000000
1!
b101 %
1'
b101 +
#885280000000
0!
0'
#885290000000
1!
b110 %
1'
b110 +
#885300000000
0!
0'
#885310000000
1!
b111 %
1'
b111 +
#885320000000
0!
0'
#885330000000
1!
0$
b1000 %
1'
0*
b1000 +
#885340000000
0!
0'
#885350000000
1!
b1001 %
1'
b1001 +
#885360000000
0!
0'
#885370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#885380000000
0!
0'
#885390000000
1!
1$
b1 %
1'
1*
b1 +
#885400000000
0!
0'
#885410000000
1!
b10 %
1'
b10 +
#885420000000
0!
0'
#885430000000
1!
b11 %
1'
b11 +
#885440000000
0!
0'
#885450000000
1!
b100 %
1'
b100 +
#885460000000
0!
0'
#885470000000
1!
b101 %
1'
b101 +
#885480000000
0!
0'
#885490000000
1!
0$
b110 %
1'
0*
b110 +
#885500000000
0!
0'
#885510000000
1!
b111 %
1'
b111 +
#885520000000
0!
0'
#885530000000
1!
b1000 %
1'
b1000 +
#885540000000
0!
0'
#885550000000
1!
b1001 %
1'
b1001 +
#885560000000
0!
0'
#885570000000
1!
b0 %
1'
b0 +
#885580000000
1"
1(
#885590000000
0!
0"
b100 &
0'
0(
b100 ,
#885600000000
1!
1$
b1 %
1'
1*
b1 +
#885610000000
0!
0'
#885620000000
1!
b10 %
1'
b10 +
#885630000000
0!
0'
#885640000000
1!
b11 %
1'
b11 +
#885650000000
0!
0'
#885660000000
1!
b100 %
1'
b100 +
#885670000000
0!
0'
#885680000000
1!
b101 %
1'
b101 +
#885690000000
0!
0'
#885700000000
1!
b110 %
1'
b110 +
#885710000000
0!
0'
#885720000000
1!
b111 %
1'
b111 +
#885730000000
0!
0'
#885740000000
1!
0$
b1000 %
1'
0*
b1000 +
#885750000000
0!
0'
#885760000000
1!
b1001 %
1'
b1001 +
#885770000000
0!
0'
#885780000000
1!
b0 %
1'
b0 +
#885790000000
0!
0'
#885800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#885810000000
0!
0'
#885820000000
1!
b10 %
1'
b10 +
#885830000000
0!
0'
#885840000000
1!
b11 %
1'
b11 +
#885850000000
0!
0'
#885860000000
1!
b100 %
1'
b100 +
#885870000000
0!
0'
#885880000000
1!
b101 %
1'
b101 +
#885890000000
0!
0'
#885900000000
1!
0$
b110 %
1'
0*
b110 +
#885910000000
0!
0'
#885920000000
1!
b111 %
1'
b111 +
#885930000000
0!
0'
#885940000000
1!
b1000 %
1'
b1000 +
#885950000000
0!
0'
#885960000000
1!
b1001 %
1'
b1001 +
#885970000000
0!
0'
#885980000000
1!
b0 %
1'
b0 +
#885990000000
0!
0'
#886000000000
1!
1$
b1 %
1'
1*
b1 +
#886010000000
1"
1(
#886020000000
0!
0"
b100 &
0'
0(
b100 ,
#886030000000
1!
b10 %
1'
b10 +
#886040000000
0!
0'
#886050000000
1!
b11 %
1'
b11 +
#886060000000
0!
0'
#886070000000
1!
b100 %
1'
b100 +
#886080000000
0!
0'
#886090000000
1!
b101 %
1'
b101 +
#886100000000
0!
0'
#886110000000
1!
b110 %
1'
b110 +
#886120000000
0!
0'
#886130000000
1!
b111 %
1'
b111 +
#886140000000
0!
0'
#886150000000
1!
0$
b1000 %
1'
0*
b1000 +
#886160000000
0!
0'
#886170000000
1!
b1001 %
1'
b1001 +
#886180000000
0!
0'
#886190000000
1!
b0 %
1'
b0 +
#886200000000
0!
0'
#886210000000
1!
1$
b1 %
1'
1*
b1 +
#886220000000
0!
0'
#886230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#886240000000
0!
0'
#886250000000
1!
b11 %
1'
b11 +
#886260000000
0!
0'
#886270000000
1!
b100 %
1'
b100 +
#886280000000
0!
0'
#886290000000
1!
b101 %
1'
b101 +
#886300000000
0!
0'
#886310000000
1!
0$
b110 %
1'
0*
b110 +
#886320000000
0!
0'
#886330000000
1!
b111 %
1'
b111 +
#886340000000
0!
0'
#886350000000
1!
b1000 %
1'
b1000 +
#886360000000
0!
0'
#886370000000
1!
b1001 %
1'
b1001 +
#886380000000
0!
0'
#886390000000
1!
b0 %
1'
b0 +
#886400000000
0!
0'
#886410000000
1!
1$
b1 %
1'
1*
b1 +
#886420000000
0!
0'
#886430000000
1!
b10 %
1'
b10 +
#886440000000
1"
1(
#886450000000
0!
0"
b100 &
0'
0(
b100 ,
#886460000000
1!
b11 %
1'
b11 +
#886470000000
0!
0'
#886480000000
1!
b100 %
1'
b100 +
#886490000000
0!
0'
#886500000000
1!
b101 %
1'
b101 +
#886510000000
0!
0'
#886520000000
1!
b110 %
1'
b110 +
#886530000000
0!
0'
#886540000000
1!
b111 %
1'
b111 +
#886550000000
0!
0'
#886560000000
1!
0$
b1000 %
1'
0*
b1000 +
#886570000000
0!
0'
#886580000000
1!
b1001 %
1'
b1001 +
#886590000000
0!
0'
#886600000000
1!
b0 %
1'
b0 +
#886610000000
0!
0'
#886620000000
1!
1$
b1 %
1'
1*
b1 +
#886630000000
0!
0'
#886640000000
1!
b10 %
1'
b10 +
#886650000000
0!
0'
#886660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#886670000000
0!
0'
#886680000000
1!
b100 %
1'
b100 +
#886690000000
0!
0'
#886700000000
1!
b101 %
1'
b101 +
#886710000000
0!
0'
#886720000000
1!
0$
b110 %
1'
0*
b110 +
#886730000000
0!
0'
#886740000000
1!
b111 %
1'
b111 +
#886750000000
0!
0'
#886760000000
1!
b1000 %
1'
b1000 +
#886770000000
0!
0'
#886780000000
1!
b1001 %
1'
b1001 +
#886790000000
0!
0'
#886800000000
1!
b0 %
1'
b0 +
#886810000000
0!
0'
#886820000000
1!
1$
b1 %
1'
1*
b1 +
#886830000000
0!
0'
#886840000000
1!
b10 %
1'
b10 +
#886850000000
0!
0'
#886860000000
1!
b11 %
1'
b11 +
#886870000000
1"
1(
#886880000000
0!
0"
b100 &
0'
0(
b100 ,
#886890000000
1!
b100 %
1'
b100 +
#886900000000
0!
0'
#886910000000
1!
b101 %
1'
b101 +
#886920000000
0!
0'
#886930000000
1!
b110 %
1'
b110 +
#886940000000
0!
0'
#886950000000
1!
b111 %
1'
b111 +
#886960000000
0!
0'
#886970000000
1!
0$
b1000 %
1'
0*
b1000 +
#886980000000
0!
0'
#886990000000
1!
b1001 %
1'
b1001 +
#887000000000
0!
0'
#887010000000
1!
b0 %
1'
b0 +
#887020000000
0!
0'
#887030000000
1!
1$
b1 %
1'
1*
b1 +
#887040000000
0!
0'
#887050000000
1!
b10 %
1'
b10 +
#887060000000
0!
0'
#887070000000
1!
b11 %
1'
b11 +
#887080000000
0!
0'
#887090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#887100000000
0!
0'
#887110000000
1!
b101 %
1'
b101 +
#887120000000
0!
0'
#887130000000
1!
0$
b110 %
1'
0*
b110 +
#887140000000
0!
0'
#887150000000
1!
b111 %
1'
b111 +
#887160000000
0!
0'
#887170000000
1!
b1000 %
1'
b1000 +
#887180000000
0!
0'
#887190000000
1!
b1001 %
1'
b1001 +
#887200000000
0!
0'
#887210000000
1!
b0 %
1'
b0 +
#887220000000
0!
0'
#887230000000
1!
1$
b1 %
1'
1*
b1 +
#887240000000
0!
0'
#887250000000
1!
b10 %
1'
b10 +
#887260000000
0!
0'
#887270000000
1!
b11 %
1'
b11 +
#887280000000
0!
0'
#887290000000
1!
b100 %
1'
b100 +
#887300000000
1"
1(
#887310000000
0!
0"
b100 &
0'
0(
b100 ,
#887320000000
1!
b101 %
1'
b101 +
#887330000000
0!
0'
#887340000000
1!
b110 %
1'
b110 +
#887350000000
0!
0'
#887360000000
1!
b111 %
1'
b111 +
#887370000000
0!
0'
#887380000000
1!
0$
b1000 %
1'
0*
b1000 +
#887390000000
0!
0'
#887400000000
1!
b1001 %
1'
b1001 +
#887410000000
0!
0'
#887420000000
1!
b0 %
1'
b0 +
#887430000000
0!
0'
#887440000000
1!
1$
b1 %
1'
1*
b1 +
#887450000000
0!
0'
#887460000000
1!
b10 %
1'
b10 +
#887470000000
0!
0'
#887480000000
1!
b11 %
1'
b11 +
#887490000000
0!
0'
#887500000000
1!
b100 %
1'
b100 +
#887510000000
0!
0'
#887520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#887530000000
0!
0'
#887540000000
1!
0$
b110 %
1'
0*
b110 +
#887550000000
0!
0'
#887560000000
1!
b111 %
1'
b111 +
#887570000000
0!
0'
#887580000000
1!
b1000 %
1'
b1000 +
#887590000000
0!
0'
#887600000000
1!
b1001 %
1'
b1001 +
#887610000000
0!
0'
#887620000000
1!
b0 %
1'
b0 +
#887630000000
0!
0'
#887640000000
1!
1$
b1 %
1'
1*
b1 +
#887650000000
0!
0'
#887660000000
1!
b10 %
1'
b10 +
#887670000000
0!
0'
#887680000000
1!
b11 %
1'
b11 +
#887690000000
0!
0'
#887700000000
1!
b100 %
1'
b100 +
#887710000000
0!
0'
#887720000000
1!
b101 %
1'
b101 +
#887730000000
1"
1(
#887740000000
0!
0"
b100 &
0'
0(
b100 ,
#887750000000
1!
b110 %
1'
b110 +
#887760000000
0!
0'
#887770000000
1!
b111 %
1'
b111 +
#887780000000
0!
0'
#887790000000
1!
0$
b1000 %
1'
0*
b1000 +
#887800000000
0!
0'
#887810000000
1!
b1001 %
1'
b1001 +
#887820000000
0!
0'
#887830000000
1!
b0 %
1'
b0 +
#887840000000
0!
0'
#887850000000
1!
1$
b1 %
1'
1*
b1 +
#887860000000
0!
0'
#887870000000
1!
b10 %
1'
b10 +
#887880000000
0!
0'
#887890000000
1!
b11 %
1'
b11 +
#887900000000
0!
0'
#887910000000
1!
b100 %
1'
b100 +
#887920000000
0!
0'
#887930000000
1!
b101 %
1'
b101 +
#887940000000
0!
0'
#887950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#887960000000
0!
0'
#887970000000
1!
b111 %
1'
b111 +
#887980000000
0!
0'
#887990000000
1!
b1000 %
1'
b1000 +
#888000000000
0!
0'
#888010000000
1!
b1001 %
1'
b1001 +
#888020000000
0!
0'
#888030000000
1!
b0 %
1'
b0 +
#888040000000
0!
0'
#888050000000
1!
1$
b1 %
1'
1*
b1 +
#888060000000
0!
0'
#888070000000
1!
b10 %
1'
b10 +
#888080000000
0!
0'
#888090000000
1!
b11 %
1'
b11 +
#888100000000
0!
0'
#888110000000
1!
b100 %
1'
b100 +
#888120000000
0!
0'
#888130000000
1!
b101 %
1'
b101 +
#888140000000
0!
0'
#888150000000
1!
0$
b110 %
1'
0*
b110 +
#888160000000
1"
1(
#888170000000
0!
0"
b100 &
0'
0(
b100 ,
#888180000000
1!
1$
b111 %
1'
1*
b111 +
#888190000000
0!
0'
#888200000000
1!
0$
b1000 %
1'
0*
b1000 +
#888210000000
0!
0'
#888220000000
1!
b1001 %
1'
b1001 +
#888230000000
0!
0'
#888240000000
1!
b0 %
1'
b0 +
#888250000000
0!
0'
#888260000000
1!
1$
b1 %
1'
1*
b1 +
#888270000000
0!
0'
#888280000000
1!
b10 %
1'
b10 +
#888290000000
0!
0'
#888300000000
1!
b11 %
1'
b11 +
#888310000000
0!
0'
#888320000000
1!
b100 %
1'
b100 +
#888330000000
0!
0'
#888340000000
1!
b101 %
1'
b101 +
#888350000000
0!
0'
#888360000000
1!
b110 %
1'
b110 +
#888370000000
0!
0'
#888380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#888390000000
0!
0'
#888400000000
1!
b1000 %
1'
b1000 +
#888410000000
0!
0'
#888420000000
1!
b1001 %
1'
b1001 +
#888430000000
0!
0'
#888440000000
1!
b0 %
1'
b0 +
#888450000000
0!
0'
#888460000000
1!
1$
b1 %
1'
1*
b1 +
#888470000000
0!
0'
#888480000000
1!
b10 %
1'
b10 +
#888490000000
0!
0'
#888500000000
1!
b11 %
1'
b11 +
#888510000000
0!
0'
#888520000000
1!
b100 %
1'
b100 +
#888530000000
0!
0'
#888540000000
1!
b101 %
1'
b101 +
#888550000000
0!
0'
#888560000000
1!
0$
b110 %
1'
0*
b110 +
#888570000000
0!
0'
#888580000000
1!
b111 %
1'
b111 +
#888590000000
1"
1(
#888600000000
0!
0"
b100 &
0'
0(
b100 ,
#888610000000
1!
b1000 %
1'
b1000 +
#888620000000
0!
0'
#888630000000
1!
b1001 %
1'
b1001 +
#888640000000
0!
0'
#888650000000
1!
b0 %
1'
b0 +
#888660000000
0!
0'
#888670000000
1!
1$
b1 %
1'
1*
b1 +
#888680000000
0!
0'
#888690000000
1!
b10 %
1'
b10 +
#888700000000
0!
0'
#888710000000
1!
b11 %
1'
b11 +
#888720000000
0!
0'
#888730000000
1!
b100 %
1'
b100 +
#888740000000
0!
0'
#888750000000
1!
b101 %
1'
b101 +
#888760000000
0!
0'
#888770000000
1!
b110 %
1'
b110 +
#888780000000
0!
0'
#888790000000
1!
b111 %
1'
b111 +
#888800000000
0!
0'
#888810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#888820000000
0!
0'
#888830000000
1!
b1001 %
1'
b1001 +
#888840000000
0!
0'
#888850000000
1!
b0 %
1'
b0 +
#888860000000
0!
0'
#888870000000
1!
1$
b1 %
1'
1*
b1 +
#888880000000
0!
0'
#888890000000
1!
b10 %
1'
b10 +
#888900000000
0!
0'
#888910000000
1!
b11 %
1'
b11 +
#888920000000
0!
0'
#888930000000
1!
b100 %
1'
b100 +
#888940000000
0!
0'
#888950000000
1!
b101 %
1'
b101 +
#888960000000
0!
0'
#888970000000
1!
0$
b110 %
1'
0*
b110 +
#888980000000
0!
0'
#888990000000
1!
b111 %
1'
b111 +
#889000000000
0!
0'
#889010000000
1!
b1000 %
1'
b1000 +
#889020000000
1"
1(
#889030000000
0!
0"
b100 &
0'
0(
b100 ,
#889040000000
1!
b1001 %
1'
b1001 +
#889050000000
0!
0'
#889060000000
1!
b0 %
1'
b0 +
#889070000000
0!
0'
#889080000000
1!
1$
b1 %
1'
1*
b1 +
#889090000000
0!
0'
#889100000000
1!
b10 %
1'
b10 +
#889110000000
0!
0'
#889120000000
1!
b11 %
1'
b11 +
#889130000000
0!
0'
#889140000000
1!
b100 %
1'
b100 +
#889150000000
0!
0'
#889160000000
1!
b101 %
1'
b101 +
#889170000000
0!
0'
#889180000000
1!
b110 %
1'
b110 +
#889190000000
0!
0'
#889200000000
1!
b111 %
1'
b111 +
#889210000000
0!
0'
#889220000000
1!
0$
b1000 %
1'
0*
b1000 +
#889230000000
0!
0'
#889240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#889250000000
0!
0'
#889260000000
1!
b0 %
1'
b0 +
#889270000000
0!
0'
#889280000000
1!
1$
b1 %
1'
1*
b1 +
#889290000000
0!
0'
#889300000000
1!
b10 %
1'
b10 +
#889310000000
0!
0'
#889320000000
1!
b11 %
1'
b11 +
#889330000000
0!
0'
#889340000000
1!
b100 %
1'
b100 +
#889350000000
0!
0'
#889360000000
1!
b101 %
1'
b101 +
#889370000000
0!
0'
#889380000000
1!
0$
b110 %
1'
0*
b110 +
#889390000000
0!
0'
#889400000000
1!
b111 %
1'
b111 +
#889410000000
0!
0'
#889420000000
1!
b1000 %
1'
b1000 +
#889430000000
0!
0'
#889440000000
1!
b1001 %
1'
b1001 +
#889450000000
1"
1(
#889460000000
0!
0"
b100 &
0'
0(
b100 ,
#889470000000
1!
b0 %
1'
b0 +
#889480000000
0!
0'
#889490000000
1!
1$
b1 %
1'
1*
b1 +
#889500000000
0!
0'
#889510000000
1!
b10 %
1'
b10 +
#889520000000
0!
0'
#889530000000
1!
b11 %
1'
b11 +
#889540000000
0!
0'
#889550000000
1!
b100 %
1'
b100 +
#889560000000
0!
0'
#889570000000
1!
b101 %
1'
b101 +
#889580000000
0!
0'
#889590000000
1!
b110 %
1'
b110 +
#889600000000
0!
0'
#889610000000
1!
b111 %
1'
b111 +
#889620000000
0!
0'
#889630000000
1!
0$
b1000 %
1'
0*
b1000 +
#889640000000
0!
0'
#889650000000
1!
b1001 %
1'
b1001 +
#889660000000
0!
0'
#889670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#889680000000
0!
0'
#889690000000
1!
1$
b1 %
1'
1*
b1 +
#889700000000
0!
0'
#889710000000
1!
b10 %
1'
b10 +
#889720000000
0!
0'
#889730000000
1!
b11 %
1'
b11 +
#889740000000
0!
0'
#889750000000
1!
b100 %
1'
b100 +
#889760000000
0!
0'
#889770000000
1!
b101 %
1'
b101 +
#889780000000
0!
0'
#889790000000
1!
0$
b110 %
1'
0*
b110 +
#889800000000
0!
0'
#889810000000
1!
b111 %
1'
b111 +
#889820000000
0!
0'
#889830000000
1!
b1000 %
1'
b1000 +
#889840000000
0!
0'
#889850000000
1!
b1001 %
1'
b1001 +
#889860000000
0!
0'
#889870000000
1!
b0 %
1'
b0 +
#889880000000
1"
1(
#889890000000
0!
0"
b100 &
0'
0(
b100 ,
#889900000000
1!
1$
b1 %
1'
1*
b1 +
#889910000000
0!
0'
#889920000000
1!
b10 %
1'
b10 +
#889930000000
0!
0'
#889940000000
1!
b11 %
1'
b11 +
#889950000000
0!
0'
#889960000000
1!
b100 %
1'
b100 +
#889970000000
0!
0'
#889980000000
1!
b101 %
1'
b101 +
#889990000000
0!
0'
#890000000000
1!
b110 %
1'
b110 +
#890010000000
0!
0'
#890020000000
1!
b111 %
1'
b111 +
#890030000000
0!
0'
#890040000000
1!
0$
b1000 %
1'
0*
b1000 +
#890050000000
0!
0'
#890060000000
1!
b1001 %
1'
b1001 +
#890070000000
0!
0'
#890080000000
1!
b0 %
1'
b0 +
#890090000000
0!
0'
#890100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#890110000000
0!
0'
#890120000000
1!
b10 %
1'
b10 +
#890130000000
0!
0'
#890140000000
1!
b11 %
1'
b11 +
#890150000000
0!
0'
#890160000000
1!
b100 %
1'
b100 +
#890170000000
0!
0'
#890180000000
1!
b101 %
1'
b101 +
#890190000000
0!
0'
#890200000000
1!
0$
b110 %
1'
0*
b110 +
#890210000000
0!
0'
#890220000000
1!
b111 %
1'
b111 +
#890230000000
0!
0'
#890240000000
1!
b1000 %
1'
b1000 +
#890250000000
0!
0'
#890260000000
1!
b1001 %
1'
b1001 +
#890270000000
0!
0'
#890280000000
1!
b0 %
1'
b0 +
#890290000000
0!
0'
#890300000000
1!
1$
b1 %
1'
1*
b1 +
#890310000000
1"
1(
#890320000000
0!
0"
b100 &
0'
0(
b100 ,
#890330000000
1!
b10 %
1'
b10 +
#890340000000
0!
0'
#890350000000
1!
b11 %
1'
b11 +
#890360000000
0!
0'
#890370000000
1!
b100 %
1'
b100 +
#890380000000
0!
0'
#890390000000
1!
b101 %
1'
b101 +
#890400000000
0!
0'
#890410000000
1!
b110 %
1'
b110 +
#890420000000
0!
0'
#890430000000
1!
b111 %
1'
b111 +
#890440000000
0!
0'
#890450000000
1!
0$
b1000 %
1'
0*
b1000 +
#890460000000
0!
0'
#890470000000
1!
b1001 %
1'
b1001 +
#890480000000
0!
0'
#890490000000
1!
b0 %
1'
b0 +
#890500000000
0!
0'
#890510000000
1!
1$
b1 %
1'
1*
b1 +
#890520000000
0!
0'
#890530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#890540000000
0!
0'
#890550000000
1!
b11 %
1'
b11 +
#890560000000
0!
0'
#890570000000
1!
b100 %
1'
b100 +
#890580000000
0!
0'
#890590000000
1!
b101 %
1'
b101 +
#890600000000
0!
0'
#890610000000
1!
0$
b110 %
1'
0*
b110 +
#890620000000
0!
0'
#890630000000
1!
b111 %
1'
b111 +
#890640000000
0!
0'
#890650000000
1!
b1000 %
1'
b1000 +
#890660000000
0!
0'
#890670000000
1!
b1001 %
1'
b1001 +
#890680000000
0!
0'
#890690000000
1!
b0 %
1'
b0 +
#890700000000
0!
0'
#890710000000
1!
1$
b1 %
1'
1*
b1 +
#890720000000
0!
0'
#890730000000
1!
b10 %
1'
b10 +
#890740000000
1"
1(
#890750000000
0!
0"
b100 &
0'
0(
b100 ,
#890760000000
1!
b11 %
1'
b11 +
#890770000000
0!
0'
#890780000000
1!
b100 %
1'
b100 +
#890790000000
0!
0'
#890800000000
1!
b101 %
1'
b101 +
#890810000000
0!
0'
#890820000000
1!
b110 %
1'
b110 +
#890830000000
0!
0'
#890840000000
1!
b111 %
1'
b111 +
#890850000000
0!
0'
#890860000000
1!
0$
b1000 %
1'
0*
b1000 +
#890870000000
0!
0'
#890880000000
1!
b1001 %
1'
b1001 +
#890890000000
0!
0'
#890900000000
1!
b0 %
1'
b0 +
#890910000000
0!
0'
#890920000000
1!
1$
b1 %
1'
1*
b1 +
#890930000000
0!
0'
#890940000000
1!
b10 %
1'
b10 +
#890950000000
0!
0'
#890960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#890970000000
0!
0'
#890980000000
1!
b100 %
1'
b100 +
#890990000000
0!
0'
#891000000000
1!
b101 %
1'
b101 +
#891010000000
0!
0'
#891020000000
1!
0$
b110 %
1'
0*
b110 +
#891030000000
0!
0'
#891040000000
1!
b111 %
1'
b111 +
#891050000000
0!
0'
#891060000000
1!
b1000 %
1'
b1000 +
#891070000000
0!
0'
#891080000000
1!
b1001 %
1'
b1001 +
#891090000000
0!
0'
#891100000000
1!
b0 %
1'
b0 +
#891110000000
0!
0'
#891120000000
1!
1$
b1 %
1'
1*
b1 +
#891130000000
0!
0'
#891140000000
1!
b10 %
1'
b10 +
#891150000000
0!
0'
#891160000000
1!
b11 %
1'
b11 +
#891170000000
1"
1(
#891180000000
0!
0"
b100 &
0'
0(
b100 ,
#891190000000
1!
b100 %
1'
b100 +
#891200000000
0!
0'
#891210000000
1!
b101 %
1'
b101 +
#891220000000
0!
0'
#891230000000
1!
b110 %
1'
b110 +
#891240000000
0!
0'
#891250000000
1!
b111 %
1'
b111 +
#891260000000
0!
0'
#891270000000
1!
0$
b1000 %
1'
0*
b1000 +
#891280000000
0!
0'
#891290000000
1!
b1001 %
1'
b1001 +
#891300000000
0!
0'
#891310000000
1!
b0 %
1'
b0 +
#891320000000
0!
0'
#891330000000
1!
1$
b1 %
1'
1*
b1 +
#891340000000
0!
0'
#891350000000
1!
b10 %
1'
b10 +
#891360000000
0!
0'
#891370000000
1!
b11 %
1'
b11 +
#891380000000
0!
0'
#891390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#891400000000
0!
0'
#891410000000
1!
b101 %
1'
b101 +
#891420000000
0!
0'
#891430000000
1!
0$
b110 %
1'
0*
b110 +
#891440000000
0!
0'
#891450000000
1!
b111 %
1'
b111 +
#891460000000
0!
0'
#891470000000
1!
b1000 %
1'
b1000 +
#891480000000
0!
0'
#891490000000
1!
b1001 %
1'
b1001 +
#891500000000
0!
0'
#891510000000
1!
b0 %
1'
b0 +
#891520000000
0!
0'
#891530000000
1!
1$
b1 %
1'
1*
b1 +
#891540000000
0!
0'
#891550000000
1!
b10 %
1'
b10 +
#891560000000
0!
0'
#891570000000
1!
b11 %
1'
b11 +
#891580000000
0!
0'
#891590000000
1!
b100 %
1'
b100 +
#891600000000
1"
1(
#891610000000
0!
0"
b100 &
0'
0(
b100 ,
#891620000000
1!
b101 %
1'
b101 +
#891630000000
0!
0'
#891640000000
1!
b110 %
1'
b110 +
#891650000000
0!
0'
#891660000000
1!
b111 %
1'
b111 +
#891670000000
0!
0'
#891680000000
1!
0$
b1000 %
1'
0*
b1000 +
#891690000000
0!
0'
#891700000000
1!
b1001 %
1'
b1001 +
#891710000000
0!
0'
#891720000000
1!
b0 %
1'
b0 +
#891730000000
0!
0'
#891740000000
1!
1$
b1 %
1'
1*
b1 +
#891750000000
0!
0'
#891760000000
1!
b10 %
1'
b10 +
#891770000000
0!
0'
#891780000000
1!
b11 %
1'
b11 +
#891790000000
0!
0'
#891800000000
1!
b100 %
1'
b100 +
#891810000000
0!
0'
#891820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#891830000000
0!
0'
#891840000000
1!
0$
b110 %
1'
0*
b110 +
#891850000000
0!
0'
#891860000000
1!
b111 %
1'
b111 +
#891870000000
0!
0'
#891880000000
1!
b1000 %
1'
b1000 +
#891890000000
0!
0'
#891900000000
1!
b1001 %
1'
b1001 +
#891910000000
0!
0'
#891920000000
1!
b0 %
1'
b0 +
#891930000000
0!
0'
#891940000000
1!
1$
b1 %
1'
1*
b1 +
#891950000000
0!
0'
#891960000000
1!
b10 %
1'
b10 +
#891970000000
0!
0'
#891980000000
1!
b11 %
1'
b11 +
#891990000000
0!
0'
#892000000000
1!
b100 %
1'
b100 +
#892010000000
0!
0'
#892020000000
1!
b101 %
1'
b101 +
#892030000000
1"
1(
#892040000000
0!
0"
b100 &
0'
0(
b100 ,
#892050000000
1!
b110 %
1'
b110 +
#892060000000
0!
0'
#892070000000
1!
b111 %
1'
b111 +
#892080000000
0!
0'
#892090000000
1!
0$
b1000 %
1'
0*
b1000 +
#892100000000
0!
0'
#892110000000
1!
b1001 %
1'
b1001 +
#892120000000
0!
0'
#892130000000
1!
b0 %
1'
b0 +
#892140000000
0!
0'
#892150000000
1!
1$
b1 %
1'
1*
b1 +
#892160000000
0!
0'
#892170000000
1!
b10 %
1'
b10 +
#892180000000
0!
0'
#892190000000
1!
b11 %
1'
b11 +
#892200000000
0!
0'
#892210000000
1!
b100 %
1'
b100 +
#892220000000
0!
0'
#892230000000
1!
b101 %
1'
b101 +
#892240000000
0!
0'
#892250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#892260000000
0!
0'
#892270000000
1!
b111 %
1'
b111 +
#892280000000
0!
0'
#892290000000
1!
b1000 %
1'
b1000 +
#892300000000
0!
0'
#892310000000
1!
b1001 %
1'
b1001 +
#892320000000
0!
0'
#892330000000
1!
b0 %
1'
b0 +
#892340000000
0!
0'
#892350000000
1!
1$
b1 %
1'
1*
b1 +
#892360000000
0!
0'
#892370000000
1!
b10 %
1'
b10 +
#892380000000
0!
0'
#892390000000
1!
b11 %
1'
b11 +
#892400000000
0!
0'
#892410000000
1!
b100 %
1'
b100 +
#892420000000
0!
0'
#892430000000
1!
b101 %
1'
b101 +
#892440000000
0!
0'
#892450000000
1!
0$
b110 %
1'
0*
b110 +
#892460000000
1"
1(
#892470000000
0!
0"
b100 &
0'
0(
b100 ,
#892480000000
1!
1$
b111 %
1'
1*
b111 +
#892490000000
0!
0'
#892500000000
1!
0$
b1000 %
1'
0*
b1000 +
#892510000000
0!
0'
#892520000000
1!
b1001 %
1'
b1001 +
#892530000000
0!
0'
#892540000000
1!
b0 %
1'
b0 +
#892550000000
0!
0'
#892560000000
1!
1$
b1 %
1'
1*
b1 +
#892570000000
0!
0'
#892580000000
1!
b10 %
1'
b10 +
#892590000000
0!
0'
#892600000000
1!
b11 %
1'
b11 +
#892610000000
0!
0'
#892620000000
1!
b100 %
1'
b100 +
#892630000000
0!
0'
#892640000000
1!
b101 %
1'
b101 +
#892650000000
0!
0'
#892660000000
1!
b110 %
1'
b110 +
#892670000000
0!
0'
#892680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#892690000000
0!
0'
#892700000000
1!
b1000 %
1'
b1000 +
#892710000000
0!
0'
#892720000000
1!
b1001 %
1'
b1001 +
#892730000000
0!
0'
#892740000000
1!
b0 %
1'
b0 +
#892750000000
0!
0'
#892760000000
1!
1$
b1 %
1'
1*
b1 +
#892770000000
0!
0'
#892780000000
1!
b10 %
1'
b10 +
#892790000000
0!
0'
#892800000000
1!
b11 %
1'
b11 +
#892810000000
0!
0'
#892820000000
1!
b100 %
1'
b100 +
#892830000000
0!
0'
#892840000000
1!
b101 %
1'
b101 +
#892850000000
0!
0'
#892860000000
1!
0$
b110 %
1'
0*
b110 +
#892870000000
0!
0'
#892880000000
1!
b111 %
1'
b111 +
#892890000000
1"
1(
#892900000000
0!
0"
b100 &
0'
0(
b100 ,
#892910000000
1!
b1000 %
1'
b1000 +
#892920000000
0!
0'
#892930000000
1!
b1001 %
1'
b1001 +
#892940000000
0!
0'
#892950000000
1!
b0 %
1'
b0 +
#892960000000
0!
0'
#892970000000
1!
1$
b1 %
1'
1*
b1 +
#892980000000
0!
0'
#892990000000
1!
b10 %
1'
b10 +
#893000000000
0!
0'
#893010000000
1!
b11 %
1'
b11 +
#893020000000
0!
0'
#893030000000
1!
b100 %
1'
b100 +
#893040000000
0!
0'
#893050000000
1!
b101 %
1'
b101 +
#893060000000
0!
0'
#893070000000
1!
b110 %
1'
b110 +
#893080000000
0!
0'
#893090000000
1!
b111 %
1'
b111 +
#893100000000
0!
0'
#893110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#893120000000
0!
0'
#893130000000
1!
b1001 %
1'
b1001 +
#893140000000
0!
0'
#893150000000
1!
b0 %
1'
b0 +
#893160000000
0!
0'
#893170000000
1!
1$
b1 %
1'
1*
b1 +
#893180000000
0!
0'
#893190000000
1!
b10 %
1'
b10 +
#893200000000
0!
0'
#893210000000
1!
b11 %
1'
b11 +
#893220000000
0!
0'
#893230000000
1!
b100 %
1'
b100 +
#893240000000
0!
0'
#893250000000
1!
b101 %
1'
b101 +
#893260000000
0!
0'
#893270000000
1!
0$
b110 %
1'
0*
b110 +
#893280000000
0!
0'
#893290000000
1!
b111 %
1'
b111 +
#893300000000
0!
0'
#893310000000
1!
b1000 %
1'
b1000 +
#893320000000
1"
1(
#893330000000
0!
0"
b100 &
0'
0(
b100 ,
#893340000000
1!
b1001 %
1'
b1001 +
#893350000000
0!
0'
#893360000000
1!
b0 %
1'
b0 +
#893370000000
0!
0'
#893380000000
1!
1$
b1 %
1'
1*
b1 +
#893390000000
0!
0'
#893400000000
1!
b10 %
1'
b10 +
#893410000000
0!
0'
#893420000000
1!
b11 %
1'
b11 +
#893430000000
0!
0'
#893440000000
1!
b100 %
1'
b100 +
#893450000000
0!
0'
#893460000000
1!
b101 %
1'
b101 +
#893470000000
0!
0'
#893480000000
1!
b110 %
1'
b110 +
#893490000000
0!
0'
#893500000000
1!
b111 %
1'
b111 +
#893510000000
0!
0'
#893520000000
1!
0$
b1000 %
1'
0*
b1000 +
#893530000000
0!
0'
#893540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#893550000000
0!
0'
#893560000000
1!
b0 %
1'
b0 +
#893570000000
0!
0'
#893580000000
1!
1$
b1 %
1'
1*
b1 +
#893590000000
0!
0'
#893600000000
1!
b10 %
1'
b10 +
#893610000000
0!
0'
#893620000000
1!
b11 %
1'
b11 +
#893630000000
0!
0'
#893640000000
1!
b100 %
1'
b100 +
#893650000000
0!
0'
#893660000000
1!
b101 %
1'
b101 +
#893670000000
0!
0'
#893680000000
1!
0$
b110 %
1'
0*
b110 +
#893690000000
0!
0'
#893700000000
1!
b111 %
1'
b111 +
#893710000000
0!
0'
#893720000000
1!
b1000 %
1'
b1000 +
#893730000000
0!
0'
#893740000000
1!
b1001 %
1'
b1001 +
#893750000000
1"
1(
#893760000000
0!
0"
b100 &
0'
0(
b100 ,
#893770000000
1!
b0 %
1'
b0 +
#893780000000
0!
0'
#893790000000
1!
1$
b1 %
1'
1*
b1 +
#893800000000
0!
0'
#893810000000
1!
b10 %
1'
b10 +
#893820000000
0!
0'
#893830000000
1!
b11 %
1'
b11 +
#893840000000
0!
0'
#893850000000
1!
b100 %
1'
b100 +
#893860000000
0!
0'
#893870000000
1!
b101 %
1'
b101 +
#893880000000
0!
0'
#893890000000
1!
b110 %
1'
b110 +
#893900000000
0!
0'
#893910000000
1!
b111 %
1'
b111 +
#893920000000
0!
0'
#893930000000
1!
0$
b1000 %
1'
0*
b1000 +
#893940000000
0!
0'
#893950000000
1!
b1001 %
1'
b1001 +
#893960000000
0!
0'
#893970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#893980000000
0!
0'
#893990000000
1!
1$
b1 %
1'
1*
b1 +
#894000000000
0!
0'
#894010000000
1!
b10 %
1'
b10 +
#894020000000
0!
0'
#894030000000
1!
b11 %
1'
b11 +
#894040000000
0!
0'
#894050000000
1!
b100 %
1'
b100 +
#894060000000
0!
0'
#894070000000
1!
b101 %
1'
b101 +
#894080000000
0!
0'
#894090000000
1!
0$
b110 %
1'
0*
b110 +
#894100000000
0!
0'
#894110000000
1!
b111 %
1'
b111 +
#894120000000
0!
0'
#894130000000
1!
b1000 %
1'
b1000 +
#894140000000
0!
0'
#894150000000
1!
b1001 %
1'
b1001 +
#894160000000
0!
0'
#894170000000
1!
b0 %
1'
b0 +
#894180000000
1"
1(
#894190000000
0!
0"
b100 &
0'
0(
b100 ,
#894200000000
1!
1$
b1 %
1'
1*
b1 +
#894210000000
0!
0'
#894220000000
1!
b10 %
1'
b10 +
#894230000000
0!
0'
#894240000000
1!
b11 %
1'
b11 +
#894250000000
0!
0'
#894260000000
1!
b100 %
1'
b100 +
#894270000000
0!
0'
#894280000000
1!
b101 %
1'
b101 +
#894290000000
0!
0'
#894300000000
1!
b110 %
1'
b110 +
#894310000000
0!
0'
#894320000000
1!
b111 %
1'
b111 +
#894330000000
0!
0'
#894340000000
1!
0$
b1000 %
1'
0*
b1000 +
#894350000000
0!
0'
#894360000000
1!
b1001 %
1'
b1001 +
#894370000000
0!
0'
#894380000000
1!
b0 %
1'
b0 +
#894390000000
0!
0'
#894400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#894410000000
0!
0'
#894420000000
1!
b10 %
1'
b10 +
#894430000000
0!
0'
#894440000000
1!
b11 %
1'
b11 +
#894450000000
0!
0'
#894460000000
1!
b100 %
1'
b100 +
#894470000000
0!
0'
#894480000000
1!
b101 %
1'
b101 +
#894490000000
0!
0'
#894500000000
1!
0$
b110 %
1'
0*
b110 +
#894510000000
0!
0'
#894520000000
1!
b111 %
1'
b111 +
#894530000000
0!
0'
#894540000000
1!
b1000 %
1'
b1000 +
#894550000000
0!
0'
#894560000000
1!
b1001 %
1'
b1001 +
#894570000000
0!
0'
#894580000000
1!
b0 %
1'
b0 +
#894590000000
0!
0'
#894600000000
1!
1$
b1 %
1'
1*
b1 +
#894610000000
1"
1(
#894620000000
0!
0"
b100 &
0'
0(
b100 ,
#894630000000
1!
b10 %
1'
b10 +
#894640000000
0!
0'
#894650000000
1!
b11 %
1'
b11 +
#894660000000
0!
0'
#894670000000
1!
b100 %
1'
b100 +
#894680000000
0!
0'
#894690000000
1!
b101 %
1'
b101 +
#894700000000
0!
0'
#894710000000
1!
b110 %
1'
b110 +
#894720000000
0!
0'
#894730000000
1!
b111 %
1'
b111 +
#894740000000
0!
0'
#894750000000
1!
0$
b1000 %
1'
0*
b1000 +
#894760000000
0!
0'
#894770000000
1!
b1001 %
1'
b1001 +
#894780000000
0!
0'
#894790000000
1!
b0 %
1'
b0 +
#894800000000
0!
0'
#894810000000
1!
1$
b1 %
1'
1*
b1 +
#894820000000
0!
0'
#894830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#894840000000
0!
0'
#894850000000
1!
b11 %
1'
b11 +
#894860000000
0!
0'
#894870000000
1!
b100 %
1'
b100 +
#894880000000
0!
0'
#894890000000
1!
b101 %
1'
b101 +
#894900000000
0!
0'
#894910000000
1!
0$
b110 %
1'
0*
b110 +
#894920000000
0!
0'
#894930000000
1!
b111 %
1'
b111 +
#894940000000
0!
0'
#894950000000
1!
b1000 %
1'
b1000 +
#894960000000
0!
0'
#894970000000
1!
b1001 %
1'
b1001 +
#894980000000
0!
0'
#894990000000
1!
b0 %
1'
b0 +
#895000000000
0!
0'
#895010000000
1!
1$
b1 %
1'
1*
b1 +
#895020000000
0!
0'
#895030000000
1!
b10 %
1'
b10 +
#895040000000
1"
1(
#895050000000
0!
0"
b100 &
0'
0(
b100 ,
#895060000000
1!
b11 %
1'
b11 +
#895070000000
0!
0'
#895080000000
1!
b100 %
1'
b100 +
#895090000000
0!
0'
#895100000000
1!
b101 %
1'
b101 +
#895110000000
0!
0'
#895120000000
1!
b110 %
1'
b110 +
#895130000000
0!
0'
#895140000000
1!
b111 %
1'
b111 +
#895150000000
0!
0'
#895160000000
1!
0$
b1000 %
1'
0*
b1000 +
#895170000000
0!
0'
#895180000000
1!
b1001 %
1'
b1001 +
#895190000000
0!
0'
#895200000000
1!
b0 %
1'
b0 +
#895210000000
0!
0'
#895220000000
1!
1$
b1 %
1'
1*
b1 +
#895230000000
0!
0'
#895240000000
1!
b10 %
1'
b10 +
#895250000000
0!
0'
#895260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#895270000000
0!
0'
#895280000000
1!
b100 %
1'
b100 +
#895290000000
0!
0'
#895300000000
1!
b101 %
1'
b101 +
#895310000000
0!
0'
#895320000000
1!
0$
b110 %
1'
0*
b110 +
#895330000000
0!
0'
#895340000000
1!
b111 %
1'
b111 +
#895350000000
0!
0'
#895360000000
1!
b1000 %
1'
b1000 +
#895370000000
0!
0'
#895380000000
1!
b1001 %
1'
b1001 +
#895390000000
0!
0'
#895400000000
1!
b0 %
1'
b0 +
#895410000000
0!
0'
#895420000000
1!
1$
b1 %
1'
1*
b1 +
#895430000000
0!
0'
#895440000000
1!
b10 %
1'
b10 +
#895450000000
0!
0'
#895460000000
1!
b11 %
1'
b11 +
#895470000000
1"
1(
#895480000000
0!
0"
b100 &
0'
0(
b100 ,
#895490000000
1!
b100 %
1'
b100 +
#895500000000
0!
0'
#895510000000
1!
b101 %
1'
b101 +
#895520000000
0!
0'
#895530000000
1!
b110 %
1'
b110 +
#895540000000
0!
0'
#895550000000
1!
b111 %
1'
b111 +
#895560000000
0!
0'
#895570000000
1!
0$
b1000 %
1'
0*
b1000 +
#895580000000
0!
0'
#895590000000
1!
b1001 %
1'
b1001 +
#895600000000
0!
0'
#895610000000
1!
b0 %
1'
b0 +
#895620000000
0!
0'
#895630000000
1!
1$
b1 %
1'
1*
b1 +
#895640000000
0!
0'
#895650000000
1!
b10 %
1'
b10 +
#895660000000
0!
0'
#895670000000
1!
b11 %
1'
b11 +
#895680000000
0!
0'
#895690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#895700000000
0!
0'
#895710000000
1!
b101 %
1'
b101 +
#895720000000
0!
0'
#895730000000
1!
0$
b110 %
1'
0*
b110 +
#895740000000
0!
0'
#895750000000
1!
b111 %
1'
b111 +
#895760000000
0!
0'
#895770000000
1!
b1000 %
1'
b1000 +
#895780000000
0!
0'
#895790000000
1!
b1001 %
1'
b1001 +
#895800000000
0!
0'
#895810000000
1!
b0 %
1'
b0 +
#895820000000
0!
0'
#895830000000
1!
1$
b1 %
1'
1*
b1 +
#895840000000
0!
0'
#895850000000
1!
b10 %
1'
b10 +
#895860000000
0!
0'
#895870000000
1!
b11 %
1'
b11 +
#895880000000
0!
0'
#895890000000
1!
b100 %
1'
b100 +
#895900000000
1"
1(
#895910000000
0!
0"
b100 &
0'
0(
b100 ,
#895920000000
1!
b101 %
1'
b101 +
#895930000000
0!
0'
#895940000000
1!
b110 %
1'
b110 +
#895950000000
0!
0'
#895960000000
1!
b111 %
1'
b111 +
#895970000000
0!
0'
#895980000000
1!
0$
b1000 %
1'
0*
b1000 +
#895990000000
0!
0'
#896000000000
1!
b1001 %
1'
b1001 +
#896010000000
0!
0'
#896020000000
1!
b0 %
1'
b0 +
#896030000000
0!
0'
#896040000000
1!
1$
b1 %
1'
1*
b1 +
#896050000000
0!
0'
#896060000000
1!
b10 %
1'
b10 +
#896070000000
0!
0'
#896080000000
1!
b11 %
1'
b11 +
#896090000000
0!
0'
#896100000000
1!
b100 %
1'
b100 +
#896110000000
0!
0'
#896120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#896130000000
0!
0'
#896140000000
1!
0$
b110 %
1'
0*
b110 +
#896150000000
0!
0'
#896160000000
1!
b111 %
1'
b111 +
#896170000000
0!
0'
#896180000000
1!
b1000 %
1'
b1000 +
#896190000000
0!
0'
#896200000000
1!
b1001 %
1'
b1001 +
#896210000000
0!
0'
#896220000000
1!
b0 %
1'
b0 +
#896230000000
0!
0'
#896240000000
1!
1$
b1 %
1'
1*
b1 +
#896250000000
0!
0'
#896260000000
1!
b10 %
1'
b10 +
#896270000000
0!
0'
#896280000000
1!
b11 %
1'
b11 +
#896290000000
0!
0'
#896300000000
1!
b100 %
1'
b100 +
#896310000000
0!
0'
#896320000000
1!
b101 %
1'
b101 +
#896330000000
1"
1(
#896340000000
0!
0"
b100 &
0'
0(
b100 ,
#896350000000
1!
b110 %
1'
b110 +
#896360000000
0!
0'
#896370000000
1!
b111 %
1'
b111 +
#896380000000
0!
0'
#896390000000
1!
0$
b1000 %
1'
0*
b1000 +
#896400000000
0!
0'
#896410000000
1!
b1001 %
1'
b1001 +
#896420000000
0!
0'
#896430000000
1!
b0 %
1'
b0 +
#896440000000
0!
0'
#896450000000
1!
1$
b1 %
1'
1*
b1 +
#896460000000
0!
0'
#896470000000
1!
b10 %
1'
b10 +
#896480000000
0!
0'
#896490000000
1!
b11 %
1'
b11 +
#896500000000
0!
0'
#896510000000
1!
b100 %
1'
b100 +
#896520000000
0!
0'
#896530000000
1!
b101 %
1'
b101 +
#896540000000
0!
0'
#896550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#896560000000
0!
0'
#896570000000
1!
b111 %
1'
b111 +
#896580000000
0!
0'
#896590000000
1!
b1000 %
1'
b1000 +
#896600000000
0!
0'
#896610000000
1!
b1001 %
1'
b1001 +
#896620000000
0!
0'
#896630000000
1!
b0 %
1'
b0 +
#896640000000
0!
0'
#896650000000
1!
1$
b1 %
1'
1*
b1 +
#896660000000
0!
0'
#896670000000
1!
b10 %
1'
b10 +
#896680000000
0!
0'
#896690000000
1!
b11 %
1'
b11 +
#896700000000
0!
0'
#896710000000
1!
b100 %
1'
b100 +
#896720000000
0!
0'
#896730000000
1!
b101 %
1'
b101 +
#896740000000
0!
0'
#896750000000
1!
0$
b110 %
1'
0*
b110 +
#896760000000
1"
1(
#896770000000
0!
0"
b100 &
0'
0(
b100 ,
#896780000000
1!
1$
b111 %
1'
1*
b111 +
#896790000000
0!
0'
#896800000000
1!
0$
b1000 %
1'
0*
b1000 +
#896810000000
0!
0'
#896820000000
1!
b1001 %
1'
b1001 +
#896830000000
0!
0'
#896840000000
1!
b0 %
1'
b0 +
#896850000000
0!
0'
#896860000000
1!
1$
b1 %
1'
1*
b1 +
#896870000000
0!
0'
#896880000000
1!
b10 %
1'
b10 +
#896890000000
0!
0'
#896900000000
1!
b11 %
1'
b11 +
#896910000000
0!
0'
#896920000000
1!
b100 %
1'
b100 +
#896930000000
0!
0'
#896940000000
1!
b101 %
1'
b101 +
#896950000000
0!
0'
#896960000000
1!
b110 %
1'
b110 +
#896970000000
0!
0'
#896980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#896990000000
0!
0'
#897000000000
1!
b1000 %
1'
b1000 +
#897010000000
0!
0'
#897020000000
1!
b1001 %
1'
b1001 +
#897030000000
0!
0'
#897040000000
1!
b0 %
1'
b0 +
#897050000000
0!
0'
#897060000000
1!
1$
b1 %
1'
1*
b1 +
#897070000000
0!
0'
#897080000000
1!
b10 %
1'
b10 +
#897090000000
0!
0'
#897100000000
1!
b11 %
1'
b11 +
#897110000000
0!
0'
#897120000000
1!
b100 %
1'
b100 +
#897130000000
0!
0'
#897140000000
1!
b101 %
1'
b101 +
#897150000000
0!
0'
#897160000000
1!
0$
b110 %
1'
0*
b110 +
#897170000000
0!
0'
#897180000000
1!
b111 %
1'
b111 +
#897190000000
1"
1(
#897200000000
0!
0"
b100 &
0'
0(
b100 ,
#897210000000
1!
b1000 %
1'
b1000 +
#897220000000
0!
0'
#897230000000
1!
b1001 %
1'
b1001 +
#897240000000
0!
0'
#897250000000
1!
b0 %
1'
b0 +
#897260000000
0!
0'
#897270000000
1!
1$
b1 %
1'
1*
b1 +
#897280000000
0!
0'
#897290000000
1!
b10 %
1'
b10 +
#897300000000
0!
0'
#897310000000
1!
b11 %
1'
b11 +
#897320000000
0!
0'
#897330000000
1!
b100 %
1'
b100 +
#897340000000
0!
0'
#897350000000
1!
b101 %
1'
b101 +
#897360000000
0!
0'
#897370000000
1!
b110 %
1'
b110 +
#897380000000
0!
0'
#897390000000
1!
b111 %
1'
b111 +
#897400000000
0!
0'
#897410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#897420000000
0!
0'
#897430000000
1!
b1001 %
1'
b1001 +
#897440000000
0!
0'
#897450000000
1!
b0 %
1'
b0 +
#897460000000
0!
0'
#897470000000
1!
1$
b1 %
1'
1*
b1 +
#897480000000
0!
0'
#897490000000
1!
b10 %
1'
b10 +
#897500000000
0!
0'
#897510000000
1!
b11 %
1'
b11 +
#897520000000
0!
0'
#897530000000
1!
b100 %
1'
b100 +
#897540000000
0!
0'
#897550000000
1!
b101 %
1'
b101 +
#897560000000
0!
0'
#897570000000
1!
0$
b110 %
1'
0*
b110 +
#897580000000
0!
0'
#897590000000
1!
b111 %
1'
b111 +
#897600000000
0!
0'
#897610000000
1!
b1000 %
1'
b1000 +
#897620000000
1"
1(
#897630000000
0!
0"
b100 &
0'
0(
b100 ,
#897640000000
1!
b1001 %
1'
b1001 +
#897650000000
0!
0'
#897660000000
1!
b0 %
1'
b0 +
#897670000000
0!
0'
#897680000000
1!
1$
b1 %
1'
1*
b1 +
#897690000000
0!
0'
#897700000000
1!
b10 %
1'
b10 +
#897710000000
0!
0'
#897720000000
1!
b11 %
1'
b11 +
#897730000000
0!
0'
#897740000000
1!
b100 %
1'
b100 +
#897750000000
0!
0'
#897760000000
1!
b101 %
1'
b101 +
#897770000000
0!
0'
#897780000000
1!
b110 %
1'
b110 +
#897790000000
0!
0'
#897800000000
1!
b111 %
1'
b111 +
#897810000000
0!
0'
#897820000000
1!
0$
b1000 %
1'
0*
b1000 +
#897830000000
0!
0'
#897840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#897850000000
0!
0'
#897860000000
1!
b0 %
1'
b0 +
#897870000000
0!
0'
#897880000000
1!
1$
b1 %
1'
1*
b1 +
#897890000000
0!
0'
#897900000000
1!
b10 %
1'
b10 +
#897910000000
0!
0'
#897920000000
1!
b11 %
1'
b11 +
#897930000000
0!
0'
#897940000000
1!
b100 %
1'
b100 +
#897950000000
0!
0'
#897960000000
1!
b101 %
1'
b101 +
#897970000000
0!
0'
#897980000000
1!
0$
b110 %
1'
0*
b110 +
#897990000000
0!
0'
#898000000000
1!
b111 %
1'
b111 +
#898010000000
0!
0'
#898020000000
1!
b1000 %
1'
b1000 +
#898030000000
0!
0'
#898040000000
1!
b1001 %
1'
b1001 +
#898050000000
1"
1(
#898060000000
0!
0"
b100 &
0'
0(
b100 ,
#898070000000
1!
b0 %
1'
b0 +
#898080000000
0!
0'
#898090000000
1!
1$
b1 %
1'
1*
b1 +
#898100000000
0!
0'
#898110000000
1!
b10 %
1'
b10 +
#898120000000
0!
0'
#898130000000
1!
b11 %
1'
b11 +
#898140000000
0!
0'
#898150000000
1!
b100 %
1'
b100 +
#898160000000
0!
0'
#898170000000
1!
b101 %
1'
b101 +
#898180000000
0!
0'
#898190000000
1!
b110 %
1'
b110 +
#898200000000
0!
0'
#898210000000
1!
b111 %
1'
b111 +
#898220000000
0!
0'
#898230000000
1!
0$
b1000 %
1'
0*
b1000 +
#898240000000
0!
0'
#898250000000
1!
b1001 %
1'
b1001 +
#898260000000
0!
0'
#898270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#898280000000
0!
0'
#898290000000
1!
1$
b1 %
1'
1*
b1 +
#898300000000
0!
0'
#898310000000
1!
b10 %
1'
b10 +
#898320000000
0!
0'
#898330000000
1!
b11 %
1'
b11 +
#898340000000
0!
0'
#898350000000
1!
b100 %
1'
b100 +
#898360000000
0!
0'
#898370000000
1!
b101 %
1'
b101 +
#898380000000
0!
0'
#898390000000
1!
0$
b110 %
1'
0*
b110 +
#898400000000
0!
0'
#898410000000
1!
b111 %
1'
b111 +
#898420000000
0!
0'
#898430000000
1!
b1000 %
1'
b1000 +
#898440000000
0!
0'
#898450000000
1!
b1001 %
1'
b1001 +
#898460000000
0!
0'
#898470000000
1!
b0 %
1'
b0 +
#898480000000
1"
1(
#898490000000
0!
0"
b100 &
0'
0(
b100 ,
#898500000000
1!
1$
b1 %
1'
1*
b1 +
#898510000000
0!
0'
#898520000000
1!
b10 %
1'
b10 +
#898530000000
0!
0'
#898540000000
1!
b11 %
1'
b11 +
#898550000000
0!
0'
#898560000000
1!
b100 %
1'
b100 +
#898570000000
0!
0'
#898580000000
1!
b101 %
1'
b101 +
#898590000000
0!
0'
#898600000000
1!
b110 %
1'
b110 +
#898610000000
0!
0'
#898620000000
1!
b111 %
1'
b111 +
#898630000000
0!
0'
#898640000000
1!
0$
b1000 %
1'
0*
b1000 +
#898650000000
0!
0'
#898660000000
1!
b1001 %
1'
b1001 +
#898670000000
0!
0'
#898680000000
1!
b0 %
1'
b0 +
#898690000000
0!
0'
#898700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#898710000000
0!
0'
#898720000000
1!
b10 %
1'
b10 +
#898730000000
0!
0'
#898740000000
1!
b11 %
1'
b11 +
#898750000000
0!
0'
#898760000000
1!
b100 %
1'
b100 +
#898770000000
0!
0'
#898780000000
1!
b101 %
1'
b101 +
#898790000000
0!
0'
#898800000000
1!
0$
b110 %
1'
0*
b110 +
#898810000000
0!
0'
#898820000000
1!
b111 %
1'
b111 +
#898830000000
0!
0'
#898840000000
1!
b1000 %
1'
b1000 +
#898850000000
0!
0'
#898860000000
1!
b1001 %
1'
b1001 +
#898870000000
0!
0'
#898880000000
1!
b0 %
1'
b0 +
#898890000000
0!
0'
#898900000000
1!
1$
b1 %
1'
1*
b1 +
#898910000000
1"
1(
#898920000000
0!
0"
b100 &
0'
0(
b100 ,
#898930000000
1!
b10 %
1'
b10 +
#898940000000
0!
0'
#898950000000
1!
b11 %
1'
b11 +
#898960000000
0!
0'
#898970000000
1!
b100 %
1'
b100 +
#898980000000
0!
0'
#898990000000
1!
b101 %
1'
b101 +
#899000000000
0!
0'
#899010000000
1!
b110 %
1'
b110 +
#899020000000
0!
0'
#899030000000
1!
b111 %
1'
b111 +
#899040000000
0!
0'
#899050000000
1!
0$
b1000 %
1'
0*
b1000 +
#899060000000
0!
0'
#899070000000
1!
b1001 %
1'
b1001 +
#899080000000
0!
0'
#899090000000
1!
b0 %
1'
b0 +
#899100000000
0!
0'
#899110000000
1!
1$
b1 %
1'
1*
b1 +
#899120000000
0!
0'
#899130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#899140000000
0!
0'
#899150000000
1!
b11 %
1'
b11 +
#899160000000
0!
0'
#899170000000
1!
b100 %
1'
b100 +
#899180000000
0!
0'
#899190000000
1!
b101 %
1'
b101 +
#899200000000
0!
0'
#899210000000
1!
0$
b110 %
1'
0*
b110 +
#899220000000
0!
0'
#899230000000
1!
b111 %
1'
b111 +
#899240000000
0!
0'
#899250000000
1!
b1000 %
1'
b1000 +
#899260000000
0!
0'
#899270000000
1!
b1001 %
1'
b1001 +
#899280000000
0!
0'
#899290000000
1!
b0 %
1'
b0 +
#899300000000
0!
0'
#899310000000
1!
1$
b1 %
1'
1*
b1 +
#899320000000
0!
0'
#899330000000
1!
b10 %
1'
b10 +
#899340000000
1"
1(
#899350000000
0!
0"
b100 &
0'
0(
b100 ,
#899360000000
1!
b11 %
1'
b11 +
#899370000000
0!
0'
#899380000000
1!
b100 %
1'
b100 +
#899390000000
0!
0'
#899400000000
1!
b101 %
1'
b101 +
#899410000000
0!
0'
#899420000000
1!
b110 %
1'
b110 +
#899430000000
0!
0'
#899440000000
1!
b111 %
1'
b111 +
#899450000000
0!
0'
#899460000000
1!
0$
b1000 %
1'
0*
b1000 +
#899470000000
0!
0'
#899480000000
1!
b1001 %
1'
b1001 +
#899490000000
0!
0'
#899500000000
1!
b0 %
1'
b0 +
#899510000000
0!
0'
#899520000000
1!
1$
b1 %
1'
1*
b1 +
#899530000000
0!
0'
#899540000000
1!
b10 %
1'
b10 +
#899550000000
0!
0'
#899560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#899570000000
0!
0'
#899580000000
1!
b100 %
1'
b100 +
#899590000000
0!
0'
#899600000000
1!
b101 %
1'
b101 +
#899610000000
0!
0'
#899620000000
1!
0$
b110 %
1'
0*
b110 +
#899630000000
0!
0'
#899640000000
1!
b111 %
1'
b111 +
#899650000000
0!
0'
#899660000000
1!
b1000 %
1'
b1000 +
#899670000000
0!
0'
#899680000000
1!
b1001 %
1'
b1001 +
#899690000000
0!
0'
#899700000000
1!
b0 %
1'
b0 +
#899710000000
0!
0'
#899720000000
1!
1$
b1 %
1'
1*
b1 +
#899730000000
0!
0'
#899740000000
1!
b10 %
1'
b10 +
#899750000000
0!
0'
#899760000000
1!
b11 %
1'
b11 +
#899770000000
1"
1(
#899780000000
0!
0"
b100 &
0'
0(
b100 ,
#899790000000
1!
b100 %
1'
b100 +
#899800000000
0!
0'
#899810000000
1!
b101 %
1'
b101 +
#899820000000
0!
0'
#899830000000
1!
b110 %
1'
b110 +
#899840000000
0!
0'
#899850000000
1!
b111 %
1'
b111 +
#899860000000
0!
0'
#899870000000
1!
0$
b1000 %
1'
0*
b1000 +
#899880000000
0!
0'
#899890000000
1!
b1001 %
1'
b1001 +
#899900000000
0!
0'
#899910000000
1!
b0 %
1'
b0 +
#899920000000
0!
0'
#899930000000
1!
1$
b1 %
1'
1*
b1 +
#899940000000
0!
0'
#899950000000
1!
b10 %
1'
b10 +
#899960000000
0!
0'
#899970000000
1!
b11 %
1'
b11 +
#899980000000
0!
0'
#899990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#900000000000
0!
0'
#900010000000
1!
b101 %
1'
b101 +
#900020000000
0!
0'
#900030000000
1!
0$
b110 %
1'
0*
b110 +
#900040000000
0!
0'
#900050000000
1!
b111 %
1'
b111 +
#900060000000
0!
0'
#900070000000
1!
b1000 %
1'
b1000 +
#900080000000
0!
0'
#900090000000
1!
b1001 %
1'
b1001 +
#900100000000
0!
0'
#900110000000
1!
b0 %
1'
b0 +
#900120000000
0!
0'
#900130000000
1!
1$
b1 %
1'
1*
b1 +
#900140000000
0!
0'
#900150000000
1!
b10 %
1'
b10 +
#900160000000
0!
0'
#900170000000
1!
b11 %
1'
b11 +
#900180000000
0!
0'
#900190000000
1!
b100 %
1'
b100 +
#900200000000
1"
1(
#900210000000
0!
0"
b100 &
0'
0(
b100 ,
#900220000000
1!
b101 %
1'
b101 +
#900230000000
0!
0'
#900240000000
1!
b110 %
1'
b110 +
#900250000000
0!
0'
#900260000000
1!
b111 %
1'
b111 +
#900270000000
0!
0'
#900280000000
1!
0$
b1000 %
1'
0*
b1000 +
#900290000000
0!
0'
#900300000000
1!
b1001 %
1'
b1001 +
#900310000000
0!
0'
#900320000000
1!
b0 %
1'
b0 +
#900330000000
0!
0'
#900340000000
1!
1$
b1 %
1'
1*
b1 +
#900350000000
0!
0'
#900360000000
1!
b10 %
1'
b10 +
#900370000000
0!
0'
#900380000000
1!
b11 %
1'
b11 +
#900390000000
0!
0'
#900400000000
1!
b100 %
1'
b100 +
#900410000000
0!
0'
#900420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#900430000000
0!
0'
#900440000000
1!
0$
b110 %
1'
0*
b110 +
#900450000000
0!
0'
#900460000000
1!
b111 %
1'
b111 +
#900470000000
0!
0'
#900480000000
1!
b1000 %
1'
b1000 +
#900490000000
0!
0'
#900500000000
1!
b1001 %
1'
b1001 +
#900510000000
0!
0'
#900520000000
1!
b0 %
1'
b0 +
#900530000000
0!
0'
#900540000000
1!
1$
b1 %
1'
1*
b1 +
#900550000000
0!
0'
#900560000000
1!
b10 %
1'
b10 +
#900570000000
0!
0'
#900580000000
1!
b11 %
1'
b11 +
#900590000000
0!
0'
#900600000000
1!
b100 %
1'
b100 +
#900610000000
0!
0'
#900620000000
1!
b101 %
1'
b101 +
#900630000000
1"
1(
#900640000000
0!
0"
b100 &
0'
0(
b100 ,
#900650000000
1!
b110 %
1'
b110 +
#900660000000
0!
0'
#900670000000
1!
b111 %
1'
b111 +
#900680000000
0!
0'
#900690000000
1!
0$
b1000 %
1'
0*
b1000 +
#900700000000
0!
0'
#900710000000
1!
b1001 %
1'
b1001 +
#900720000000
0!
0'
#900730000000
1!
b0 %
1'
b0 +
#900740000000
0!
0'
#900750000000
1!
1$
b1 %
1'
1*
b1 +
#900760000000
0!
0'
#900770000000
1!
b10 %
1'
b10 +
#900780000000
0!
0'
#900790000000
1!
b11 %
1'
b11 +
#900800000000
0!
0'
#900810000000
1!
b100 %
1'
b100 +
#900820000000
0!
0'
#900830000000
1!
b101 %
1'
b101 +
#900840000000
0!
0'
#900850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#900860000000
0!
0'
#900870000000
1!
b111 %
1'
b111 +
#900880000000
0!
0'
#900890000000
1!
b1000 %
1'
b1000 +
#900900000000
0!
0'
#900910000000
1!
b1001 %
1'
b1001 +
#900920000000
0!
0'
#900930000000
1!
b0 %
1'
b0 +
#900940000000
0!
0'
#900950000000
1!
1$
b1 %
1'
1*
b1 +
#900960000000
0!
0'
#900970000000
1!
b10 %
1'
b10 +
#900980000000
0!
0'
#900990000000
1!
b11 %
1'
b11 +
#901000000000
0!
0'
#901010000000
1!
b100 %
1'
b100 +
#901020000000
0!
0'
#901030000000
1!
b101 %
1'
b101 +
#901040000000
0!
0'
#901050000000
1!
0$
b110 %
1'
0*
b110 +
#901060000000
1"
1(
#901070000000
0!
0"
b100 &
0'
0(
b100 ,
#901080000000
1!
1$
b111 %
1'
1*
b111 +
#901090000000
0!
0'
#901100000000
1!
0$
b1000 %
1'
0*
b1000 +
#901110000000
0!
0'
#901120000000
1!
b1001 %
1'
b1001 +
#901130000000
0!
0'
#901140000000
1!
b0 %
1'
b0 +
#901150000000
0!
0'
#901160000000
1!
1$
b1 %
1'
1*
b1 +
#901170000000
0!
0'
#901180000000
1!
b10 %
1'
b10 +
#901190000000
0!
0'
#901200000000
1!
b11 %
1'
b11 +
#901210000000
0!
0'
#901220000000
1!
b100 %
1'
b100 +
#901230000000
0!
0'
#901240000000
1!
b101 %
1'
b101 +
#901250000000
0!
0'
#901260000000
1!
b110 %
1'
b110 +
#901270000000
0!
0'
#901280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#901290000000
0!
0'
#901300000000
1!
b1000 %
1'
b1000 +
#901310000000
0!
0'
#901320000000
1!
b1001 %
1'
b1001 +
#901330000000
0!
0'
#901340000000
1!
b0 %
1'
b0 +
#901350000000
0!
0'
#901360000000
1!
1$
b1 %
1'
1*
b1 +
#901370000000
0!
0'
#901380000000
1!
b10 %
1'
b10 +
#901390000000
0!
0'
#901400000000
1!
b11 %
1'
b11 +
#901410000000
0!
0'
#901420000000
1!
b100 %
1'
b100 +
#901430000000
0!
0'
#901440000000
1!
b101 %
1'
b101 +
#901450000000
0!
0'
#901460000000
1!
0$
b110 %
1'
0*
b110 +
#901470000000
0!
0'
#901480000000
1!
b111 %
1'
b111 +
#901490000000
1"
1(
#901500000000
0!
0"
b100 &
0'
0(
b100 ,
#901510000000
1!
b1000 %
1'
b1000 +
#901520000000
0!
0'
#901530000000
1!
b1001 %
1'
b1001 +
#901540000000
0!
0'
#901550000000
1!
b0 %
1'
b0 +
#901560000000
0!
0'
#901570000000
1!
1$
b1 %
1'
1*
b1 +
#901580000000
0!
0'
#901590000000
1!
b10 %
1'
b10 +
#901600000000
0!
0'
#901610000000
1!
b11 %
1'
b11 +
#901620000000
0!
0'
#901630000000
1!
b100 %
1'
b100 +
#901640000000
0!
0'
#901650000000
1!
b101 %
1'
b101 +
#901660000000
0!
0'
#901670000000
1!
b110 %
1'
b110 +
#901680000000
0!
0'
#901690000000
1!
b111 %
1'
b111 +
#901700000000
0!
0'
#901710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#901720000000
0!
0'
#901730000000
1!
b1001 %
1'
b1001 +
#901740000000
0!
0'
#901750000000
1!
b0 %
1'
b0 +
#901760000000
0!
0'
#901770000000
1!
1$
b1 %
1'
1*
b1 +
#901780000000
0!
0'
#901790000000
1!
b10 %
1'
b10 +
#901800000000
0!
0'
#901810000000
1!
b11 %
1'
b11 +
#901820000000
0!
0'
#901830000000
1!
b100 %
1'
b100 +
#901840000000
0!
0'
#901850000000
1!
b101 %
1'
b101 +
#901860000000
0!
0'
#901870000000
1!
0$
b110 %
1'
0*
b110 +
#901880000000
0!
0'
#901890000000
1!
b111 %
1'
b111 +
#901900000000
0!
0'
#901910000000
1!
b1000 %
1'
b1000 +
#901920000000
1"
1(
#901930000000
0!
0"
b100 &
0'
0(
b100 ,
#901940000000
1!
b1001 %
1'
b1001 +
#901950000000
0!
0'
#901960000000
1!
b0 %
1'
b0 +
#901970000000
0!
0'
#901980000000
1!
1$
b1 %
1'
1*
b1 +
#901990000000
0!
0'
#902000000000
1!
b10 %
1'
b10 +
#902010000000
0!
0'
#902020000000
1!
b11 %
1'
b11 +
#902030000000
0!
0'
#902040000000
1!
b100 %
1'
b100 +
#902050000000
0!
0'
#902060000000
1!
b101 %
1'
b101 +
#902070000000
0!
0'
#902080000000
1!
b110 %
1'
b110 +
#902090000000
0!
0'
#902100000000
1!
b111 %
1'
b111 +
#902110000000
0!
0'
#902120000000
1!
0$
b1000 %
1'
0*
b1000 +
#902130000000
0!
0'
#902140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#902150000000
0!
0'
#902160000000
1!
b0 %
1'
b0 +
#902170000000
0!
0'
#902180000000
1!
1$
b1 %
1'
1*
b1 +
#902190000000
0!
0'
#902200000000
1!
b10 %
1'
b10 +
#902210000000
0!
0'
#902220000000
1!
b11 %
1'
b11 +
#902230000000
0!
0'
#902240000000
1!
b100 %
1'
b100 +
#902250000000
0!
0'
#902260000000
1!
b101 %
1'
b101 +
#902270000000
0!
0'
#902280000000
1!
0$
b110 %
1'
0*
b110 +
#902290000000
0!
0'
#902300000000
1!
b111 %
1'
b111 +
#902310000000
0!
0'
#902320000000
1!
b1000 %
1'
b1000 +
#902330000000
0!
0'
#902340000000
1!
b1001 %
1'
b1001 +
#902350000000
1"
1(
#902360000000
0!
0"
b100 &
0'
0(
b100 ,
#902370000000
1!
b0 %
1'
b0 +
#902380000000
0!
0'
#902390000000
1!
1$
b1 %
1'
1*
b1 +
#902400000000
0!
0'
#902410000000
1!
b10 %
1'
b10 +
#902420000000
0!
0'
#902430000000
1!
b11 %
1'
b11 +
#902440000000
0!
0'
#902450000000
1!
b100 %
1'
b100 +
#902460000000
0!
0'
#902470000000
1!
b101 %
1'
b101 +
#902480000000
0!
0'
#902490000000
1!
b110 %
1'
b110 +
#902500000000
0!
0'
#902510000000
1!
b111 %
1'
b111 +
#902520000000
0!
0'
#902530000000
1!
0$
b1000 %
1'
0*
b1000 +
#902540000000
0!
0'
#902550000000
1!
b1001 %
1'
b1001 +
#902560000000
0!
0'
#902570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#902580000000
0!
0'
#902590000000
1!
1$
b1 %
1'
1*
b1 +
#902600000000
0!
0'
#902610000000
1!
b10 %
1'
b10 +
#902620000000
0!
0'
#902630000000
1!
b11 %
1'
b11 +
#902640000000
0!
0'
#902650000000
1!
b100 %
1'
b100 +
#902660000000
0!
0'
#902670000000
1!
b101 %
1'
b101 +
#902680000000
0!
0'
#902690000000
1!
0$
b110 %
1'
0*
b110 +
#902700000000
0!
0'
#902710000000
1!
b111 %
1'
b111 +
#902720000000
0!
0'
#902730000000
1!
b1000 %
1'
b1000 +
#902740000000
0!
0'
#902750000000
1!
b1001 %
1'
b1001 +
#902760000000
0!
0'
#902770000000
1!
b0 %
1'
b0 +
#902780000000
1"
1(
#902790000000
0!
0"
b100 &
0'
0(
b100 ,
#902800000000
1!
1$
b1 %
1'
1*
b1 +
#902810000000
0!
0'
#902820000000
1!
b10 %
1'
b10 +
#902830000000
0!
0'
#902840000000
1!
b11 %
1'
b11 +
#902850000000
0!
0'
#902860000000
1!
b100 %
1'
b100 +
#902870000000
0!
0'
#902880000000
1!
b101 %
1'
b101 +
#902890000000
0!
0'
#902900000000
1!
b110 %
1'
b110 +
#902910000000
0!
0'
#902920000000
1!
b111 %
1'
b111 +
#902930000000
0!
0'
#902940000000
1!
0$
b1000 %
1'
0*
b1000 +
#902950000000
0!
0'
#902960000000
1!
b1001 %
1'
b1001 +
#902970000000
0!
0'
#902980000000
1!
b0 %
1'
b0 +
#902990000000
0!
0'
#903000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#903010000000
0!
0'
#903020000000
1!
b10 %
1'
b10 +
#903030000000
0!
0'
#903040000000
1!
b11 %
1'
b11 +
#903050000000
0!
0'
#903060000000
1!
b100 %
1'
b100 +
#903070000000
0!
0'
#903080000000
1!
b101 %
1'
b101 +
#903090000000
0!
0'
#903100000000
1!
0$
b110 %
1'
0*
b110 +
#903110000000
0!
0'
#903120000000
1!
b111 %
1'
b111 +
#903130000000
0!
0'
#903140000000
1!
b1000 %
1'
b1000 +
#903150000000
0!
0'
#903160000000
1!
b1001 %
1'
b1001 +
#903170000000
0!
0'
#903180000000
1!
b0 %
1'
b0 +
#903190000000
0!
0'
#903200000000
1!
1$
b1 %
1'
1*
b1 +
#903210000000
1"
1(
#903220000000
0!
0"
b100 &
0'
0(
b100 ,
#903230000000
1!
b10 %
1'
b10 +
#903240000000
0!
0'
#903250000000
1!
b11 %
1'
b11 +
#903260000000
0!
0'
#903270000000
1!
b100 %
1'
b100 +
#903280000000
0!
0'
#903290000000
1!
b101 %
1'
b101 +
#903300000000
0!
0'
#903310000000
1!
b110 %
1'
b110 +
#903320000000
0!
0'
#903330000000
1!
b111 %
1'
b111 +
#903340000000
0!
0'
#903350000000
1!
0$
b1000 %
1'
0*
b1000 +
#903360000000
0!
0'
#903370000000
1!
b1001 %
1'
b1001 +
#903380000000
0!
0'
#903390000000
1!
b0 %
1'
b0 +
#903400000000
0!
0'
#903410000000
1!
1$
b1 %
1'
1*
b1 +
#903420000000
0!
0'
#903430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#903440000000
0!
0'
#903450000000
1!
b11 %
1'
b11 +
#903460000000
0!
0'
#903470000000
1!
b100 %
1'
b100 +
#903480000000
0!
0'
#903490000000
1!
b101 %
1'
b101 +
#903500000000
0!
0'
#903510000000
1!
0$
b110 %
1'
0*
b110 +
#903520000000
0!
0'
#903530000000
1!
b111 %
1'
b111 +
#903540000000
0!
0'
#903550000000
1!
b1000 %
1'
b1000 +
#903560000000
0!
0'
#903570000000
1!
b1001 %
1'
b1001 +
#903580000000
0!
0'
#903590000000
1!
b0 %
1'
b0 +
#903600000000
0!
0'
#903610000000
1!
1$
b1 %
1'
1*
b1 +
#903620000000
0!
0'
#903630000000
1!
b10 %
1'
b10 +
#903640000000
1"
1(
#903650000000
0!
0"
b100 &
0'
0(
b100 ,
#903660000000
1!
b11 %
1'
b11 +
#903670000000
0!
0'
#903680000000
1!
b100 %
1'
b100 +
#903690000000
0!
0'
#903700000000
1!
b101 %
1'
b101 +
#903710000000
0!
0'
#903720000000
1!
b110 %
1'
b110 +
#903730000000
0!
0'
#903740000000
1!
b111 %
1'
b111 +
#903750000000
0!
0'
#903760000000
1!
0$
b1000 %
1'
0*
b1000 +
#903770000000
0!
0'
#903780000000
1!
b1001 %
1'
b1001 +
#903790000000
0!
0'
#903800000000
1!
b0 %
1'
b0 +
#903810000000
0!
0'
#903820000000
1!
1$
b1 %
1'
1*
b1 +
#903830000000
0!
0'
#903840000000
1!
b10 %
1'
b10 +
#903850000000
0!
0'
#903860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#903870000000
0!
0'
#903880000000
1!
b100 %
1'
b100 +
#903890000000
0!
0'
#903900000000
1!
b101 %
1'
b101 +
#903910000000
0!
0'
#903920000000
1!
0$
b110 %
1'
0*
b110 +
#903930000000
0!
0'
#903940000000
1!
b111 %
1'
b111 +
#903950000000
0!
0'
#903960000000
1!
b1000 %
1'
b1000 +
#903970000000
0!
0'
#903980000000
1!
b1001 %
1'
b1001 +
#903990000000
0!
0'
#904000000000
1!
b0 %
1'
b0 +
#904010000000
0!
0'
#904020000000
1!
1$
b1 %
1'
1*
b1 +
#904030000000
0!
0'
#904040000000
1!
b10 %
1'
b10 +
#904050000000
0!
0'
#904060000000
1!
b11 %
1'
b11 +
#904070000000
1"
1(
#904080000000
0!
0"
b100 &
0'
0(
b100 ,
#904090000000
1!
b100 %
1'
b100 +
#904100000000
0!
0'
#904110000000
1!
b101 %
1'
b101 +
#904120000000
0!
0'
#904130000000
1!
b110 %
1'
b110 +
#904140000000
0!
0'
#904150000000
1!
b111 %
1'
b111 +
#904160000000
0!
0'
#904170000000
1!
0$
b1000 %
1'
0*
b1000 +
#904180000000
0!
0'
#904190000000
1!
b1001 %
1'
b1001 +
#904200000000
0!
0'
#904210000000
1!
b0 %
1'
b0 +
#904220000000
0!
0'
#904230000000
1!
1$
b1 %
1'
1*
b1 +
#904240000000
0!
0'
#904250000000
1!
b10 %
1'
b10 +
#904260000000
0!
0'
#904270000000
1!
b11 %
1'
b11 +
#904280000000
0!
0'
#904290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#904300000000
0!
0'
#904310000000
1!
b101 %
1'
b101 +
#904320000000
0!
0'
#904330000000
1!
0$
b110 %
1'
0*
b110 +
#904340000000
0!
0'
#904350000000
1!
b111 %
1'
b111 +
#904360000000
0!
0'
#904370000000
1!
b1000 %
1'
b1000 +
#904380000000
0!
0'
#904390000000
1!
b1001 %
1'
b1001 +
#904400000000
0!
0'
#904410000000
1!
b0 %
1'
b0 +
#904420000000
0!
0'
#904430000000
1!
1$
b1 %
1'
1*
b1 +
#904440000000
0!
0'
#904450000000
1!
b10 %
1'
b10 +
#904460000000
0!
0'
#904470000000
1!
b11 %
1'
b11 +
#904480000000
0!
0'
#904490000000
1!
b100 %
1'
b100 +
#904500000000
1"
1(
#904510000000
0!
0"
b100 &
0'
0(
b100 ,
#904520000000
1!
b101 %
1'
b101 +
#904530000000
0!
0'
#904540000000
1!
b110 %
1'
b110 +
#904550000000
0!
0'
#904560000000
1!
b111 %
1'
b111 +
#904570000000
0!
0'
#904580000000
1!
0$
b1000 %
1'
0*
b1000 +
#904590000000
0!
0'
#904600000000
1!
b1001 %
1'
b1001 +
#904610000000
0!
0'
#904620000000
1!
b0 %
1'
b0 +
#904630000000
0!
0'
#904640000000
1!
1$
b1 %
1'
1*
b1 +
#904650000000
0!
0'
#904660000000
1!
b10 %
1'
b10 +
#904670000000
0!
0'
#904680000000
1!
b11 %
1'
b11 +
#904690000000
0!
0'
#904700000000
1!
b100 %
1'
b100 +
#904710000000
0!
0'
#904720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#904730000000
0!
0'
#904740000000
1!
0$
b110 %
1'
0*
b110 +
#904750000000
0!
0'
#904760000000
1!
b111 %
1'
b111 +
#904770000000
0!
0'
#904780000000
1!
b1000 %
1'
b1000 +
#904790000000
0!
0'
#904800000000
1!
b1001 %
1'
b1001 +
#904810000000
0!
0'
#904820000000
1!
b0 %
1'
b0 +
#904830000000
0!
0'
#904840000000
1!
1$
b1 %
1'
1*
b1 +
#904850000000
0!
0'
#904860000000
1!
b10 %
1'
b10 +
#904870000000
0!
0'
#904880000000
1!
b11 %
1'
b11 +
#904890000000
0!
0'
#904900000000
1!
b100 %
1'
b100 +
#904910000000
0!
0'
#904920000000
1!
b101 %
1'
b101 +
#904930000000
1"
1(
#904940000000
0!
0"
b100 &
0'
0(
b100 ,
#904950000000
1!
b110 %
1'
b110 +
#904960000000
0!
0'
#904970000000
1!
b111 %
1'
b111 +
#904980000000
0!
0'
#904990000000
1!
0$
b1000 %
1'
0*
b1000 +
#905000000000
0!
0'
#905010000000
1!
b1001 %
1'
b1001 +
#905020000000
0!
0'
#905030000000
1!
b0 %
1'
b0 +
#905040000000
0!
0'
#905050000000
1!
1$
b1 %
1'
1*
b1 +
#905060000000
0!
0'
#905070000000
1!
b10 %
1'
b10 +
#905080000000
0!
0'
#905090000000
1!
b11 %
1'
b11 +
#905100000000
0!
0'
#905110000000
1!
b100 %
1'
b100 +
#905120000000
0!
0'
#905130000000
1!
b101 %
1'
b101 +
#905140000000
0!
0'
#905150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#905160000000
0!
0'
#905170000000
1!
b111 %
1'
b111 +
#905180000000
0!
0'
#905190000000
1!
b1000 %
1'
b1000 +
#905200000000
0!
0'
#905210000000
1!
b1001 %
1'
b1001 +
#905220000000
0!
0'
#905230000000
1!
b0 %
1'
b0 +
#905240000000
0!
0'
#905250000000
1!
1$
b1 %
1'
1*
b1 +
#905260000000
0!
0'
#905270000000
1!
b10 %
1'
b10 +
#905280000000
0!
0'
#905290000000
1!
b11 %
1'
b11 +
#905300000000
0!
0'
#905310000000
1!
b100 %
1'
b100 +
#905320000000
0!
0'
#905330000000
1!
b101 %
1'
b101 +
#905340000000
0!
0'
#905350000000
1!
0$
b110 %
1'
0*
b110 +
#905360000000
1"
1(
#905370000000
0!
0"
b100 &
0'
0(
b100 ,
#905380000000
1!
1$
b111 %
1'
1*
b111 +
#905390000000
0!
0'
#905400000000
1!
0$
b1000 %
1'
0*
b1000 +
#905410000000
0!
0'
#905420000000
1!
b1001 %
1'
b1001 +
#905430000000
0!
0'
#905440000000
1!
b0 %
1'
b0 +
#905450000000
0!
0'
#905460000000
1!
1$
b1 %
1'
1*
b1 +
#905470000000
0!
0'
#905480000000
1!
b10 %
1'
b10 +
#905490000000
0!
0'
#905500000000
1!
b11 %
1'
b11 +
#905510000000
0!
0'
#905520000000
1!
b100 %
1'
b100 +
#905530000000
0!
0'
#905540000000
1!
b101 %
1'
b101 +
#905550000000
0!
0'
#905560000000
1!
b110 %
1'
b110 +
#905570000000
0!
0'
#905580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#905590000000
0!
0'
#905600000000
1!
b1000 %
1'
b1000 +
#905610000000
0!
0'
#905620000000
1!
b1001 %
1'
b1001 +
#905630000000
0!
0'
#905640000000
1!
b0 %
1'
b0 +
#905650000000
0!
0'
#905660000000
1!
1$
b1 %
1'
1*
b1 +
#905670000000
0!
0'
#905680000000
1!
b10 %
1'
b10 +
#905690000000
0!
0'
#905700000000
1!
b11 %
1'
b11 +
#905710000000
0!
0'
#905720000000
1!
b100 %
1'
b100 +
#905730000000
0!
0'
#905740000000
1!
b101 %
1'
b101 +
#905750000000
0!
0'
#905760000000
1!
0$
b110 %
1'
0*
b110 +
#905770000000
0!
0'
#905780000000
1!
b111 %
1'
b111 +
#905790000000
1"
1(
#905800000000
0!
0"
b100 &
0'
0(
b100 ,
#905810000000
1!
b1000 %
1'
b1000 +
#905820000000
0!
0'
#905830000000
1!
b1001 %
1'
b1001 +
#905840000000
0!
0'
#905850000000
1!
b0 %
1'
b0 +
#905860000000
0!
0'
#905870000000
1!
1$
b1 %
1'
1*
b1 +
#905880000000
0!
0'
#905890000000
1!
b10 %
1'
b10 +
#905900000000
0!
0'
#905910000000
1!
b11 %
1'
b11 +
#905920000000
0!
0'
#905930000000
1!
b100 %
1'
b100 +
#905940000000
0!
0'
#905950000000
1!
b101 %
1'
b101 +
#905960000000
0!
0'
#905970000000
1!
b110 %
1'
b110 +
#905980000000
0!
0'
#905990000000
1!
b111 %
1'
b111 +
#906000000000
0!
0'
#906010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#906020000000
0!
0'
#906030000000
1!
b1001 %
1'
b1001 +
#906040000000
0!
0'
#906050000000
1!
b0 %
1'
b0 +
#906060000000
0!
0'
#906070000000
1!
1$
b1 %
1'
1*
b1 +
#906080000000
0!
0'
#906090000000
1!
b10 %
1'
b10 +
#906100000000
0!
0'
#906110000000
1!
b11 %
1'
b11 +
#906120000000
0!
0'
#906130000000
1!
b100 %
1'
b100 +
#906140000000
0!
0'
#906150000000
1!
b101 %
1'
b101 +
#906160000000
0!
0'
#906170000000
1!
0$
b110 %
1'
0*
b110 +
#906180000000
0!
0'
#906190000000
1!
b111 %
1'
b111 +
#906200000000
0!
0'
#906210000000
1!
b1000 %
1'
b1000 +
#906220000000
1"
1(
#906230000000
0!
0"
b100 &
0'
0(
b100 ,
#906240000000
1!
b1001 %
1'
b1001 +
#906250000000
0!
0'
#906260000000
1!
b0 %
1'
b0 +
#906270000000
0!
0'
#906280000000
1!
1$
b1 %
1'
1*
b1 +
#906290000000
0!
0'
#906300000000
1!
b10 %
1'
b10 +
#906310000000
0!
0'
#906320000000
1!
b11 %
1'
b11 +
#906330000000
0!
0'
#906340000000
1!
b100 %
1'
b100 +
#906350000000
0!
0'
#906360000000
1!
b101 %
1'
b101 +
#906370000000
0!
0'
#906380000000
1!
b110 %
1'
b110 +
#906390000000
0!
0'
#906400000000
1!
b111 %
1'
b111 +
#906410000000
0!
0'
#906420000000
1!
0$
b1000 %
1'
0*
b1000 +
#906430000000
0!
0'
#906440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#906450000000
0!
0'
#906460000000
1!
b0 %
1'
b0 +
#906470000000
0!
0'
#906480000000
1!
1$
b1 %
1'
1*
b1 +
#906490000000
0!
0'
#906500000000
1!
b10 %
1'
b10 +
#906510000000
0!
0'
#906520000000
1!
b11 %
1'
b11 +
#906530000000
0!
0'
#906540000000
1!
b100 %
1'
b100 +
#906550000000
0!
0'
#906560000000
1!
b101 %
1'
b101 +
#906570000000
0!
0'
#906580000000
1!
0$
b110 %
1'
0*
b110 +
#906590000000
0!
0'
#906600000000
1!
b111 %
1'
b111 +
#906610000000
0!
0'
#906620000000
1!
b1000 %
1'
b1000 +
#906630000000
0!
0'
#906640000000
1!
b1001 %
1'
b1001 +
#906650000000
1"
1(
#906660000000
0!
0"
b100 &
0'
0(
b100 ,
#906670000000
1!
b0 %
1'
b0 +
#906680000000
0!
0'
#906690000000
1!
1$
b1 %
1'
1*
b1 +
#906700000000
0!
0'
#906710000000
1!
b10 %
1'
b10 +
#906720000000
0!
0'
#906730000000
1!
b11 %
1'
b11 +
#906740000000
0!
0'
#906750000000
1!
b100 %
1'
b100 +
#906760000000
0!
0'
#906770000000
1!
b101 %
1'
b101 +
#906780000000
0!
0'
#906790000000
1!
b110 %
1'
b110 +
#906800000000
0!
0'
#906810000000
1!
b111 %
1'
b111 +
#906820000000
0!
0'
#906830000000
1!
0$
b1000 %
1'
0*
b1000 +
#906840000000
0!
0'
#906850000000
1!
b1001 %
1'
b1001 +
#906860000000
0!
0'
#906870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#906880000000
0!
0'
#906890000000
1!
1$
b1 %
1'
1*
b1 +
#906900000000
0!
0'
#906910000000
1!
b10 %
1'
b10 +
#906920000000
0!
0'
#906930000000
1!
b11 %
1'
b11 +
#906940000000
0!
0'
#906950000000
1!
b100 %
1'
b100 +
#906960000000
0!
0'
#906970000000
1!
b101 %
1'
b101 +
#906980000000
0!
0'
#906990000000
1!
0$
b110 %
1'
0*
b110 +
#907000000000
0!
0'
#907010000000
1!
b111 %
1'
b111 +
#907020000000
0!
0'
#907030000000
1!
b1000 %
1'
b1000 +
#907040000000
0!
0'
#907050000000
1!
b1001 %
1'
b1001 +
#907060000000
0!
0'
#907070000000
1!
b0 %
1'
b0 +
#907080000000
1"
1(
#907090000000
0!
0"
b100 &
0'
0(
b100 ,
#907100000000
1!
1$
b1 %
1'
1*
b1 +
#907110000000
0!
0'
#907120000000
1!
b10 %
1'
b10 +
#907130000000
0!
0'
#907140000000
1!
b11 %
1'
b11 +
#907150000000
0!
0'
#907160000000
1!
b100 %
1'
b100 +
#907170000000
0!
0'
#907180000000
1!
b101 %
1'
b101 +
#907190000000
0!
0'
#907200000000
1!
b110 %
1'
b110 +
#907210000000
0!
0'
#907220000000
1!
b111 %
1'
b111 +
#907230000000
0!
0'
#907240000000
1!
0$
b1000 %
1'
0*
b1000 +
#907250000000
0!
0'
#907260000000
1!
b1001 %
1'
b1001 +
#907270000000
0!
0'
#907280000000
1!
b0 %
1'
b0 +
#907290000000
0!
0'
#907300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#907310000000
0!
0'
#907320000000
1!
b10 %
1'
b10 +
#907330000000
0!
0'
#907340000000
1!
b11 %
1'
b11 +
#907350000000
0!
0'
#907360000000
1!
b100 %
1'
b100 +
#907370000000
0!
0'
#907380000000
1!
b101 %
1'
b101 +
#907390000000
0!
0'
#907400000000
1!
0$
b110 %
1'
0*
b110 +
#907410000000
0!
0'
#907420000000
1!
b111 %
1'
b111 +
#907430000000
0!
0'
#907440000000
1!
b1000 %
1'
b1000 +
#907450000000
0!
0'
#907460000000
1!
b1001 %
1'
b1001 +
#907470000000
0!
0'
#907480000000
1!
b0 %
1'
b0 +
#907490000000
0!
0'
#907500000000
1!
1$
b1 %
1'
1*
b1 +
#907510000000
1"
1(
#907520000000
0!
0"
b100 &
0'
0(
b100 ,
#907530000000
1!
b10 %
1'
b10 +
#907540000000
0!
0'
#907550000000
1!
b11 %
1'
b11 +
#907560000000
0!
0'
#907570000000
1!
b100 %
1'
b100 +
#907580000000
0!
0'
#907590000000
1!
b101 %
1'
b101 +
#907600000000
0!
0'
#907610000000
1!
b110 %
1'
b110 +
#907620000000
0!
0'
#907630000000
1!
b111 %
1'
b111 +
#907640000000
0!
0'
#907650000000
1!
0$
b1000 %
1'
0*
b1000 +
#907660000000
0!
0'
#907670000000
1!
b1001 %
1'
b1001 +
#907680000000
0!
0'
#907690000000
1!
b0 %
1'
b0 +
#907700000000
0!
0'
#907710000000
1!
1$
b1 %
1'
1*
b1 +
#907720000000
0!
0'
#907730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#907740000000
0!
0'
#907750000000
1!
b11 %
1'
b11 +
#907760000000
0!
0'
#907770000000
1!
b100 %
1'
b100 +
#907780000000
0!
0'
#907790000000
1!
b101 %
1'
b101 +
#907800000000
0!
0'
#907810000000
1!
0$
b110 %
1'
0*
b110 +
#907820000000
0!
0'
#907830000000
1!
b111 %
1'
b111 +
#907840000000
0!
0'
#907850000000
1!
b1000 %
1'
b1000 +
#907860000000
0!
0'
#907870000000
1!
b1001 %
1'
b1001 +
#907880000000
0!
0'
#907890000000
1!
b0 %
1'
b0 +
#907900000000
0!
0'
#907910000000
1!
1$
b1 %
1'
1*
b1 +
#907920000000
0!
0'
#907930000000
1!
b10 %
1'
b10 +
#907940000000
1"
1(
#907950000000
0!
0"
b100 &
0'
0(
b100 ,
#907960000000
1!
b11 %
1'
b11 +
#907970000000
0!
0'
#907980000000
1!
b100 %
1'
b100 +
#907990000000
0!
0'
#908000000000
1!
b101 %
1'
b101 +
#908010000000
0!
0'
#908020000000
1!
b110 %
1'
b110 +
#908030000000
0!
0'
#908040000000
1!
b111 %
1'
b111 +
#908050000000
0!
0'
#908060000000
1!
0$
b1000 %
1'
0*
b1000 +
#908070000000
0!
0'
#908080000000
1!
b1001 %
1'
b1001 +
#908090000000
0!
0'
#908100000000
1!
b0 %
1'
b0 +
#908110000000
0!
0'
#908120000000
1!
1$
b1 %
1'
1*
b1 +
#908130000000
0!
0'
#908140000000
1!
b10 %
1'
b10 +
#908150000000
0!
0'
#908160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#908170000000
0!
0'
#908180000000
1!
b100 %
1'
b100 +
#908190000000
0!
0'
#908200000000
1!
b101 %
1'
b101 +
#908210000000
0!
0'
#908220000000
1!
0$
b110 %
1'
0*
b110 +
#908230000000
0!
0'
#908240000000
1!
b111 %
1'
b111 +
#908250000000
0!
0'
#908260000000
1!
b1000 %
1'
b1000 +
#908270000000
0!
0'
#908280000000
1!
b1001 %
1'
b1001 +
#908290000000
0!
0'
#908300000000
1!
b0 %
1'
b0 +
#908310000000
0!
0'
#908320000000
1!
1$
b1 %
1'
1*
b1 +
#908330000000
0!
0'
#908340000000
1!
b10 %
1'
b10 +
#908350000000
0!
0'
#908360000000
1!
b11 %
1'
b11 +
#908370000000
1"
1(
#908380000000
0!
0"
b100 &
0'
0(
b100 ,
#908390000000
1!
b100 %
1'
b100 +
#908400000000
0!
0'
#908410000000
1!
b101 %
1'
b101 +
#908420000000
0!
0'
#908430000000
1!
b110 %
1'
b110 +
#908440000000
0!
0'
#908450000000
1!
b111 %
1'
b111 +
#908460000000
0!
0'
#908470000000
1!
0$
b1000 %
1'
0*
b1000 +
#908480000000
0!
0'
#908490000000
1!
b1001 %
1'
b1001 +
#908500000000
0!
0'
#908510000000
1!
b0 %
1'
b0 +
#908520000000
0!
0'
#908530000000
1!
1$
b1 %
1'
1*
b1 +
#908540000000
0!
0'
#908550000000
1!
b10 %
1'
b10 +
#908560000000
0!
0'
#908570000000
1!
b11 %
1'
b11 +
#908580000000
0!
0'
#908590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#908600000000
0!
0'
#908610000000
1!
b101 %
1'
b101 +
#908620000000
0!
0'
#908630000000
1!
0$
b110 %
1'
0*
b110 +
#908640000000
0!
0'
#908650000000
1!
b111 %
1'
b111 +
#908660000000
0!
0'
#908670000000
1!
b1000 %
1'
b1000 +
#908680000000
0!
0'
#908690000000
1!
b1001 %
1'
b1001 +
#908700000000
0!
0'
#908710000000
1!
b0 %
1'
b0 +
#908720000000
0!
0'
#908730000000
1!
1$
b1 %
1'
1*
b1 +
#908740000000
0!
0'
#908750000000
1!
b10 %
1'
b10 +
#908760000000
0!
0'
#908770000000
1!
b11 %
1'
b11 +
#908780000000
0!
0'
#908790000000
1!
b100 %
1'
b100 +
#908800000000
1"
1(
#908810000000
0!
0"
b100 &
0'
0(
b100 ,
#908820000000
1!
b101 %
1'
b101 +
#908830000000
0!
0'
#908840000000
1!
b110 %
1'
b110 +
#908850000000
0!
0'
#908860000000
1!
b111 %
1'
b111 +
#908870000000
0!
0'
#908880000000
1!
0$
b1000 %
1'
0*
b1000 +
#908890000000
0!
0'
#908900000000
1!
b1001 %
1'
b1001 +
#908910000000
0!
0'
#908920000000
1!
b0 %
1'
b0 +
#908930000000
0!
0'
#908940000000
1!
1$
b1 %
1'
1*
b1 +
#908950000000
0!
0'
#908960000000
1!
b10 %
1'
b10 +
#908970000000
0!
0'
#908980000000
1!
b11 %
1'
b11 +
#908990000000
0!
0'
#909000000000
1!
b100 %
1'
b100 +
#909010000000
0!
0'
#909020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#909030000000
0!
0'
#909040000000
1!
0$
b110 %
1'
0*
b110 +
#909050000000
0!
0'
#909060000000
1!
b111 %
1'
b111 +
#909070000000
0!
0'
#909080000000
1!
b1000 %
1'
b1000 +
#909090000000
0!
0'
#909100000000
1!
b1001 %
1'
b1001 +
#909110000000
0!
0'
#909120000000
1!
b0 %
1'
b0 +
#909130000000
0!
0'
#909140000000
1!
1$
b1 %
1'
1*
b1 +
#909150000000
0!
0'
#909160000000
1!
b10 %
1'
b10 +
#909170000000
0!
0'
#909180000000
1!
b11 %
1'
b11 +
#909190000000
0!
0'
#909200000000
1!
b100 %
1'
b100 +
#909210000000
0!
0'
#909220000000
1!
b101 %
1'
b101 +
#909230000000
1"
1(
#909240000000
0!
0"
b100 &
0'
0(
b100 ,
#909250000000
1!
b110 %
1'
b110 +
#909260000000
0!
0'
#909270000000
1!
b111 %
1'
b111 +
#909280000000
0!
0'
#909290000000
1!
0$
b1000 %
1'
0*
b1000 +
#909300000000
0!
0'
#909310000000
1!
b1001 %
1'
b1001 +
#909320000000
0!
0'
#909330000000
1!
b0 %
1'
b0 +
#909340000000
0!
0'
#909350000000
1!
1$
b1 %
1'
1*
b1 +
#909360000000
0!
0'
#909370000000
1!
b10 %
1'
b10 +
#909380000000
0!
0'
#909390000000
1!
b11 %
1'
b11 +
#909400000000
0!
0'
#909410000000
1!
b100 %
1'
b100 +
#909420000000
0!
0'
#909430000000
1!
b101 %
1'
b101 +
#909440000000
0!
0'
#909450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#909460000000
0!
0'
#909470000000
1!
b111 %
1'
b111 +
#909480000000
0!
0'
#909490000000
1!
b1000 %
1'
b1000 +
#909500000000
0!
0'
#909510000000
1!
b1001 %
1'
b1001 +
#909520000000
0!
0'
#909530000000
1!
b0 %
1'
b0 +
#909540000000
0!
0'
#909550000000
1!
1$
b1 %
1'
1*
b1 +
#909560000000
0!
0'
#909570000000
1!
b10 %
1'
b10 +
#909580000000
0!
0'
#909590000000
1!
b11 %
1'
b11 +
#909600000000
0!
0'
#909610000000
1!
b100 %
1'
b100 +
#909620000000
0!
0'
#909630000000
1!
b101 %
1'
b101 +
#909640000000
0!
0'
#909650000000
1!
0$
b110 %
1'
0*
b110 +
#909660000000
1"
1(
#909670000000
0!
0"
b100 &
0'
0(
b100 ,
#909680000000
1!
1$
b111 %
1'
1*
b111 +
#909690000000
0!
0'
#909700000000
1!
0$
b1000 %
1'
0*
b1000 +
#909710000000
0!
0'
#909720000000
1!
b1001 %
1'
b1001 +
#909730000000
0!
0'
#909740000000
1!
b0 %
1'
b0 +
#909750000000
0!
0'
#909760000000
1!
1$
b1 %
1'
1*
b1 +
#909770000000
0!
0'
#909780000000
1!
b10 %
1'
b10 +
#909790000000
0!
0'
#909800000000
1!
b11 %
1'
b11 +
#909810000000
0!
0'
#909820000000
1!
b100 %
1'
b100 +
#909830000000
0!
0'
#909840000000
1!
b101 %
1'
b101 +
#909850000000
0!
0'
#909860000000
1!
b110 %
1'
b110 +
#909870000000
0!
0'
#909880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#909890000000
0!
0'
#909900000000
1!
b1000 %
1'
b1000 +
#909910000000
0!
0'
#909920000000
1!
b1001 %
1'
b1001 +
#909930000000
0!
0'
#909940000000
1!
b0 %
1'
b0 +
#909950000000
0!
0'
#909960000000
1!
1$
b1 %
1'
1*
b1 +
#909970000000
0!
0'
#909980000000
1!
b10 %
1'
b10 +
#909990000000
0!
0'
#910000000000
1!
b11 %
1'
b11 +
#910010000000
0!
0'
#910020000000
1!
b100 %
1'
b100 +
#910030000000
0!
0'
#910040000000
1!
b101 %
1'
b101 +
#910050000000
0!
0'
#910060000000
1!
0$
b110 %
1'
0*
b110 +
#910070000000
0!
0'
#910080000000
1!
b111 %
1'
b111 +
#910090000000
1"
1(
#910100000000
0!
0"
b100 &
0'
0(
b100 ,
#910110000000
1!
b1000 %
1'
b1000 +
#910120000000
0!
0'
#910130000000
1!
b1001 %
1'
b1001 +
#910140000000
0!
0'
#910150000000
1!
b0 %
1'
b0 +
#910160000000
0!
0'
#910170000000
1!
1$
b1 %
1'
1*
b1 +
#910180000000
0!
0'
#910190000000
1!
b10 %
1'
b10 +
#910200000000
0!
0'
#910210000000
1!
b11 %
1'
b11 +
#910220000000
0!
0'
#910230000000
1!
b100 %
1'
b100 +
#910240000000
0!
0'
#910250000000
1!
b101 %
1'
b101 +
#910260000000
0!
0'
#910270000000
1!
b110 %
1'
b110 +
#910280000000
0!
0'
#910290000000
1!
b111 %
1'
b111 +
#910300000000
0!
0'
#910310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#910320000000
0!
0'
#910330000000
1!
b1001 %
1'
b1001 +
#910340000000
0!
0'
#910350000000
1!
b0 %
1'
b0 +
#910360000000
0!
0'
#910370000000
1!
1$
b1 %
1'
1*
b1 +
#910380000000
0!
0'
#910390000000
1!
b10 %
1'
b10 +
#910400000000
0!
0'
#910410000000
1!
b11 %
1'
b11 +
#910420000000
0!
0'
#910430000000
1!
b100 %
1'
b100 +
#910440000000
0!
0'
#910450000000
1!
b101 %
1'
b101 +
#910460000000
0!
0'
#910470000000
1!
0$
b110 %
1'
0*
b110 +
#910480000000
0!
0'
#910490000000
1!
b111 %
1'
b111 +
#910500000000
0!
0'
#910510000000
1!
b1000 %
1'
b1000 +
#910520000000
1"
1(
#910530000000
0!
0"
b100 &
0'
0(
b100 ,
#910540000000
1!
b1001 %
1'
b1001 +
#910550000000
0!
0'
#910560000000
1!
b0 %
1'
b0 +
#910570000000
0!
0'
#910580000000
1!
1$
b1 %
1'
1*
b1 +
#910590000000
0!
0'
#910600000000
1!
b10 %
1'
b10 +
#910610000000
0!
0'
#910620000000
1!
b11 %
1'
b11 +
#910630000000
0!
0'
#910640000000
1!
b100 %
1'
b100 +
#910650000000
0!
0'
#910660000000
1!
b101 %
1'
b101 +
#910670000000
0!
0'
#910680000000
1!
b110 %
1'
b110 +
#910690000000
0!
0'
#910700000000
1!
b111 %
1'
b111 +
#910710000000
0!
0'
#910720000000
1!
0$
b1000 %
1'
0*
b1000 +
#910730000000
0!
0'
#910740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#910750000000
0!
0'
#910760000000
1!
b0 %
1'
b0 +
#910770000000
0!
0'
#910780000000
1!
1$
b1 %
1'
1*
b1 +
#910790000000
0!
0'
#910800000000
1!
b10 %
1'
b10 +
#910810000000
0!
0'
#910820000000
1!
b11 %
1'
b11 +
#910830000000
0!
0'
#910840000000
1!
b100 %
1'
b100 +
#910850000000
0!
0'
#910860000000
1!
b101 %
1'
b101 +
#910870000000
0!
0'
#910880000000
1!
0$
b110 %
1'
0*
b110 +
#910890000000
0!
0'
#910900000000
1!
b111 %
1'
b111 +
#910910000000
0!
0'
#910920000000
1!
b1000 %
1'
b1000 +
#910930000000
0!
0'
#910940000000
1!
b1001 %
1'
b1001 +
#910950000000
1"
1(
#910960000000
0!
0"
b100 &
0'
0(
b100 ,
#910970000000
1!
b0 %
1'
b0 +
#910980000000
0!
0'
#910990000000
1!
1$
b1 %
1'
1*
b1 +
#911000000000
0!
0'
#911010000000
1!
b10 %
1'
b10 +
#911020000000
0!
0'
#911030000000
1!
b11 %
1'
b11 +
#911040000000
0!
0'
#911050000000
1!
b100 %
1'
b100 +
#911060000000
0!
0'
#911070000000
1!
b101 %
1'
b101 +
#911080000000
0!
0'
#911090000000
1!
b110 %
1'
b110 +
#911100000000
0!
0'
#911110000000
1!
b111 %
1'
b111 +
#911120000000
0!
0'
#911130000000
1!
0$
b1000 %
1'
0*
b1000 +
#911140000000
0!
0'
#911150000000
1!
b1001 %
1'
b1001 +
#911160000000
0!
0'
#911170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#911180000000
0!
0'
#911190000000
1!
1$
b1 %
1'
1*
b1 +
#911200000000
0!
0'
#911210000000
1!
b10 %
1'
b10 +
#911220000000
0!
0'
#911230000000
1!
b11 %
1'
b11 +
#911240000000
0!
0'
#911250000000
1!
b100 %
1'
b100 +
#911260000000
0!
0'
#911270000000
1!
b101 %
1'
b101 +
#911280000000
0!
0'
#911290000000
1!
0$
b110 %
1'
0*
b110 +
#911300000000
0!
0'
#911310000000
1!
b111 %
1'
b111 +
#911320000000
0!
0'
#911330000000
1!
b1000 %
1'
b1000 +
#911340000000
0!
0'
#911350000000
1!
b1001 %
1'
b1001 +
#911360000000
0!
0'
#911370000000
1!
b0 %
1'
b0 +
#911380000000
1"
1(
#911390000000
0!
0"
b100 &
0'
0(
b100 ,
#911400000000
1!
1$
b1 %
1'
1*
b1 +
#911410000000
0!
0'
#911420000000
1!
b10 %
1'
b10 +
#911430000000
0!
0'
#911440000000
1!
b11 %
1'
b11 +
#911450000000
0!
0'
#911460000000
1!
b100 %
1'
b100 +
#911470000000
0!
0'
#911480000000
1!
b101 %
1'
b101 +
#911490000000
0!
0'
#911500000000
1!
b110 %
1'
b110 +
#911510000000
0!
0'
#911520000000
1!
b111 %
1'
b111 +
#911530000000
0!
0'
#911540000000
1!
0$
b1000 %
1'
0*
b1000 +
#911550000000
0!
0'
#911560000000
1!
b1001 %
1'
b1001 +
#911570000000
0!
0'
#911580000000
1!
b0 %
1'
b0 +
#911590000000
0!
0'
#911600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#911610000000
0!
0'
#911620000000
1!
b10 %
1'
b10 +
#911630000000
0!
0'
#911640000000
1!
b11 %
1'
b11 +
#911650000000
0!
0'
#911660000000
1!
b100 %
1'
b100 +
#911670000000
0!
0'
#911680000000
1!
b101 %
1'
b101 +
#911690000000
0!
0'
#911700000000
1!
0$
b110 %
1'
0*
b110 +
#911710000000
0!
0'
#911720000000
1!
b111 %
1'
b111 +
#911730000000
0!
0'
#911740000000
1!
b1000 %
1'
b1000 +
#911750000000
0!
0'
#911760000000
1!
b1001 %
1'
b1001 +
#911770000000
0!
0'
#911780000000
1!
b0 %
1'
b0 +
#911790000000
0!
0'
#911800000000
1!
1$
b1 %
1'
1*
b1 +
#911810000000
1"
1(
#911820000000
0!
0"
b100 &
0'
0(
b100 ,
#911830000000
1!
b10 %
1'
b10 +
#911840000000
0!
0'
#911850000000
1!
b11 %
1'
b11 +
#911860000000
0!
0'
#911870000000
1!
b100 %
1'
b100 +
#911880000000
0!
0'
#911890000000
1!
b101 %
1'
b101 +
#911900000000
0!
0'
#911910000000
1!
b110 %
1'
b110 +
#911920000000
0!
0'
#911930000000
1!
b111 %
1'
b111 +
#911940000000
0!
0'
#911950000000
1!
0$
b1000 %
1'
0*
b1000 +
#911960000000
0!
0'
#911970000000
1!
b1001 %
1'
b1001 +
#911980000000
0!
0'
#911990000000
1!
b0 %
1'
b0 +
#912000000000
0!
0'
#912010000000
1!
1$
b1 %
1'
1*
b1 +
#912020000000
0!
0'
#912030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#912040000000
0!
0'
#912050000000
1!
b11 %
1'
b11 +
#912060000000
0!
0'
#912070000000
1!
b100 %
1'
b100 +
#912080000000
0!
0'
#912090000000
1!
b101 %
1'
b101 +
#912100000000
0!
0'
#912110000000
1!
0$
b110 %
1'
0*
b110 +
#912120000000
0!
0'
#912130000000
1!
b111 %
1'
b111 +
#912140000000
0!
0'
#912150000000
1!
b1000 %
1'
b1000 +
#912160000000
0!
0'
#912170000000
1!
b1001 %
1'
b1001 +
#912180000000
0!
0'
#912190000000
1!
b0 %
1'
b0 +
#912200000000
0!
0'
#912210000000
1!
1$
b1 %
1'
1*
b1 +
#912220000000
0!
0'
#912230000000
1!
b10 %
1'
b10 +
#912240000000
1"
1(
#912250000000
0!
0"
b100 &
0'
0(
b100 ,
#912260000000
1!
b11 %
1'
b11 +
#912270000000
0!
0'
#912280000000
1!
b100 %
1'
b100 +
#912290000000
0!
0'
#912300000000
1!
b101 %
1'
b101 +
#912310000000
0!
0'
#912320000000
1!
b110 %
1'
b110 +
#912330000000
0!
0'
#912340000000
1!
b111 %
1'
b111 +
#912350000000
0!
0'
#912360000000
1!
0$
b1000 %
1'
0*
b1000 +
#912370000000
0!
0'
#912380000000
1!
b1001 %
1'
b1001 +
#912390000000
0!
0'
#912400000000
1!
b0 %
1'
b0 +
#912410000000
0!
0'
#912420000000
1!
1$
b1 %
1'
1*
b1 +
#912430000000
0!
0'
#912440000000
1!
b10 %
1'
b10 +
#912450000000
0!
0'
#912460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#912470000000
0!
0'
#912480000000
1!
b100 %
1'
b100 +
#912490000000
0!
0'
#912500000000
1!
b101 %
1'
b101 +
#912510000000
0!
0'
#912520000000
1!
0$
b110 %
1'
0*
b110 +
#912530000000
0!
0'
#912540000000
1!
b111 %
1'
b111 +
#912550000000
0!
0'
#912560000000
1!
b1000 %
1'
b1000 +
#912570000000
0!
0'
#912580000000
1!
b1001 %
1'
b1001 +
#912590000000
0!
0'
#912600000000
1!
b0 %
1'
b0 +
#912610000000
0!
0'
#912620000000
1!
1$
b1 %
1'
1*
b1 +
#912630000000
0!
0'
#912640000000
1!
b10 %
1'
b10 +
#912650000000
0!
0'
#912660000000
1!
b11 %
1'
b11 +
#912670000000
1"
1(
#912680000000
0!
0"
b100 &
0'
0(
b100 ,
#912690000000
1!
b100 %
1'
b100 +
#912700000000
0!
0'
#912710000000
1!
b101 %
1'
b101 +
#912720000000
0!
0'
#912730000000
1!
b110 %
1'
b110 +
#912740000000
0!
0'
#912750000000
1!
b111 %
1'
b111 +
#912760000000
0!
0'
#912770000000
1!
0$
b1000 %
1'
0*
b1000 +
#912780000000
0!
0'
#912790000000
1!
b1001 %
1'
b1001 +
#912800000000
0!
0'
#912810000000
1!
b0 %
1'
b0 +
#912820000000
0!
0'
#912830000000
1!
1$
b1 %
1'
1*
b1 +
#912840000000
0!
0'
#912850000000
1!
b10 %
1'
b10 +
#912860000000
0!
0'
#912870000000
1!
b11 %
1'
b11 +
#912880000000
0!
0'
#912890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#912900000000
0!
0'
#912910000000
1!
b101 %
1'
b101 +
#912920000000
0!
0'
#912930000000
1!
0$
b110 %
1'
0*
b110 +
#912940000000
0!
0'
#912950000000
1!
b111 %
1'
b111 +
#912960000000
0!
0'
#912970000000
1!
b1000 %
1'
b1000 +
#912980000000
0!
0'
#912990000000
1!
b1001 %
1'
b1001 +
#913000000000
0!
0'
#913010000000
1!
b0 %
1'
b0 +
#913020000000
0!
0'
#913030000000
1!
1$
b1 %
1'
1*
b1 +
#913040000000
0!
0'
#913050000000
1!
b10 %
1'
b10 +
#913060000000
0!
0'
#913070000000
1!
b11 %
1'
b11 +
#913080000000
0!
0'
#913090000000
1!
b100 %
1'
b100 +
#913100000000
1"
1(
#913110000000
0!
0"
b100 &
0'
0(
b100 ,
#913120000000
1!
b101 %
1'
b101 +
#913130000000
0!
0'
#913140000000
1!
b110 %
1'
b110 +
#913150000000
0!
0'
#913160000000
1!
b111 %
1'
b111 +
#913170000000
0!
0'
#913180000000
1!
0$
b1000 %
1'
0*
b1000 +
#913190000000
0!
0'
#913200000000
1!
b1001 %
1'
b1001 +
#913210000000
0!
0'
#913220000000
1!
b0 %
1'
b0 +
#913230000000
0!
0'
#913240000000
1!
1$
b1 %
1'
1*
b1 +
#913250000000
0!
0'
#913260000000
1!
b10 %
1'
b10 +
#913270000000
0!
0'
#913280000000
1!
b11 %
1'
b11 +
#913290000000
0!
0'
#913300000000
1!
b100 %
1'
b100 +
#913310000000
0!
0'
#913320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#913330000000
0!
0'
#913340000000
1!
0$
b110 %
1'
0*
b110 +
#913350000000
0!
0'
#913360000000
1!
b111 %
1'
b111 +
#913370000000
0!
0'
#913380000000
1!
b1000 %
1'
b1000 +
#913390000000
0!
0'
#913400000000
1!
b1001 %
1'
b1001 +
#913410000000
0!
0'
#913420000000
1!
b0 %
1'
b0 +
#913430000000
0!
0'
#913440000000
1!
1$
b1 %
1'
1*
b1 +
#913450000000
0!
0'
#913460000000
1!
b10 %
1'
b10 +
#913470000000
0!
0'
#913480000000
1!
b11 %
1'
b11 +
#913490000000
0!
0'
#913500000000
1!
b100 %
1'
b100 +
#913510000000
0!
0'
#913520000000
1!
b101 %
1'
b101 +
#913530000000
1"
1(
#913540000000
0!
0"
b100 &
0'
0(
b100 ,
#913550000000
1!
b110 %
1'
b110 +
#913560000000
0!
0'
#913570000000
1!
b111 %
1'
b111 +
#913580000000
0!
0'
#913590000000
1!
0$
b1000 %
1'
0*
b1000 +
#913600000000
0!
0'
#913610000000
1!
b1001 %
1'
b1001 +
#913620000000
0!
0'
#913630000000
1!
b0 %
1'
b0 +
#913640000000
0!
0'
#913650000000
1!
1$
b1 %
1'
1*
b1 +
#913660000000
0!
0'
#913670000000
1!
b10 %
1'
b10 +
#913680000000
0!
0'
#913690000000
1!
b11 %
1'
b11 +
#913700000000
0!
0'
#913710000000
1!
b100 %
1'
b100 +
#913720000000
0!
0'
#913730000000
1!
b101 %
1'
b101 +
#913740000000
0!
0'
#913750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#913760000000
0!
0'
#913770000000
1!
b111 %
1'
b111 +
#913780000000
0!
0'
#913790000000
1!
b1000 %
1'
b1000 +
#913800000000
0!
0'
#913810000000
1!
b1001 %
1'
b1001 +
#913820000000
0!
0'
#913830000000
1!
b0 %
1'
b0 +
#913840000000
0!
0'
#913850000000
1!
1$
b1 %
1'
1*
b1 +
#913860000000
0!
0'
#913870000000
1!
b10 %
1'
b10 +
#913880000000
0!
0'
#913890000000
1!
b11 %
1'
b11 +
#913900000000
0!
0'
#913910000000
1!
b100 %
1'
b100 +
#913920000000
0!
0'
#913930000000
1!
b101 %
1'
b101 +
#913940000000
0!
0'
#913950000000
1!
0$
b110 %
1'
0*
b110 +
#913960000000
1"
1(
#913970000000
0!
0"
b100 &
0'
0(
b100 ,
#913980000000
1!
1$
b111 %
1'
1*
b111 +
#913990000000
0!
0'
#914000000000
1!
0$
b1000 %
1'
0*
b1000 +
#914010000000
0!
0'
#914020000000
1!
b1001 %
1'
b1001 +
#914030000000
0!
0'
#914040000000
1!
b0 %
1'
b0 +
#914050000000
0!
0'
#914060000000
1!
1$
b1 %
1'
1*
b1 +
#914070000000
0!
0'
#914080000000
1!
b10 %
1'
b10 +
#914090000000
0!
0'
#914100000000
1!
b11 %
1'
b11 +
#914110000000
0!
0'
#914120000000
1!
b100 %
1'
b100 +
#914130000000
0!
0'
#914140000000
1!
b101 %
1'
b101 +
#914150000000
0!
0'
#914160000000
1!
b110 %
1'
b110 +
#914170000000
0!
0'
#914180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#914190000000
0!
0'
#914200000000
1!
b1000 %
1'
b1000 +
#914210000000
0!
0'
#914220000000
1!
b1001 %
1'
b1001 +
#914230000000
0!
0'
#914240000000
1!
b0 %
1'
b0 +
#914250000000
0!
0'
#914260000000
1!
1$
b1 %
1'
1*
b1 +
#914270000000
0!
0'
#914280000000
1!
b10 %
1'
b10 +
#914290000000
0!
0'
#914300000000
1!
b11 %
1'
b11 +
#914310000000
0!
0'
#914320000000
1!
b100 %
1'
b100 +
#914330000000
0!
0'
#914340000000
1!
b101 %
1'
b101 +
#914350000000
0!
0'
#914360000000
1!
0$
b110 %
1'
0*
b110 +
#914370000000
0!
0'
#914380000000
1!
b111 %
1'
b111 +
#914390000000
1"
1(
#914400000000
0!
0"
b100 &
0'
0(
b100 ,
#914410000000
1!
b1000 %
1'
b1000 +
#914420000000
0!
0'
#914430000000
1!
b1001 %
1'
b1001 +
#914440000000
0!
0'
#914450000000
1!
b0 %
1'
b0 +
#914460000000
0!
0'
#914470000000
1!
1$
b1 %
1'
1*
b1 +
#914480000000
0!
0'
#914490000000
1!
b10 %
1'
b10 +
#914500000000
0!
0'
#914510000000
1!
b11 %
1'
b11 +
#914520000000
0!
0'
#914530000000
1!
b100 %
1'
b100 +
#914540000000
0!
0'
#914550000000
1!
b101 %
1'
b101 +
#914560000000
0!
0'
#914570000000
1!
b110 %
1'
b110 +
#914580000000
0!
0'
#914590000000
1!
b111 %
1'
b111 +
#914600000000
0!
0'
#914610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#914620000000
0!
0'
#914630000000
1!
b1001 %
1'
b1001 +
#914640000000
0!
0'
#914650000000
1!
b0 %
1'
b0 +
#914660000000
0!
0'
#914670000000
1!
1$
b1 %
1'
1*
b1 +
#914680000000
0!
0'
#914690000000
1!
b10 %
1'
b10 +
#914700000000
0!
0'
#914710000000
1!
b11 %
1'
b11 +
#914720000000
0!
0'
#914730000000
1!
b100 %
1'
b100 +
#914740000000
0!
0'
#914750000000
1!
b101 %
1'
b101 +
#914760000000
0!
0'
#914770000000
1!
0$
b110 %
1'
0*
b110 +
#914780000000
0!
0'
#914790000000
1!
b111 %
1'
b111 +
#914800000000
0!
0'
#914810000000
1!
b1000 %
1'
b1000 +
#914820000000
1"
1(
#914830000000
0!
0"
b100 &
0'
0(
b100 ,
#914840000000
1!
b1001 %
1'
b1001 +
#914850000000
0!
0'
#914860000000
1!
b0 %
1'
b0 +
#914870000000
0!
0'
#914880000000
1!
1$
b1 %
1'
1*
b1 +
#914890000000
0!
0'
#914900000000
1!
b10 %
1'
b10 +
#914910000000
0!
0'
#914920000000
1!
b11 %
1'
b11 +
#914930000000
0!
0'
#914940000000
1!
b100 %
1'
b100 +
#914950000000
0!
0'
#914960000000
1!
b101 %
1'
b101 +
#914970000000
0!
0'
#914980000000
1!
b110 %
1'
b110 +
#914990000000
0!
0'
#915000000000
1!
b111 %
1'
b111 +
#915010000000
0!
0'
#915020000000
1!
0$
b1000 %
1'
0*
b1000 +
#915030000000
0!
0'
#915040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#915050000000
0!
0'
#915060000000
1!
b0 %
1'
b0 +
#915070000000
0!
0'
#915080000000
1!
1$
b1 %
1'
1*
b1 +
#915090000000
0!
0'
#915100000000
1!
b10 %
1'
b10 +
#915110000000
0!
0'
#915120000000
1!
b11 %
1'
b11 +
#915130000000
0!
0'
#915140000000
1!
b100 %
1'
b100 +
#915150000000
0!
0'
#915160000000
1!
b101 %
1'
b101 +
#915170000000
0!
0'
#915180000000
1!
0$
b110 %
1'
0*
b110 +
#915190000000
0!
0'
#915200000000
1!
b111 %
1'
b111 +
#915210000000
0!
0'
#915220000000
1!
b1000 %
1'
b1000 +
#915230000000
0!
0'
#915240000000
1!
b1001 %
1'
b1001 +
#915250000000
1"
1(
#915260000000
0!
0"
b100 &
0'
0(
b100 ,
#915270000000
1!
b0 %
1'
b0 +
#915280000000
0!
0'
#915290000000
1!
1$
b1 %
1'
1*
b1 +
#915300000000
0!
0'
#915310000000
1!
b10 %
1'
b10 +
#915320000000
0!
0'
#915330000000
1!
b11 %
1'
b11 +
#915340000000
0!
0'
#915350000000
1!
b100 %
1'
b100 +
#915360000000
0!
0'
#915370000000
1!
b101 %
1'
b101 +
#915380000000
0!
0'
#915390000000
1!
b110 %
1'
b110 +
#915400000000
0!
0'
#915410000000
1!
b111 %
1'
b111 +
#915420000000
0!
0'
#915430000000
1!
0$
b1000 %
1'
0*
b1000 +
#915440000000
0!
0'
#915450000000
1!
b1001 %
1'
b1001 +
#915460000000
0!
0'
#915470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#915480000000
0!
0'
#915490000000
1!
1$
b1 %
1'
1*
b1 +
#915500000000
0!
0'
#915510000000
1!
b10 %
1'
b10 +
#915520000000
0!
0'
#915530000000
1!
b11 %
1'
b11 +
#915540000000
0!
0'
#915550000000
1!
b100 %
1'
b100 +
#915560000000
0!
0'
#915570000000
1!
b101 %
1'
b101 +
#915580000000
0!
0'
#915590000000
1!
0$
b110 %
1'
0*
b110 +
#915600000000
0!
0'
#915610000000
1!
b111 %
1'
b111 +
#915620000000
0!
0'
#915630000000
1!
b1000 %
1'
b1000 +
#915640000000
0!
0'
#915650000000
1!
b1001 %
1'
b1001 +
#915660000000
0!
0'
#915670000000
1!
b0 %
1'
b0 +
#915680000000
1"
1(
#915690000000
0!
0"
b100 &
0'
0(
b100 ,
#915700000000
1!
1$
b1 %
1'
1*
b1 +
#915710000000
0!
0'
#915720000000
1!
b10 %
1'
b10 +
#915730000000
0!
0'
#915740000000
1!
b11 %
1'
b11 +
#915750000000
0!
0'
#915760000000
1!
b100 %
1'
b100 +
#915770000000
0!
0'
#915780000000
1!
b101 %
1'
b101 +
#915790000000
0!
0'
#915800000000
1!
b110 %
1'
b110 +
#915810000000
0!
0'
#915820000000
1!
b111 %
1'
b111 +
#915830000000
0!
0'
#915840000000
1!
0$
b1000 %
1'
0*
b1000 +
#915850000000
0!
0'
#915860000000
1!
b1001 %
1'
b1001 +
#915870000000
0!
0'
#915880000000
1!
b0 %
1'
b0 +
#915890000000
0!
0'
#915900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#915910000000
0!
0'
#915920000000
1!
b10 %
1'
b10 +
#915930000000
0!
0'
#915940000000
1!
b11 %
1'
b11 +
#915950000000
0!
0'
#915960000000
1!
b100 %
1'
b100 +
#915970000000
0!
0'
#915980000000
1!
b101 %
1'
b101 +
#915990000000
0!
0'
#916000000000
1!
0$
b110 %
1'
0*
b110 +
#916010000000
0!
0'
#916020000000
1!
b111 %
1'
b111 +
#916030000000
0!
0'
#916040000000
1!
b1000 %
1'
b1000 +
#916050000000
0!
0'
#916060000000
1!
b1001 %
1'
b1001 +
#916070000000
0!
0'
#916080000000
1!
b0 %
1'
b0 +
#916090000000
0!
0'
#916100000000
1!
1$
b1 %
1'
1*
b1 +
#916110000000
1"
1(
#916120000000
0!
0"
b100 &
0'
0(
b100 ,
#916130000000
1!
b10 %
1'
b10 +
#916140000000
0!
0'
#916150000000
1!
b11 %
1'
b11 +
#916160000000
0!
0'
#916170000000
1!
b100 %
1'
b100 +
#916180000000
0!
0'
#916190000000
1!
b101 %
1'
b101 +
#916200000000
0!
0'
#916210000000
1!
b110 %
1'
b110 +
#916220000000
0!
0'
#916230000000
1!
b111 %
1'
b111 +
#916240000000
0!
0'
#916250000000
1!
0$
b1000 %
1'
0*
b1000 +
#916260000000
0!
0'
#916270000000
1!
b1001 %
1'
b1001 +
#916280000000
0!
0'
#916290000000
1!
b0 %
1'
b0 +
#916300000000
0!
0'
#916310000000
1!
1$
b1 %
1'
1*
b1 +
#916320000000
0!
0'
#916330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#916340000000
0!
0'
#916350000000
1!
b11 %
1'
b11 +
#916360000000
0!
0'
#916370000000
1!
b100 %
1'
b100 +
#916380000000
0!
0'
#916390000000
1!
b101 %
1'
b101 +
#916400000000
0!
0'
#916410000000
1!
0$
b110 %
1'
0*
b110 +
#916420000000
0!
0'
#916430000000
1!
b111 %
1'
b111 +
#916440000000
0!
0'
#916450000000
1!
b1000 %
1'
b1000 +
#916460000000
0!
0'
#916470000000
1!
b1001 %
1'
b1001 +
#916480000000
0!
0'
#916490000000
1!
b0 %
1'
b0 +
#916500000000
0!
0'
#916510000000
1!
1$
b1 %
1'
1*
b1 +
#916520000000
0!
0'
#916530000000
1!
b10 %
1'
b10 +
#916540000000
1"
1(
#916550000000
0!
0"
b100 &
0'
0(
b100 ,
#916560000000
1!
b11 %
1'
b11 +
#916570000000
0!
0'
#916580000000
1!
b100 %
1'
b100 +
#916590000000
0!
0'
#916600000000
1!
b101 %
1'
b101 +
#916610000000
0!
0'
#916620000000
1!
b110 %
1'
b110 +
#916630000000
0!
0'
#916640000000
1!
b111 %
1'
b111 +
#916650000000
0!
0'
#916660000000
1!
0$
b1000 %
1'
0*
b1000 +
#916670000000
0!
0'
#916680000000
1!
b1001 %
1'
b1001 +
#916690000000
0!
0'
#916700000000
1!
b0 %
1'
b0 +
#916710000000
0!
0'
#916720000000
1!
1$
b1 %
1'
1*
b1 +
#916730000000
0!
0'
#916740000000
1!
b10 %
1'
b10 +
#916750000000
0!
0'
#916760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#916770000000
0!
0'
#916780000000
1!
b100 %
1'
b100 +
#916790000000
0!
0'
#916800000000
1!
b101 %
1'
b101 +
#916810000000
0!
0'
#916820000000
1!
0$
b110 %
1'
0*
b110 +
#916830000000
0!
0'
#916840000000
1!
b111 %
1'
b111 +
#916850000000
0!
0'
#916860000000
1!
b1000 %
1'
b1000 +
#916870000000
0!
0'
#916880000000
1!
b1001 %
1'
b1001 +
#916890000000
0!
0'
#916900000000
1!
b0 %
1'
b0 +
#916910000000
0!
0'
#916920000000
1!
1$
b1 %
1'
1*
b1 +
#916930000000
0!
0'
#916940000000
1!
b10 %
1'
b10 +
#916950000000
0!
0'
#916960000000
1!
b11 %
1'
b11 +
#916970000000
1"
1(
#916980000000
0!
0"
b100 &
0'
0(
b100 ,
#916990000000
1!
b100 %
1'
b100 +
#917000000000
0!
0'
#917010000000
1!
b101 %
1'
b101 +
#917020000000
0!
0'
#917030000000
1!
b110 %
1'
b110 +
#917040000000
0!
0'
#917050000000
1!
b111 %
1'
b111 +
#917060000000
0!
0'
#917070000000
1!
0$
b1000 %
1'
0*
b1000 +
#917080000000
0!
0'
#917090000000
1!
b1001 %
1'
b1001 +
#917100000000
0!
0'
#917110000000
1!
b0 %
1'
b0 +
#917120000000
0!
0'
#917130000000
1!
1$
b1 %
1'
1*
b1 +
#917140000000
0!
0'
#917150000000
1!
b10 %
1'
b10 +
#917160000000
0!
0'
#917170000000
1!
b11 %
1'
b11 +
#917180000000
0!
0'
#917190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#917200000000
0!
0'
#917210000000
1!
b101 %
1'
b101 +
#917220000000
0!
0'
#917230000000
1!
0$
b110 %
1'
0*
b110 +
#917240000000
0!
0'
#917250000000
1!
b111 %
1'
b111 +
#917260000000
0!
0'
#917270000000
1!
b1000 %
1'
b1000 +
#917280000000
0!
0'
#917290000000
1!
b1001 %
1'
b1001 +
#917300000000
0!
0'
#917310000000
1!
b0 %
1'
b0 +
#917320000000
0!
0'
#917330000000
1!
1$
b1 %
1'
1*
b1 +
#917340000000
0!
0'
#917350000000
1!
b10 %
1'
b10 +
#917360000000
0!
0'
#917370000000
1!
b11 %
1'
b11 +
#917380000000
0!
0'
#917390000000
1!
b100 %
1'
b100 +
#917400000000
1"
1(
#917410000000
0!
0"
b100 &
0'
0(
b100 ,
#917420000000
1!
b101 %
1'
b101 +
#917430000000
0!
0'
#917440000000
1!
b110 %
1'
b110 +
#917450000000
0!
0'
#917460000000
1!
b111 %
1'
b111 +
#917470000000
0!
0'
#917480000000
1!
0$
b1000 %
1'
0*
b1000 +
#917490000000
0!
0'
#917500000000
1!
b1001 %
1'
b1001 +
#917510000000
0!
0'
#917520000000
1!
b0 %
1'
b0 +
#917530000000
0!
0'
#917540000000
1!
1$
b1 %
1'
1*
b1 +
#917550000000
0!
0'
#917560000000
1!
b10 %
1'
b10 +
#917570000000
0!
0'
#917580000000
1!
b11 %
1'
b11 +
#917590000000
0!
0'
#917600000000
1!
b100 %
1'
b100 +
#917610000000
0!
0'
#917620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#917630000000
0!
0'
#917640000000
1!
0$
b110 %
1'
0*
b110 +
#917650000000
0!
0'
#917660000000
1!
b111 %
1'
b111 +
#917670000000
0!
0'
#917680000000
1!
b1000 %
1'
b1000 +
#917690000000
0!
0'
#917700000000
1!
b1001 %
1'
b1001 +
#917710000000
0!
0'
#917720000000
1!
b0 %
1'
b0 +
#917730000000
0!
0'
#917740000000
1!
1$
b1 %
1'
1*
b1 +
#917750000000
0!
0'
#917760000000
1!
b10 %
1'
b10 +
#917770000000
0!
0'
#917780000000
1!
b11 %
1'
b11 +
#917790000000
0!
0'
#917800000000
1!
b100 %
1'
b100 +
#917810000000
0!
0'
#917820000000
1!
b101 %
1'
b101 +
#917830000000
1"
1(
#917840000000
0!
0"
b100 &
0'
0(
b100 ,
#917850000000
1!
b110 %
1'
b110 +
#917860000000
0!
0'
#917870000000
1!
b111 %
1'
b111 +
#917880000000
0!
0'
#917890000000
1!
0$
b1000 %
1'
0*
b1000 +
#917900000000
0!
0'
#917910000000
1!
b1001 %
1'
b1001 +
#917920000000
0!
0'
#917930000000
1!
b0 %
1'
b0 +
#917940000000
0!
0'
#917950000000
1!
1$
b1 %
1'
1*
b1 +
#917960000000
0!
0'
#917970000000
1!
b10 %
1'
b10 +
#917980000000
0!
0'
#917990000000
1!
b11 %
1'
b11 +
#918000000000
0!
0'
#918010000000
1!
b100 %
1'
b100 +
#918020000000
0!
0'
#918030000000
1!
b101 %
1'
b101 +
#918040000000
0!
0'
#918050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#918060000000
0!
0'
#918070000000
1!
b111 %
1'
b111 +
#918080000000
0!
0'
#918090000000
1!
b1000 %
1'
b1000 +
#918100000000
0!
0'
#918110000000
1!
b1001 %
1'
b1001 +
#918120000000
0!
0'
#918130000000
1!
b0 %
1'
b0 +
#918140000000
0!
0'
#918150000000
1!
1$
b1 %
1'
1*
b1 +
#918160000000
0!
0'
#918170000000
1!
b10 %
1'
b10 +
#918180000000
0!
0'
#918190000000
1!
b11 %
1'
b11 +
#918200000000
0!
0'
#918210000000
1!
b100 %
1'
b100 +
#918220000000
0!
0'
#918230000000
1!
b101 %
1'
b101 +
#918240000000
0!
0'
#918250000000
1!
0$
b110 %
1'
0*
b110 +
#918260000000
1"
1(
#918270000000
0!
0"
b100 &
0'
0(
b100 ,
#918280000000
1!
1$
b111 %
1'
1*
b111 +
#918290000000
0!
0'
#918300000000
1!
0$
b1000 %
1'
0*
b1000 +
#918310000000
0!
0'
#918320000000
1!
b1001 %
1'
b1001 +
#918330000000
0!
0'
#918340000000
1!
b0 %
1'
b0 +
#918350000000
0!
0'
#918360000000
1!
1$
b1 %
1'
1*
b1 +
#918370000000
0!
0'
#918380000000
1!
b10 %
1'
b10 +
#918390000000
0!
0'
#918400000000
1!
b11 %
1'
b11 +
#918410000000
0!
0'
#918420000000
1!
b100 %
1'
b100 +
#918430000000
0!
0'
#918440000000
1!
b101 %
1'
b101 +
#918450000000
0!
0'
#918460000000
1!
b110 %
1'
b110 +
#918470000000
0!
0'
#918480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#918490000000
0!
0'
#918500000000
1!
b1000 %
1'
b1000 +
#918510000000
0!
0'
#918520000000
1!
b1001 %
1'
b1001 +
#918530000000
0!
0'
#918540000000
1!
b0 %
1'
b0 +
#918550000000
0!
0'
#918560000000
1!
1$
b1 %
1'
1*
b1 +
#918570000000
0!
0'
#918580000000
1!
b10 %
1'
b10 +
#918590000000
0!
0'
#918600000000
1!
b11 %
1'
b11 +
#918610000000
0!
0'
#918620000000
1!
b100 %
1'
b100 +
#918630000000
0!
0'
#918640000000
1!
b101 %
1'
b101 +
#918650000000
0!
0'
#918660000000
1!
0$
b110 %
1'
0*
b110 +
#918670000000
0!
0'
#918680000000
1!
b111 %
1'
b111 +
#918690000000
1"
1(
#918700000000
0!
0"
b100 &
0'
0(
b100 ,
#918710000000
1!
b1000 %
1'
b1000 +
#918720000000
0!
0'
#918730000000
1!
b1001 %
1'
b1001 +
#918740000000
0!
0'
#918750000000
1!
b0 %
1'
b0 +
#918760000000
0!
0'
#918770000000
1!
1$
b1 %
1'
1*
b1 +
#918780000000
0!
0'
#918790000000
1!
b10 %
1'
b10 +
#918800000000
0!
0'
#918810000000
1!
b11 %
1'
b11 +
#918820000000
0!
0'
#918830000000
1!
b100 %
1'
b100 +
#918840000000
0!
0'
#918850000000
1!
b101 %
1'
b101 +
#918860000000
0!
0'
#918870000000
1!
b110 %
1'
b110 +
#918880000000
0!
0'
#918890000000
1!
b111 %
1'
b111 +
#918900000000
0!
0'
#918910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#918920000000
0!
0'
#918930000000
1!
b1001 %
1'
b1001 +
#918940000000
0!
0'
#918950000000
1!
b0 %
1'
b0 +
#918960000000
0!
0'
#918970000000
1!
1$
b1 %
1'
1*
b1 +
#918980000000
0!
0'
#918990000000
1!
b10 %
1'
b10 +
#919000000000
0!
0'
#919010000000
1!
b11 %
1'
b11 +
#919020000000
0!
0'
#919030000000
1!
b100 %
1'
b100 +
#919040000000
0!
0'
#919050000000
1!
b101 %
1'
b101 +
#919060000000
0!
0'
#919070000000
1!
0$
b110 %
1'
0*
b110 +
#919080000000
0!
0'
#919090000000
1!
b111 %
1'
b111 +
#919100000000
0!
0'
#919110000000
1!
b1000 %
1'
b1000 +
#919120000000
1"
1(
#919130000000
0!
0"
b100 &
0'
0(
b100 ,
#919140000000
1!
b1001 %
1'
b1001 +
#919150000000
0!
0'
#919160000000
1!
b0 %
1'
b0 +
#919170000000
0!
0'
#919180000000
1!
1$
b1 %
1'
1*
b1 +
#919190000000
0!
0'
#919200000000
1!
b10 %
1'
b10 +
#919210000000
0!
0'
#919220000000
1!
b11 %
1'
b11 +
#919230000000
0!
0'
#919240000000
1!
b100 %
1'
b100 +
#919250000000
0!
0'
#919260000000
1!
b101 %
1'
b101 +
#919270000000
0!
0'
#919280000000
1!
b110 %
1'
b110 +
#919290000000
0!
0'
#919300000000
1!
b111 %
1'
b111 +
#919310000000
0!
0'
#919320000000
1!
0$
b1000 %
1'
0*
b1000 +
#919330000000
0!
0'
#919340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#919350000000
0!
0'
#919360000000
1!
b0 %
1'
b0 +
#919370000000
0!
0'
#919380000000
1!
1$
b1 %
1'
1*
b1 +
#919390000000
0!
0'
#919400000000
1!
b10 %
1'
b10 +
#919410000000
0!
0'
#919420000000
1!
b11 %
1'
b11 +
#919430000000
0!
0'
#919440000000
1!
b100 %
1'
b100 +
#919450000000
0!
0'
#919460000000
1!
b101 %
1'
b101 +
#919470000000
0!
0'
#919480000000
1!
0$
b110 %
1'
0*
b110 +
#919490000000
0!
0'
#919500000000
1!
b111 %
1'
b111 +
#919510000000
0!
0'
#919520000000
1!
b1000 %
1'
b1000 +
#919530000000
0!
0'
#919540000000
1!
b1001 %
1'
b1001 +
#919550000000
1"
1(
#919560000000
0!
0"
b100 &
0'
0(
b100 ,
#919570000000
1!
b0 %
1'
b0 +
#919580000000
0!
0'
#919590000000
1!
1$
b1 %
1'
1*
b1 +
#919600000000
0!
0'
#919610000000
1!
b10 %
1'
b10 +
#919620000000
0!
0'
#919630000000
1!
b11 %
1'
b11 +
#919640000000
0!
0'
#919650000000
1!
b100 %
1'
b100 +
#919660000000
0!
0'
#919670000000
1!
b101 %
1'
b101 +
#919680000000
0!
0'
#919690000000
1!
b110 %
1'
b110 +
#919700000000
0!
0'
#919710000000
1!
b111 %
1'
b111 +
#919720000000
0!
0'
#919730000000
1!
0$
b1000 %
1'
0*
b1000 +
#919740000000
0!
0'
#919750000000
1!
b1001 %
1'
b1001 +
#919760000000
0!
0'
#919770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#919780000000
0!
0'
#919790000000
1!
1$
b1 %
1'
1*
b1 +
#919800000000
0!
0'
#919810000000
1!
b10 %
1'
b10 +
#919820000000
0!
0'
#919830000000
1!
b11 %
1'
b11 +
#919840000000
0!
0'
#919850000000
1!
b100 %
1'
b100 +
#919860000000
0!
0'
#919870000000
1!
b101 %
1'
b101 +
#919880000000
0!
0'
#919890000000
1!
0$
b110 %
1'
0*
b110 +
#919900000000
0!
0'
#919910000000
1!
b111 %
1'
b111 +
#919920000000
0!
0'
#919930000000
1!
b1000 %
1'
b1000 +
#919940000000
0!
0'
#919950000000
1!
b1001 %
1'
b1001 +
#919960000000
0!
0'
#919970000000
1!
b0 %
1'
b0 +
#919980000000
1"
1(
#919990000000
0!
0"
b100 &
0'
0(
b100 ,
#920000000000
1!
1$
b1 %
1'
1*
b1 +
#920010000000
0!
0'
#920020000000
1!
b10 %
1'
b10 +
#920030000000
0!
0'
#920040000000
1!
b11 %
1'
b11 +
#920050000000
0!
0'
#920060000000
1!
b100 %
1'
b100 +
#920070000000
0!
0'
#920080000000
1!
b101 %
1'
b101 +
#920090000000
0!
0'
#920100000000
1!
b110 %
1'
b110 +
#920110000000
0!
0'
#920120000000
1!
b111 %
1'
b111 +
#920130000000
0!
0'
#920140000000
1!
0$
b1000 %
1'
0*
b1000 +
#920150000000
0!
0'
#920160000000
1!
b1001 %
1'
b1001 +
#920170000000
0!
0'
#920180000000
1!
b0 %
1'
b0 +
#920190000000
0!
0'
#920200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#920210000000
0!
0'
#920220000000
1!
b10 %
1'
b10 +
#920230000000
0!
0'
#920240000000
1!
b11 %
1'
b11 +
#920250000000
0!
0'
#920260000000
1!
b100 %
1'
b100 +
#920270000000
0!
0'
#920280000000
1!
b101 %
1'
b101 +
#920290000000
0!
0'
#920300000000
1!
0$
b110 %
1'
0*
b110 +
#920310000000
0!
0'
#920320000000
1!
b111 %
1'
b111 +
#920330000000
0!
0'
#920340000000
1!
b1000 %
1'
b1000 +
#920350000000
0!
0'
#920360000000
1!
b1001 %
1'
b1001 +
#920370000000
0!
0'
#920380000000
1!
b0 %
1'
b0 +
#920390000000
0!
0'
#920400000000
1!
1$
b1 %
1'
1*
b1 +
#920410000000
1"
1(
#920420000000
0!
0"
b100 &
0'
0(
b100 ,
#920430000000
1!
b10 %
1'
b10 +
#920440000000
0!
0'
#920450000000
1!
b11 %
1'
b11 +
#920460000000
0!
0'
#920470000000
1!
b100 %
1'
b100 +
#920480000000
0!
0'
#920490000000
1!
b101 %
1'
b101 +
#920500000000
0!
0'
#920510000000
1!
b110 %
1'
b110 +
#920520000000
0!
0'
#920530000000
1!
b111 %
1'
b111 +
#920540000000
0!
0'
#920550000000
1!
0$
b1000 %
1'
0*
b1000 +
#920560000000
0!
0'
#920570000000
1!
b1001 %
1'
b1001 +
#920580000000
0!
0'
#920590000000
1!
b0 %
1'
b0 +
#920600000000
0!
0'
#920610000000
1!
1$
b1 %
1'
1*
b1 +
#920620000000
0!
0'
#920630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#920640000000
0!
0'
#920650000000
1!
b11 %
1'
b11 +
#920660000000
0!
0'
#920670000000
1!
b100 %
1'
b100 +
#920680000000
0!
0'
#920690000000
1!
b101 %
1'
b101 +
#920700000000
0!
0'
#920710000000
1!
0$
b110 %
1'
0*
b110 +
#920720000000
0!
0'
#920730000000
1!
b111 %
1'
b111 +
#920740000000
0!
0'
#920750000000
1!
b1000 %
1'
b1000 +
#920760000000
0!
0'
#920770000000
1!
b1001 %
1'
b1001 +
#920780000000
0!
0'
#920790000000
1!
b0 %
1'
b0 +
#920800000000
0!
0'
#920810000000
1!
1$
b1 %
1'
1*
b1 +
#920820000000
0!
0'
#920830000000
1!
b10 %
1'
b10 +
#920840000000
1"
1(
#920850000000
0!
0"
b100 &
0'
0(
b100 ,
#920860000000
1!
b11 %
1'
b11 +
#920870000000
0!
0'
#920880000000
1!
b100 %
1'
b100 +
#920890000000
0!
0'
#920900000000
1!
b101 %
1'
b101 +
#920910000000
0!
0'
#920920000000
1!
b110 %
1'
b110 +
#920930000000
0!
0'
#920940000000
1!
b111 %
1'
b111 +
#920950000000
0!
0'
#920960000000
1!
0$
b1000 %
1'
0*
b1000 +
#920970000000
0!
0'
#920980000000
1!
b1001 %
1'
b1001 +
#920990000000
0!
0'
#921000000000
1!
b0 %
1'
b0 +
#921010000000
0!
0'
#921020000000
1!
1$
b1 %
1'
1*
b1 +
#921030000000
0!
0'
#921040000000
1!
b10 %
1'
b10 +
#921050000000
0!
0'
#921060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#921070000000
0!
0'
#921080000000
1!
b100 %
1'
b100 +
#921090000000
0!
0'
#921100000000
1!
b101 %
1'
b101 +
#921110000000
0!
0'
#921120000000
1!
0$
b110 %
1'
0*
b110 +
#921130000000
0!
0'
#921140000000
1!
b111 %
1'
b111 +
#921150000000
0!
0'
#921160000000
1!
b1000 %
1'
b1000 +
#921170000000
0!
0'
#921180000000
1!
b1001 %
1'
b1001 +
#921190000000
0!
0'
#921200000000
1!
b0 %
1'
b0 +
#921210000000
0!
0'
#921220000000
1!
1$
b1 %
1'
1*
b1 +
#921230000000
0!
0'
#921240000000
1!
b10 %
1'
b10 +
#921250000000
0!
0'
#921260000000
1!
b11 %
1'
b11 +
#921270000000
1"
1(
#921280000000
0!
0"
b100 &
0'
0(
b100 ,
#921290000000
1!
b100 %
1'
b100 +
#921300000000
0!
0'
#921310000000
1!
b101 %
1'
b101 +
#921320000000
0!
0'
#921330000000
1!
b110 %
1'
b110 +
#921340000000
0!
0'
#921350000000
1!
b111 %
1'
b111 +
#921360000000
0!
0'
#921370000000
1!
0$
b1000 %
1'
0*
b1000 +
#921380000000
0!
0'
#921390000000
1!
b1001 %
1'
b1001 +
#921400000000
0!
0'
#921410000000
1!
b0 %
1'
b0 +
#921420000000
0!
0'
#921430000000
1!
1$
b1 %
1'
1*
b1 +
#921440000000
0!
0'
#921450000000
1!
b10 %
1'
b10 +
#921460000000
0!
0'
#921470000000
1!
b11 %
1'
b11 +
#921480000000
0!
0'
#921490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#921500000000
0!
0'
#921510000000
1!
b101 %
1'
b101 +
#921520000000
0!
0'
#921530000000
1!
0$
b110 %
1'
0*
b110 +
#921540000000
0!
0'
#921550000000
1!
b111 %
1'
b111 +
#921560000000
0!
0'
#921570000000
1!
b1000 %
1'
b1000 +
#921580000000
0!
0'
#921590000000
1!
b1001 %
1'
b1001 +
#921600000000
0!
0'
#921610000000
1!
b0 %
1'
b0 +
#921620000000
0!
0'
#921630000000
1!
1$
b1 %
1'
1*
b1 +
#921640000000
0!
0'
#921650000000
1!
b10 %
1'
b10 +
#921660000000
0!
0'
#921670000000
1!
b11 %
1'
b11 +
#921680000000
0!
0'
#921690000000
1!
b100 %
1'
b100 +
#921700000000
1"
1(
#921710000000
0!
0"
b100 &
0'
0(
b100 ,
#921720000000
1!
b101 %
1'
b101 +
#921730000000
0!
0'
#921740000000
1!
b110 %
1'
b110 +
#921750000000
0!
0'
#921760000000
1!
b111 %
1'
b111 +
#921770000000
0!
0'
#921780000000
1!
0$
b1000 %
1'
0*
b1000 +
#921790000000
0!
0'
#921800000000
1!
b1001 %
1'
b1001 +
#921810000000
0!
0'
#921820000000
1!
b0 %
1'
b0 +
#921830000000
0!
0'
#921840000000
1!
1$
b1 %
1'
1*
b1 +
#921850000000
0!
0'
#921860000000
1!
b10 %
1'
b10 +
#921870000000
0!
0'
#921880000000
1!
b11 %
1'
b11 +
#921890000000
0!
0'
#921900000000
1!
b100 %
1'
b100 +
#921910000000
0!
0'
#921920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#921930000000
0!
0'
#921940000000
1!
0$
b110 %
1'
0*
b110 +
#921950000000
0!
0'
#921960000000
1!
b111 %
1'
b111 +
#921970000000
0!
0'
#921980000000
1!
b1000 %
1'
b1000 +
#921990000000
0!
0'
#922000000000
1!
b1001 %
1'
b1001 +
#922010000000
0!
0'
#922020000000
1!
b0 %
1'
b0 +
#922030000000
0!
0'
#922040000000
1!
1$
b1 %
1'
1*
b1 +
#922050000000
0!
0'
#922060000000
1!
b10 %
1'
b10 +
#922070000000
0!
0'
#922080000000
1!
b11 %
1'
b11 +
#922090000000
0!
0'
#922100000000
1!
b100 %
1'
b100 +
#922110000000
0!
0'
#922120000000
1!
b101 %
1'
b101 +
#922130000000
1"
1(
#922140000000
0!
0"
b100 &
0'
0(
b100 ,
#922150000000
1!
b110 %
1'
b110 +
#922160000000
0!
0'
#922170000000
1!
b111 %
1'
b111 +
#922180000000
0!
0'
#922190000000
1!
0$
b1000 %
1'
0*
b1000 +
#922200000000
0!
0'
#922210000000
1!
b1001 %
1'
b1001 +
#922220000000
0!
0'
#922230000000
1!
b0 %
1'
b0 +
#922240000000
0!
0'
#922250000000
1!
1$
b1 %
1'
1*
b1 +
#922260000000
0!
0'
#922270000000
1!
b10 %
1'
b10 +
#922280000000
0!
0'
#922290000000
1!
b11 %
1'
b11 +
#922300000000
0!
0'
#922310000000
1!
b100 %
1'
b100 +
#922320000000
0!
0'
#922330000000
1!
b101 %
1'
b101 +
#922340000000
0!
0'
#922350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#922360000000
0!
0'
#922370000000
1!
b111 %
1'
b111 +
#922380000000
0!
0'
#922390000000
1!
b1000 %
1'
b1000 +
#922400000000
0!
0'
#922410000000
1!
b1001 %
1'
b1001 +
#922420000000
0!
0'
#922430000000
1!
b0 %
1'
b0 +
#922440000000
0!
0'
#922450000000
1!
1$
b1 %
1'
1*
b1 +
#922460000000
0!
0'
#922470000000
1!
b10 %
1'
b10 +
#922480000000
0!
0'
#922490000000
1!
b11 %
1'
b11 +
#922500000000
0!
0'
#922510000000
1!
b100 %
1'
b100 +
#922520000000
0!
0'
#922530000000
1!
b101 %
1'
b101 +
#922540000000
0!
0'
#922550000000
1!
0$
b110 %
1'
0*
b110 +
#922560000000
1"
1(
#922570000000
0!
0"
b100 &
0'
0(
b100 ,
#922580000000
1!
1$
b111 %
1'
1*
b111 +
#922590000000
0!
0'
#922600000000
1!
0$
b1000 %
1'
0*
b1000 +
#922610000000
0!
0'
#922620000000
1!
b1001 %
1'
b1001 +
#922630000000
0!
0'
#922640000000
1!
b0 %
1'
b0 +
#922650000000
0!
0'
#922660000000
1!
1$
b1 %
1'
1*
b1 +
#922670000000
0!
0'
#922680000000
1!
b10 %
1'
b10 +
#922690000000
0!
0'
#922700000000
1!
b11 %
1'
b11 +
#922710000000
0!
0'
#922720000000
1!
b100 %
1'
b100 +
#922730000000
0!
0'
#922740000000
1!
b101 %
1'
b101 +
#922750000000
0!
0'
#922760000000
1!
b110 %
1'
b110 +
#922770000000
0!
0'
#922780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#922790000000
0!
0'
#922800000000
1!
b1000 %
1'
b1000 +
#922810000000
0!
0'
#922820000000
1!
b1001 %
1'
b1001 +
#922830000000
0!
0'
#922840000000
1!
b0 %
1'
b0 +
#922850000000
0!
0'
#922860000000
1!
1$
b1 %
1'
1*
b1 +
#922870000000
0!
0'
#922880000000
1!
b10 %
1'
b10 +
#922890000000
0!
0'
#922900000000
1!
b11 %
1'
b11 +
#922910000000
0!
0'
#922920000000
1!
b100 %
1'
b100 +
#922930000000
0!
0'
#922940000000
1!
b101 %
1'
b101 +
#922950000000
0!
0'
#922960000000
1!
0$
b110 %
1'
0*
b110 +
#922970000000
0!
0'
#922980000000
1!
b111 %
1'
b111 +
#922990000000
1"
1(
#923000000000
0!
0"
b100 &
0'
0(
b100 ,
#923010000000
1!
b1000 %
1'
b1000 +
#923020000000
0!
0'
#923030000000
1!
b1001 %
1'
b1001 +
#923040000000
0!
0'
#923050000000
1!
b0 %
1'
b0 +
#923060000000
0!
0'
#923070000000
1!
1$
b1 %
1'
1*
b1 +
#923080000000
0!
0'
#923090000000
1!
b10 %
1'
b10 +
#923100000000
0!
0'
#923110000000
1!
b11 %
1'
b11 +
#923120000000
0!
0'
#923130000000
1!
b100 %
1'
b100 +
#923140000000
0!
0'
#923150000000
1!
b101 %
1'
b101 +
#923160000000
0!
0'
#923170000000
1!
b110 %
1'
b110 +
#923180000000
0!
0'
#923190000000
1!
b111 %
1'
b111 +
#923200000000
0!
0'
#923210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#923220000000
0!
0'
#923230000000
1!
b1001 %
1'
b1001 +
#923240000000
0!
0'
#923250000000
1!
b0 %
1'
b0 +
#923260000000
0!
0'
#923270000000
1!
1$
b1 %
1'
1*
b1 +
#923280000000
0!
0'
#923290000000
1!
b10 %
1'
b10 +
#923300000000
0!
0'
#923310000000
1!
b11 %
1'
b11 +
#923320000000
0!
0'
#923330000000
1!
b100 %
1'
b100 +
#923340000000
0!
0'
#923350000000
1!
b101 %
1'
b101 +
#923360000000
0!
0'
#923370000000
1!
0$
b110 %
1'
0*
b110 +
#923380000000
0!
0'
#923390000000
1!
b111 %
1'
b111 +
#923400000000
0!
0'
#923410000000
1!
b1000 %
1'
b1000 +
#923420000000
1"
1(
#923430000000
0!
0"
b100 &
0'
0(
b100 ,
#923440000000
1!
b1001 %
1'
b1001 +
#923450000000
0!
0'
#923460000000
1!
b0 %
1'
b0 +
#923470000000
0!
0'
#923480000000
1!
1$
b1 %
1'
1*
b1 +
#923490000000
0!
0'
#923500000000
1!
b10 %
1'
b10 +
#923510000000
0!
0'
#923520000000
1!
b11 %
1'
b11 +
#923530000000
0!
0'
#923540000000
1!
b100 %
1'
b100 +
#923550000000
0!
0'
#923560000000
1!
b101 %
1'
b101 +
#923570000000
0!
0'
#923580000000
1!
b110 %
1'
b110 +
#923590000000
0!
0'
#923600000000
1!
b111 %
1'
b111 +
#923610000000
0!
0'
#923620000000
1!
0$
b1000 %
1'
0*
b1000 +
#923630000000
0!
0'
#923640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#923650000000
0!
0'
#923660000000
1!
b0 %
1'
b0 +
#923670000000
0!
0'
#923680000000
1!
1$
b1 %
1'
1*
b1 +
#923690000000
0!
0'
#923700000000
1!
b10 %
1'
b10 +
#923710000000
0!
0'
#923720000000
1!
b11 %
1'
b11 +
#923730000000
0!
0'
#923740000000
1!
b100 %
1'
b100 +
#923750000000
0!
0'
#923760000000
1!
b101 %
1'
b101 +
#923770000000
0!
0'
#923780000000
1!
0$
b110 %
1'
0*
b110 +
#923790000000
0!
0'
#923800000000
1!
b111 %
1'
b111 +
#923810000000
0!
0'
#923820000000
1!
b1000 %
1'
b1000 +
#923830000000
0!
0'
#923840000000
1!
b1001 %
1'
b1001 +
#923850000000
1"
1(
#923860000000
0!
0"
b100 &
0'
0(
b100 ,
#923870000000
1!
b0 %
1'
b0 +
#923880000000
0!
0'
#923890000000
1!
1$
b1 %
1'
1*
b1 +
#923900000000
0!
0'
#923910000000
1!
b10 %
1'
b10 +
#923920000000
0!
0'
#923930000000
1!
b11 %
1'
b11 +
#923940000000
0!
0'
#923950000000
1!
b100 %
1'
b100 +
#923960000000
0!
0'
#923970000000
1!
b101 %
1'
b101 +
#923980000000
0!
0'
#923990000000
1!
b110 %
1'
b110 +
#924000000000
0!
0'
#924010000000
1!
b111 %
1'
b111 +
#924020000000
0!
0'
#924030000000
1!
0$
b1000 %
1'
0*
b1000 +
#924040000000
0!
0'
#924050000000
1!
b1001 %
1'
b1001 +
#924060000000
0!
0'
#924070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#924080000000
0!
0'
#924090000000
1!
1$
b1 %
1'
1*
b1 +
#924100000000
0!
0'
#924110000000
1!
b10 %
1'
b10 +
#924120000000
0!
0'
#924130000000
1!
b11 %
1'
b11 +
#924140000000
0!
0'
#924150000000
1!
b100 %
1'
b100 +
#924160000000
0!
0'
#924170000000
1!
b101 %
1'
b101 +
#924180000000
0!
0'
#924190000000
1!
0$
b110 %
1'
0*
b110 +
#924200000000
0!
0'
#924210000000
1!
b111 %
1'
b111 +
#924220000000
0!
0'
#924230000000
1!
b1000 %
1'
b1000 +
#924240000000
0!
0'
#924250000000
1!
b1001 %
1'
b1001 +
#924260000000
0!
0'
#924270000000
1!
b0 %
1'
b0 +
#924280000000
1"
1(
#924290000000
0!
0"
b100 &
0'
0(
b100 ,
#924300000000
1!
1$
b1 %
1'
1*
b1 +
#924310000000
0!
0'
#924320000000
1!
b10 %
1'
b10 +
#924330000000
0!
0'
#924340000000
1!
b11 %
1'
b11 +
#924350000000
0!
0'
#924360000000
1!
b100 %
1'
b100 +
#924370000000
0!
0'
#924380000000
1!
b101 %
1'
b101 +
#924390000000
0!
0'
#924400000000
1!
b110 %
1'
b110 +
#924410000000
0!
0'
#924420000000
1!
b111 %
1'
b111 +
#924430000000
0!
0'
#924440000000
1!
0$
b1000 %
1'
0*
b1000 +
#924450000000
0!
0'
#924460000000
1!
b1001 %
1'
b1001 +
#924470000000
0!
0'
#924480000000
1!
b0 %
1'
b0 +
#924490000000
0!
0'
#924500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#924510000000
0!
0'
#924520000000
1!
b10 %
1'
b10 +
#924530000000
0!
0'
#924540000000
1!
b11 %
1'
b11 +
#924550000000
0!
0'
#924560000000
1!
b100 %
1'
b100 +
#924570000000
0!
0'
#924580000000
1!
b101 %
1'
b101 +
#924590000000
0!
0'
#924600000000
1!
0$
b110 %
1'
0*
b110 +
#924610000000
0!
0'
#924620000000
1!
b111 %
1'
b111 +
#924630000000
0!
0'
#924640000000
1!
b1000 %
1'
b1000 +
#924650000000
0!
0'
#924660000000
1!
b1001 %
1'
b1001 +
#924670000000
0!
0'
#924680000000
1!
b0 %
1'
b0 +
#924690000000
0!
0'
#924700000000
1!
1$
b1 %
1'
1*
b1 +
#924710000000
1"
1(
#924720000000
0!
0"
b100 &
0'
0(
b100 ,
#924730000000
1!
b10 %
1'
b10 +
#924740000000
0!
0'
#924750000000
1!
b11 %
1'
b11 +
#924760000000
0!
0'
#924770000000
1!
b100 %
1'
b100 +
#924780000000
0!
0'
#924790000000
1!
b101 %
1'
b101 +
#924800000000
0!
0'
#924810000000
1!
b110 %
1'
b110 +
#924820000000
0!
0'
#924830000000
1!
b111 %
1'
b111 +
#924840000000
0!
0'
#924850000000
1!
0$
b1000 %
1'
0*
b1000 +
#924860000000
0!
0'
#924870000000
1!
b1001 %
1'
b1001 +
#924880000000
0!
0'
#924890000000
1!
b0 %
1'
b0 +
#924900000000
0!
0'
#924910000000
1!
1$
b1 %
1'
1*
b1 +
#924920000000
0!
0'
#924930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#924940000000
0!
0'
#924950000000
1!
b11 %
1'
b11 +
#924960000000
0!
0'
#924970000000
1!
b100 %
1'
b100 +
#924980000000
0!
0'
#924990000000
1!
b101 %
1'
b101 +
#925000000000
0!
0'
#925010000000
1!
0$
b110 %
1'
0*
b110 +
#925020000000
0!
0'
#925030000000
1!
b111 %
1'
b111 +
#925040000000
0!
0'
#925050000000
1!
b1000 %
1'
b1000 +
#925060000000
0!
0'
#925070000000
1!
b1001 %
1'
b1001 +
#925080000000
0!
0'
#925090000000
1!
b0 %
1'
b0 +
#925100000000
0!
0'
#925110000000
1!
1$
b1 %
1'
1*
b1 +
#925120000000
0!
0'
#925130000000
1!
b10 %
1'
b10 +
#925140000000
1"
1(
#925150000000
0!
0"
b100 &
0'
0(
b100 ,
#925160000000
1!
b11 %
1'
b11 +
#925170000000
0!
0'
#925180000000
1!
b100 %
1'
b100 +
#925190000000
0!
0'
#925200000000
1!
b101 %
1'
b101 +
#925210000000
0!
0'
#925220000000
1!
b110 %
1'
b110 +
#925230000000
0!
0'
#925240000000
1!
b111 %
1'
b111 +
#925250000000
0!
0'
#925260000000
1!
0$
b1000 %
1'
0*
b1000 +
#925270000000
0!
0'
#925280000000
1!
b1001 %
1'
b1001 +
#925290000000
0!
0'
#925300000000
1!
b0 %
1'
b0 +
#925310000000
0!
0'
#925320000000
1!
1$
b1 %
1'
1*
b1 +
#925330000000
0!
0'
#925340000000
1!
b10 %
1'
b10 +
#925350000000
0!
0'
#925360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#925370000000
0!
0'
#925380000000
1!
b100 %
1'
b100 +
#925390000000
0!
0'
#925400000000
1!
b101 %
1'
b101 +
#925410000000
0!
0'
#925420000000
1!
0$
b110 %
1'
0*
b110 +
#925430000000
0!
0'
#925440000000
1!
b111 %
1'
b111 +
#925450000000
0!
0'
#925460000000
1!
b1000 %
1'
b1000 +
#925470000000
0!
0'
#925480000000
1!
b1001 %
1'
b1001 +
#925490000000
0!
0'
#925500000000
1!
b0 %
1'
b0 +
#925510000000
0!
0'
#925520000000
1!
1$
b1 %
1'
1*
b1 +
#925530000000
0!
0'
#925540000000
1!
b10 %
1'
b10 +
#925550000000
0!
0'
#925560000000
1!
b11 %
1'
b11 +
#925570000000
1"
1(
#925580000000
0!
0"
b100 &
0'
0(
b100 ,
#925590000000
1!
b100 %
1'
b100 +
#925600000000
0!
0'
#925610000000
1!
b101 %
1'
b101 +
#925620000000
0!
0'
#925630000000
1!
b110 %
1'
b110 +
#925640000000
0!
0'
#925650000000
1!
b111 %
1'
b111 +
#925660000000
0!
0'
#925670000000
1!
0$
b1000 %
1'
0*
b1000 +
#925680000000
0!
0'
#925690000000
1!
b1001 %
1'
b1001 +
#925700000000
0!
0'
#925710000000
1!
b0 %
1'
b0 +
#925720000000
0!
0'
#925730000000
1!
1$
b1 %
1'
1*
b1 +
#925740000000
0!
0'
#925750000000
1!
b10 %
1'
b10 +
#925760000000
0!
0'
#925770000000
1!
b11 %
1'
b11 +
#925780000000
0!
0'
#925790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#925800000000
0!
0'
#925810000000
1!
b101 %
1'
b101 +
#925820000000
0!
0'
#925830000000
1!
0$
b110 %
1'
0*
b110 +
#925840000000
0!
0'
#925850000000
1!
b111 %
1'
b111 +
#925860000000
0!
0'
#925870000000
1!
b1000 %
1'
b1000 +
#925880000000
0!
0'
#925890000000
1!
b1001 %
1'
b1001 +
#925900000000
0!
0'
#925910000000
1!
b0 %
1'
b0 +
#925920000000
0!
0'
#925930000000
1!
1$
b1 %
1'
1*
b1 +
#925940000000
0!
0'
#925950000000
1!
b10 %
1'
b10 +
#925960000000
0!
0'
#925970000000
1!
b11 %
1'
b11 +
#925980000000
0!
0'
#925990000000
1!
b100 %
1'
b100 +
#926000000000
1"
1(
#926010000000
0!
0"
b100 &
0'
0(
b100 ,
#926020000000
1!
b101 %
1'
b101 +
#926030000000
0!
0'
#926040000000
1!
b110 %
1'
b110 +
#926050000000
0!
0'
#926060000000
1!
b111 %
1'
b111 +
#926070000000
0!
0'
#926080000000
1!
0$
b1000 %
1'
0*
b1000 +
#926090000000
0!
0'
#926100000000
1!
b1001 %
1'
b1001 +
#926110000000
0!
0'
#926120000000
1!
b0 %
1'
b0 +
#926130000000
0!
0'
#926140000000
1!
1$
b1 %
1'
1*
b1 +
#926150000000
0!
0'
#926160000000
1!
b10 %
1'
b10 +
#926170000000
0!
0'
#926180000000
1!
b11 %
1'
b11 +
#926190000000
0!
0'
#926200000000
1!
b100 %
1'
b100 +
#926210000000
0!
0'
#926220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#926230000000
0!
0'
#926240000000
1!
0$
b110 %
1'
0*
b110 +
#926250000000
0!
0'
#926260000000
1!
b111 %
1'
b111 +
#926270000000
0!
0'
#926280000000
1!
b1000 %
1'
b1000 +
#926290000000
0!
0'
#926300000000
1!
b1001 %
1'
b1001 +
#926310000000
0!
0'
#926320000000
1!
b0 %
1'
b0 +
#926330000000
0!
0'
#926340000000
1!
1$
b1 %
1'
1*
b1 +
#926350000000
0!
0'
#926360000000
1!
b10 %
1'
b10 +
#926370000000
0!
0'
#926380000000
1!
b11 %
1'
b11 +
#926390000000
0!
0'
#926400000000
1!
b100 %
1'
b100 +
#926410000000
0!
0'
#926420000000
1!
b101 %
1'
b101 +
#926430000000
1"
1(
#926440000000
0!
0"
b100 &
0'
0(
b100 ,
#926450000000
1!
b110 %
1'
b110 +
#926460000000
0!
0'
#926470000000
1!
b111 %
1'
b111 +
#926480000000
0!
0'
#926490000000
1!
0$
b1000 %
1'
0*
b1000 +
#926500000000
0!
0'
#926510000000
1!
b1001 %
1'
b1001 +
#926520000000
0!
0'
#926530000000
1!
b0 %
1'
b0 +
#926540000000
0!
0'
#926550000000
1!
1$
b1 %
1'
1*
b1 +
#926560000000
0!
0'
#926570000000
1!
b10 %
1'
b10 +
#926580000000
0!
0'
#926590000000
1!
b11 %
1'
b11 +
#926600000000
0!
0'
#926610000000
1!
b100 %
1'
b100 +
#926620000000
0!
0'
#926630000000
1!
b101 %
1'
b101 +
#926640000000
0!
0'
#926650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#926660000000
0!
0'
#926670000000
1!
b111 %
1'
b111 +
#926680000000
0!
0'
#926690000000
1!
b1000 %
1'
b1000 +
#926700000000
0!
0'
#926710000000
1!
b1001 %
1'
b1001 +
#926720000000
0!
0'
#926730000000
1!
b0 %
1'
b0 +
#926740000000
0!
0'
#926750000000
1!
1$
b1 %
1'
1*
b1 +
#926760000000
0!
0'
#926770000000
1!
b10 %
1'
b10 +
#926780000000
0!
0'
#926790000000
1!
b11 %
1'
b11 +
#926800000000
0!
0'
#926810000000
1!
b100 %
1'
b100 +
#926820000000
0!
0'
#926830000000
1!
b101 %
1'
b101 +
#926840000000
0!
0'
#926850000000
1!
0$
b110 %
1'
0*
b110 +
#926860000000
1"
1(
#926870000000
0!
0"
b100 &
0'
0(
b100 ,
#926880000000
1!
1$
b111 %
1'
1*
b111 +
#926890000000
0!
0'
#926900000000
1!
0$
b1000 %
1'
0*
b1000 +
#926910000000
0!
0'
#926920000000
1!
b1001 %
1'
b1001 +
#926930000000
0!
0'
#926940000000
1!
b0 %
1'
b0 +
#926950000000
0!
0'
#926960000000
1!
1$
b1 %
1'
1*
b1 +
#926970000000
0!
0'
#926980000000
1!
b10 %
1'
b10 +
#926990000000
0!
0'
#927000000000
1!
b11 %
1'
b11 +
#927010000000
0!
0'
#927020000000
1!
b100 %
1'
b100 +
#927030000000
0!
0'
#927040000000
1!
b101 %
1'
b101 +
#927050000000
0!
0'
#927060000000
1!
b110 %
1'
b110 +
#927070000000
0!
0'
#927080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#927090000000
0!
0'
#927100000000
1!
b1000 %
1'
b1000 +
#927110000000
0!
0'
#927120000000
1!
b1001 %
1'
b1001 +
#927130000000
0!
0'
#927140000000
1!
b0 %
1'
b0 +
#927150000000
0!
0'
#927160000000
1!
1$
b1 %
1'
1*
b1 +
#927170000000
0!
0'
#927180000000
1!
b10 %
1'
b10 +
#927190000000
0!
0'
#927200000000
1!
b11 %
1'
b11 +
#927210000000
0!
0'
#927220000000
1!
b100 %
1'
b100 +
#927230000000
0!
0'
#927240000000
1!
b101 %
1'
b101 +
#927250000000
0!
0'
#927260000000
1!
0$
b110 %
1'
0*
b110 +
#927270000000
0!
0'
#927280000000
1!
b111 %
1'
b111 +
#927290000000
1"
1(
#927300000000
0!
0"
b100 &
0'
0(
b100 ,
#927310000000
1!
b1000 %
1'
b1000 +
#927320000000
0!
0'
#927330000000
1!
b1001 %
1'
b1001 +
#927340000000
0!
0'
#927350000000
1!
b0 %
1'
b0 +
#927360000000
0!
0'
#927370000000
1!
1$
b1 %
1'
1*
b1 +
#927380000000
0!
0'
#927390000000
1!
b10 %
1'
b10 +
#927400000000
0!
0'
#927410000000
1!
b11 %
1'
b11 +
#927420000000
0!
0'
#927430000000
1!
b100 %
1'
b100 +
#927440000000
0!
0'
#927450000000
1!
b101 %
1'
b101 +
#927460000000
0!
0'
#927470000000
1!
b110 %
1'
b110 +
#927480000000
0!
0'
#927490000000
1!
b111 %
1'
b111 +
#927500000000
0!
0'
#927510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#927520000000
0!
0'
#927530000000
1!
b1001 %
1'
b1001 +
#927540000000
0!
0'
#927550000000
1!
b0 %
1'
b0 +
#927560000000
0!
0'
#927570000000
1!
1$
b1 %
1'
1*
b1 +
#927580000000
0!
0'
#927590000000
1!
b10 %
1'
b10 +
#927600000000
0!
0'
#927610000000
1!
b11 %
1'
b11 +
#927620000000
0!
0'
#927630000000
1!
b100 %
1'
b100 +
#927640000000
0!
0'
#927650000000
1!
b101 %
1'
b101 +
#927660000000
0!
0'
#927670000000
1!
0$
b110 %
1'
0*
b110 +
#927680000000
0!
0'
#927690000000
1!
b111 %
1'
b111 +
#927700000000
0!
0'
#927710000000
1!
b1000 %
1'
b1000 +
#927720000000
1"
1(
#927730000000
0!
0"
b100 &
0'
0(
b100 ,
#927740000000
1!
b1001 %
1'
b1001 +
#927750000000
0!
0'
#927760000000
1!
b0 %
1'
b0 +
#927770000000
0!
0'
#927780000000
1!
1$
b1 %
1'
1*
b1 +
#927790000000
0!
0'
#927800000000
1!
b10 %
1'
b10 +
#927810000000
0!
0'
#927820000000
1!
b11 %
1'
b11 +
#927830000000
0!
0'
#927840000000
1!
b100 %
1'
b100 +
#927850000000
0!
0'
#927860000000
1!
b101 %
1'
b101 +
#927870000000
0!
0'
#927880000000
1!
b110 %
1'
b110 +
#927890000000
0!
0'
#927900000000
1!
b111 %
1'
b111 +
#927910000000
0!
0'
#927920000000
1!
0$
b1000 %
1'
0*
b1000 +
#927930000000
0!
0'
#927940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#927950000000
0!
0'
#927960000000
1!
b0 %
1'
b0 +
#927970000000
0!
0'
#927980000000
1!
1$
b1 %
1'
1*
b1 +
#927990000000
0!
0'
#928000000000
1!
b10 %
1'
b10 +
#928010000000
0!
0'
#928020000000
1!
b11 %
1'
b11 +
#928030000000
0!
0'
#928040000000
1!
b100 %
1'
b100 +
#928050000000
0!
0'
#928060000000
1!
b101 %
1'
b101 +
#928070000000
0!
0'
#928080000000
1!
0$
b110 %
1'
0*
b110 +
#928090000000
0!
0'
#928100000000
1!
b111 %
1'
b111 +
#928110000000
0!
0'
#928120000000
1!
b1000 %
1'
b1000 +
#928130000000
0!
0'
#928140000000
1!
b1001 %
1'
b1001 +
#928150000000
1"
1(
#928160000000
0!
0"
b100 &
0'
0(
b100 ,
#928170000000
1!
b0 %
1'
b0 +
#928180000000
0!
0'
#928190000000
1!
1$
b1 %
1'
1*
b1 +
#928200000000
0!
0'
#928210000000
1!
b10 %
1'
b10 +
#928220000000
0!
0'
#928230000000
1!
b11 %
1'
b11 +
#928240000000
0!
0'
#928250000000
1!
b100 %
1'
b100 +
#928260000000
0!
0'
#928270000000
1!
b101 %
1'
b101 +
#928280000000
0!
0'
#928290000000
1!
b110 %
1'
b110 +
#928300000000
0!
0'
#928310000000
1!
b111 %
1'
b111 +
#928320000000
0!
0'
#928330000000
1!
0$
b1000 %
1'
0*
b1000 +
#928340000000
0!
0'
#928350000000
1!
b1001 %
1'
b1001 +
#928360000000
0!
0'
#928370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#928380000000
0!
0'
#928390000000
1!
1$
b1 %
1'
1*
b1 +
#928400000000
0!
0'
#928410000000
1!
b10 %
1'
b10 +
#928420000000
0!
0'
#928430000000
1!
b11 %
1'
b11 +
#928440000000
0!
0'
#928450000000
1!
b100 %
1'
b100 +
#928460000000
0!
0'
#928470000000
1!
b101 %
1'
b101 +
#928480000000
0!
0'
#928490000000
1!
0$
b110 %
1'
0*
b110 +
#928500000000
0!
0'
#928510000000
1!
b111 %
1'
b111 +
#928520000000
0!
0'
#928530000000
1!
b1000 %
1'
b1000 +
#928540000000
0!
0'
#928550000000
1!
b1001 %
1'
b1001 +
#928560000000
0!
0'
#928570000000
1!
b0 %
1'
b0 +
#928580000000
1"
1(
#928590000000
0!
0"
b100 &
0'
0(
b100 ,
#928600000000
1!
1$
b1 %
1'
1*
b1 +
#928610000000
0!
0'
#928620000000
1!
b10 %
1'
b10 +
#928630000000
0!
0'
#928640000000
1!
b11 %
1'
b11 +
#928650000000
0!
0'
#928660000000
1!
b100 %
1'
b100 +
#928670000000
0!
0'
#928680000000
1!
b101 %
1'
b101 +
#928690000000
0!
0'
#928700000000
1!
b110 %
1'
b110 +
#928710000000
0!
0'
#928720000000
1!
b111 %
1'
b111 +
#928730000000
0!
0'
#928740000000
1!
0$
b1000 %
1'
0*
b1000 +
#928750000000
0!
0'
#928760000000
1!
b1001 %
1'
b1001 +
#928770000000
0!
0'
#928780000000
1!
b0 %
1'
b0 +
#928790000000
0!
0'
#928800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#928810000000
0!
0'
#928820000000
1!
b10 %
1'
b10 +
#928830000000
0!
0'
#928840000000
1!
b11 %
1'
b11 +
#928850000000
0!
0'
#928860000000
1!
b100 %
1'
b100 +
#928870000000
0!
0'
#928880000000
1!
b101 %
1'
b101 +
#928890000000
0!
0'
#928900000000
1!
0$
b110 %
1'
0*
b110 +
#928910000000
0!
0'
#928920000000
1!
b111 %
1'
b111 +
#928930000000
0!
0'
#928940000000
1!
b1000 %
1'
b1000 +
#928950000000
0!
0'
#928960000000
1!
b1001 %
1'
b1001 +
#928970000000
0!
0'
#928980000000
1!
b0 %
1'
b0 +
#928990000000
0!
0'
#929000000000
1!
1$
b1 %
1'
1*
b1 +
#929010000000
1"
1(
#929020000000
0!
0"
b100 &
0'
0(
b100 ,
#929030000000
1!
b10 %
1'
b10 +
#929040000000
0!
0'
#929050000000
1!
b11 %
1'
b11 +
#929060000000
0!
0'
#929070000000
1!
b100 %
1'
b100 +
#929080000000
0!
0'
#929090000000
1!
b101 %
1'
b101 +
#929100000000
0!
0'
#929110000000
1!
b110 %
1'
b110 +
#929120000000
0!
0'
#929130000000
1!
b111 %
1'
b111 +
#929140000000
0!
0'
#929150000000
1!
0$
b1000 %
1'
0*
b1000 +
#929160000000
0!
0'
#929170000000
1!
b1001 %
1'
b1001 +
#929180000000
0!
0'
#929190000000
1!
b0 %
1'
b0 +
#929200000000
0!
0'
#929210000000
1!
1$
b1 %
1'
1*
b1 +
#929220000000
0!
0'
#929230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#929240000000
0!
0'
#929250000000
1!
b11 %
1'
b11 +
#929260000000
0!
0'
#929270000000
1!
b100 %
1'
b100 +
#929280000000
0!
0'
#929290000000
1!
b101 %
1'
b101 +
#929300000000
0!
0'
#929310000000
1!
0$
b110 %
1'
0*
b110 +
#929320000000
0!
0'
#929330000000
1!
b111 %
1'
b111 +
#929340000000
0!
0'
#929350000000
1!
b1000 %
1'
b1000 +
#929360000000
0!
0'
#929370000000
1!
b1001 %
1'
b1001 +
#929380000000
0!
0'
#929390000000
1!
b0 %
1'
b0 +
#929400000000
0!
0'
#929410000000
1!
1$
b1 %
1'
1*
b1 +
#929420000000
0!
0'
#929430000000
1!
b10 %
1'
b10 +
#929440000000
1"
1(
#929450000000
0!
0"
b100 &
0'
0(
b100 ,
#929460000000
1!
b11 %
1'
b11 +
#929470000000
0!
0'
#929480000000
1!
b100 %
1'
b100 +
#929490000000
0!
0'
#929500000000
1!
b101 %
1'
b101 +
#929510000000
0!
0'
#929520000000
1!
b110 %
1'
b110 +
#929530000000
0!
0'
#929540000000
1!
b111 %
1'
b111 +
#929550000000
0!
0'
#929560000000
1!
0$
b1000 %
1'
0*
b1000 +
#929570000000
0!
0'
#929580000000
1!
b1001 %
1'
b1001 +
#929590000000
0!
0'
#929600000000
1!
b0 %
1'
b0 +
#929610000000
0!
0'
#929620000000
1!
1$
b1 %
1'
1*
b1 +
#929630000000
0!
0'
#929640000000
1!
b10 %
1'
b10 +
#929650000000
0!
0'
#929660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#929670000000
0!
0'
#929680000000
1!
b100 %
1'
b100 +
#929690000000
0!
0'
#929700000000
1!
b101 %
1'
b101 +
#929710000000
0!
0'
#929720000000
1!
0$
b110 %
1'
0*
b110 +
#929730000000
0!
0'
#929740000000
1!
b111 %
1'
b111 +
#929750000000
0!
0'
#929760000000
1!
b1000 %
1'
b1000 +
#929770000000
0!
0'
#929780000000
1!
b1001 %
1'
b1001 +
#929790000000
0!
0'
#929800000000
1!
b0 %
1'
b0 +
#929810000000
0!
0'
#929820000000
1!
1$
b1 %
1'
1*
b1 +
#929830000000
0!
0'
#929840000000
1!
b10 %
1'
b10 +
#929850000000
0!
0'
#929860000000
1!
b11 %
1'
b11 +
#929870000000
1"
1(
#929880000000
0!
0"
b100 &
0'
0(
b100 ,
#929890000000
1!
b100 %
1'
b100 +
#929900000000
0!
0'
#929910000000
1!
b101 %
1'
b101 +
#929920000000
0!
0'
#929930000000
1!
b110 %
1'
b110 +
#929940000000
0!
0'
#929950000000
1!
b111 %
1'
b111 +
#929960000000
0!
0'
#929970000000
1!
0$
b1000 %
1'
0*
b1000 +
#929980000000
0!
0'
#929990000000
1!
b1001 %
1'
b1001 +
#930000000000
0!
0'
#930010000000
1!
b0 %
1'
b0 +
#930020000000
0!
0'
#930030000000
1!
1$
b1 %
1'
1*
b1 +
#930040000000
0!
0'
#930050000000
1!
b10 %
1'
b10 +
#930060000000
0!
0'
#930070000000
1!
b11 %
1'
b11 +
#930080000000
0!
0'
#930090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#930100000000
0!
0'
#930110000000
1!
b101 %
1'
b101 +
#930120000000
0!
0'
#930130000000
1!
0$
b110 %
1'
0*
b110 +
#930140000000
0!
0'
#930150000000
1!
b111 %
1'
b111 +
#930160000000
0!
0'
#930170000000
1!
b1000 %
1'
b1000 +
#930180000000
0!
0'
#930190000000
1!
b1001 %
1'
b1001 +
#930200000000
0!
0'
#930210000000
1!
b0 %
1'
b0 +
#930220000000
0!
0'
#930230000000
1!
1$
b1 %
1'
1*
b1 +
#930240000000
0!
0'
#930250000000
1!
b10 %
1'
b10 +
#930260000000
0!
0'
#930270000000
1!
b11 %
1'
b11 +
#930280000000
0!
0'
#930290000000
1!
b100 %
1'
b100 +
#930300000000
1"
1(
#930310000000
0!
0"
b100 &
0'
0(
b100 ,
#930320000000
1!
b101 %
1'
b101 +
#930330000000
0!
0'
#930340000000
1!
b110 %
1'
b110 +
#930350000000
0!
0'
#930360000000
1!
b111 %
1'
b111 +
#930370000000
0!
0'
#930380000000
1!
0$
b1000 %
1'
0*
b1000 +
#930390000000
0!
0'
#930400000000
1!
b1001 %
1'
b1001 +
#930410000000
0!
0'
#930420000000
1!
b0 %
1'
b0 +
#930430000000
0!
0'
#930440000000
1!
1$
b1 %
1'
1*
b1 +
#930450000000
0!
0'
#930460000000
1!
b10 %
1'
b10 +
#930470000000
0!
0'
#930480000000
1!
b11 %
1'
b11 +
#930490000000
0!
0'
#930500000000
1!
b100 %
1'
b100 +
#930510000000
0!
0'
#930520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#930530000000
0!
0'
#930540000000
1!
0$
b110 %
1'
0*
b110 +
#930550000000
0!
0'
#930560000000
1!
b111 %
1'
b111 +
#930570000000
0!
0'
#930580000000
1!
b1000 %
1'
b1000 +
#930590000000
0!
0'
#930600000000
1!
b1001 %
1'
b1001 +
#930610000000
0!
0'
#930620000000
1!
b0 %
1'
b0 +
#930630000000
0!
0'
#930640000000
1!
1$
b1 %
1'
1*
b1 +
#930650000000
0!
0'
#930660000000
1!
b10 %
1'
b10 +
#930670000000
0!
0'
#930680000000
1!
b11 %
1'
b11 +
#930690000000
0!
0'
#930700000000
1!
b100 %
1'
b100 +
#930710000000
0!
0'
#930720000000
1!
b101 %
1'
b101 +
#930730000000
1"
1(
#930740000000
0!
0"
b100 &
0'
0(
b100 ,
#930750000000
1!
b110 %
1'
b110 +
#930760000000
0!
0'
#930770000000
1!
b111 %
1'
b111 +
#930780000000
0!
0'
#930790000000
1!
0$
b1000 %
1'
0*
b1000 +
#930800000000
0!
0'
#930810000000
1!
b1001 %
1'
b1001 +
#930820000000
0!
0'
#930830000000
1!
b0 %
1'
b0 +
#930840000000
0!
0'
#930850000000
1!
1$
b1 %
1'
1*
b1 +
#930860000000
0!
0'
#930870000000
1!
b10 %
1'
b10 +
#930880000000
0!
0'
#930890000000
1!
b11 %
1'
b11 +
#930900000000
0!
0'
#930910000000
1!
b100 %
1'
b100 +
#930920000000
0!
0'
#930930000000
1!
b101 %
1'
b101 +
#930940000000
0!
0'
#930950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#930960000000
0!
0'
#930970000000
1!
b111 %
1'
b111 +
#930980000000
0!
0'
#930990000000
1!
b1000 %
1'
b1000 +
#931000000000
0!
0'
#931010000000
1!
b1001 %
1'
b1001 +
#931020000000
0!
0'
#931030000000
1!
b0 %
1'
b0 +
#931040000000
0!
0'
#931050000000
1!
1$
b1 %
1'
1*
b1 +
#931060000000
0!
0'
#931070000000
1!
b10 %
1'
b10 +
#931080000000
0!
0'
#931090000000
1!
b11 %
1'
b11 +
#931100000000
0!
0'
#931110000000
1!
b100 %
1'
b100 +
#931120000000
0!
0'
#931130000000
1!
b101 %
1'
b101 +
#931140000000
0!
0'
#931150000000
1!
0$
b110 %
1'
0*
b110 +
#931160000000
1"
1(
#931170000000
0!
0"
b100 &
0'
0(
b100 ,
#931180000000
1!
1$
b111 %
1'
1*
b111 +
#931190000000
0!
0'
#931200000000
1!
0$
b1000 %
1'
0*
b1000 +
#931210000000
0!
0'
#931220000000
1!
b1001 %
1'
b1001 +
#931230000000
0!
0'
#931240000000
1!
b0 %
1'
b0 +
#931250000000
0!
0'
#931260000000
1!
1$
b1 %
1'
1*
b1 +
#931270000000
0!
0'
#931280000000
1!
b10 %
1'
b10 +
#931290000000
0!
0'
#931300000000
1!
b11 %
1'
b11 +
#931310000000
0!
0'
#931320000000
1!
b100 %
1'
b100 +
#931330000000
0!
0'
#931340000000
1!
b101 %
1'
b101 +
#931350000000
0!
0'
#931360000000
1!
b110 %
1'
b110 +
#931370000000
0!
0'
#931380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#931390000000
0!
0'
#931400000000
1!
b1000 %
1'
b1000 +
#931410000000
0!
0'
#931420000000
1!
b1001 %
1'
b1001 +
#931430000000
0!
0'
#931440000000
1!
b0 %
1'
b0 +
#931450000000
0!
0'
#931460000000
1!
1$
b1 %
1'
1*
b1 +
#931470000000
0!
0'
#931480000000
1!
b10 %
1'
b10 +
#931490000000
0!
0'
#931500000000
1!
b11 %
1'
b11 +
#931510000000
0!
0'
#931520000000
1!
b100 %
1'
b100 +
#931530000000
0!
0'
#931540000000
1!
b101 %
1'
b101 +
#931550000000
0!
0'
#931560000000
1!
0$
b110 %
1'
0*
b110 +
#931570000000
0!
0'
#931580000000
1!
b111 %
1'
b111 +
#931590000000
1"
1(
#931600000000
0!
0"
b100 &
0'
0(
b100 ,
#931610000000
1!
b1000 %
1'
b1000 +
#931620000000
0!
0'
#931630000000
1!
b1001 %
1'
b1001 +
#931640000000
0!
0'
#931650000000
1!
b0 %
1'
b0 +
#931660000000
0!
0'
#931670000000
1!
1$
b1 %
1'
1*
b1 +
#931680000000
0!
0'
#931690000000
1!
b10 %
1'
b10 +
#931700000000
0!
0'
#931710000000
1!
b11 %
1'
b11 +
#931720000000
0!
0'
#931730000000
1!
b100 %
1'
b100 +
#931740000000
0!
0'
#931750000000
1!
b101 %
1'
b101 +
#931760000000
0!
0'
#931770000000
1!
b110 %
1'
b110 +
#931780000000
0!
0'
#931790000000
1!
b111 %
1'
b111 +
#931800000000
0!
0'
#931810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#931820000000
0!
0'
#931830000000
1!
b1001 %
1'
b1001 +
#931840000000
0!
0'
#931850000000
1!
b0 %
1'
b0 +
#931860000000
0!
0'
#931870000000
1!
1$
b1 %
1'
1*
b1 +
#931880000000
0!
0'
#931890000000
1!
b10 %
1'
b10 +
#931900000000
0!
0'
#931910000000
1!
b11 %
1'
b11 +
#931920000000
0!
0'
#931930000000
1!
b100 %
1'
b100 +
#931940000000
0!
0'
#931950000000
1!
b101 %
1'
b101 +
#931960000000
0!
0'
#931970000000
1!
0$
b110 %
1'
0*
b110 +
#931980000000
0!
0'
#931990000000
1!
b111 %
1'
b111 +
#932000000000
0!
0'
#932010000000
1!
b1000 %
1'
b1000 +
#932020000000
1"
1(
#932030000000
0!
0"
b100 &
0'
0(
b100 ,
#932040000000
1!
b1001 %
1'
b1001 +
#932050000000
0!
0'
#932060000000
1!
b0 %
1'
b0 +
#932070000000
0!
0'
#932080000000
1!
1$
b1 %
1'
1*
b1 +
#932090000000
0!
0'
#932100000000
1!
b10 %
1'
b10 +
#932110000000
0!
0'
#932120000000
1!
b11 %
1'
b11 +
#932130000000
0!
0'
#932140000000
1!
b100 %
1'
b100 +
#932150000000
0!
0'
#932160000000
1!
b101 %
1'
b101 +
#932170000000
0!
0'
#932180000000
1!
b110 %
1'
b110 +
#932190000000
0!
0'
#932200000000
1!
b111 %
1'
b111 +
#932210000000
0!
0'
#932220000000
1!
0$
b1000 %
1'
0*
b1000 +
#932230000000
0!
0'
#932240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#932250000000
0!
0'
#932260000000
1!
b0 %
1'
b0 +
#932270000000
0!
0'
#932280000000
1!
1$
b1 %
1'
1*
b1 +
#932290000000
0!
0'
#932300000000
1!
b10 %
1'
b10 +
#932310000000
0!
0'
#932320000000
1!
b11 %
1'
b11 +
#932330000000
0!
0'
#932340000000
1!
b100 %
1'
b100 +
#932350000000
0!
0'
#932360000000
1!
b101 %
1'
b101 +
#932370000000
0!
0'
#932380000000
1!
0$
b110 %
1'
0*
b110 +
#932390000000
0!
0'
#932400000000
1!
b111 %
1'
b111 +
#932410000000
0!
0'
#932420000000
1!
b1000 %
1'
b1000 +
#932430000000
0!
0'
#932440000000
1!
b1001 %
1'
b1001 +
#932450000000
1"
1(
#932460000000
0!
0"
b100 &
0'
0(
b100 ,
#932470000000
1!
b0 %
1'
b0 +
#932480000000
0!
0'
#932490000000
1!
1$
b1 %
1'
1*
b1 +
#932500000000
0!
0'
#932510000000
1!
b10 %
1'
b10 +
#932520000000
0!
0'
#932530000000
1!
b11 %
1'
b11 +
#932540000000
0!
0'
#932550000000
1!
b100 %
1'
b100 +
#932560000000
0!
0'
#932570000000
1!
b101 %
1'
b101 +
#932580000000
0!
0'
#932590000000
1!
b110 %
1'
b110 +
#932600000000
0!
0'
#932610000000
1!
b111 %
1'
b111 +
#932620000000
0!
0'
#932630000000
1!
0$
b1000 %
1'
0*
b1000 +
#932640000000
0!
0'
#932650000000
1!
b1001 %
1'
b1001 +
#932660000000
0!
0'
#932670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#932680000000
0!
0'
#932690000000
1!
1$
b1 %
1'
1*
b1 +
#932700000000
0!
0'
#932710000000
1!
b10 %
1'
b10 +
#932720000000
0!
0'
#932730000000
1!
b11 %
1'
b11 +
#932740000000
0!
0'
#932750000000
1!
b100 %
1'
b100 +
#932760000000
0!
0'
#932770000000
1!
b101 %
1'
b101 +
#932780000000
0!
0'
#932790000000
1!
0$
b110 %
1'
0*
b110 +
#932800000000
0!
0'
#932810000000
1!
b111 %
1'
b111 +
#932820000000
0!
0'
#932830000000
1!
b1000 %
1'
b1000 +
#932840000000
0!
0'
#932850000000
1!
b1001 %
1'
b1001 +
#932860000000
0!
0'
#932870000000
1!
b0 %
1'
b0 +
#932880000000
1"
1(
#932890000000
0!
0"
b100 &
0'
0(
b100 ,
#932900000000
1!
1$
b1 %
1'
1*
b1 +
#932910000000
0!
0'
#932920000000
1!
b10 %
1'
b10 +
#932930000000
0!
0'
#932940000000
1!
b11 %
1'
b11 +
#932950000000
0!
0'
#932960000000
1!
b100 %
1'
b100 +
#932970000000
0!
0'
#932980000000
1!
b101 %
1'
b101 +
#932990000000
0!
0'
#933000000000
1!
b110 %
1'
b110 +
#933010000000
0!
0'
#933020000000
1!
b111 %
1'
b111 +
#933030000000
0!
0'
#933040000000
1!
0$
b1000 %
1'
0*
b1000 +
#933050000000
0!
0'
#933060000000
1!
b1001 %
1'
b1001 +
#933070000000
0!
0'
#933080000000
1!
b0 %
1'
b0 +
#933090000000
0!
0'
#933100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#933110000000
0!
0'
#933120000000
1!
b10 %
1'
b10 +
#933130000000
0!
0'
#933140000000
1!
b11 %
1'
b11 +
#933150000000
0!
0'
#933160000000
1!
b100 %
1'
b100 +
#933170000000
0!
0'
#933180000000
1!
b101 %
1'
b101 +
#933190000000
0!
0'
#933200000000
1!
0$
b110 %
1'
0*
b110 +
#933210000000
0!
0'
#933220000000
1!
b111 %
1'
b111 +
#933230000000
0!
0'
#933240000000
1!
b1000 %
1'
b1000 +
#933250000000
0!
0'
#933260000000
1!
b1001 %
1'
b1001 +
#933270000000
0!
0'
#933280000000
1!
b0 %
1'
b0 +
#933290000000
0!
0'
#933300000000
1!
1$
b1 %
1'
1*
b1 +
#933310000000
1"
1(
#933320000000
0!
0"
b100 &
0'
0(
b100 ,
#933330000000
1!
b10 %
1'
b10 +
#933340000000
0!
0'
#933350000000
1!
b11 %
1'
b11 +
#933360000000
0!
0'
#933370000000
1!
b100 %
1'
b100 +
#933380000000
0!
0'
#933390000000
1!
b101 %
1'
b101 +
#933400000000
0!
0'
#933410000000
1!
b110 %
1'
b110 +
#933420000000
0!
0'
#933430000000
1!
b111 %
1'
b111 +
#933440000000
0!
0'
#933450000000
1!
0$
b1000 %
1'
0*
b1000 +
#933460000000
0!
0'
#933470000000
1!
b1001 %
1'
b1001 +
#933480000000
0!
0'
#933490000000
1!
b0 %
1'
b0 +
#933500000000
0!
0'
#933510000000
1!
1$
b1 %
1'
1*
b1 +
#933520000000
0!
0'
#933530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#933540000000
0!
0'
#933550000000
1!
b11 %
1'
b11 +
#933560000000
0!
0'
#933570000000
1!
b100 %
1'
b100 +
#933580000000
0!
0'
#933590000000
1!
b101 %
1'
b101 +
#933600000000
0!
0'
#933610000000
1!
0$
b110 %
1'
0*
b110 +
#933620000000
0!
0'
#933630000000
1!
b111 %
1'
b111 +
#933640000000
0!
0'
#933650000000
1!
b1000 %
1'
b1000 +
#933660000000
0!
0'
#933670000000
1!
b1001 %
1'
b1001 +
#933680000000
0!
0'
#933690000000
1!
b0 %
1'
b0 +
#933700000000
0!
0'
#933710000000
1!
1$
b1 %
1'
1*
b1 +
#933720000000
0!
0'
#933730000000
1!
b10 %
1'
b10 +
#933740000000
1"
1(
#933750000000
0!
0"
b100 &
0'
0(
b100 ,
#933760000000
1!
b11 %
1'
b11 +
#933770000000
0!
0'
#933780000000
1!
b100 %
1'
b100 +
#933790000000
0!
0'
#933800000000
1!
b101 %
1'
b101 +
#933810000000
0!
0'
#933820000000
1!
b110 %
1'
b110 +
#933830000000
0!
0'
#933840000000
1!
b111 %
1'
b111 +
#933850000000
0!
0'
#933860000000
1!
0$
b1000 %
1'
0*
b1000 +
#933870000000
0!
0'
#933880000000
1!
b1001 %
1'
b1001 +
#933890000000
0!
0'
#933900000000
1!
b0 %
1'
b0 +
#933910000000
0!
0'
#933920000000
1!
1$
b1 %
1'
1*
b1 +
#933930000000
0!
0'
#933940000000
1!
b10 %
1'
b10 +
#933950000000
0!
0'
#933960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#933970000000
0!
0'
#933980000000
1!
b100 %
1'
b100 +
#933990000000
0!
0'
#934000000000
1!
b101 %
1'
b101 +
#934010000000
0!
0'
#934020000000
1!
0$
b110 %
1'
0*
b110 +
#934030000000
0!
0'
#934040000000
1!
b111 %
1'
b111 +
#934050000000
0!
0'
#934060000000
1!
b1000 %
1'
b1000 +
#934070000000
0!
0'
#934080000000
1!
b1001 %
1'
b1001 +
#934090000000
0!
0'
#934100000000
1!
b0 %
1'
b0 +
#934110000000
0!
0'
#934120000000
1!
1$
b1 %
1'
1*
b1 +
#934130000000
0!
0'
#934140000000
1!
b10 %
1'
b10 +
#934150000000
0!
0'
#934160000000
1!
b11 %
1'
b11 +
#934170000000
1"
1(
#934180000000
0!
0"
b100 &
0'
0(
b100 ,
#934190000000
1!
b100 %
1'
b100 +
#934200000000
0!
0'
#934210000000
1!
b101 %
1'
b101 +
#934220000000
0!
0'
#934230000000
1!
b110 %
1'
b110 +
#934240000000
0!
0'
#934250000000
1!
b111 %
1'
b111 +
#934260000000
0!
0'
#934270000000
1!
0$
b1000 %
1'
0*
b1000 +
#934280000000
0!
0'
#934290000000
1!
b1001 %
1'
b1001 +
#934300000000
0!
0'
#934310000000
1!
b0 %
1'
b0 +
#934320000000
0!
0'
#934330000000
1!
1$
b1 %
1'
1*
b1 +
#934340000000
0!
0'
#934350000000
1!
b10 %
1'
b10 +
#934360000000
0!
0'
#934370000000
1!
b11 %
1'
b11 +
#934380000000
0!
0'
#934390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#934400000000
0!
0'
#934410000000
1!
b101 %
1'
b101 +
#934420000000
0!
0'
#934430000000
1!
0$
b110 %
1'
0*
b110 +
#934440000000
0!
0'
#934450000000
1!
b111 %
1'
b111 +
#934460000000
0!
0'
#934470000000
1!
b1000 %
1'
b1000 +
#934480000000
0!
0'
#934490000000
1!
b1001 %
1'
b1001 +
#934500000000
0!
0'
#934510000000
1!
b0 %
1'
b0 +
#934520000000
0!
0'
#934530000000
1!
1$
b1 %
1'
1*
b1 +
#934540000000
0!
0'
#934550000000
1!
b10 %
1'
b10 +
#934560000000
0!
0'
#934570000000
1!
b11 %
1'
b11 +
#934580000000
0!
0'
#934590000000
1!
b100 %
1'
b100 +
#934600000000
1"
1(
#934610000000
0!
0"
b100 &
0'
0(
b100 ,
#934620000000
1!
b101 %
1'
b101 +
#934630000000
0!
0'
#934640000000
1!
b110 %
1'
b110 +
#934650000000
0!
0'
#934660000000
1!
b111 %
1'
b111 +
#934670000000
0!
0'
#934680000000
1!
0$
b1000 %
1'
0*
b1000 +
#934690000000
0!
0'
#934700000000
1!
b1001 %
1'
b1001 +
#934710000000
0!
0'
#934720000000
1!
b0 %
1'
b0 +
#934730000000
0!
0'
#934740000000
1!
1$
b1 %
1'
1*
b1 +
#934750000000
0!
0'
#934760000000
1!
b10 %
1'
b10 +
#934770000000
0!
0'
#934780000000
1!
b11 %
1'
b11 +
#934790000000
0!
0'
#934800000000
1!
b100 %
1'
b100 +
#934810000000
0!
0'
#934820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#934830000000
0!
0'
#934840000000
1!
0$
b110 %
1'
0*
b110 +
#934850000000
0!
0'
#934860000000
1!
b111 %
1'
b111 +
#934870000000
0!
0'
#934880000000
1!
b1000 %
1'
b1000 +
#934890000000
0!
0'
#934900000000
1!
b1001 %
1'
b1001 +
#934910000000
0!
0'
#934920000000
1!
b0 %
1'
b0 +
#934930000000
0!
0'
#934940000000
1!
1$
b1 %
1'
1*
b1 +
#934950000000
0!
0'
#934960000000
1!
b10 %
1'
b10 +
#934970000000
0!
0'
#934980000000
1!
b11 %
1'
b11 +
#934990000000
0!
0'
#935000000000
1!
b100 %
1'
b100 +
#935010000000
0!
0'
#935020000000
1!
b101 %
1'
b101 +
#935030000000
1"
1(
#935040000000
0!
0"
b100 &
0'
0(
b100 ,
#935050000000
1!
b110 %
1'
b110 +
#935060000000
0!
0'
#935070000000
1!
b111 %
1'
b111 +
#935080000000
0!
0'
#935090000000
1!
0$
b1000 %
1'
0*
b1000 +
#935100000000
0!
0'
#935110000000
1!
b1001 %
1'
b1001 +
#935120000000
0!
0'
#935130000000
1!
b0 %
1'
b0 +
#935140000000
0!
0'
#935150000000
1!
1$
b1 %
1'
1*
b1 +
#935160000000
0!
0'
#935170000000
1!
b10 %
1'
b10 +
#935180000000
0!
0'
#935190000000
1!
b11 %
1'
b11 +
#935200000000
0!
0'
#935210000000
1!
b100 %
1'
b100 +
#935220000000
0!
0'
#935230000000
1!
b101 %
1'
b101 +
#935240000000
0!
0'
#935250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#935260000000
0!
0'
#935270000000
1!
b111 %
1'
b111 +
#935280000000
0!
0'
#935290000000
1!
b1000 %
1'
b1000 +
#935300000000
0!
0'
#935310000000
1!
b1001 %
1'
b1001 +
#935320000000
0!
0'
#935330000000
1!
b0 %
1'
b0 +
#935340000000
0!
0'
#935350000000
1!
1$
b1 %
1'
1*
b1 +
#935360000000
0!
0'
#935370000000
1!
b10 %
1'
b10 +
#935380000000
0!
0'
#935390000000
1!
b11 %
1'
b11 +
#935400000000
0!
0'
#935410000000
1!
b100 %
1'
b100 +
#935420000000
0!
0'
#935430000000
1!
b101 %
1'
b101 +
#935440000000
0!
0'
#935450000000
1!
0$
b110 %
1'
0*
b110 +
#935460000000
1"
1(
#935470000000
0!
0"
b100 &
0'
0(
b100 ,
#935480000000
1!
1$
b111 %
1'
1*
b111 +
#935490000000
0!
0'
#935500000000
1!
0$
b1000 %
1'
0*
b1000 +
#935510000000
0!
0'
#935520000000
1!
b1001 %
1'
b1001 +
#935530000000
0!
0'
#935540000000
1!
b0 %
1'
b0 +
#935550000000
0!
0'
#935560000000
1!
1$
b1 %
1'
1*
b1 +
#935570000000
0!
0'
#935580000000
1!
b10 %
1'
b10 +
#935590000000
0!
0'
#935600000000
1!
b11 %
1'
b11 +
#935610000000
0!
0'
#935620000000
1!
b100 %
1'
b100 +
#935630000000
0!
0'
#935640000000
1!
b101 %
1'
b101 +
#935650000000
0!
0'
#935660000000
1!
b110 %
1'
b110 +
#935670000000
0!
0'
#935680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#935690000000
0!
0'
#935700000000
1!
b1000 %
1'
b1000 +
#935710000000
0!
0'
#935720000000
1!
b1001 %
1'
b1001 +
#935730000000
0!
0'
#935740000000
1!
b0 %
1'
b0 +
#935750000000
0!
0'
#935760000000
1!
1$
b1 %
1'
1*
b1 +
#935770000000
0!
0'
#935780000000
1!
b10 %
1'
b10 +
#935790000000
0!
0'
#935800000000
1!
b11 %
1'
b11 +
#935810000000
0!
0'
#935820000000
1!
b100 %
1'
b100 +
#935830000000
0!
0'
#935840000000
1!
b101 %
1'
b101 +
#935850000000
0!
0'
#935860000000
1!
0$
b110 %
1'
0*
b110 +
#935870000000
0!
0'
#935880000000
1!
b111 %
1'
b111 +
#935890000000
1"
1(
#935900000000
0!
0"
b100 &
0'
0(
b100 ,
#935910000000
1!
b1000 %
1'
b1000 +
#935920000000
0!
0'
#935930000000
1!
b1001 %
1'
b1001 +
#935940000000
0!
0'
#935950000000
1!
b0 %
1'
b0 +
#935960000000
0!
0'
#935970000000
1!
1$
b1 %
1'
1*
b1 +
#935980000000
0!
0'
#935990000000
1!
b10 %
1'
b10 +
#936000000000
0!
0'
#936010000000
1!
b11 %
1'
b11 +
#936020000000
0!
0'
#936030000000
1!
b100 %
1'
b100 +
#936040000000
0!
0'
#936050000000
1!
b101 %
1'
b101 +
#936060000000
0!
0'
#936070000000
1!
b110 %
1'
b110 +
#936080000000
0!
0'
#936090000000
1!
b111 %
1'
b111 +
#936100000000
0!
0'
#936110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#936120000000
0!
0'
#936130000000
1!
b1001 %
1'
b1001 +
#936140000000
0!
0'
#936150000000
1!
b0 %
1'
b0 +
#936160000000
0!
0'
#936170000000
1!
1$
b1 %
1'
1*
b1 +
#936180000000
0!
0'
#936190000000
1!
b10 %
1'
b10 +
#936200000000
0!
0'
#936210000000
1!
b11 %
1'
b11 +
#936220000000
0!
0'
#936230000000
1!
b100 %
1'
b100 +
#936240000000
0!
0'
#936250000000
1!
b101 %
1'
b101 +
#936260000000
0!
0'
#936270000000
1!
0$
b110 %
1'
0*
b110 +
#936280000000
0!
0'
#936290000000
1!
b111 %
1'
b111 +
#936300000000
0!
0'
#936310000000
1!
b1000 %
1'
b1000 +
#936320000000
1"
1(
#936330000000
0!
0"
b100 &
0'
0(
b100 ,
#936340000000
1!
b1001 %
1'
b1001 +
#936350000000
0!
0'
#936360000000
1!
b0 %
1'
b0 +
#936370000000
0!
0'
#936380000000
1!
1$
b1 %
1'
1*
b1 +
#936390000000
0!
0'
#936400000000
1!
b10 %
1'
b10 +
#936410000000
0!
0'
#936420000000
1!
b11 %
1'
b11 +
#936430000000
0!
0'
#936440000000
1!
b100 %
1'
b100 +
#936450000000
0!
0'
#936460000000
1!
b101 %
1'
b101 +
#936470000000
0!
0'
#936480000000
1!
b110 %
1'
b110 +
#936490000000
0!
0'
#936500000000
1!
b111 %
1'
b111 +
#936510000000
0!
0'
#936520000000
1!
0$
b1000 %
1'
0*
b1000 +
#936530000000
0!
0'
#936540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#936550000000
0!
0'
#936560000000
1!
b0 %
1'
b0 +
#936570000000
0!
0'
#936580000000
1!
1$
b1 %
1'
1*
b1 +
#936590000000
0!
0'
#936600000000
1!
b10 %
1'
b10 +
#936610000000
0!
0'
#936620000000
1!
b11 %
1'
b11 +
#936630000000
0!
0'
#936640000000
1!
b100 %
1'
b100 +
#936650000000
0!
0'
#936660000000
1!
b101 %
1'
b101 +
#936670000000
0!
0'
#936680000000
1!
0$
b110 %
1'
0*
b110 +
#936690000000
0!
0'
#936700000000
1!
b111 %
1'
b111 +
#936710000000
0!
0'
#936720000000
1!
b1000 %
1'
b1000 +
#936730000000
0!
0'
#936740000000
1!
b1001 %
1'
b1001 +
#936750000000
1"
1(
#936760000000
0!
0"
b100 &
0'
0(
b100 ,
#936770000000
1!
b0 %
1'
b0 +
#936780000000
0!
0'
#936790000000
1!
1$
b1 %
1'
1*
b1 +
#936800000000
0!
0'
#936810000000
1!
b10 %
1'
b10 +
#936820000000
0!
0'
#936830000000
1!
b11 %
1'
b11 +
#936840000000
0!
0'
#936850000000
1!
b100 %
1'
b100 +
#936860000000
0!
0'
#936870000000
1!
b101 %
1'
b101 +
#936880000000
0!
0'
#936890000000
1!
b110 %
1'
b110 +
#936900000000
0!
0'
#936910000000
1!
b111 %
1'
b111 +
#936920000000
0!
0'
#936930000000
1!
0$
b1000 %
1'
0*
b1000 +
#936940000000
0!
0'
#936950000000
1!
b1001 %
1'
b1001 +
#936960000000
0!
0'
#936970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#936980000000
0!
0'
#936990000000
1!
1$
b1 %
1'
1*
b1 +
#937000000000
0!
0'
#937010000000
1!
b10 %
1'
b10 +
#937020000000
0!
0'
#937030000000
1!
b11 %
1'
b11 +
#937040000000
0!
0'
#937050000000
1!
b100 %
1'
b100 +
#937060000000
0!
0'
#937070000000
1!
b101 %
1'
b101 +
#937080000000
0!
0'
#937090000000
1!
0$
b110 %
1'
0*
b110 +
#937100000000
0!
0'
#937110000000
1!
b111 %
1'
b111 +
#937120000000
0!
0'
#937130000000
1!
b1000 %
1'
b1000 +
#937140000000
0!
0'
#937150000000
1!
b1001 %
1'
b1001 +
#937160000000
0!
0'
#937170000000
1!
b0 %
1'
b0 +
#937180000000
1"
1(
#937190000000
0!
0"
b100 &
0'
0(
b100 ,
#937200000000
1!
1$
b1 %
1'
1*
b1 +
#937210000000
0!
0'
#937220000000
1!
b10 %
1'
b10 +
#937230000000
0!
0'
#937240000000
1!
b11 %
1'
b11 +
#937250000000
0!
0'
#937260000000
1!
b100 %
1'
b100 +
#937270000000
0!
0'
#937280000000
1!
b101 %
1'
b101 +
#937290000000
0!
0'
#937300000000
1!
b110 %
1'
b110 +
#937310000000
0!
0'
#937320000000
1!
b111 %
1'
b111 +
#937330000000
0!
0'
#937340000000
1!
0$
b1000 %
1'
0*
b1000 +
#937350000000
0!
0'
#937360000000
1!
b1001 %
1'
b1001 +
#937370000000
0!
0'
#937380000000
1!
b0 %
1'
b0 +
#937390000000
0!
0'
#937400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#937410000000
0!
0'
#937420000000
1!
b10 %
1'
b10 +
#937430000000
0!
0'
#937440000000
1!
b11 %
1'
b11 +
#937450000000
0!
0'
#937460000000
1!
b100 %
1'
b100 +
#937470000000
0!
0'
#937480000000
1!
b101 %
1'
b101 +
#937490000000
0!
0'
#937500000000
1!
0$
b110 %
1'
0*
b110 +
#937510000000
0!
0'
#937520000000
1!
b111 %
1'
b111 +
#937530000000
0!
0'
#937540000000
1!
b1000 %
1'
b1000 +
#937550000000
0!
0'
#937560000000
1!
b1001 %
1'
b1001 +
#937570000000
0!
0'
#937580000000
1!
b0 %
1'
b0 +
#937590000000
0!
0'
#937600000000
1!
1$
b1 %
1'
1*
b1 +
#937610000000
1"
1(
#937620000000
0!
0"
b100 &
0'
0(
b100 ,
#937630000000
1!
b10 %
1'
b10 +
#937640000000
0!
0'
#937650000000
1!
b11 %
1'
b11 +
#937660000000
0!
0'
#937670000000
1!
b100 %
1'
b100 +
#937680000000
0!
0'
#937690000000
1!
b101 %
1'
b101 +
#937700000000
0!
0'
#937710000000
1!
b110 %
1'
b110 +
#937720000000
0!
0'
#937730000000
1!
b111 %
1'
b111 +
#937740000000
0!
0'
#937750000000
1!
0$
b1000 %
1'
0*
b1000 +
#937760000000
0!
0'
#937770000000
1!
b1001 %
1'
b1001 +
#937780000000
0!
0'
#937790000000
1!
b0 %
1'
b0 +
#937800000000
0!
0'
#937810000000
1!
1$
b1 %
1'
1*
b1 +
#937820000000
0!
0'
#937830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#937840000000
0!
0'
#937850000000
1!
b11 %
1'
b11 +
#937860000000
0!
0'
#937870000000
1!
b100 %
1'
b100 +
#937880000000
0!
0'
#937890000000
1!
b101 %
1'
b101 +
#937900000000
0!
0'
#937910000000
1!
0$
b110 %
1'
0*
b110 +
#937920000000
0!
0'
#937930000000
1!
b111 %
1'
b111 +
#937940000000
0!
0'
#937950000000
1!
b1000 %
1'
b1000 +
#937960000000
0!
0'
#937970000000
1!
b1001 %
1'
b1001 +
#937980000000
0!
0'
#937990000000
1!
b0 %
1'
b0 +
#938000000000
0!
0'
#938010000000
1!
1$
b1 %
1'
1*
b1 +
#938020000000
0!
0'
#938030000000
1!
b10 %
1'
b10 +
#938040000000
1"
1(
#938050000000
0!
0"
b100 &
0'
0(
b100 ,
#938060000000
1!
b11 %
1'
b11 +
#938070000000
0!
0'
#938080000000
1!
b100 %
1'
b100 +
#938090000000
0!
0'
#938100000000
1!
b101 %
1'
b101 +
#938110000000
0!
0'
#938120000000
1!
b110 %
1'
b110 +
#938130000000
0!
0'
#938140000000
1!
b111 %
1'
b111 +
#938150000000
0!
0'
#938160000000
1!
0$
b1000 %
1'
0*
b1000 +
#938170000000
0!
0'
#938180000000
1!
b1001 %
1'
b1001 +
#938190000000
0!
0'
#938200000000
1!
b0 %
1'
b0 +
#938210000000
0!
0'
#938220000000
1!
1$
b1 %
1'
1*
b1 +
#938230000000
0!
0'
#938240000000
1!
b10 %
1'
b10 +
#938250000000
0!
0'
#938260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#938270000000
0!
0'
#938280000000
1!
b100 %
1'
b100 +
#938290000000
0!
0'
#938300000000
1!
b101 %
1'
b101 +
#938310000000
0!
0'
#938320000000
1!
0$
b110 %
1'
0*
b110 +
#938330000000
0!
0'
#938340000000
1!
b111 %
1'
b111 +
#938350000000
0!
0'
#938360000000
1!
b1000 %
1'
b1000 +
#938370000000
0!
0'
#938380000000
1!
b1001 %
1'
b1001 +
#938390000000
0!
0'
#938400000000
1!
b0 %
1'
b0 +
#938410000000
0!
0'
#938420000000
1!
1$
b1 %
1'
1*
b1 +
#938430000000
0!
0'
#938440000000
1!
b10 %
1'
b10 +
#938450000000
0!
0'
#938460000000
1!
b11 %
1'
b11 +
#938470000000
1"
1(
#938480000000
0!
0"
b100 &
0'
0(
b100 ,
#938490000000
1!
b100 %
1'
b100 +
#938500000000
0!
0'
#938510000000
1!
b101 %
1'
b101 +
#938520000000
0!
0'
#938530000000
1!
b110 %
1'
b110 +
#938540000000
0!
0'
#938550000000
1!
b111 %
1'
b111 +
#938560000000
0!
0'
#938570000000
1!
0$
b1000 %
1'
0*
b1000 +
#938580000000
0!
0'
#938590000000
1!
b1001 %
1'
b1001 +
#938600000000
0!
0'
#938610000000
1!
b0 %
1'
b0 +
#938620000000
0!
0'
#938630000000
1!
1$
b1 %
1'
1*
b1 +
#938640000000
0!
0'
#938650000000
1!
b10 %
1'
b10 +
#938660000000
0!
0'
#938670000000
1!
b11 %
1'
b11 +
#938680000000
0!
0'
#938690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#938700000000
0!
0'
#938710000000
1!
b101 %
1'
b101 +
#938720000000
0!
0'
#938730000000
1!
0$
b110 %
1'
0*
b110 +
#938740000000
0!
0'
#938750000000
1!
b111 %
1'
b111 +
#938760000000
0!
0'
#938770000000
1!
b1000 %
1'
b1000 +
#938780000000
0!
0'
#938790000000
1!
b1001 %
1'
b1001 +
#938800000000
0!
0'
#938810000000
1!
b0 %
1'
b0 +
#938820000000
0!
0'
#938830000000
1!
1$
b1 %
1'
1*
b1 +
#938840000000
0!
0'
#938850000000
1!
b10 %
1'
b10 +
#938860000000
0!
0'
#938870000000
1!
b11 %
1'
b11 +
#938880000000
0!
0'
#938890000000
1!
b100 %
1'
b100 +
#938900000000
1"
1(
#938910000000
0!
0"
b100 &
0'
0(
b100 ,
#938920000000
1!
b101 %
1'
b101 +
#938930000000
0!
0'
#938940000000
1!
b110 %
1'
b110 +
#938950000000
0!
0'
#938960000000
1!
b111 %
1'
b111 +
#938970000000
0!
0'
#938980000000
1!
0$
b1000 %
1'
0*
b1000 +
#938990000000
0!
0'
#939000000000
1!
b1001 %
1'
b1001 +
#939010000000
0!
0'
#939020000000
1!
b0 %
1'
b0 +
#939030000000
0!
0'
#939040000000
1!
1$
b1 %
1'
1*
b1 +
#939050000000
0!
0'
#939060000000
1!
b10 %
1'
b10 +
#939070000000
0!
0'
#939080000000
1!
b11 %
1'
b11 +
#939090000000
0!
0'
#939100000000
1!
b100 %
1'
b100 +
#939110000000
0!
0'
#939120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#939130000000
0!
0'
#939140000000
1!
0$
b110 %
1'
0*
b110 +
#939150000000
0!
0'
#939160000000
1!
b111 %
1'
b111 +
#939170000000
0!
0'
#939180000000
1!
b1000 %
1'
b1000 +
#939190000000
0!
0'
#939200000000
1!
b1001 %
1'
b1001 +
#939210000000
0!
0'
#939220000000
1!
b0 %
1'
b0 +
#939230000000
0!
0'
#939240000000
1!
1$
b1 %
1'
1*
b1 +
#939250000000
0!
0'
#939260000000
1!
b10 %
1'
b10 +
#939270000000
0!
0'
#939280000000
1!
b11 %
1'
b11 +
#939290000000
0!
0'
#939300000000
1!
b100 %
1'
b100 +
#939310000000
0!
0'
#939320000000
1!
b101 %
1'
b101 +
#939330000000
1"
1(
#939340000000
0!
0"
b100 &
0'
0(
b100 ,
#939350000000
1!
b110 %
1'
b110 +
#939360000000
0!
0'
#939370000000
1!
b111 %
1'
b111 +
#939380000000
0!
0'
#939390000000
1!
0$
b1000 %
1'
0*
b1000 +
#939400000000
0!
0'
#939410000000
1!
b1001 %
1'
b1001 +
#939420000000
0!
0'
#939430000000
1!
b0 %
1'
b0 +
#939440000000
0!
0'
#939450000000
1!
1$
b1 %
1'
1*
b1 +
#939460000000
0!
0'
#939470000000
1!
b10 %
1'
b10 +
#939480000000
0!
0'
#939490000000
1!
b11 %
1'
b11 +
#939500000000
0!
0'
#939510000000
1!
b100 %
1'
b100 +
#939520000000
0!
0'
#939530000000
1!
b101 %
1'
b101 +
#939540000000
0!
0'
#939550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#939560000000
0!
0'
#939570000000
1!
b111 %
1'
b111 +
#939580000000
0!
0'
#939590000000
1!
b1000 %
1'
b1000 +
#939600000000
0!
0'
#939610000000
1!
b1001 %
1'
b1001 +
#939620000000
0!
0'
#939630000000
1!
b0 %
1'
b0 +
#939640000000
0!
0'
#939650000000
1!
1$
b1 %
1'
1*
b1 +
#939660000000
0!
0'
#939670000000
1!
b10 %
1'
b10 +
#939680000000
0!
0'
#939690000000
1!
b11 %
1'
b11 +
#939700000000
0!
0'
#939710000000
1!
b100 %
1'
b100 +
#939720000000
0!
0'
#939730000000
1!
b101 %
1'
b101 +
#939740000000
0!
0'
#939750000000
1!
0$
b110 %
1'
0*
b110 +
#939760000000
1"
1(
#939770000000
0!
0"
b100 &
0'
0(
b100 ,
#939780000000
1!
1$
b111 %
1'
1*
b111 +
#939790000000
0!
0'
#939800000000
1!
0$
b1000 %
1'
0*
b1000 +
#939810000000
0!
0'
#939820000000
1!
b1001 %
1'
b1001 +
#939830000000
0!
0'
#939840000000
1!
b0 %
1'
b0 +
#939850000000
0!
0'
#939860000000
1!
1$
b1 %
1'
1*
b1 +
#939870000000
0!
0'
#939880000000
1!
b10 %
1'
b10 +
#939890000000
0!
0'
#939900000000
1!
b11 %
1'
b11 +
#939910000000
0!
0'
#939920000000
1!
b100 %
1'
b100 +
#939930000000
0!
0'
#939940000000
1!
b101 %
1'
b101 +
#939950000000
0!
0'
#939960000000
1!
b110 %
1'
b110 +
#939970000000
0!
0'
#939980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#939990000000
0!
0'
#940000000000
1!
b1000 %
1'
b1000 +
#940010000000
0!
0'
#940020000000
1!
b1001 %
1'
b1001 +
#940030000000
0!
0'
#940040000000
1!
b0 %
1'
b0 +
#940050000000
0!
0'
#940060000000
1!
1$
b1 %
1'
1*
b1 +
#940070000000
0!
0'
#940080000000
1!
b10 %
1'
b10 +
#940090000000
0!
0'
#940100000000
1!
b11 %
1'
b11 +
#940110000000
0!
0'
#940120000000
1!
b100 %
1'
b100 +
#940130000000
0!
0'
#940140000000
1!
b101 %
1'
b101 +
#940150000000
0!
0'
#940160000000
1!
0$
b110 %
1'
0*
b110 +
#940170000000
0!
0'
#940180000000
1!
b111 %
1'
b111 +
#940190000000
1"
1(
#940200000000
0!
0"
b100 &
0'
0(
b100 ,
#940210000000
1!
b1000 %
1'
b1000 +
#940220000000
0!
0'
#940230000000
1!
b1001 %
1'
b1001 +
#940240000000
0!
0'
#940250000000
1!
b0 %
1'
b0 +
#940260000000
0!
0'
#940270000000
1!
1$
b1 %
1'
1*
b1 +
#940280000000
0!
0'
#940290000000
1!
b10 %
1'
b10 +
#940300000000
0!
0'
#940310000000
1!
b11 %
1'
b11 +
#940320000000
0!
0'
#940330000000
1!
b100 %
1'
b100 +
#940340000000
0!
0'
#940350000000
1!
b101 %
1'
b101 +
#940360000000
0!
0'
#940370000000
1!
b110 %
1'
b110 +
#940380000000
0!
0'
#940390000000
1!
b111 %
1'
b111 +
#940400000000
0!
0'
#940410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#940420000000
0!
0'
#940430000000
1!
b1001 %
1'
b1001 +
#940440000000
0!
0'
#940450000000
1!
b0 %
1'
b0 +
#940460000000
0!
0'
#940470000000
1!
1$
b1 %
1'
1*
b1 +
#940480000000
0!
0'
#940490000000
1!
b10 %
1'
b10 +
#940500000000
0!
0'
#940510000000
1!
b11 %
1'
b11 +
#940520000000
0!
0'
#940530000000
1!
b100 %
1'
b100 +
#940540000000
0!
0'
#940550000000
1!
b101 %
1'
b101 +
#940560000000
0!
0'
#940570000000
1!
0$
b110 %
1'
0*
b110 +
#940580000000
0!
0'
#940590000000
1!
b111 %
1'
b111 +
#940600000000
0!
0'
#940610000000
1!
b1000 %
1'
b1000 +
#940620000000
1"
1(
#940630000000
0!
0"
b100 &
0'
0(
b100 ,
#940640000000
1!
b1001 %
1'
b1001 +
#940650000000
0!
0'
#940660000000
1!
b0 %
1'
b0 +
#940670000000
0!
0'
#940680000000
1!
1$
b1 %
1'
1*
b1 +
#940690000000
0!
0'
#940700000000
1!
b10 %
1'
b10 +
#940710000000
0!
0'
#940720000000
1!
b11 %
1'
b11 +
#940730000000
0!
0'
#940740000000
1!
b100 %
1'
b100 +
#940750000000
0!
0'
#940760000000
1!
b101 %
1'
b101 +
#940770000000
0!
0'
#940780000000
1!
b110 %
1'
b110 +
#940790000000
0!
0'
#940800000000
1!
b111 %
1'
b111 +
#940810000000
0!
0'
#940820000000
1!
0$
b1000 %
1'
0*
b1000 +
#940830000000
0!
0'
#940840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#940850000000
0!
0'
#940860000000
1!
b0 %
1'
b0 +
#940870000000
0!
0'
#940880000000
1!
1$
b1 %
1'
1*
b1 +
#940890000000
0!
0'
#940900000000
1!
b10 %
1'
b10 +
#940910000000
0!
0'
#940920000000
1!
b11 %
1'
b11 +
#940930000000
0!
0'
#940940000000
1!
b100 %
1'
b100 +
#940950000000
0!
0'
#940960000000
1!
b101 %
1'
b101 +
#940970000000
0!
0'
#940980000000
1!
0$
b110 %
1'
0*
b110 +
#940990000000
0!
0'
#941000000000
1!
b111 %
1'
b111 +
#941010000000
0!
0'
#941020000000
1!
b1000 %
1'
b1000 +
#941030000000
0!
0'
#941040000000
1!
b1001 %
1'
b1001 +
#941050000000
1"
1(
#941060000000
0!
0"
b100 &
0'
0(
b100 ,
#941070000000
1!
b0 %
1'
b0 +
#941080000000
0!
0'
#941090000000
1!
1$
b1 %
1'
1*
b1 +
#941100000000
0!
0'
#941110000000
1!
b10 %
1'
b10 +
#941120000000
0!
0'
#941130000000
1!
b11 %
1'
b11 +
#941140000000
0!
0'
#941150000000
1!
b100 %
1'
b100 +
#941160000000
0!
0'
#941170000000
1!
b101 %
1'
b101 +
#941180000000
0!
0'
#941190000000
1!
b110 %
1'
b110 +
#941200000000
0!
0'
#941210000000
1!
b111 %
1'
b111 +
#941220000000
0!
0'
#941230000000
1!
0$
b1000 %
1'
0*
b1000 +
#941240000000
0!
0'
#941250000000
1!
b1001 %
1'
b1001 +
#941260000000
0!
0'
#941270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#941280000000
0!
0'
#941290000000
1!
1$
b1 %
1'
1*
b1 +
#941300000000
0!
0'
#941310000000
1!
b10 %
1'
b10 +
#941320000000
0!
0'
#941330000000
1!
b11 %
1'
b11 +
#941340000000
0!
0'
#941350000000
1!
b100 %
1'
b100 +
#941360000000
0!
0'
#941370000000
1!
b101 %
1'
b101 +
#941380000000
0!
0'
#941390000000
1!
0$
b110 %
1'
0*
b110 +
#941400000000
0!
0'
#941410000000
1!
b111 %
1'
b111 +
#941420000000
0!
0'
#941430000000
1!
b1000 %
1'
b1000 +
#941440000000
0!
0'
#941450000000
1!
b1001 %
1'
b1001 +
#941460000000
0!
0'
#941470000000
1!
b0 %
1'
b0 +
#941480000000
1"
1(
#941490000000
0!
0"
b100 &
0'
0(
b100 ,
#941500000000
1!
1$
b1 %
1'
1*
b1 +
#941510000000
0!
0'
#941520000000
1!
b10 %
1'
b10 +
#941530000000
0!
0'
#941540000000
1!
b11 %
1'
b11 +
#941550000000
0!
0'
#941560000000
1!
b100 %
1'
b100 +
#941570000000
0!
0'
#941580000000
1!
b101 %
1'
b101 +
#941590000000
0!
0'
#941600000000
1!
b110 %
1'
b110 +
#941610000000
0!
0'
#941620000000
1!
b111 %
1'
b111 +
#941630000000
0!
0'
#941640000000
1!
0$
b1000 %
1'
0*
b1000 +
#941650000000
0!
0'
#941660000000
1!
b1001 %
1'
b1001 +
#941670000000
0!
0'
#941680000000
1!
b0 %
1'
b0 +
#941690000000
0!
0'
#941700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#941710000000
0!
0'
#941720000000
1!
b10 %
1'
b10 +
#941730000000
0!
0'
#941740000000
1!
b11 %
1'
b11 +
#941750000000
0!
0'
#941760000000
1!
b100 %
1'
b100 +
#941770000000
0!
0'
#941780000000
1!
b101 %
1'
b101 +
#941790000000
0!
0'
#941800000000
1!
0$
b110 %
1'
0*
b110 +
#941810000000
0!
0'
#941820000000
1!
b111 %
1'
b111 +
#941830000000
0!
0'
#941840000000
1!
b1000 %
1'
b1000 +
#941850000000
0!
0'
#941860000000
1!
b1001 %
1'
b1001 +
#941870000000
0!
0'
#941880000000
1!
b0 %
1'
b0 +
#941890000000
0!
0'
#941900000000
1!
1$
b1 %
1'
1*
b1 +
#941910000000
1"
1(
#941920000000
0!
0"
b100 &
0'
0(
b100 ,
#941930000000
1!
b10 %
1'
b10 +
#941940000000
0!
0'
#941950000000
1!
b11 %
1'
b11 +
#941960000000
0!
0'
#941970000000
1!
b100 %
1'
b100 +
#941980000000
0!
0'
#941990000000
1!
b101 %
1'
b101 +
#942000000000
0!
0'
#942010000000
1!
b110 %
1'
b110 +
#942020000000
0!
0'
#942030000000
1!
b111 %
1'
b111 +
#942040000000
0!
0'
#942050000000
1!
0$
b1000 %
1'
0*
b1000 +
#942060000000
0!
0'
#942070000000
1!
b1001 %
1'
b1001 +
#942080000000
0!
0'
#942090000000
1!
b0 %
1'
b0 +
#942100000000
0!
0'
#942110000000
1!
1$
b1 %
1'
1*
b1 +
#942120000000
0!
0'
#942130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#942140000000
0!
0'
#942150000000
1!
b11 %
1'
b11 +
#942160000000
0!
0'
#942170000000
1!
b100 %
1'
b100 +
#942180000000
0!
0'
#942190000000
1!
b101 %
1'
b101 +
#942200000000
0!
0'
#942210000000
1!
0$
b110 %
1'
0*
b110 +
#942220000000
0!
0'
#942230000000
1!
b111 %
1'
b111 +
#942240000000
0!
0'
#942250000000
1!
b1000 %
1'
b1000 +
#942260000000
0!
0'
#942270000000
1!
b1001 %
1'
b1001 +
#942280000000
0!
0'
#942290000000
1!
b0 %
1'
b0 +
#942300000000
0!
0'
#942310000000
1!
1$
b1 %
1'
1*
b1 +
#942320000000
0!
0'
#942330000000
1!
b10 %
1'
b10 +
#942340000000
1"
1(
#942350000000
0!
0"
b100 &
0'
0(
b100 ,
#942360000000
1!
b11 %
1'
b11 +
#942370000000
0!
0'
#942380000000
1!
b100 %
1'
b100 +
#942390000000
0!
0'
#942400000000
1!
b101 %
1'
b101 +
#942410000000
0!
0'
#942420000000
1!
b110 %
1'
b110 +
#942430000000
0!
0'
#942440000000
1!
b111 %
1'
b111 +
#942450000000
0!
0'
#942460000000
1!
0$
b1000 %
1'
0*
b1000 +
#942470000000
0!
0'
#942480000000
1!
b1001 %
1'
b1001 +
#942490000000
0!
0'
#942500000000
1!
b0 %
1'
b0 +
#942510000000
0!
0'
#942520000000
1!
1$
b1 %
1'
1*
b1 +
#942530000000
0!
0'
#942540000000
1!
b10 %
1'
b10 +
#942550000000
0!
0'
#942560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#942570000000
0!
0'
#942580000000
1!
b100 %
1'
b100 +
#942590000000
0!
0'
#942600000000
1!
b101 %
1'
b101 +
#942610000000
0!
0'
#942620000000
1!
0$
b110 %
1'
0*
b110 +
#942630000000
0!
0'
#942640000000
1!
b111 %
1'
b111 +
#942650000000
0!
0'
#942660000000
1!
b1000 %
1'
b1000 +
#942670000000
0!
0'
#942680000000
1!
b1001 %
1'
b1001 +
#942690000000
0!
0'
#942700000000
1!
b0 %
1'
b0 +
#942710000000
0!
0'
#942720000000
1!
1$
b1 %
1'
1*
b1 +
#942730000000
0!
0'
#942740000000
1!
b10 %
1'
b10 +
#942750000000
0!
0'
#942760000000
1!
b11 %
1'
b11 +
#942770000000
1"
1(
#942780000000
0!
0"
b100 &
0'
0(
b100 ,
#942790000000
1!
b100 %
1'
b100 +
#942800000000
0!
0'
#942810000000
1!
b101 %
1'
b101 +
#942820000000
0!
0'
#942830000000
1!
b110 %
1'
b110 +
#942840000000
0!
0'
#942850000000
1!
b111 %
1'
b111 +
#942860000000
0!
0'
#942870000000
1!
0$
b1000 %
1'
0*
b1000 +
#942880000000
0!
0'
#942890000000
1!
b1001 %
1'
b1001 +
#942900000000
0!
0'
#942910000000
1!
b0 %
1'
b0 +
#942920000000
0!
0'
#942930000000
1!
1$
b1 %
1'
1*
b1 +
#942940000000
0!
0'
#942950000000
1!
b10 %
1'
b10 +
#942960000000
0!
0'
#942970000000
1!
b11 %
1'
b11 +
#942980000000
0!
0'
#942990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#943000000000
0!
0'
#943010000000
1!
b101 %
1'
b101 +
#943020000000
0!
0'
#943030000000
1!
0$
b110 %
1'
0*
b110 +
#943040000000
0!
0'
#943050000000
1!
b111 %
1'
b111 +
#943060000000
0!
0'
#943070000000
1!
b1000 %
1'
b1000 +
#943080000000
0!
0'
#943090000000
1!
b1001 %
1'
b1001 +
#943100000000
0!
0'
#943110000000
1!
b0 %
1'
b0 +
#943120000000
0!
0'
#943130000000
1!
1$
b1 %
1'
1*
b1 +
#943140000000
0!
0'
#943150000000
1!
b10 %
1'
b10 +
#943160000000
0!
0'
#943170000000
1!
b11 %
1'
b11 +
#943180000000
0!
0'
#943190000000
1!
b100 %
1'
b100 +
#943200000000
1"
1(
#943210000000
0!
0"
b100 &
0'
0(
b100 ,
#943220000000
1!
b101 %
1'
b101 +
#943230000000
0!
0'
#943240000000
1!
b110 %
1'
b110 +
#943250000000
0!
0'
#943260000000
1!
b111 %
1'
b111 +
#943270000000
0!
0'
#943280000000
1!
0$
b1000 %
1'
0*
b1000 +
#943290000000
0!
0'
#943300000000
1!
b1001 %
1'
b1001 +
#943310000000
0!
0'
#943320000000
1!
b0 %
1'
b0 +
#943330000000
0!
0'
#943340000000
1!
1$
b1 %
1'
1*
b1 +
#943350000000
0!
0'
#943360000000
1!
b10 %
1'
b10 +
#943370000000
0!
0'
#943380000000
1!
b11 %
1'
b11 +
#943390000000
0!
0'
#943400000000
1!
b100 %
1'
b100 +
#943410000000
0!
0'
#943420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#943430000000
0!
0'
#943440000000
1!
0$
b110 %
1'
0*
b110 +
#943450000000
0!
0'
#943460000000
1!
b111 %
1'
b111 +
#943470000000
0!
0'
#943480000000
1!
b1000 %
1'
b1000 +
#943490000000
0!
0'
#943500000000
1!
b1001 %
1'
b1001 +
#943510000000
0!
0'
#943520000000
1!
b0 %
1'
b0 +
#943530000000
0!
0'
#943540000000
1!
1$
b1 %
1'
1*
b1 +
#943550000000
0!
0'
#943560000000
1!
b10 %
1'
b10 +
#943570000000
0!
0'
#943580000000
1!
b11 %
1'
b11 +
#943590000000
0!
0'
#943600000000
1!
b100 %
1'
b100 +
#943610000000
0!
0'
#943620000000
1!
b101 %
1'
b101 +
#943630000000
1"
1(
#943640000000
0!
0"
b100 &
0'
0(
b100 ,
#943650000000
1!
b110 %
1'
b110 +
#943660000000
0!
0'
#943670000000
1!
b111 %
1'
b111 +
#943680000000
0!
0'
#943690000000
1!
0$
b1000 %
1'
0*
b1000 +
#943700000000
0!
0'
#943710000000
1!
b1001 %
1'
b1001 +
#943720000000
0!
0'
#943730000000
1!
b0 %
1'
b0 +
#943740000000
0!
0'
#943750000000
1!
1$
b1 %
1'
1*
b1 +
#943760000000
0!
0'
#943770000000
1!
b10 %
1'
b10 +
#943780000000
0!
0'
#943790000000
1!
b11 %
1'
b11 +
#943800000000
0!
0'
#943810000000
1!
b100 %
1'
b100 +
#943820000000
0!
0'
#943830000000
1!
b101 %
1'
b101 +
#943840000000
0!
0'
#943850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#943860000000
0!
0'
#943870000000
1!
b111 %
1'
b111 +
#943880000000
0!
0'
#943890000000
1!
b1000 %
1'
b1000 +
#943900000000
0!
0'
#943910000000
1!
b1001 %
1'
b1001 +
#943920000000
0!
0'
#943930000000
1!
b0 %
1'
b0 +
#943940000000
0!
0'
#943950000000
1!
1$
b1 %
1'
1*
b1 +
#943960000000
0!
0'
#943970000000
1!
b10 %
1'
b10 +
#943980000000
0!
0'
#943990000000
1!
b11 %
1'
b11 +
#944000000000
0!
0'
#944010000000
1!
b100 %
1'
b100 +
#944020000000
0!
0'
#944030000000
1!
b101 %
1'
b101 +
#944040000000
0!
0'
#944050000000
1!
0$
b110 %
1'
0*
b110 +
#944060000000
1"
1(
#944070000000
0!
0"
b100 &
0'
0(
b100 ,
#944080000000
1!
1$
b111 %
1'
1*
b111 +
#944090000000
0!
0'
#944100000000
1!
0$
b1000 %
1'
0*
b1000 +
#944110000000
0!
0'
#944120000000
1!
b1001 %
1'
b1001 +
#944130000000
0!
0'
#944140000000
1!
b0 %
1'
b0 +
#944150000000
0!
0'
#944160000000
1!
1$
b1 %
1'
1*
b1 +
#944170000000
0!
0'
#944180000000
1!
b10 %
1'
b10 +
#944190000000
0!
0'
#944200000000
1!
b11 %
1'
b11 +
#944210000000
0!
0'
#944220000000
1!
b100 %
1'
b100 +
#944230000000
0!
0'
#944240000000
1!
b101 %
1'
b101 +
#944250000000
0!
0'
#944260000000
1!
b110 %
1'
b110 +
#944270000000
0!
0'
#944280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#944290000000
0!
0'
#944300000000
1!
b1000 %
1'
b1000 +
#944310000000
0!
0'
#944320000000
1!
b1001 %
1'
b1001 +
#944330000000
0!
0'
#944340000000
1!
b0 %
1'
b0 +
#944350000000
0!
0'
#944360000000
1!
1$
b1 %
1'
1*
b1 +
#944370000000
0!
0'
#944380000000
1!
b10 %
1'
b10 +
#944390000000
0!
0'
#944400000000
1!
b11 %
1'
b11 +
#944410000000
0!
0'
#944420000000
1!
b100 %
1'
b100 +
#944430000000
0!
0'
#944440000000
1!
b101 %
1'
b101 +
#944450000000
0!
0'
#944460000000
1!
0$
b110 %
1'
0*
b110 +
#944470000000
0!
0'
#944480000000
1!
b111 %
1'
b111 +
#944490000000
1"
1(
#944500000000
0!
0"
b100 &
0'
0(
b100 ,
#944510000000
1!
b1000 %
1'
b1000 +
#944520000000
0!
0'
#944530000000
1!
b1001 %
1'
b1001 +
#944540000000
0!
0'
#944550000000
1!
b0 %
1'
b0 +
#944560000000
0!
0'
#944570000000
1!
1$
b1 %
1'
1*
b1 +
#944580000000
0!
0'
#944590000000
1!
b10 %
1'
b10 +
#944600000000
0!
0'
#944610000000
1!
b11 %
1'
b11 +
#944620000000
0!
0'
#944630000000
1!
b100 %
1'
b100 +
#944640000000
0!
0'
#944650000000
1!
b101 %
1'
b101 +
#944660000000
0!
0'
#944670000000
1!
b110 %
1'
b110 +
#944680000000
0!
0'
#944690000000
1!
b111 %
1'
b111 +
#944700000000
0!
0'
#944710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#944720000000
0!
0'
#944730000000
1!
b1001 %
1'
b1001 +
#944740000000
0!
0'
#944750000000
1!
b0 %
1'
b0 +
#944760000000
0!
0'
#944770000000
1!
1$
b1 %
1'
1*
b1 +
#944780000000
0!
0'
#944790000000
1!
b10 %
1'
b10 +
#944800000000
0!
0'
#944810000000
1!
b11 %
1'
b11 +
#944820000000
0!
0'
#944830000000
1!
b100 %
1'
b100 +
#944840000000
0!
0'
#944850000000
1!
b101 %
1'
b101 +
#944860000000
0!
0'
#944870000000
1!
0$
b110 %
1'
0*
b110 +
#944880000000
0!
0'
#944890000000
1!
b111 %
1'
b111 +
#944900000000
0!
0'
#944910000000
1!
b1000 %
1'
b1000 +
#944920000000
1"
1(
#944930000000
0!
0"
b100 &
0'
0(
b100 ,
#944940000000
1!
b1001 %
1'
b1001 +
#944950000000
0!
0'
#944960000000
1!
b0 %
1'
b0 +
#944970000000
0!
0'
#944980000000
1!
1$
b1 %
1'
1*
b1 +
#944990000000
0!
0'
#945000000000
1!
b10 %
1'
b10 +
#945010000000
0!
0'
#945020000000
1!
b11 %
1'
b11 +
#945030000000
0!
0'
#945040000000
1!
b100 %
1'
b100 +
#945050000000
0!
0'
#945060000000
1!
b101 %
1'
b101 +
#945070000000
0!
0'
#945080000000
1!
b110 %
1'
b110 +
#945090000000
0!
0'
#945100000000
1!
b111 %
1'
b111 +
#945110000000
0!
0'
#945120000000
1!
0$
b1000 %
1'
0*
b1000 +
#945130000000
0!
0'
#945140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#945150000000
0!
0'
#945160000000
1!
b0 %
1'
b0 +
#945170000000
0!
0'
#945180000000
1!
1$
b1 %
1'
1*
b1 +
#945190000000
0!
0'
#945200000000
1!
b10 %
1'
b10 +
#945210000000
0!
0'
#945220000000
1!
b11 %
1'
b11 +
#945230000000
0!
0'
#945240000000
1!
b100 %
1'
b100 +
#945250000000
0!
0'
#945260000000
1!
b101 %
1'
b101 +
#945270000000
0!
0'
#945280000000
1!
0$
b110 %
1'
0*
b110 +
#945290000000
0!
0'
#945300000000
1!
b111 %
1'
b111 +
#945310000000
0!
0'
#945320000000
1!
b1000 %
1'
b1000 +
#945330000000
0!
0'
#945340000000
1!
b1001 %
1'
b1001 +
#945350000000
1"
1(
#945360000000
0!
0"
b100 &
0'
0(
b100 ,
#945370000000
1!
b0 %
1'
b0 +
#945380000000
0!
0'
#945390000000
1!
1$
b1 %
1'
1*
b1 +
#945400000000
0!
0'
#945410000000
1!
b10 %
1'
b10 +
#945420000000
0!
0'
#945430000000
1!
b11 %
1'
b11 +
#945440000000
0!
0'
#945450000000
1!
b100 %
1'
b100 +
#945460000000
0!
0'
#945470000000
1!
b101 %
1'
b101 +
#945480000000
0!
0'
#945490000000
1!
b110 %
1'
b110 +
#945500000000
0!
0'
#945510000000
1!
b111 %
1'
b111 +
#945520000000
0!
0'
#945530000000
1!
0$
b1000 %
1'
0*
b1000 +
#945540000000
0!
0'
#945550000000
1!
b1001 %
1'
b1001 +
#945560000000
0!
0'
#945570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#945580000000
0!
0'
#945590000000
1!
1$
b1 %
1'
1*
b1 +
#945600000000
0!
0'
#945610000000
1!
b10 %
1'
b10 +
#945620000000
0!
0'
#945630000000
1!
b11 %
1'
b11 +
#945640000000
0!
0'
#945650000000
1!
b100 %
1'
b100 +
#945660000000
0!
0'
#945670000000
1!
b101 %
1'
b101 +
#945680000000
0!
0'
#945690000000
1!
0$
b110 %
1'
0*
b110 +
#945700000000
0!
0'
#945710000000
1!
b111 %
1'
b111 +
#945720000000
0!
0'
#945730000000
1!
b1000 %
1'
b1000 +
#945740000000
0!
0'
#945750000000
1!
b1001 %
1'
b1001 +
#945760000000
0!
0'
#945770000000
1!
b0 %
1'
b0 +
#945780000000
1"
1(
#945790000000
0!
0"
b100 &
0'
0(
b100 ,
#945800000000
1!
1$
b1 %
1'
1*
b1 +
#945810000000
0!
0'
#945820000000
1!
b10 %
1'
b10 +
#945830000000
0!
0'
#945840000000
1!
b11 %
1'
b11 +
#945850000000
0!
0'
#945860000000
1!
b100 %
1'
b100 +
#945870000000
0!
0'
#945880000000
1!
b101 %
1'
b101 +
#945890000000
0!
0'
#945900000000
1!
b110 %
1'
b110 +
#945910000000
0!
0'
#945920000000
1!
b111 %
1'
b111 +
#945930000000
0!
0'
#945940000000
1!
0$
b1000 %
1'
0*
b1000 +
#945950000000
0!
0'
#945960000000
1!
b1001 %
1'
b1001 +
#945970000000
0!
0'
#945980000000
1!
b0 %
1'
b0 +
#945990000000
0!
0'
#946000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#946010000000
0!
0'
#946020000000
1!
b10 %
1'
b10 +
#946030000000
0!
0'
#946040000000
1!
b11 %
1'
b11 +
#946050000000
0!
0'
#946060000000
1!
b100 %
1'
b100 +
#946070000000
0!
0'
#946080000000
1!
b101 %
1'
b101 +
#946090000000
0!
0'
#946100000000
1!
0$
b110 %
1'
0*
b110 +
#946110000000
0!
0'
#946120000000
1!
b111 %
1'
b111 +
#946130000000
0!
0'
#946140000000
1!
b1000 %
1'
b1000 +
#946150000000
0!
0'
#946160000000
1!
b1001 %
1'
b1001 +
#946170000000
0!
0'
#946180000000
1!
b0 %
1'
b0 +
#946190000000
0!
0'
#946200000000
1!
1$
b1 %
1'
1*
b1 +
#946210000000
1"
1(
#946220000000
0!
0"
b100 &
0'
0(
b100 ,
#946230000000
1!
b10 %
1'
b10 +
#946240000000
0!
0'
#946250000000
1!
b11 %
1'
b11 +
#946260000000
0!
0'
#946270000000
1!
b100 %
1'
b100 +
#946280000000
0!
0'
#946290000000
1!
b101 %
1'
b101 +
#946300000000
0!
0'
#946310000000
1!
b110 %
1'
b110 +
#946320000000
0!
0'
#946330000000
1!
b111 %
1'
b111 +
#946340000000
0!
0'
#946350000000
1!
0$
b1000 %
1'
0*
b1000 +
#946360000000
0!
0'
#946370000000
1!
b1001 %
1'
b1001 +
#946380000000
0!
0'
#946390000000
1!
b0 %
1'
b0 +
#946400000000
0!
0'
#946410000000
1!
1$
b1 %
1'
1*
b1 +
#946420000000
0!
0'
#946430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#946440000000
0!
0'
#946450000000
1!
b11 %
1'
b11 +
#946460000000
0!
0'
#946470000000
1!
b100 %
1'
b100 +
#946480000000
0!
0'
#946490000000
1!
b101 %
1'
b101 +
#946500000000
0!
0'
#946510000000
1!
0$
b110 %
1'
0*
b110 +
#946520000000
0!
0'
#946530000000
1!
b111 %
1'
b111 +
#946540000000
0!
0'
#946550000000
1!
b1000 %
1'
b1000 +
#946560000000
0!
0'
#946570000000
1!
b1001 %
1'
b1001 +
#946580000000
0!
0'
#946590000000
1!
b0 %
1'
b0 +
#946600000000
0!
0'
#946610000000
1!
1$
b1 %
1'
1*
b1 +
#946620000000
0!
0'
#946630000000
1!
b10 %
1'
b10 +
#946640000000
1"
1(
#946650000000
0!
0"
b100 &
0'
0(
b100 ,
#946660000000
1!
b11 %
1'
b11 +
#946670000000
0!
0'
#946680000000
1!
b100 %
1'
b100 +
#946690000000
0!
0'
#946700000000
1!
b101 %
1'
b101 +
#946710000000
0!
0'
#946720000000
1!
b110 %
1'
b110 +
#946730000000
0!
0'
#946740000000
1!
b111 %
1'
b111 +
#946750000000
0!
0'
#946760000000
1!
0$
b1000 %
1'
0*
b1000 +
#946770000000
0!
0'
#946780000000
1!
b1001 %
1'
b1001 +
#946790000000
0!
0'
#946800000000
1!
b0 %
1'
b0 +
#946810000000
0!
0'
#946820000000
1!
1$
b1 %
1'
1*
b1 +
#946830000000
0!
0'
#946840000000
1!
b10 %
1'
b10 +
#946850000000
0!
0'
#946860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#946870000000
0!
0'
#946880000000
1!
b100 %
1'
b100 +
#946890000000
0!
0'
#946900000000
1!
b101 %
1'
b101 +
#946910000000
0!
0'
#946920000000
1!
0$
b110 %
1'
0*
b110 +
#946930000000
0!
0'
#946940000000
1!
b111 %
1'
b111 +
#946950000000
0!
0'
#946960000000
1!
b1000 %
1'
b1000 +
#946970000000
0!
0'
#946980000000
1!
b1001 %
1'
b1001 +
#946990000000
0!
0'
#947000000000
1!
b0 %
1'
b0 +
#947010000000
0!
0'
#947020000000
1!
1$
b1 %
1'
1*
b1 +
#947030000000
0!
0'
#947040000000
1!
b10 %
1'
b10 +
#947050000000
0!
0'
#947060000000
1!
b11 %
1'
b11 +
#947070000000
1"
1(
#947080000000
0!
0"
b100 &
0'
0(
b100 ,
#947090000000
1!
b100 %
1'
b100 +
#947100000000
0!
0'
#947110000000
1!
b101 %
1'
b101 +
#947120000000
0!
0'
#947130000000
1!
b110 %
1'
b110 +
#947140000000
0!
0'
#947150000000
1!
b111 %
1'
b111 +
#947160000000
0!
0'
#947170000000
1!
0$
b1000 %
1'
0*
b1000 +
#947180000000
0!
0'
#947190000000
1!
b1001 %
1'
b1001 +
#947200000000
0!
0'
#947210000000
1!
b0 %
1'
b0 +
#947220000000
0!
0'
#947230000000
1!
1$
b1 %
1'
1*
b1 +
#947240000000
0!
0'
#947250000000
1!
b10 %
1'
b10 +
#947260000000
0!
0'
#947270000000
1!
b11 %
1'
b11 +
#947280000000
0!
0'
#947290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#947300000000
0!
0'
#947310000000
1!
b101 %
1'
b101 +
#947320000000
0!
0'
#947330000000
1!
0$
b110 %
1'
0*
b110 +
#947340000000
0!
0'
#947350000000
1!
b111 %
1'
b111 +
#947360000000
0!
0'
#947370000000
1!
b1000 %
1'
b1000 +
#947380000000
0!
0'
#947390000000
1!
b1001 %
1'
b1001 +
#947400000000
0!
0'
#947410000000
1!
b0 %
1'
b0 +
#947420000000
0!
0'
#947430000000
1!
1$
b1 %
1'
1*
b1 +
#947440000000
0!
0'
#947450000000
1!
b10 %
1'
b10 +
#947460000000
0!
0'
#947470000000
1!
b11 %
1'
b11 +
#947480000000
0!
0'
#947490000000
1!
b100 %
1'
b100 +
#947500000000
1"
1(
#947510000000
0!
0"
b100 &
0'
0(
b100 ,
#947520000000
1!
b101 %
1'
b101 +
#947530000000
0!
0'
#947540000000
1!
b110 %
1'
b110 +
#947550000000
0!
0'
#947560000000
1!
b111 %
1'
b111 +
#947570000000
0!
0'
#947580000000
1!
0$
b1000 %
1'
0*
b1000 +
#947590000000
0!
0'
#947600000000
1!
b1001 %
1'
b1001 +
#947610000000
0!
0'
#947620000000
1!
b0 %
1'
b0 +
#947630000000
0!
0'
#947640000000
1!
1$
b1 %
1'
1*
b1 +
#947650000000
0!
0'
#947660000000
1!
b10 %
1'
b10 +
#947670000000
0!
0'
#947680000000
1!
b11 %
1'
b11 +
#947690000000
0!
0'
#947700000000
1!
b100 %
1'
b100 +
#947710000000
0!
0'
#947720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#947730000000
0!
0'
#947740000000
1!
0$
b110 %
1'
0*
b110 +
#947750000000
0!
0'
#947760000000
1!
b111 %
1'
b111 +
#947770000000
0!
0'
#947780000000
1!
b1000 %
1'
b1000 +
#947790000000
0!
0'
#947800000000
1!
b1001 %
1'
b1001 +
#947810000000
0!
0'
#947820000000
1!
b0 %
1'
b0 +
#947830000000
0!
0'
#947840000000
1!
1$
b1 %
1'
1*
b1 +
#947850000000
0!
0'
#947860000000
1!
b10 %
1'
b10 +
#947870000000
0!
0'
#947880000000
1!
b11 %
1'
b11 +
#947890000000
0!
0'
#947900000000
1!
b100 %
1'
b100 +
#947910000000
0!
0'
#947920000000
1!
b101 %
1'
b101 +
#947930000000
1"
1(
#947940000000
0!
0"
b100 &
0'
0(
b100 ,
#947950000000
1!
b110 %
1'
b110 +
#947960000000
0!
0'
#947970000000
1!
b111 %
1'
b111 +
#947980000000
0!
0'
#947990000000
1!
0$
b1000 %
1'
0*
b1000 +
#948000000000
0!
0'
#948010000000
1!
b1001 %
1'
b1001 +
#948020000000
0!
0'
#948030000000
1!
b0 %
1'
b0 +
#948040000000
0!
0'
#948050000000
1!
1$
b1 %
1'
1*
b1 +
#948060000000
0!
0'
#948070000000
1!
b10 %
1'
b10 +
#948080000000
0!
0'
#948090000000
1!
b11 %
1'
b11 +
#948100000000
0!
0'
#948110000000
1!
b100 %
1'
b100 +
#948120000000
0!
0'
#948130000000
1!
b101 %
1'
b101 +
#948140000000
0!
0'
#948150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#948160000000
0!
0'
#948170000000
1!
b111 %
1'
b111 +
#948180000000
0!
0'
#948190000000
1!
b1000 %
1'
b1000 +
#948200000000
0!
0'
#948210000000
1!
b1001 %
1'
b1001 +
#948220000000
0!
0'
#948230000000
1!
b0 %
1'
b0 +
#948240000000
0!
0'
#948250000000
1!
1$
b1 %
1'
1*
b1 +
#948260000000
0!
0'
#948270000000
1!
b10 %
1'
b10 +
#948280000000
0!
0'
#948290000000
1!
b11 %
1'
b11 +
#948300000000
0!
0'
#948310000000
1!
b100 %
1'
b100 +
#948320000000
0!
0'
#948330000000
1!
b101 %
1'
b101 +
#948340000000
0!
0'
#948350000000
1!
0$
b110 %
1'
0*
b110 +
#948360000000
1"
1(
#948370000000
0!
0"
b100 &
0'
0(
b100 ,
#948380000000
1!
1$
b111 %
1'
1*
b111 +
#948390000000
0!
0'
#948400000000
1!
0$
b1000 %
1'
0*
b1000 +
#948410000000
0!
0'
#948420000000
1!
b1001 %
1'
b1001 +
#948430000000
0!
0'
#948440000000
1!
b0 %
1'
b0 +
#948450000000
0!
0'
#948460000000
1!
1$
b1 %
1'
1*
b1 +
#948470000000
0!
0'
#948480000000
1!
b10 %
1'
b10 +
#948490000000
0!
0'
#948500000000
1!
b11 %
1'
b11 +
#948510000000
0!
0'
#948520000000
1!
b100 %
1'
b100 +
#948530000000
0!
0'
#948540000000
1!
b101 %
1'
b101 +
#948550000000
0!
0'
#948560000000
1!
b110 %
1'
b110 +
#948570000000
0!
0'
#948580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#948590000000
0!
0'
#948600000000
1!
b1000 %
1'
b1000 +
#948610000000
0!
0'
#948620000000
1!
b1001 %
1'
b1001 +
#948630000000
0!
0'
#948640000000
1!
b0 %
1'
b0 +
#948650000000
0!
0'
#948660000000
1!
1$
b1 %
1'
1*
b1 +
#948670000000
0!
0'
#948680000000
1!
b10 %
1'
b10 +
#948690000000
0!
0'
#948700000000
1!
b11 %
1'
b11 +
#948710000000
0!
0'
#948720000000
1!
b100 %
1'
b100 +
#948730000000
0!
0'
#948740000000
1!
b101 %
1'
b101 +
#948750000000
0!
0'
#948760000000
1!
0$
b110 %
1'
0*
b110 +
#948770000000
0!
0'
#948780000000
1!
b111 %
1'
b111 +
#948790000000
1"
1(
#948800000000
0!
0"
b100 &
0'
0(
b100 ,
#948810000000
1!
b1000 %
1'
b1000 +
#948820000000
0!
0'
#948830000000
1!
b1001 %
1'
b1001 +
#948840000000
0!
0'
#948850000000
1!
b0 %
1'
b0 +
#948860000000
0!
0'
#948870000000
1!
1$
b1 %
1'
1*
b1 +
#948880000000
0!
0'
#948890000000
1!
b10 %
1'
b10 +
#948900000000
0!
0'
#948910000000
1!
b11 %
1'
b11 +
#948920000000
0!
0'
#948930000000
1!
b100 %
1'
b100 +
#948940000000
0!
0'
#948950000000
1!
b101 %
1'
b101 +
#948960000000
0!
0'
#948970000000
1!
b110 %
1'
b110 +
#948980000000
0!
0'
#948990000000
1!
b111 %
1'
b111 +
#949000000000
0!
0'
#949010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#949020000000
0!
0'
#949030000000
1!
b1001 %
1'
b1001 +
#949040000000
0!
0'
#949050000000
1!
b0 %
1'
b0 +
#949060000000
0!
0'
#949070000000
1!
1$
b1 %
1'
1*
b1 +
#949080000000
0!
0'
#949090000000
1!
b10 %
1'
b10 +
#949100000000
0!
0'
#949110000000
1!
b11 %
1'
b11 +
#949120000000
0!
0'
#949130000000
1!
b100 %
1'
b100 +
#949140000000
0!
0'
#949150000000
1!
b101 %
1'
b101 +
#949160000000
0!
0'
#949170000000
1!
0$
b110 %
1'
0*
b110 +
#949180000000
0!
0'
#949190000000
1!
b111 %
1'
b111 +
#949200000000
0!
0'
#949210000000
1!
b1000 %
1'
b1000 +
#949220000000
1"
1(
#949230000000
0!
0"
b100 &
0'
0(
b100 ,
#949240000000
1!
b1001 %
1'
b1001 +
#949250000000
0!
0'
#949260000000
1!
b0 %
1'
b0 +
#949270000000
0!
0'
#949280000000
1!
1$
b1 %
1'
1*
b1 +
#949290000000
0!
0'
#949300000000
1!
b10 %
1'
b10 +
#949310000000
0!
0'
#949320000000
1!
b11 %
1'
b11 +
#949330000000
0!
0'
#949340000000
1!
b100 %
1'
b100 +
#949350000000
0!
0'
#949360000000
1!
b101 %
1'
b101 +
#949370000000
0!
0'
#949380000000
1!
b110 %
1'
b110 +
#949390000000
0!
0'
#949400000000
1!
b111 %
1'
b111 +
#949410000000
0!
0'
#949420000000
1!
0$
b1000 %
1'
0*
b1000 +
#949430000000
0!
0'
#949440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#949450000000
0!
0'
#949460000000
1!
b0 %
1'
b0 +
#949470000000
0!
0'
#949480000000
1!
1$
b1 %
1'
1*
b1 +
#949490000000
0!
0'
#949500000000
1!
b10 %
1'
b10 +
#949510000000
0!
0'
#949520000000
1!
b11 %
1'
b11 +
#949530000000
0!
0'
#949540000000
1!
b100 %
1'
b100 +
#949550000000
0!
0'
#949560000000
1!
b101 %
1'
b101 +
#949570000000
0!
0'
#949580000000
1!
0$
b110 %
1'
0*
b110 +
#949590000000
0!
0'
#949600000000
1!
b111 %
1'
b111 +
#949610000000
0!
0'
#949620000000
1!
b1000 %
1'
b1000 +
#949630000000
0!
0'
#949640000000
1!
b1001 %
1'
b1001 +
#949650000000
1"
1(
#949660000000
0!
0"
b100 &
0'
0(
b100 ,
#949670000000
1!
b0 %
1'
b0 +
#949680000000
0!
0'
#949690000000
1!
1$
b1 %
1'
1*
b1 +
#949700000000
0!
0'
#949710000000
1!
b10 %
1'
b10 +
#949720000000
0!
0'
#949730000000
1!
b11 %
1'
b11 +
#949740000000
0!
0'
#949750000000
1!
b100 %
1'
b100 +
#949760000000
0!
0'
#949770000000
1!
b101 %
1'
b101 +
#949780000000
0!
0'
#949790000000
1!
b110 %
1'
b110 +
#949800000000
0!
0'
#949810000000
1!
b111 %
1'
b111 +
#949820000000
0!
0'
#949830000000
1!
0$
b1000 %
1'
0*
b1000 +
#949840000000
0!
0'
#949850000000
1!
b1001 %
1'
b1001 +
#949860000000
0!
0'
#949870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#949880000000
0!
0'
#949890000000
1!
1$
b1 %
1'
1*
b1 +
#949900000000
0!
0'
#949910000000
1!
b10 %
1'
b10 +
#949920000000
0!
0'
#949930000000
1!
b11 %
1'
b11 +
#949940000000
0!
0'
#949950000000
1!
b100 %
1'
b100 +
#949960000000
0!
0'
#949970000000
1!
b101 %
1'
b101 +
#949980000000
0!
0'
#949990000000
1!
0$
b110 %
1'
0*
b110 +
#950000000000
0!
0'
#950010000000
1!
b111 %
1'
b111 +
#950020000000
0!
0'
#950030000000
1!
b1000 %
1'
b1000 +
#950040000000
0!
0'
#950050000000
1!
b1001 %
1'
b1001 +
#950060000000
0!
0'
#950070000000
1!
b0 %
1'
b0 +
#950080000000
1"
1(
#950090000000
0!
0"
b100 &
0'
0(
b100 ,
#950100000000
1!
1$
b1 %
1'
1*
b1 +
#950110000000
0!
0'
#950120000000
1!
b10 %
1'
b10 +
#950130000000
0!
0'
#950140000000
1!
b11 %
1'
b11 +
#950150000000
0!
0'
#950160000000
1!
b100 %
1'
b100 +
#950170000000
0!
0'
#950180000000
1!
b101 %
1'
b101 +
#950190000000
0!
0'
#950200000000
1!
b110 %
1'
b110 +
#950210000000
0!
0'
#950220000000
1!
b111 %
1'
b111 +
#950230000000
0!
0'
#950240000000
1!
0$
b1000 %
1'
0*
b1000 +
#950250000000
0!
0'
#950260000000
1!
b1001 %
1'
b1001 +
#950270000000
0!
0'
#950280000000
1!
b0 %
1'
b0 +
#950290000000
0!
0'
#950300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#950310000000
0!
0'
#950320000000
1!
b10 %
1'
b10 +
#950330000000
0!
0'
#950340000000
1!
b11 %
1'
b11 +
#950350000000
0!
0'
#950360000000
1!
b100 %
1'
b100 +
#950370000000
0!
0'
#950380000000
1!
b101 %
1'
b101 +
#950390000000
0!
0'
#950400000000
1!
0$
b110 %
1'
0*
b110 +
#950410000000
0!
0'
#950420000000
1!
b111 %
1'
b111 +
#950430000000
0!
0'
#950440000000
1!
b1000 %
1'
b1000 +
#950450000000
0!
0'
#950460000000
1!
b1001 %
1'
b1001 +
#950470000000
0!
0'
#950480000000
1!
b0 %
1'
b0 +
#950490000000
0!
0'
#950500000000
1!
1$
b1 %
1'
1*
b1 +
#950510000000
1"
1(
#950520000000
0!
0"
b100 &
0'
0(
b100 ,
#950530000000
1!
b10 %
1'
b10 +
#950540000000
0!
0'
#950550000000
1!
b11 %
1'
b11 +
#950560000000
0!
0'
#950570000000
1!
b100 %
1'
b100 +
#950580000000
0!
0'
#950590000000
1!
b101 %
1'
b101 +
#950600000000
0!
0'
#950610000000
1!
b110 %
1'
b110 +
#950620000000
0!
0'
#950630000000
1!
b111 %
1'
b111 +
#950640000000
0!
0'
#950650000000
1!
0$
b1000 %
1'
0*
b1000 +
#950660000000
0!
0'
#950670000000
1!
b1001 %
1'
b1001 +
#950680000000
0!
0'
#950690000000
1!
b0 %
1'
b0 +
#950700000000
0!
0'
#950710000000
1!
1$
b1 %
1'
1*
b1 +
#950720000000
0!
0'
#950730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#950740000000
0!
0'
#950750000000
1!
b11 %
1'
b11 +
#950760000000
0!
0'
#950770000000
1!
b100 %
1'
b100 +
#950780000000
0!
0'
#950790000000
1!
b101 %
1'
b101 +
#950800000000
0!
0'
#950810000000
1!
0$
b110 %
1'
0*
b110 +
#950820000000
0!
0'
#950830000000
1!
b111 %
1'
b111 +
#950840000000
0!
0'
#950850000000
1!
b1000 %
1'
b1000 +
#950860000000
0!
0'
#950870000000
1!
b1001 %
1'
b1001 +
#950880000000
0!
0'
#950890000000
1!
b0 %
1'
b0 +
#950900000000
0!
0'
#950910000000
1!
1$
b1 %
1'
1*
b1 +
#950920000000
0!
0'
#950930000000
1!
b10 %
1'
b10 +
#950940000000
1"
1(
#950950000000
0!
0"
b100 &
0'
0(
b100 ,
#950960000000
1!
b11 %
1'
b11 +
#950970000000
0!
0'
#950980000000
1!
b100 %
1'
b100 +
#950990000000
0!
0'
#951000000000
1!
b101 %
1'
b101 +
#951010000000
0!
0'
#951020000000
1!
b110 %
1'
b110 +
#951030000000
0!
0'
#951040000000
1!
b111 %
1'
b111 +
#951050000000
0!
0'
#951060000000
1!
0$
b1000 %
1'
0*
b1000 +
#951070000000
0!
0'
#951080000000
1!
b1001 %
1'
b1001 +
#951090000000
0!
0'
#951100000000
1!
b0 %
1'
b0 +
#951110000000
0!
0'
#951120000000
1!
1$
b1 %
1'
1*
b1 +
#951130000000
0!
0'
#951140000000
1!
b10 %
1'
b10 +
#951150000000
0!
0'
#951160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#951170000000
0!
0'
#951180000000
1!
b100 %
1'
b100 +
#951190000000
0!
0'
#951200000000
1!
b101 %
1'
b101 +
#951210000000
0!
0'
#951220000000
1!
0$
b110 %
1'
0*
b110 +
#951230000000
0!
0'
#951240000000
1!
b111 %
1'
b111 +
#951250000000
0!
0'
#951260000000
1!
b1000 %
1'
b1000 +
#951270000000
0!
0'
#951280000000
1!
b1001 %
1'
b1001 +
#951290000000
0!
0'
#951300000000
1!
b0 %
1'
b0 +
#951310000000
0!
0'
#951320000000
1!
1$
b1 %
1'
1*
b1 +
#951330000000
0!
0'
#951340000000
1!
b10 %
1'
b10 +
#951350000000
0!
0'
#951360000000
1!
b11 %
1'
b11 +
#951370000000
1"
1(
#951380000000
0!
0"
b100 &
0'
0(
b100 ,
#951390000000
1!
b100 %
1'
b100 +
#951400000000
0!
0'
#951410000000
1!
b101 %
1'
b101 +
#951420000000
0!
0'
#951430000000
1!
b110 %
1'
b110 +
#951440000000
0!
0'
#951450000000
1!
b111 %
1'
b111 +
#951460000000
0!
0'
#951470000000
1!
0$
b1000 %
1'
0*
b1000 +
#951480000000
0!
0'
#951490000000
1!
b1001 %
1'
b1001 +
#951500000000
0!
0'
#951510000000
1!
b0 %
1'
b0 +
#951520000000
0!
0'
#951530000000
1!
1$
b1 %
1'
1*
b1 +
#951540000000
0!
0'
#951550000000
1!
b10 %
1'
b10 +
#951560000000
0!
0'
#951570000000
1!
b11 %
1'
b11 +
#951580000000
0!
0'
#951590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#951600000000
0!
0'
#951610000000
1!
b101 %
1'
b101 +
#951620000000
0!
0'
#951630000000
1!
0$
b110 %
1'
0*
b110 +
#951640000000
0!
0'
#951650000000
1!
b111 %
1'
b111 +
#951660000000
0!
0'
#951670000000
1!
b1000 %
1'
b1000 +
#951680000000
0!
0'
#951690000000
1!
b1001 %
1'
b1001 +
#951700000000
0!
0'
#951710000000
1!
b0 %
1'
b0 +
#951720000000
0!
0'
#951730000000
1!
1$
b1 %
1'
1*
b1 +
#951740000000
0!
0'
#951750000000
1!
b10 %
1'
b10 +
#951760000000
0!
0'
#951770000000
1!
b11 %
1'
b11 +
#951780000000
0!
0'
#951790000000
1!
b100 %
1'
b100 +
#951800000000
1"
1(
#951810000000
0!
0"
b100 &
0'
0(
b100 ,
#951820000000
1!
b101 %
1'
b101 +
#951830000000
0!
0'
#951840000000
1!
b110 %
1'
b110 +
#951850000000
0!
0'
#951860000000
1!
b111 %
1'
b111 +
#951870000000
0!
0'
#951880000000
1!
0$
b1000 %
1'
0*
b1000 +
#951890000000
0!
0'
#951900000000
1!
b1001 %
1'
b1001 +
#951910000000
0!
0'
#951920000000
1!
b0 %
1'
b0 +
#951930000000
0!
0'
#951940000000
1!
1$
b1 %
1'
1*
b1 +
#951950000000
0!
0'
#951960000000
1!
b10 %
1'
b10 +
#951970000000
0!
0'
#951980000000
1!
b11 %
1'
b11 +
#951990000000
0!
0'
#952000000000
1!
b100 %
1'
b100 +
#952010000000
0!
0'
#952020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#952030000000
0!
0'
#952040000000
1!
0$
b110 %
1'
0*
b110 +
#952050000000
0!
0'
#952060000000
1!
b111 %
1'
b111 +
#952070000000
0!
0'
#952080000000
1!
b1000 %
1'
b1000 +
#952090000000
0!
0'
#952100000000
1!
b1001 %
1'
b1001 +
#952110000000
0!
0'
#952120000000
1!
b0 %
1'
b0 +
#952130000000
0!
0'
#952140000000
1!
1$
b1 %
1'
1*
b1 +
#952150000000
0!
0'
#952160000000
1!
b10 %
1'
b10 +
#952170000000
0!
0'
#952180000000
1!
b11 %
1'
b11 +
#952190000000
0!
0'
#952200000000
1!
b100 %
1'
b100 +
#952210000000
0!
0'
#952220000000
1!
b101 %
1'
b101 +
#952230000000
1"
1(
#952240000000
0!
0"
b100 &
0'
0(
b100 ,
#952250000000
1!
b110 %
1'
b110 +
#952260000000
0!
0'
#952270000000
1!
b111 %
1'
b111 +
#952280000000
0!
0'
#952290000000
1!
0$
b1000 %
1'
0*
b1000 +
#952300000000
0!
0'
#952310000000
1!
b1001 %
1'
b1001 +
#952320000000
0!
0'
#952330000000
1!
b0 %
1'
b0 +
#952340000000
0!
0'
#952350000000
1!
1$
b1 %
1'
1*
b1 +
#952360000000
0!
0'
#952370000000
1!
b10 %
1'
b10 +
#952380000000
0!
0'
#952390000000
1!
b11 %
1'
b11 +
#952400000000
0!
0'
#952410000000
1!
b100 %
1'
b100 +
#952420000000
0!
0'
#952430000000
1!
b101 %
1'
b101 +
#952440000000
0!
0'
#952450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#952460000000
0!
0'
#952470000000
1!
b111 %
1'
b111 +
#952480000000
0!
0'
#952490000000
1!
b1000 %
1'
b1000 +
#952500000000
0!
0'
#952510000000
1!
b1001 %
1'
b1001 +
#952520000000
0!
0'
#952530000000
1!
b0 %
1'
b0 +
#952540000000
0!
0'
#952550000000
1!
1$
b1 %
1'
1*
b1 +
#952560000000
0!
0'
#952570000000
1!
b10 %
1'
b10 +
#952580000000
0!
0'
#952590000000
1!
b11 %
1'
b11 +
#952600000000
0!
0'
#952610000000
1!
b100 %
1'
b100 +
#952620000000
0!
0'
#952630000000
1!
b101 %
1'
b101 +
#952640000000
0!
0'
#952650000000
1!
0$
b110 %
1'
0*
b110 +
#952660000000
1"
1(
#952670000000
0!
0"
b100 &
0'
0(
b100 ,
#952680000000
1!
1$
b111 %
1'
1*
b111 +
#952690000000
0!
0'
#952700000000
1!
0$
b1000 %
1'
0*
b1000 +
#952710000000
0!
0'
#952720000000
1!
b1001 %
1'
b1001 +
#952730000000
0!
0'
#952740000000
1!
b0 %
1'
b0 +
#952750000000
0!
0'
#952760000000
1!
1$
b1 %
1'
1*
b1 +
#952770000000
0!
0'
#952780000000
1!
b10 %
1'
b10 +
#952790000000
0!
0'
#952800000000
1!
b11 %
1'
b11 +
#952810000000
0!
0'
#952820000000
1!
b100 %
1'
b100 +
#952830000000
0!
0'
#952840000000
1!
b101 %
1'
b101 +
#952850000000
0!
0'
#952860000000
1!
b110 %
1'
b110 +
#952870000000
0!
0'
#952880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#952890000000
0!
0'
#952900000000
1!
b1000 %
1'
b1000 +
#952910000000
0!
0'
#952920000000
1!
b1001 %
1'
b1001 +
#952930000000
0!
0'
#952940000000
1!
b0 %
1'
b0 +
#952950000000
0!
0'
#952960000000
1!
1$
b1 %
1'
1*
b1 +
#952970000000
0!
0'
#952980000000
1!
b10 %
1'
b10 +
#952990000000
0!
0'
#953000000000
1!
b11 %
1'
b11 +
#953010000000
0!
0'
#953020000000
1!
b100 %
1'
b100 +
#953030000000
0!
0'
#953040000000
1!
b101 %
1'
b101 +
#953050000000
0!
0'
#953060000000
1!
0$
b110 %
1'
0*
b110 +
#953070000000
0!
0'
#953080000000
1!
b111 %
1'
b111 +
#953090000000
1"
1(
#953100000000
0!
0"
b100 &
0'
0(
b100 ,
#953110000000
1!
b1000 %
1'
b1000 +
#953120000000
0!
0'
#953130000000
1!
b1001 %
1'
b1001 +
#953140000000
0!
0'
#953150000000
1!
b0 %
1'
b0 +
#953160000000
0!
0'
#953170000000
1!
1$
b1 %
1'
1*
b1 +
#953180000000
0!
0'
#953190000000
1!
b10 %
1'
b10 +
#953200000000
0!
0'
#953210000000
1!
b11 %
1'
b11 +
#953220000000
0!
0'
#953230000000
1!
b100 %
1'
b100 +
#953240000000
0!
0'
#953250000000
1!
b101 %
1'
b101 +
#953260000000
0!
0'
#953270000000
1!
b110 %
1'
b110 +
#953280000000
0!
0'
#953290000000
1!
b111 %
1'
b111 +
#953300000000
0!
0'
#953310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#953320000000
0!
0'
#953330000000
1!
b1001 %
1'
b1001 +
#953340000000
0!
0'
#953350000000
1!
b0 %
1'
b0 +
#953360000000
0!
0'
#953370000000
1!
1$
b1 %
1'
1*
b1 +
#953380000000
0!
0'
#953390000000
1!
b10 %
1'
b10 +
#953400000000
0!
0'
#953410000000
1!
b11 %
1'
b11 +
#953420000000
0!
0'
#953430000000
1!
b100 %
1'
b100 +
#953440000000
0!
0'
#953450000000
1!
b101 %
1'
b101 +
#953460000000
0!
0'
#953470000000
1!
0$
b110 %
1'
0*
b110 +
#953480000000
0!
0'
#953490000000
1!
b111 %
1'
b111 +
#953500000000
0!
0'
#953510000000
1!
b1000 %
1'
b1000 +
#953520000000
1"
1(
#953530000000
0!
0"
b100 &
0'
0(
b100 ,
#953540000000
1!
b1001 %
1'
b1001 +
#953550000000
0!
0'
#953560000000
1!
b0 %
1'
b0 +
#953570000000
0!
0'
#953580000000
1!
1$
b1 %
1'
1*
b1 +
#953590000000
0!
0'
#953600000000
1!
b10 %
1'
b10 +
#953610000000
0!
0'
#953620000000
1!
b11 %
1'
b11 +
#953630000000
0!
0'
#953640000000
1!
b100 %
1'
b100 +
#953650000000
0!
0'
#953660000000
1!
b101 %
1'
b101 +
#953670000000
0!
0'
#953680000000
1!
b110 %
1'
b110 +
#953690000000
0!
0'
#953700000000
1!
b111 %
1'
b111 +
#953710000000
0!
0'
#953720000000
1!
0$
b1000 %
1'
0*
b1000 +
#953730000000
0!
0'
#953740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#953750000000
0!
0'
#953760000000
1!
b0 %
1'
b0 +
#953770000000
0!
0'
#953780000000
1!
1$
b1 %
1'
1*
b1 +
#953790000000
0!
0'
#953800000000
1!
b10 %
1'
b10 +
#953810000000
0!
0'
#953820000000
1!
b11 %
1'
b11 +
#953830000000
0!
0'
#953840000000
1!
b100 %
1'
b100 +
#953850000000
0!
0'
#953860000000
1!
b101 %
1'
b101 +
#953870000000
0!
0'
#953880000000
1!
0$
b110 %
1'
0*
b110 +
#953890000000
0!
0'
#953900000000
1!
b111 %
1'
b111 +
#953910000000
0!
0'
#953920000000
1!
b1000 %
1'
b1000 +
#953930000000
0!
0'
#953940000000
1!
b1001 %
1'
b1001 +
#953950000000
1"
1(
#953960000000
0!
0"
b100 &
0'
0(
b100 ,
#953970000000
1!
b0 %
1'
b0 +
#953980000000
0!
0'
#953990000000
1!
1$
b1 %
1'
1*
b1 +
#954000000000
0!
0'
#954010000000
1!
b10 %
1'
b10 +
#954020000000
0!
0'
#954030000000
1!
b11 %
1'
b11 +
#954040000000
0!
0'
#954050000000
1!
b100 %
1'
b100 +
#954060000000
0!
0'
#954070000000
1!
b101 %
1'
b101 +
#954080000000
0!
0'
#954090000000
1!
b110 %
1'
b110 +
#954100000000
0!
0'
#954110000000
1!
b111 %
1'
b111 +
#954120000000
0!
0'
#954130000000
1!
0$
b1000 %
1'
0*
b1000 +
#954140000000
0!
0'
#954150000000
1!
b1001 %
1'
b1001 +
#954160000000
0!
0'
#954170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#954180000000
0!
0'
#954190000000
1!
1$
b1 %
1'
1*
b1 +
#954200000000
0!
0'
#954210000000
1!
b10 %
1'
b10 +
#954220000000
0!
0'
#954230000000
1!
b11 %
1'
b11 +
#954240000000
0!
0'
#954250000000
1!
b100 %
1'
b100 +
#954260000000
0!
0'
#954270000000
1!
b101 %
1'
b101 +
#954280000000
0!
0'
#954290000000
1!
0$
b110 %
1'
0*
b110 +
#954300000000
0!
0'
#954310000000
1!
b111 %
1'
b111 +
#954320000000
0!
0'
#954330000000
1!
b1000 %
1'
b1000 +
#954340000000
0!
0'
#954350000000
1!
b1001 %
1'
b1001 +
#954360000000
0!
0'
#954370000000
1!
b0 %
1'
b0 +
#954380000000
1"
1(
#954390000000
0!
0"
b100 &
0'
0(
b100 ,
#954400000000
1!
1$
b1 %
1'
1*
b1 +
#954410000000
0!
0'
#954420000000
1!
b10 %
1'
b10 +
#954430000000
0!
0'
#954440000000
1!
b11 %
1'
b11 +
#954450000000
0!
0'
#954460000000
1!
b100 %
1'
b100 +
#954470000000
0!
0'
#954480000000
1!
b101 %
1'
b101 +
#954490000000
0!
0'
#954500000000
1!
b110 %
1'
b110 +
#954510000000
0!
0'
#954520000000
1!
b111 %
1'
b111 +
#954530000000
0!
0'
#954540000000
1!
0$
b1000 %
1'
0*
b1000 +
#954550000000
0!
0'
#954560000000
1!
b1001 %
1'
b1001 +
#954570000000
0!
0'
#954580000000
1!
b0 %
1'
b0 +
#954590000000
0!
0'
#954600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#954610000000
0!
0'
#954620000000
1!
b10 %
1'
b10 +
#954630000000
0!
0'
#954640000000
1!
b11 %
1'
b11 +
#954650000000
0!
0'
#954660000000
1!
b100 %
1'
b100 +
#954670000000
0!
0'
#954680000000
1!
b101 %
1'
b101 +
#954690000000
0!
0'
#954700000000
1!
0$
b110 %
1'
0*
b110 +
#954710000000
0!
0'
#954720000000
1!
b111 %
1'
b111 +
#954730000000
0!
0'
#954740000000
1!
b1000 %
1'
b1000 +
#954750000000
0!
0'
#954760000000
1!
b1001 %
1'
b1001 +
#954770000000
0!
0'
#954780000000
1!
b0 %
1'
b0 +
#954790000000
0!
0'
#954800000000
1!
1$
b1 %
1'
1*
b1 +
#954810000000
1"
1(
#954820000000
0!
0"
b100 &
0'
0(
b100 ,
#954830000000
1!
b10 %
1'
b10 +
#954840000000
0!
0'
#954850000000
1!
b11 %
1'
b11 +
#954860000000
0!
0'
#954870000000
1!
b100 %
1'
b100 +
#954880000000
0!
0'
#954890000000
1!
b101 %
1'
b101 +
#954900000000
0!
0'
#954910000000
1!
b110 %
1'
b110 +
#954920000000
0!
0'
#954930000000
1!
b111 %
1'
b111 +
#954940000000
0!
0'
#954950000000
1!
0$
b1000 %
1'
0*
b1000 +
#954960000000
0!
0'
#954970000000
1!
b1001 %
1'
b1001 +
#954980000000
0!
0'
#954990000000
1!
b0 %
1'
b0 +
#955000000000
0!
0'
#955010000000
1!
1$
b1 %
1'
1*
b1 +
#955020000000
0!
0'
#955030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#955040000000
0!
0'
#955050000000
1!
b11 %
1'
b11 +
#955060000000
0!
0'
#955070000000
1!
b100 %
1'
b100 +
#955080000000
0!
0'
#955090000000
1!
b101 %
1'
b101 +
#955100000000
0!
0'
#955110000000
1!
0$
b110 %
1'
0*
b110 +
#955120000000
0!
0'
#955130000000
1!
b111 %
1'
b111 +
#955140000000
0!
0'
#955150000000
1!
b1000 %
1'
b1000 +
#955160000000
0!
0'
#955170000000
1!
b1001 %
1'
b1001 +
#955180000000
0!
0'
#955190000000
1!
b0 %
1'
b0 +
#955200000000
0!
0'
#955210000000
1!
1$
b1 %
1'
1*
b1 +
#955220000000
0!
0'
#955230000000
1!
b10 %
1'
b10 +
#955240000000
1"
1(
#955250000000
0!
0"
b100 &
0'
0(
b100 ,
#955260000000
1!
b11 %
1'
b11 +
#955270000000
0!
0'
#955280000000
1!
b100 %
1'
b100 +
#955290000000
0!
0'
#955300000000
1!
b101 %
1'
b101 +
#955310000000
0!
0'
#955320000000
1!
b110 %
1'
b110 +
#955330000000
0!
0'
#955340000000
1!
b111 %
1'
b111 +
#955350000000
0!
0'
#955360000000
1!
0$
b1000 %
1'
0*
b1000 +
#955370000000
0!
0'
#955380000000
1!
b1001 %
1'
b1001 +
#955390000000
0!
0'
#955400000000
1!
b0 %
1'
b0 +
#955410000000
0!
0'
#955420000000
1!
1$
b1 %
1'
1*
b1 +
#955430000000
0!
0'
#955440000000
1!
b10 %
1'
b10 +
#955450000000
0!
0'
#955460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#955470000000
0!
0'
#955480000000
1!
b100 %
1'
b100 +
#955490000000
0!
0'
#955500000000
1!
b101 %
1'
b101 +
#955510000000
0!
0'
#955520000000
1!
0$
b110 %
1'
0*
b110 +
#955530000000
0!
0'
#955540000000
1!
b111 %
1'
b111 +
#955550000000
0!
0'
#955560000000
1!
b1000 %
1'
b1000 +
#955570000000
0!
0'
#955580000000
1!
b1001 %
1'
b1001 +
#955590000000
0!
0'
#955600000000
1!
b0 %
1'
b0 +
#955610000000
0!
0'
#955620000000
1!
1$
b1 %
1'
1*
b1 +
#955630000000
0!
0'
#955640000000
1!
b10 %
1'
b10 +
#955650000000
0!
0'
#955660000000
1!
b11 %
1'
b11 +
#955670000000
1"
1(
#955680000000
0!
0"
b100 &
0'
0(
b100 ,
#955690000000
1!
b100 %
1'
b100 +
#955700000000
0!
0'
#955710000000
1!
b101 %
1'
b101 +
#955720000000
0!
0'
#955730000000
1!
b110 %
1'
b110 +
#955740000000
0!
0'
#955750000000
1!
b111 %
1'
b111 +
#955760000000
0!
0'
#955770000000
1!
0$
b1000 %
1'
0*
b1000 +
#955780000000
0!
0'
#955790000000
1!
b1001 %
1'
b1001 +
#955800000000
0!
0'
#955810000000
1!
b0 %
1'
b0 +
#955820000000
0!
0'
#955830000000
1!
1$
b1 %
1'
1*
b1 +
#955840000000
0!
0'
#955850000000
1!
b10 %
1'
b10 +
#955860000000
0!
0'
#955870000000
1!
b11 %
1'
b11 +
#955880000000
0!
0'
#955890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#955900000000
0!
0'
#955910000000
1!
b101 %
1'
b101 +
#955920000000
0!
0'
#955930000000
1!
0$
b110 %
1'
0*
b110 +
#955940000000
0!
0'
#955950000000
1!
b111 %
1'
b111 +
#955960000000
0!
0'
#955970000000
1!
b1000 %
1'
b1000 +
#955980000000
0!
0'
#955990000000
1!
b1001 %
1'
b1001 +
#956000000000
0!
0'
#956010000000
1!
b0 %
1'
b0 +
#956020000000
0!
0'
#956030000000
1!
1$
b1 %
1'
1*
b1 +
#956040000000
0!
0'
#956050000000
1!
b10 %
1'
b10 +
#956060000000
0!
0'
#956070000000
1!
b11 %
1'
b11 +
#956080000000
0!
0'
#956090000000
1!
b100 %
1'
b100 +
#956100000000
1"
1(
#956110000000
0!
0"
b100 &
0'
0(
b100 ,
#956120000000
1!
b101 %
1'
b101 +
#956130000000
0!
0'
#956140000000
1!
b110 %
1'
b110 +
#956150000000
0!
0'
#956160000000
1!
b111 %
1'
b111 +
#956170000000
0!
0'
#956180000000
1!
0$
b1000 %
1'
0*
b1000 +
#956190000000
0!
0'
#956200000000
1!
b1001 %
1'
b1001 +
#956210000000
0!
0'
#956220000000
1!
b0 %
1'
b0 +
#956230000000
0!
0'
#956240000000
1!
1$
b1 %
1'
1*
b1 +
#956250000000
0!
0'
#956260000000
1!
b10 %
1'
b10 +
#956270000000
0!
0'
#956280000000
1!
b11 %
1'
b11 +
#956290000000
0!
0'
#956300000000
1!
b100 %
1'
b100 +
#956310000000
0!
0'
#956320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#956330000000
0!
0'
#956340000000
1!
0$
b110 %
1'
0*
b110 +
#956350000000
0!
0'
#956360000000
1!
b111 %
1'
b111 +
#956370000000
0!
0'
#956380000000
1!
b1000 %
1'
b1000 +
#956390000000
0!
0'
#956400000000
1!
b1001 %
1'
b1001 +
#956410000000
0!
0'
#956420000000
1!
b0 %
1'
b0 +
#956430000000
0!
0'
#956440000000
1!
1$
b1 %
1'
1*
b1 +
#956450000000
0!
0'
#956460000000
1!
b10 %
1'
b10 +
#956470000000
0!
0'
#956480000000
1!
b11 %
1'
b11 +
#956490000000
0!
0'
#956500000000
1!
b100 %
1'
b100 +
#956510000000
0!
0'
#956520000000
1!
b101 %
1'
b101 +
#956530000000
1"
1(
#956540000000
0!
0"
b100 &
0'
0(
b100 ,
#956550000000
1!
b110 %
1'
b110 +
#956560000000
0!
0'
#956570000000
1!
b111 %
1'
b111 +
#956580000000
0!
0'
#956590000000
1!
0$
b1000 %
1'
0*
b1000 +
#956600000000
0!
0'
#956610000000
1!
b1001 %
1'
b1001 +
#956620000000
0!
0'
#956630000000
1!
b0 %
1'
b0 +
#956640000000
0!
0'
#956650000000
1!
1$
b1 %
1'
1*
b1 +
#956660000000
0!
0'
#956670000000
1!
b10 %
1'
b10 +
#956680000000
0!
0'
#956690000000
1!
b11 %
1'
b11 +
#956700000000
0!
0'
#956710000000
1!
b100 %
1'
b100 +
#956720000000
0!
0'
#956730000000
1!
b101 %
1'
b101 +
#956740000000
0!
0'
#956750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#956760000000
0!
0'
#956770000000
1!
b111 %
1'
b111 +
#956780000000
0!
0'
#956790000000
1!
b1000 %
1'
b1000 +
#956800000000
0!
0'
#956810000000
1!
b1001 %
1'
b1001 +
#956820000000
0!
0'
#956830000000
1!
b0 %
1'
b0 +
#956840000000
0!
0'
#956850000000
1!
1$
b1 %
1'
1*
b1 +
#956860000000
0!
0'
#956870000000
1!
b10 %
1'
b10 +
#956880000000
0!
0'
#956890000000
1!
b11 %
1'
b11 +
#956900000000
0!
0'
#956910000000
1!
b100 %
1'
b100 +
#956920000000
0!
0'
#956930000000
1!
b101 %
1'
b101 +
#956940000000
0!
0'
#956950000000
1!
0$
b110 %
1'
0*
b110 +
#956960000000
1"
1(
#956970000000
0!
0"
b100 &
0'
0(
b100 ,
#956980000000
1!
1$
b111 %
1'
1*
b111 +
#956990000000
0!
0'
#957000000000
1!
0$
b1000 %
1'
0*
b1000 +
#957010000000
0!
0'
#957020000000
1!
b1001 %
1'
b1001 +
#957030000000
0!
0'
#957040000000
1!
b0 %
1'
b0 +
#957050000000
0!
0'
#957060000000
1!
1$
b1 %
1'
1*
b1 +
#957070000000
0!
0'
#957080000000
1!
b10 %
1'
b10 +
#957090000000
0!
0'
#957100000000
1!
b11 %
1'
b11 +
#957110000000
0!
0'
#957120000000
1!
b100 %
1'
b100 +
#957130000000
0!
0'
#957140000000
1!
b101 %
1'
b101 +
#957150000000
0!
0'
#957160000000
1!
b110 %
1'
b110 +
#957170000000
0!
0'
#957180000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#957190000000
0!
0'
#957200000000
1!
b1000 %
1'
b1000 +
#957210000000
0!
0'
#957220000000
1!
b1001 %
1'
b1001 +
#957230000000
0!
0'
#957240000000
1!
b0 %
1'
b0 +
#957250000000
0!
0'
#957260000000
1!
1$
b1 %
1'
1*
b1 +
#957270000000
0!
0'
#957280000000
1!
b10 %
1'
b10 +
#957290000000
0!
0'
#957300000000
1!
b11 %
1'
b11 +
#957310000000
0!
0'
#957320000000
1!
b100 %
1'
b100 +
#957330000000
0!
0'
#957340000000
1!
b101 %
1'
b101 +
#957350000000
0!
0'
#957360000000
1!
0$
b110 %
1'
0*
b110 +
#957370000000
0!
0'
#957380000000
1!
b111 %
1'
b111 +
#957390000000
1"
1(
#957400000000
0!
0"
b100 &
0'
0(
b100 ,
#957410000000
1!
b1000 %
1'
b1000 +
#957420000000
0!
0'
#957430000000
1!
b1001 %
1'
b1001 +
#957440000000
0!
0'
#957450000000
1!
b0 %
1'
b0 +
#957460000000
0!
0'
#957470000000
1!
1$
b1 %
1'
1*
b1 +
#957480000000
0!
0'
#957490000000
1!
b10 %
1'
b10 +
#957500000000
0!
0'
#957510000000
1!
b11 %
1'
b11 +
#957520000000
0!
0'
#957530000000
1!
b100 %
1'
b100 +
#957540000000
0!
0'
#957550000000
1!
b101 %
1'
b101 +
#957560000000
0!
0'
#957570000000
1!
b110 %
1'
b110 +
#957580000000
0!
0'
#957590000000
1!
b111 %
1'
b111 +
#957600000000
0!
0'
#957610000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#957620000000
0!
0'
#957630000000
1!
b1001 %
1'
b1001 +
#957640000000
0!
0'
#957650000000
1!
b0 %
1'
b0 +
#957660000000
0!
0'
#957670000000
1!
1$
b1 %
1'
1*
b1 +
#957680000000
0!
0'
#957690000000
1!
b10 %
1'
b10 +
#957700000000
0!
0'
#957710000000
1!
b11 %
1'
b11 +
#957720000000
0!
0'
#957730000000
1!
b100 %
1'
b100 +
#957740000000
0!
0'
#957750000000
1!
b101 %
1'
b101 +
#957760000000
0!
0'
#957770000000
1!
0$
b110 %
1'
0*
b110 +
#957780000000
0!
0'
#957790000000
1!
b111 %
1'
b111 +
#957800000000
0!
0'
#957810000000
1!
b1000 %
1'
b1000 +
#957820000000
1"
1(
#957830000000
0!
0"
b100 &
0'
0(
b100 ,
#957840000000
1!
b1001 %
1'
b1001 +
#957850000000
0!
0'
#957860000000
1!
b0 %
1'
b0 +
#957870000000
0!
0'
#957880000000
1!
1$
b1 %
1'
1*
b1 +
#957890000000
0!
0'
#957900000000
1!
b10 %
1'
b10 +
#957910000000
0!
0'
#957920000000
1!
b11 %
1'
b11 +
#957930000000
0!
0'
#957940000000
1!
b100 %
1'
b100 +
#957950000000
0!
0'
#957960000000
1!
b101 %
1'
b101 +
#957970000000
0!
0'
#957980000000
1!
b110 %
1'
b110 +
#957990000000
0!
0'
#958000000000
1!
b111 %
1'
b111 +
#958010000000
0!
0'
#958020000000
1!
0$
b1000 %
1'
0*
b1000 +
#958030000000
0!
0'
#958040000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#958050000000
0!
0'
#958060000000
1!
b0 %
1'
b0 +
#958070000000
0!
0'
#958080000000
1!
1$
b1 %
1'
1*
b1 +
#958090000000
0!
0'
#958100000000
1!
b10 %
1'
b10 +
#958110000000
0!
0'
#958120000000
1!
b11 %
1'
b11 +
#958130000000
0!
0'
#958140000000
1!
b100 %
1'
b100 +
#958150000000
0!
0'
#958160000000
1!
b101 %
1'
b101 +
#958170000000
0!
0'
#958180000000
1!
0$
b110 %
1'
0*
b110 +
#958190000000
0!
0'
#958200000000
1!
b111 %
1'
b111 +
#958210000000
0!
0'
#958220000000
1!
b1000 %
1'
b1000 +
#958230000000
0!
0'
#958240000000
1!
b1001 %
1'
b1001 +
#958250000000
1"
1(
#958260000000
0!
0"
b100 &
0'
0(
b100 ,
#958270000000
1!
b0 %
1'
b0 +
#958280000000
0!
0'
#958290000000
1!
1$
b1 %
1'
1*
b1 +
#958300000000
0!
0'
#958310000000
1!
b10 %
1'
b10 +
#958320000000
0!
0'
#958330000000
1!
b11 %
1'
b11 +
#958340000000
0!
0'
#958350000000
1!
b100 %
1'
b100 +
#958360000000
0!
0'
#958370000000
1!
b101 %
1'
b101 +
#958380000000
0!
0'
#958390000000
1!
b110 %
1'
b110 +
#958400000000
0!
0'
#958410000000
1!
b111 %
1'
b111 +
#958420000000
0!
0'
#958430000000
1!
0$
b1000 %
1'
0*
b1000 +
#958440000000
0!
0'
#958450000000
1!
b1001 %
1'
b1001 +
#958460000000
0!
0'
#958470000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#958480000000
0!
0'
#958490000000
1!
1$
b1 %
1'
1*
b1 +
#958500000000
0!
0'
#958510000000
1!
b10 %
1'
b10 +
#958520000000
0!
0'
#958530000000
1!
b11 %
1'
b11 +
#958540000000
0!
0'
#958550000000
1!
b100 %
1'
b100 +
#958560000000
0!
0'
#958570000000
1!
b101 %
1'
b101 +
#958580000000
0!
0'
#958590000000
1!
0$
b110 %
1'
0*
b110 +
#958600000000
0!
0'
#958610000000
1!
b111 %
1'
b111 +
#958620000000
0!
0'
#958630000000
1!
b1000 %
1'
b1000 +
#958640000000
0!
0'
#958650000000
1!
b1001 %
1'
b1001 +
#958660000000
0!
0'
#958670000000
1!
b0 %
1'
b0 +
#958680000000
1"
1(
#958690000000
0!
0"
b100 &
0'
0(
b100 ,
#958700000000
1!
1$
b1 %
1'
1*
b1 +
#958710000000
0!
0'
#958720000000
1!
b10 %
1'
b10 +
#958730000000
0!
0'
#958740000000
1!
b11 %
1'
b11 +
#958750000000
0!
0'
#958760000000
1!
b100 %
1'
b100 +
#958770000000
0!
0'
#958780000000
1!
b101 %
1'
b101 +
#958790000000
0!
0'
#958800000000
1!
b110 %
1'
b110 +
#958810000000
0!
0'
#958820000000
1!
b111 %
1'
b111 +
#958830000000
0!
0'
#958840000000
1!
0$
b1000 %
1'
0*
b1000 +
#958850000000
0!
0'
#958860000000
1!
b1001 %
1'
b1001 +
#958870000000
0!
0'
#958880000000
1!
b0 %
1'
b0 +
#958890000000
0!
0'
#958900000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#958910000000
0!
0'
#958920000000
1!
b10 %
1'
b10 +
#958930000000
0!
0'
#958940000000
1!
b11 %
1'
b11 +
#958950000000
0!
0'
#958960000000
1!
b100 %
1'
b100 +
#958970000000
0!
0'
#958980000000
1!
b101 %
1'
b101 +
#958990000000
0!
0'
#959000000000
1!
0$
b110 %
1'
0*
b110 +
#959010000000
0!
0'
#959020000000
1!
b111 %
1'
b111 +
#959030000000
0!
0'
#959040000000
1!
b1000 %
1'
b1000 +
#959050000000
0!
0'
#959060000000
1!
b1001 %
1'
b1001 +
#959070000000
0!
0'
#959080000000
1!
b0 %
1'
b0 +
#959090000000
0!
0'
#959100000000
1!
1$
b1 %
1'
1*
b1 +
#959110000000
1"
1(
#959120000000
0!
0"
b100 &
0'
0(
b100 ,
#959130000000
1!
b10 %
1'
b10 +
#959140000000
0!
0'
#959150000000
1!
b11 %
1'
b11 +
#959160000000
0!
0'
#959170000000
1!
b100 %
1'
b100 +
#959180000000
0!
0'
#959190000000
1!
b101 %
1'
b101 +
#959200000000
0!
0'
#959210000000
1!
b110 %
1'
b110 +
#959220000000
0!
0'
#959230000000
1!
b111 %
1'
b111 +
#959240000000
0!
0'
#959250000000
1!
0$
b1000 %
1'
0*
b1000 +
#959260000000
0!
0'
#959270000000
1!
b1001 %
1'
b1001 +
#959280000000
0!
0'
#959290000000
1!
b0 %
1'
b0 +
#959300000000
0!
0'
#959310000000
1!
1$
b1 %
1'
1*
b1 +
#959320000000
0!
0'
#959330000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#959340000000
0!
0'
#959350000000
1!
b11 %
1'
b11 +
#959360000000
0!
0'
#959370000000
1!
b100 %
1'
b100 +
#959380000000
0!
0'
#959390000000
1!
b101 %
1'
b101 +
#959400000000
0!
0'
#959410000000
1!
0$
b110 %
1'
0*
b110 +
#959420000000
0!
0'
#959430000000
1!
b111 %
1'
b111 +
#959440000000
0!
0'
#959450000000
1!
b1000 %
1'
b1000 +
#959460000000
0!
0'
#959470000000
1!
b1001 %
1'
b1001 +
#959480000000
0!
0'
#959490000000
1!
b0 %
1'
b0 +
#959500000000
0!
0'
#959510000000
1!
1$
b1 %
1'
1*
b1 +
#959520000000
0!
0'
#959530000000
1!
b10 %
1'
b10 +
#959540000000
1"
1(
#959550000000
0!
0"
b100 &
0'
0(
b100 ,
#959560000000
1!
b11 %
1'
b11 +
#959570000000
0!
0'
#959580000000
1!
b100 %
1'
b100 +
#959590000000
0!
0'
#959600000000
1!
b101 %
1'
b101 +
#959610000000
0!
0'
#959620000000
1!
b110 %
1'
b110 +
#959630000000
0!
0'
#959640000000
1!
b111 %
1'
b111 +
#959650000000
0!
0'
#959660000000
1!
0$
b1000 %
1'
0*
b1000 +
#959670000000
0!
0'
#959680000000
1!
b1001 %
1'
b1001 +
#959690000000
0!
0'
#959700000000
1!
b0 %
1'
b0 +
#959710000000
0!
0'
#959720000000
1!
1$
b1 %
1'
1*
b1 +
#959730000000
0!
0'
#959740000000
1!
b10 %
1'
b10 +
#959750000000
0!
0'
#959760000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#959770000000
0!
0'
#959780000000
1!
b100 %
1'
b100 +
#959790000000
0!
0'
#959800000000
1!
b101 %
1'
b101 +
#959810000000
0!
0'
#959820000000
1!
0$
b110 %
1'
0*
b110 +
#959830000000
0!
0'
#959840000000
1!
b111 %
1'
b111 +
#959850000000
0!
0'
#959860000000
1!
b1000 %
1'
b1000 +
#959870000000
0!
0'
#959880000000
1!
b1001 %
1'
b1001 +
#959890000000
0!
0'
#959900000000
1!
b0 %
1'
b0 +
#959910000000
0!
0'
#959920000000
1!
1$
b1 %
1'
1*
b1 +
#959930000000
0!
0'
#959940000000
1!
b10 %
1'
b10 +
#959950000000
0!
0'
#959960000000
1!
b11 %
1'
b11 +
#959970000000
1"
1(
#959980000000
0!
0"
b100 &
0'
0(
b100 ,
#959990000000
1!
b100 %
1'
b100 +
#960000000000
0!
0'
#960010000000
1!
b101 %
1'
b101 +
#960020000000
0!
0'
#960030000000
1!
b110 %
1'
b110 +
#960040000000
0!
0'
#960050000000
1!
b111 %
1'
b111 +
#960060000000
0!
0'
#960070000000
1!
0$
b1000 %
1'
0*
b1000 +
#960080000000
0!
0'
#960090000000
1!
b1001 %
1'
b1001 +
#960100000000
0!
0'
#960110000000
1!
b0 %
1'
b0 +
#960120000000
0!
0'
#960130000000
1!
1$
b1 %
1'
1*
b1 +
#960140000000
0!
0'
#960150000000
1!
b10 %
1'
b10 +
#960160000000
0!
0'
#960170000000
1!
b11 %
1'
b11 +
#960180000000
0!
0'
#960190000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#960200000000
0!
0'
#960210000000
1!
b101 %
1'
b101 +
#960220000000
0!
0'
#960230000000
1!
0$
b110 %
1'
0*
b110 +
#960240000000
0!
0'
#960250000000
1!
b111 %
1'
b111 +
#960260000000
0!
0'
#960270000000
1!
b1000 %
1'
b1000 +
#960280000000
0!
0'
#960290000000
1!
b1001 %
1'
b1001 +
#960300000000
0!
0'
#960310000000
1!
b0 %
1'
b0 +
#960320000000
0!
0'
#960330000000
1!
1$
b1 %
1'
1*
b1 +
#960340000000
0!
0'
#960350000000
1!
b10 %
1'
b10 +
#960360000000
0!
0'
#960370000000
1!
b11 %
1'
b11 +
#960380000000
0!
0'
#960390000000
1!
b100 %
1'
b100 +
#960400000000
1"
1(
#960410000000
0!
0"
b100 &
0'
0(
b100 ,
#960420000000
1!
b101 %
1'
b101 +
#960430000000
0!
0'
#960440000000
1!
b110 %
1'
b110 +
#960450000000
0!
0'
#960460000000
1!
b111 %
1'
b111 +
#960470000000
0!
0'
#960480000000
1!
0$
b1000 %
1'
0*
b1000 +
#960490000000
0!
0'
#960500000000
1!
b1001 %
1'
b1001 +
#960510000000
0!
0'
#960520000000
1!
b0 %
1'
b0 +
#960530000000
0!
0'
#960540000000
1!
1$
b1 %
1'
1*
b1 +
#960550000000
0!
0'
#960560000000
1!
b10 %
1'
b10 +
#960570000000
0!
0'
#960580000000
1!
b11 %
1'
b11 +
#960590000000
0!
0'
#960600000000
1!
b100 %
1'
b100 +
#960610000000
0!
0'
#960620000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#960630000000
0!
0'
#960640000000
1!
0$
b110 %
1'
0*
b110 +
#960650000000
0!
0'
#960660000000
1!
b111 %
1'
b111 +
#960670000000
0!
0'
#960680000000
1!
b1000 %
1'
b1000 +
#960690000000
0!
0'
#960700000000
1!
b1001 %
1'
b1001 +
#960710000000
0!
0'
#960720000000
1!
b0 %
1'
b0 +
#960730000000
0!
0'
#960740000000
1!
1$
b1 %
1'
1*
b1 +
#960750000000
0!
0'
#960760000000
1!
b10 %
1'
b10 +
#960770000000
0!
0'
#960780000000
1!
b11 %
1'
b11 +
#960790000000
0!
0'
#960800000000
1!
b100 %
1'
b100 +
#960810000000
0!
0'
#960820000000
1!
b101 %
1'
b101 +
#960830000000
1"
1(
#960840000000
0!
0"
b100 &
0'
0(
b100 ,
#960850000000
1!
b110 %
1'
b110 +
#960860000000
0!
0'
#960870000000
1!
b111 %
1'
b111 +
#960880000000
0!
0'
#960890000000
1!
0$
b1000 %
1'
0*
b1000 +
#960900000000
0!
0'
#960910000000
1!
b1001 %
1'
b1001 +
#960920000000
0!
0'
#960930000000
1!
b0 %
1'
b0 +
#960940000000
0!
0'
#960950000000
1!
1$
b1 %
1'
1*
b1 +
#960960000000
0!
0'
#960970000000
1!
b10 %
1'
b10 +
#960980000000
0!
0'
#960990000000
1!
b11 %
1'
b11 +
#961000000000
0!
0'
#961010000000
1!
b100 %
1'
b100 +
#961020000000
0!
0'
#961030000000
1!
b101 %
1'
b101 +
#961040000000
0!
0'
#961050000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#961060000000
0!
0'
#961070000000
1!
b111 %
1'
b111 +
#961080000000
0!
0'
#961090000000
1!
b1000 %
1'
b1000 +
#961100000000
0!
0'
#961110000000
1!
b1001 %
1'
b1001 +
#961120000000
0!
0'
#961130000000
1!
b0 %
1'
b0 +
#961140000000
0!
0'
#961150000000
1!
1$
b1 %
1'
1*
b1 +
#961160000000
0!
0'
#961170000000
1!
b10 %
1'
b10 +
#961180000000
0!
0'
#961190000000
1!
b11 %
1'
b11 +
#961200000000
0!
0'
#961210000000
1!
b100 %
1'
b100 +
#961220000000
0!
0'
#961230000000
1!
b101 %
1'
b101 +
#961240000000
0!
0'
#961250000000
1!
0$
b110 %
1'
0*
b110 +
#961260000000
1"
1(
#961270000000
0!
0"
b100 &
0'
0(
b100 ,
#961280000000
1!
1$
b111 %
1'
1*
b111 +
#961290000000
0!
0'
#961300000000
1!
0$
b1000 %
1'
0*
b1000 +
#961310000000
0!
0'
#961320000000
1!
b1001 %
1'
b1001 +
#961330000000
0!
0'
#961340000000
1!
b0 %
1'
b0 +
#961350000000
0!
0'
#961360000000
1!
1$
b1 %
1'
1*
b1 +
#961370000000
0!
0'
#961380000000
1!
b10 %
1'
b10 +
#961390000000
0!
0'
#961400000000
1!
b11 %
1'
b11 +
#961410000000
0!
0'
#961420000000
1!
b100 %
1'
b100 +
#961430000000
0!
0'
#961440000000
1!
b101 %
1'
b101 +
#961450000000
0!
0'
#961460000000
1!
b110 %
1'
b110 +
#961470000000
0!
0'
#961480000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#961490000000
0!
0'
#961500000000
1!
b1000 %
1'
b1000 +
#961510000000
0!
0'
#961520000000
1!
b1001 %
1'
b1001 +
#961530000000
0!
0'
#961540000000
1!
b0 %
1'
b0 +
#961550000000
0!
0'
#961560000000
1!
1$
b1 %
1'
1*
b1 +
#961570000000
0!
0'
#961580000000
1!
b10 %
1'
b10 +
#961590000000
0!
0'
#961600000000
1!
b11 %
1'
b11 +
#961610000000
0!
0'
#961620000000
1!
b100 %
1'
b100 +
#961630000000
0!
0'
#961640000000
1!
b101 %
1'
b101 +
#961650000000
0!
0'
#961660000000
1!
0$
b110 %
1'
0*
b110 +
#961670000000
0!
0'
#961680000000
1!
b111 %
1'
b111 +
#961690000000
1"
1(
#961700000000
0!
0"
b100 &
0'
0(
b100 ,
#961710000000
1!
b1000 %
1'
b1000 +
#961720000000
0!
0'
#961730000000
1!
b1001 %
1'
b1001 +
#961740000000
0!
0'
#961750000000
1!
b0 %
1'
b0 +
#961760000000
0!
0'
#961770000000
1!
1$
b1 %
1'
1*
b1 +
#961780000000
0!
0'
#961790000000
1!
b10 %
1'
b10 +
#961800000000
0!
0'
#961810000000
1!
b11 %
1'
b11 +
#961820000000
0!
0'
#961830000000
1!
b100 %
1'
b100 +
#961840000000
0!
0'
#961850000000
1!
b101 %
1'
b101 +
#961860000000
0!
0'
#961870000000
1!
b110 %
1'
b110 +
#961880000000
0!
0'
#961890000000
1!
b111 %
1'
b111 +
#961900000000
0!
0'
#961910000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#961920000000
0!
0'
#961930000000
1!
b1001 %
1'
b1001 +
#961940000000
0!
0'
#961950000000
1!
b0 %
1'
b0 +
#961960000000
0!
0'
#961970000000
1!
1$
b1 %
1'
1*
b1 +
#961980000000
0!
0'
#961990000000
1!
b10 %
1'
b10 +
#962000000000
0!
0'
#962010000000
1!
b11 %
1'
b11 +
#962020000000
0!
0'
#962030000000
1!
b100 %
1'
b100 +
#962040000000
0!
0'
#962050000000
1!
b101 %
1'
b101 +
#962060000000
0!
0'
#962070000000
1!
0$
b110 %
1'
0*
b110 +
#962080000000
0!
0'
#962090000000
1!
b111 %
1'
b111 +
#962100000000
0!
0'
#962110000000
1!
b1000 %
1'
b1000 +
#962120000000
1"
1(
#962130000000
0!
0"
b100 &
0'
0(
b100 ,
#962140000000
1!
b1001 %
1'
b1001 +
#962150000000
0!
0'
#962160000000
1!
b0 %
1'
b0 +
#962170000000
0!
0'
#962180000000
1!
1$
b1 %
1'
1*
b1 +
#962190000000
0!
0'
#962200000000
1!
b10 %
1'
b10 +
#962210000000
0!
0'
#962220000000
1!
b11 %
1'
b11 +
#962230000000
0!
0'
#962240000000
1!
b100 %
1'
b100 +
#962250000000
0!
0'
#962260000000
1!
b101 %
1'
b101 +
#962270000000
0!
0'
#962280000000
1!
b110 %
1'
b110 +
#962290000000
0!
0'
#962300000000
1!
b111 %
1'
b111 +
#962310000000
0!
0'
#962320000000
1!
0$
b1000 %
1'
0*
b1000 +
#962330000000
0!
0'
#962340000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#962350000000
0!
0'
#962360000000
1!
b0 %
1'
b0 +
#962370000000
0!
0'
#962380000000
1!
1$
b1 %
1'
1*
b1 +
#962390000000
0!
0'
#962400000000
1!
b10 %
1'
b10 +
#962410000000
0!
0'
#962420000000
1!
b11 %
1'
b11 +
#962430000000
0!
0'
#962440000000
1!
b100 %
1'
b100 +
#962450000000
0!
0'
#962460000000
1!
b101 %
1'
b101 +
#962470000000
0!
0'
#962480000000
1!
0$
b110 %
1'
0*
b110 +
#962490000000
0!
0'
#962500000000
1!
b111 %
1'
b111 +
#962510000000
0!
0'
#962520000000
1!
b1000 %
1'
b1000 +
#962530000000
0!
0'
#962540000000
1!
b1001 %
1'
b1001 +
#962550000000
1"
1(
#962560000000
0!
0"
b100 &
0'
0(
b100 ,
#962570000000
1!
b0 %
1'
b0 +
#962580000000
0!
0'
#962590000000
1!
1$
b1 %
1'
1*
b1 +
#962600000000
0!
0'
#962610000000
1!
b10 %
1'
b10 +
#962620000000
0!
0'
#962630000000
1!
b11 %
1'
b11 +
#962640000000
0!
0'
#962650000000
1!
b100 %
1'
b100 +
#962660000000
0!
0'
#962670000000
1!
b101 %
1'
b101 +
#962680000000
0!
0'
#962690000000
1!
b110 %
1'
b110 +
#962700000000
0!
0'
#962710000000
1!
b111 %
1'
b111 +
#962720000000
0!
0'
#962730000000
1!
0$
b1000 %
1'
0*
b1000 +
#962740000000
0!
0'
#962750000000
1!
b1001 %
1'
b1001 +
#962760000000
0!
0'
#962770000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#962780000000
0!
0'
#962790000000
1!
1$
b1 %
1'
1*
b1 +
#962800000000
0!
0'
#962810000000
1!
b10 %
1'
b10 +
#962820000000
0!
0'
#962830000000
1!
b11 %
1'
b11 +
#962840000000
0!
0'
#962850000000
1!
b100 %
1'
b100 +
#962860000000
0!
0'
#962870000000
1!
b101 %
1'
b101 +
#962880000000
0!
0'
#962890000000
1!
0$
b110 %
1'
0*
b110 +
#962900000000
0!
0'
#962910000000
1!
b111 %
1'
b111 +
#962920000000
0!
0'
#962930000000
1!
b1000 %
1'
b1000 +
#962940000000
0!
0'
#962950000000
1!
b1001 %
1'
b1001 +
#962960000000
0!
0'
#962970000000
1!
b0 %
1'
b0 +
#962980000000
1"
1(
#962990000000
0!
0"
b100 &
0'
0(
b100 ,
#963000000000
1!
1$
b1 %
1'
1*
b1 +
#963010000000
0!
0'
#963020000000
1!
b10 %
1'
b10 +
#963030000000
0!
0'
#963040000000
1!
b11 %
1'
b11 +
#963050000000
0!
0'
#963060000000
1!
b100 %
1'
b100 +
#963070000000
0!
0'
#963080000000
1!
b101 %
1'
b101 +
#963090000000
0!
0'
#963100000000
1!
b110 %
1'
b110 +
#963110000000
0!
0'
#963120000000
1!
b111 %
1'
b111 +
#963130000000
0!
0'
#963140000000
1!
0$
b1000 %
1'
0*
b1000 +
#963150000000
0!
0'
#963160000000
1!
b1001 %
1'
b1001 +
#963170000000
0!
0'
#963180000000
1!
b0 %
1'
b0 +
#963190000000
0!
0'
#963200000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#963210000000
0!
0'
#963220000000
1!
b10 %
1'
b10 +
#963230000000
0!
0'
#963240000000
1!
b11 %
1'
b11 +
#963250000000
0!
0'
#963260000000
1!
b100 %
1'
b100 +
#963270000000
0!
0'
#963280000000
1!
b101 %
1'
b101 +
#963290000000
0!
0'
#963300000000
1!
0$
b110 %
1'
0*
b110 +
#963310000000
0!
0'
#963320000000
1!
b111 %
1'
b111 +
#963330000000
0!
0'
#963340000000
1!
b1000 %
1'
b1000 +
#963350000000
0!
0'
#963360000000
1!
b1001 %
1'
b1001 +
#963370000000
0!
0'
#963380000000
1!
b0 %
1'
b0 +
#963390000000
0!
0'
#963400000000
1!
1$
b1 %
1'
1*
b1 +
#963410000000
1"
1(
#963420000000
0!
0"
b100 &
0'
0(
b100 ,
#963430000000
1!
b10 %
1'
b10 +
#963440000000
0!
0'
#963450000000
1!
b11 %
1'
b11 +
#963460000000
0!
0'
#963470000000
1!
b100 %
1'
b100 +
#963480000000
0!
0'
#963490000000
1!
b101 %
1'
b101 +
#963500000000
0!
0'
#963510000000
1!
b110 %
1'
b110 +
#963520000000
0!
0'
#963530000000
1!
b111 %
1'
b111 +
#963540000000
0!
0'
#963550000000
1!
0$
b1000 %
1'
0*
b1000 +
#963560000000
0!
0'
#963570000000
1!
b1001 %
1'
b1001 +
#963580000000
0!
0'
#963590000000
1!
b0 %
1'
b0 +
#963600000000
0!
0'
#963610000000
1!
1$
b1 %
1'
1*
b1 +
#963620000000
0!
0'
#963630000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#963640000000
0!
0'
#963650000000
1!
b11 %
1'
b11 +
#963660000000
0!
0'
#963670000000
1!
b100 %
1'
b100 +
#963680000000
0!
0'
#963690000000
1!
b101 %
1'
b101 +
#963700000000
0!
0'
#963710000000
1!
0$
b110 %
1'
0*
b110 +
#963720000000
0!
0'
#963730000000
1!
b111 %
1'
b111 +
#963740000000
0!
0'
#963750000000
1!
b1000 %
1'
b1000 +
#963760000000
0!
0'
#963770000000
1!
b1001 %
1'
b1001 +
#963780000000
0!
0'
#963790000000
1!
b0 %
1'
b0 +
#963800000000
0!
0'
#963810000000
1!
1$
b1 %
1'
1*
b1 +
#963820000000
0!
0'
#963830000000
1!
b10 %
1'
b10 +
#963840000000
1"
1(
#963850000000
0!
0"
b100 &
0'
0(
b100 ,
#963860000000
1!
b11 %
1'
b11 +
#963870000000
0!
0'
#963880000000
1!
b100 %
1'
b100 +
#963890000000
0!
0'
#963900000000
1!
b101 %
1'
b101 +
#963910000000
0!
0'
#963920000000
1!
b110 %
1'
b110 +
#963930000000
0!
0'
#963940000000
1!
b111 %
1'
b111 +
#963950000000
0!
0'
#963960000000
1!
0$
b1000 %
1'
0*
b1000 +
#963970000000
0!
0'
#963980000000
1!
b1001 %
1'
b1001 +
#963990000000
0!
0'
#964000000000
1!
b0 %
1'
b0 +
#964010000000
0!
0'
#964020000000
1!
1$
b1 %
1'
1*
b1 +
#964030000000
0!
0'
#964040000000
1!
b10 %
1'
b10 +
#964050000000
0!
0'
#964060000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#964070000000
0!
0'
#964080000000
1!
b100 %
1'
b100 +
#964090000000
0!
0'
#964100000000
1!
b101 %
1'
b101 +
#964110000000
0!
0'
#964120000000
1!
0$
b110 %
1'
0*
b110 +
#964130000000
0!
0'
#964140000000
1!
b111 %
1'
b111 +
#964150000000
0!
0'
#964160000000
1!
b1000 %
1'
b1000 +
#964170000000
0!
0'
#964180000000
1!
b1001 %
1'
b1001 +
#964190000000
0!
0'
#964200000000
1!
b0 %
1'
b0 +
#964210000000
0!
0'
#964220000000
1!
1$
b1 %
1'
1*
b1 +
#964230000000
0!
0'
#964240000000
1!
b10 %
1'
b10 +
#964250000000
0!
0'
#964260000000
1!
b11 %
1'
b11 +
#964270000000
1"
1(
#964280000000
0!
0"
b100 &
0'
0(
b100 ,
#964290000000
1!
b100 %
1'
b100 +
#964300000000
0!
0'
#964310000000
1!
b101 %
1'
b101 +
#964320000000
0!
0'
#964330000000
1!
b110 %
1'
b110 +
#964340000000
0!
0'
#964350000000
1!
b111 %
1'
b111 +
#964360000000
0!
0'
#964370000000
1!
0$
b1000 %
1'
0*
b1000 +
#964380000000
0!
0'
#964390000000
1!
b1001 %
1'
b1001 +
#964400000000
0!
0'
#964410000000
1!
b0 %
1'
b0 +
#964420000000
0!
0'
#964430000000
1!
1$
b1 %
1'
1*
b1 +
#964440000000
0!
0'
#964450000000
1!
b10 %
1'
b10 +
#964460000000
0!
0'
#964470000000
1!
b11 %
1'
b11 +
#964480000000
0!
0'
#964490000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#964500000000
0!
0'
#964510000000
1!
b101 %
1'
b101 +
#964520000000
0!
0'
#964530000000
1!
0$
b110 %
1'
0*
b110 +
#964540000000
0!
0'
#964550000000
1!
b111 %
1'
b111 +
#964560000000
0!
0'
#964570000000
1!
b1000 %
1'
b1000 +
#964580000000
0!
0'
#964590000000
1!
b1001 %
1'
b1001 +
#964600000000
0!
0'
#964610000000
1!
b0 %
1'
b0 +
#964620000000
0!
0'
#964630000000
1!
1$
b1 %
1'
1*
b1 +
#964640000000
0!
0'
#964650000000
1!
b10 %
1'
b10 +
#964660000000
0!
0'
#964670000000
1!
b11 %
1'
b11 +
#964680000000
0!
0'
#964690000000
1!
b100 %
1'
b100 +
#964700000000
1"
1(
#964710000000
0!
0"
b100 &
0'
0(
b100 ,
#964720000000
1!
b101 %
1'
b101 +
#964730000000
0!
0'
#964740000000
1!
b110 %
1'
b110 +
#964750000000
0!
0'
#964760000000
1!
b111 %
1'
b111 +
#964770000000
0!
0'
#964780000000
1!
0$
b1000 %
1'
0*
b1000 +
#964790000000
0!
0'
#964800000000
1!
b1001 %
1'
b1001 +
#964810000000
0!
0'
#964820000000
1!
b0 %
1'
b0 +
#964830000000
0!
0'
#964840000000
1!
1$
b1 %
1'
1*
b1 +
#964850000000
0!
0'
#964860000000
1!
b10 %
1'
b10 +
#964870000000
0!
0'
#964880000000
1!
b11 %
1'
b11 +
#964890000000
0!
0'
#964900000000
1!
b100 %
1'
b100 +
#964910000000
0!
0'
#964920000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#964930000000
0!
0'
#964940000000
1!
0$
b110 %
1'
0*
b110 +
#964950000000
0!
0'
#964960000000
1!
b111 %
1'
b111 +
#964970000000
0!
0'
#964980000000
1!
b1000 %
1'
b1000 +
#964990000000
0!
0'
#965000000000
1!
b1001 %
1'
b1001 +
#965010000000
0!
0'
#965020000000
1!
b0 %
1'
b0 +
#965030000000
0!
0'
#965040000000
1!
1$
b1 %
1'
1*
b1 +
#965050000000
0!
0'
#965060000000
1!
b10 %
1'
b10 +
#965070000000
0!
0'
#965080000000
1!
b11 %
1'
b11 +
#965090000000
0!
0'
#965100000000
1!
b100 %
1'
b100 +
#965110000000
0!
0'
#965120000000
1!
b101 %
1'
b101 +
#965130000000
1"
1(
#965140000000
0!
0"
b100 &
0'
0(
b100 ,
#965150000000
1!
b110 %
1'
b110 +
#965160000000
0!
0'
#965170000000
1!
b111 %
1'
b111 +
#965180000000
0!
0'
#965190000000
1!
0$
b1000 %
1'
0*
b1000 +
#965200000000
0!
0'
#965210000000
1!
b1001 %
1'
b1001 +
#965220000000
0!
0'
#965230000000
1!
b0 %
1'
b0 +
#965240000000
0!
0'
#965250000000
1!
1$
b1 %
1'
1*
b1 +
#965260000000
0!
0'
#965270000000
1!
b10 %
1'
b10 +
#965280000000
0!
0'
#965290000000
1!
b11 %
1'
b11 +
#965300000000
0!
0'
#965310000000
1!
b100 %
1'
b100 +
#965320000000
0!
0'
#965330000000
1!
b101 %
1'
b101 +
#965340000000
0!
0'
#965350000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#965360000000
0!
0'
#965370000000
1!
b111 %
1'
b111 +
#965380000000
0!
0'
#965390000000
1!
b1000 %
1'
b1000 +
#965400000000
0!
0'
#965410000000
1!
b1001 %
1'
b1001 +
#965420000000
0!
0'
#965430000000
1!
b0 %
1'
b0 +
#965440000000
0!
0'
#965450000000
1!
1$
b1 %
1'
1*
b1 +
#965460000000
0!
0'
#965470000000
1!
b10 %
1'
b10 +
#965480000000
0!
0'
#965490000000
1!
b11 %
1'
b11 +
#965500000000
0!
0'
#965510000000
1!
b100 %
1'
b100 +
#965520000000
0!
0'
#965530000000
1!
b101 %
1'
b101 +
#965540000000
0!
0'
#965550000000
1!
0$
b110 %
1'
0*
b110 +
#965560000000
1"
1(
#965570000000
0!
0"
b100 &
0'
0(
b100 ,
#965580000000
1!
1$
b111 %
1'
1*
b111 +
#965590000000
0!
0'
#965600000000
1!
0$
b1000 %
1'
0*
b1000 +
#965610000000
0!
0'
#965620000000
1!
b1001 %
1'
b1001 +
#965630000000
0!
0'
#965640000000
1!
b0 %
1'
b0 +
#965650000000
0!
0'
#965660000000
1!
1$
b1 %
1'
1*
b1 +
#965670000000
0!
0'
#965680000000
1!
b10 %
1'
b10 +
#965690000000
0!
0'
#965700000000
1!
b11 %
1'
b11 +
#965710000000
0!
0'
#965720000000
1!
b100 %
1'
b100 +
#965730000000
0!
0'
#965740000000
1!
b101 %
1'
b101 +
#965750000000
0!
0'
#965760000000
1!
b110 %
1'
b110 +
#965770000000
0!
0'
#965780000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#965790000000
0!
0'
#965800000000
1!
b1000 %
1'
b1000 +
#965810000000
0!
0'
#965820000000
1!
b1001 %
1'
b1001 +
#965830000000
0!
0'
#965840000000
1!
b0 %
1'
b0 +
#965850000000
0!
0'
#965860000000
1!
1$
b1 %
1'
1*
b1 +
#965870000000
0!
0'
#965880000000
1!
b10 %
1'
b10 +
#965890000000
0!
0'
#965900000000
1!
b11 %
1'
b11 +
#965910000000
0!
0'
#965920000000
1!
b100 %
1'
b100 +
#965930000000
0!
0'
#965940000000
1!
b101 %
1'
b101 +
#965950000000
0!
0'
#965960000000
1!
0$
b110 %
1'
0*
b110 +
#965970000000
0!
0'
#965980000000
1!
b111 %
1'
b111 +
#965990000000
1"
1(
#966000000000
0!
0"
b100 &
0'
0(
b100 ,
#966010000000
1!
b1000 %
1'
b1000 +
#966020000000
0!
0'
#966030000000
1!
b1001 %
1'
b1001 +
#966040000000
0!
0'
#966050000000
1!
b0 %
1'
b0 +
#966060000000
0!
0'
#966070000000
1!
1$
b1 %
1'
1*
b1 +
#966080000000
0!
0'
#966090000000
1!
b10 %
1'
b10 +
#966100000000
0!
0'
#966110000000
1!
b11 %
1'
b11 +
#966120000000
0!
0'
#966130000000
1!
b100 %
1'
b100 +
#966140000000
0!
0'
#966150000000
1!
b101 %
1'
b101 +
#966160000000
0!
0'
#966170000000
1!
b110 %
1'
b110 +
#966180000000
0!
0'
#966190000000
1!
b111 %
1'
b111 +
#966200000000
0!
0'
#966210000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#966220000000
0!
0'
#966230000000
1!
b1001 %
1'
b1001 +
#966240000000
0!
0'
#966250000000
1!
b0 %
1'
b0 +
#966260000000
0!
0'
#966270000000
1!
1$
b1 %
1'
1*
b1 +
#966280000000
0!
0'
#966290000000
1!
b10 %
1'
b10 +
#966300000000
0!
0'
#966310000000
1!
b11 %
1'
b11 +
#966320000000
0!
0'
#966330000000
1!
b100 %
1'
b100 +
#966340000000
0!
0'
#966350000000
1!
b101 %
1'
b101 +
#966360000000
0!
0'
#966370000000
1!
0$
b110 %
1'
0*
b110 +
#966380000000
0!
0'
#966390000000
1!
b111 %
1'
b111 +
#966400000000
0!
0'
#966410000000
1!
b1000 %
1'
b1000 +
#966420000000
1"
1(
#966430000000
0!
0"
b100 &
0'
0(
b100 ,
#966440000000
1!
b1001 %
1'
b1001 +
#966450000000
0!
0'
#966460000000
1!
b0 %
1'
b0 +
#966470000000
0!
0'
#966480000000
1!
1$
b1 %
1'
1*
b1 +
#966490000000
0!
0'
#966500000000
1!
b10 %
1'
b10 +
#966510000000
0!
0'
#966520000000
1!
b11 %
1'
b11 +
#966530000000
0!
0'
#966540000000
1!
b100 %
1'
b100 +
#966550000000
0!
0'
#966560000000
1!
b101 %
1'
b101 +
#966570000000
0!
0'
#966580000000
1!
b110 %
1'
b110 +
#966590000000
0!
0'
#966600000000
1!
b111 %
1'
b111 +
#966610000000
0!
0'
#966620000000
1!
0$
b1000 %
1'
0*
b1000 +
#966630000000
0!
0'
#966640000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#966650000000
0!
0'
#966660000000
1!
b0 %
1'
b0 +
#966670000000
0!
0'
#966680000000
1!
1$
b1 %
1'
1*
b1 +
#966690000000
0!
0'
#966700000000
1!
b10 %
1'
b10 +
#966710000000
0!
0'
#966720000000
1!
b11 %
1'
b11 +
#966730000000
0!
0'
#966740000000
1!
b100 %
1'
b100 +
#966750000000
0!
0'
#966760000000
1!
b101 %
1'
b101 +
#966770000000
0!
0'
#966780000000
1!
0$
b110 %
1'
0*
b110 +
#966790000000
0!
0'
#966800000000
1!
b111 %
1'
b111 +
#966810000000
0!
0'
#966820000000
1!
b1000 %
1'
b1000 +
#966830000000
0!
0'
#966840000000
1!
b1001 %
1'
b1001 +
#966850000000
1"
1(
#966860000000
0!
0"
b100 &
0'
0(
b100 ,
#966870000000
1!
b0 %
1'
b0 +
#966880000000
0!
0'
#966890000000
1!
1$
b1 %
1'
1*
b1 +
#966900000000
0!
0'
#966910000000
1!
b10 %
1'
b10 +
#966920000000
0!
0'
#966930000000
1!
b11 %
1'
b11 +
#966940000000
0!
0'
#966950000000
1!
b100 %
1'
b100 +
#966960000000
0!
0'
#966970000000
1!
b101 %
1'
b101 +
#966980000000
0!
0'
#966990000000
1!
b110 %
1'
b110 +
#967000000000
0!
0'
#967010000000
1!
b111 %
1'
b111 +
#967020000000
0!
0'
#967030000000
1!
0$
b1000 %
1'
0*
b1000 +
#967040000000
0!
0'
#967050000000
1!
b1001 %
1'
b1001 +
#967060000000
0!
0'
#967070000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#967080000000
0!
0'
#967090000000
1!
1$
b1 %
1'
1*
b1 +
#967100000000
0!
0'
#967110000000
1!
b10 %
1'
b10 +
#967120000000
0!
0'
#967130000000
1!
b11 %
1'
b11 +
#967140000000
0!
0'
#967150000000
1!
b100 %
1'
b100 +
#967160000000
0!
0'
#967170000000
1!
b101 %
1'
b101 +
#967180000000
0!
0'
#967190000000
1!
0$
b110 %
1'
0*
b110 +
#967200000000
0!
0'
#967210000000
1!
b111 %
1'
b111 +
#967220000000
0!
0'
#967230000000
1!
b1000 %
1'
b1000 +
#967240000000
0!
0'
#967250000000
1!
b1001 %
1'
b1001 +
#967260000000
0!
0'
#967270000000
1!
b0 %
1'
b0 +
#967280000000
1"
1(
#967290000000
0!
0"
b100 &
0'
0(
b100 ,
#967300000000
1!
1$
b1 %
1'
1*
b1 +
#967310000000
0!
0'
#967320000000
1!
b10 %
1'
b10 +
#967330000000
0!
0'
#967340000000
1!
b11 %
1'
b11 +
#967350000000
0!
0'
#967360000000
1!
b100 %
1'
b100 +
#967370000000
0!
0'
#967380000000
1!
b101 %
1'
b101 +
#967390000000
0!
0'
#967400000000
1!
b110 %
1'
b110 +
#967410000000
0!
0'
#967420000000
1!
b111 %
1'
b111 +
#967430000000
0!
0'
#967440000000
1!
0$
b1000 %
1'
0*
b1000 +
#967450000000
0!
0'
#967460000000
1!
b1001 %
1'
b1001 +
#967470000000
0!
0'
#967480000000
1!
b0 %
1'
b0 +
#967490000000
0!
0'
#967500000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#967510000000
0!
0'
#967520000000
1!
b10 %
1'
b10 +
#967530000000
0!
0'
#967540000000
1!
b11 %
1'
b11 +
#967550000000
0!
0'
#967560000000
1!
b100 %
1'
b100 +
#967570000000
0!
0'
#967580000000
1!
b101 %
1'
b101 +
#967590000000
0!
0'
#967600000000
1!
0$
b110 %
1'
0*
b110 +
#967610000000
0!
0'
#967620000000
1!
b111 %
1'
b111 +
#967630000000
0!
0'
#967640000000
1!
b1000 %
1'
b1000 +
#967650000000
0!
0'
#967660000000
1!
b1001 %
1'
b1001 +
#967670000000
0!
0'
#967680000000
1!
b0 %
1'
b0 +
#967690000000
0!
0'
#967700000000
1!
1$
b1 %
1'
1*
b1 +
#967710000000
1"
1(
#967720000000
0!
0"
b100 &
0'
0(
b100 ,
#967730000000
1!
b10 %
1'
b10 +
#967740000000
0!
0'
#967750000000
1!
b11 %
1'
b11 +
#967760000000
0!
0'
#967770000000
1!
b100 %
1'
b100 +
#967780000000
0!
0'
#967790000000
1!
b101 %
1'
b101 +
#967800000000
0!
0'
#967810000000
1!
b110 %
1'
b110 +
#967820000000
0!
0'
#967830000000
1!
b111 %
1'
b111 +
#967840000000
0!
0'
#967850000000
1!
0$
b1000 %
1'
0*
b1000 +
#967860000000
0!
0'
#967870000000
1!
b1001 %
1'
b1001 +
#967880000000
0!
0'
#967890000000
1!
b0 %
1'
b0 +
#967900000000
0!
0'
#967910000000
1!
1$
b1 %
1'
1*
b1 +
#967920000000
0!
0'
#967930000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#967940000000
0!
0'
#967950000000
1!
b11 %
1'
b11 +
#967960000000
0!
0'
#967970000000
1!
b100 %
1'
b100 +
#967980000000
0!
0'
#967990000000
1!
b101 %
1'
b101 +
#968000000000
0!
0'
#968010000000
1!
0$
b110 %
1'
0*
b110 +
#968020000000
0!
0'
#968030000000
1!
b111 %
1'
b111 +
#968040000000
0!
0'
#968050000000
1!
b1000 %
1'
b1000 +
#968060000000
0!
0'
#968070000000
1!
b1001 %
1'
b1001 +
#968080000000
0!
0'
#968090000000
1!
b0 %
1'
b0 +
#968100000000
0!
0'
#968110000000
1!
1$
b1 %
1'
1*
b1 +
#968120000000
0!
0'
#968130000000
1!
b10 %
1'
b10 +
#968140000000
1"
1(
#968150000000
0!
0"
b100 &
0'
0(
b100 ,
#968160000000
1!
b11 %
1'
b11 +
#968170000000
0!
0'
#968180000000
1!
b100 %
1'
b100 +
#968190000000
0!
0'
#968200000000
1!
b101 %
1'
b101 +
#968210000000
0!
0'
#968220000000
1!
b110 %
1'
b110 +
#968230000000
0!
0'
#968240000000
1!
b111 %
1'
b111 +
#968250000000
0!
0'
#968260000000
1!
0$
b1000 %
1'
0*
b1000 +
#968270000000
0!
0'
#968280000000
1!
b1001 %
1'
b1001 +
#968290000000
0!
0'
#968300000000
1!
b0 %
1'
b0 +
#968310000000
0!
0'
#968320000000
1!
1$
b1 %
1'
1*
b1 +
#968330000000
0!
0'
#968340000000
1!
b10 %
1'
b10 +
#968350000000
0!
0'
#968360000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#968370000000
0!
0'
#968380000000
1!
b100 %
1'
b100 +
#968390000000
0!
0'
#968400000000
1!
b101 %
1'
b101 +
#968410000000
0!
0'
#968420000000
1!
0$
b110 %
1'
0*
b110 +
#968430000000
0!
0'
#968440000000
1!
b111 %
1'
b111 +
#968450000000
0!
0'
#968460000000
1!
b1000 %
1'
b1000 +
#968470000000
0!
0'
#968480000000
1!
b1001 %
1'
b1001 +
#968490000000
0!
0'
#968500000000
1!
b0 %
1'
b0 +
#968510000000
0!
0'
#968520000000
1!
1$
b1 %
1'
1*
b1 +
#968530000000
0!
0'
#968540000000
1!
b10 %
1'
b10 +
#968550000000
0!
0'
#968560000000
1!
b11 %
1'
b11 +
#968570000000
1"
1(
#968580000000
0!
0"
b100 &
0'
0(
b100 ,
#968590000000
1!
b100 %
1'
b100 +
#968600000000
0!
0'
#968610000000
1!
b101 %
1'
b101 +
#968620000000
0!
0'
#968630000000
1!
b110 %
1'
b110 +
#968640000000
0!
0'
#968650000000
1!
b111 %
1'
b111 +
#968660000000
0!
0'
#968670000000
1!
0$
b1000 %
1'
0*
b1000 +
#968680000000
0!
0'
#968690000000
1!
b1001 %
1'
b1001 +
#968700000000
0!
0'
#968710000000
1!
b0 %
1'
b0 +
#968720000000
0!
0'
#968730000000
1!
1$
b1 %
1'
1*
b1 +
#968740000000
0!
0'
#968750000000
1!
b10 %
1'
b10 +
#968760000000
0!
0'
#968770000000
1!
b11 %
1'
b11 +
#968780000000
0!
0'
#968790000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#968800000000
0!
0'
#968810000000
1!
b101 %
1'
b101 +
#968820000000
0!
0'
#968830000000
1!
0$
b110 %
1'
0*
b110 +
#968840000000
0!
0'
#968850000000
1!
b111 %
1'
b111 +
#968860000000
0!
0'
#968870000000
1!
b1000 %
1'
b1000 +
#968880000000
0!
0'
#968890000000
1!
b1001 %
1'
b1001 +
#968900000000
0!
0'
#968910000000
1!
b0 %
1'
b0 +
#968920000000
0!
0'
#968930000000
1!
1$
b1 %
1'
1*
b1 +
#968940000000
0!
0'
#968950000000
1!
b10 %
1'
b10 +
#968960000000
0!
0'
#968970000000
1!
b11 %
1'
b11 +
#968980000000
0!
0'
#968990000000
1!
b100 %
1'
b100 +
#969000000000
1"
1(
#969010000000
0!
0"
b100 &
0'
0(
b100 ,
#969020000000
1!
b101 %
1'
b101 +
#969030000000
0!
0'
#969040000000
1!
b110 %
1'
b110 +
#969050000000
0!
0'
#969060000000
1!
b111 %
1'
b111 +
#969070000000
0!
0'
#969080000000
1!
0$
b1000 %
1'
0*
b1000 +
#969090000000
0!
0'
#969100000000
1!
b1001 %
1'
b1001 +
#969110000000
0!
0'
#969120000000
1!
b0 %
1'
b0 +
#969130000000
0!
0'
#969140000000
1!
1$
b1 %
1'
1*
b1 +
#969150000000
0!
0'
#969160000000
1!
b10 %
1'
b10 +
#969170000000
0!
0'
#969180000000
1!
b11 %
1'
b11 +
#969190000000
0!
0'
#969200000000
1!
b100 %
1'
b100 +
#969210000000
0!
0'
#969220000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#969230000000
0!
0'
#969240000000
1!
0$
b110 %
1'
0*
b110 +
#969250000000
0!
0'
#969260000000
1!
b111 %
1'
b111 +
#969270000000
0!
0'
#969280000000
1!
b1000 %
1'
b1000 +
#969290000000
0!
0'
#969300000000
1!
b1001 %
1'
b1001 +
#969310000000
0!
0'
#969320000000
1!
b0 %
1'
b0 +
#969330000000
0!
0'
#969340000000
1!
1$
b1 %
1'
1*
b1 +
#969350000000
0!
0'
#969360000000
1!
b10 %
1'
b10 +
#969370000000
0!
0'
#969380000000
1!
b11 %
1'
b11 +
#969390000000
0!
0'
#969400000000
1!
b100 %
1'
b100 +
#969410000000
0!
0'
#969420000000
1!
b101 %
1'
b101 +
#969430000000
1"
1(
#969440000000
0!
0"
b100 &
0'
0(
b100 ,
#969450000000
1!
b110 %
1'
b110 +
#969460000000
0!
0'
#969470000000
1!
b111 %
1'
b111 +
#969480000000
0!
0'
#969490000000
1!
0$
b1000 %
1'
0*
b1000 +
#969500000000
0!
0'
#969510000000
1!
b1001 %
1'
b1001 +
#969520000000
0!
0'
#969530000000
1!
b0 %
1'
b0 +
#969540000000
0!
0'
#969550000000
1!
1$
b1 %
1'
1*
b1 +
#969560000000
0!
0'
#969570000000
1!
b10 %
1'
b10 +
#969580000000
0!
0'
#969590000000
1!
b11 %
1'
b11 +
#969600000000
0!
0'
#969610000000
1!
b100 %
1'
b100 +
#969620000000
0!
0'
#969630000000
1!
b101 %
1'
b101 +
#969640000000
0!
0'
#969650000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#969660000000
0!
0'
#969670000000
1!
b111 %
1'
b111 +
#969680000000
0!
0'
#969690000000
1!
b1000 %
1'
b1000 +
#969700000000
0!
0'
#969710000000
1!
b1001 %
1'
b1001 +
#969720000000
0!
0'
#969730000000
1!
b0 %
1'
b0 +
#969740000000
0!
0'
#969750000000
1!
1$
b1 %
1'
1*
b1 +
#969760000000
0!
0'
#969770000000
1!
b10 %
1'
b10 +
#969780000000
0!
0'
#969790000000
1!
b11 %
1'
b11 +
#969800000000
0!
0'
#969810000000
1!
b100 %
1'
b100 +
#969820000000
0!
0'
#969830000000
1!
b101 %
1'
b101 +
#969840000000
0!
0'
#969850000000
1!
0$
b110 %
1'
0*
b110 +
#969860000000
1"
1(
#969870000000
0!
0"
b100 &
0'
0(
b100 ,
#969880000000
1!
1$
b111 %
1'
1*
b111 +
#969890000000
0!
0'
#969900000000
1!
0$
b1000 %
1'
0*
b1000 +
#969910000000
0!
0'
#969920000000
1!
b1001 %
1'
b1001 +
#969930000000
0!
0'
#969940000000
1!
b0 %
1'
b0 +
#969950000000
0!
0'
#969960000000
1!
1$
b1 %
1'
1*
b1 +
#969970000000
0!
0'
#969980000000
1!
b10 %
1'
b10 +
#969990000000
0!
0'
#970000000000
1!
b11 %
1'
b11 +
#970010000000
0!
0'
#970020000000
1!
b100 %
1'
b100 +
#970030000000
0!
0'
#970040000000
1!
b101 %
1'
b101 +
#970050000000
0!
0'
#970060000000
1!
b110 %
1'
b110 +
#970070000000
0!
0'
#970080000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#970090000000
0!
0'
#970100000000
1!
b1000 %
1'
b1000 +
#970110000000
0!
0'
#970120000000
1!
b1001 %
1'
b1001 +
#970130000000
0!
0'
#970140000000
1!
b0 %
1'
b0 +
#970150000000
0!
0'
#970160000000
1!
1$
b1 %
1'
1*
b1 +
#970170000000
0!
0'
#970180000000
1!
b10 %
1'
b10 +
#970190000000
0!
0'
#970200000000
1!
b11 %
1'
b11 +
#970210000000
0!
0'
#970220000000
1!
b100 %
1'
b100 +
#970230000000
0!
0'
#970240000000
1!
b101 %
1'
b101 +
#970250000000
0!
0'
#970260000000
1!
0$
b110 %
1'
0*
b110 +
#970270000000
0!
0'
#970280000000
1!
b111 %
1'
b111 +
#970290000000
1"
1(
#970300000000
0!
0"
b100 &
0'
0(
b100 ,
#970310000000
1!
b1000 %
1'
b1000 +
#970320000000
0!
0'
#970330000000
1!
b1001 %
1'
b1001 +
#970340000000
0!
0'
#970350000000
1!
b0 %
1'
b0 +
#970360000000
0!
0'
#970370000000
1!
1$
b1 %
1'
1*
b1 +
#970380000000
0!
0'
#970390000000
1!
b10 %
1'
b10 +
#970400000000
0!
0'
#970410000000
1!
b11 %
1'
b11 +
#970420000000
0!
0'
#970430000000
1!
b100 %
1'
b100 +
#970440000000
0!
0'
#970450000000
1!
b101 %
1'
b101 +
#970460000000
0!
0'
#970470000000
1!
b110 %
1'
b110 +
#970480000000
0!
0'
#970490000000
1!
b111 %
1'
b111 +
#970500000000
0!
0'
#970510000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#970520000000
0!
0'
#970530000000
1!
b1001 %
1'
b1001 +
#970540000000
0!
0'
#970550000000
1!
b0 %
1'
b0 +
#970560000000
0!
0'
#970570000000
1!
1$
b1 %
1'
1*
b1 +
#970580000000
0!
0'
#970590000000
1!
b10 %
1'
b10 +
#970600000000
0!
0'
#970610000000
1!
b11 %
1'
b11 +
#970620000000
0!
0'
#970630000000
1!
b100 %
1'
b100 +
#970640000000
0!
0'
#970650000000
1!
b101 %
1'
b101 +
#970660000000
0!
0'
#970670000000
1!
0$
b110 %
1'
0*
b110 +
#970680000000
0!
0'
#970690000000
1!
b111 %
1'
b111 +
#970700000000
0!
0'
#970710000000
1!
b1000 %
1'
b1000 +
#970720000000
1"
1(
#970730000000
0!
0"
b100 &
0'
0(
b100 ,
#970740000000
1!
b1001 %
1'
b1001 +
#970750000000
0!
0'
#970760000000
1!
b0 %
1'
b0 +
#970770000000
0!
0'
#970780000000
1!
1$
b1 %
1'
1*
b1 +
#970790000000
0!
0'
#970800000000
1!
b10 %
1'
b10 +
#970810000000
0!
0'
#970820000000
1!
b11 %
1'
b11 +
#970830000000
0!
0'
#970840000000
1!
b100 %
1'
b100 +
#970850000000
0!
0'
#970860000000
1!
b101 %
1'
b101 +
#970870000000
0!
0'
#970880000000
1!
b110 %
1'
b110 +
#970890000000
0!
0'
#970900000000
1!
b111 %
1'
b111 +
#970910000000
0!
0'
#970920000000
1!
0$
b1000 %
1'
0*
b1000 +
#970930000000
0!
0'
#970940000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#970950000000
0!
0'
#970960000000
1!
b0 %
1'
b0 +
#970970000000
0!
0'
#970980000000
1!
1$
b1 %
1'
1*
b1 +
#970990000000
0!
0'
#971000000000
1!
b10 %
1'
b10 +
#971010000000
0!
0'
#971020000000
1!
b11 %
1'
b11 +
#971030000000
0!
0'
#971040000000
1!
b100 %
1'
b100 +
#971050000000
0!
0'
#971060000000
1!
b101 %
1'
b101 +
#971070000000
0!
0'
#971080000000
1!
0$
b110 %
1'
0*
b110 +
#971090000000
0!
0'
#971100000000
1!
b111 %
1'
b111 +
#971110000000
0!
0'
#971120000000
1!
b1000 %
1'
b1000 +
#971130000000
0!
0'
#971140000000
1!
b1001 %
1'
b1001 +
#971150000000
1"
1(
#971160000000
0!
0"
b100 &
0'
0(
b100 ,
#971170000000
1!
b0 %
1'
b0 +
#971180000000
0!
0'
#971190000000
1!
1$
b1 %
1'
1*
b1 +
#971200000000
0!
0'
#971210000000
1!
b10 %
1'
b10 +
#971220000000
0!
0'
#971230000000
1!
b11 %
1'
b11 +
#971240000000
0!
0'
#971250000000
1!
b100 %
1'
b100 +
#971260000000
0!
0'
#971270000000
1!
b101 %
1'
b101 +
#971280000000
0!
0'
#971290000000
1!
b110 %
1'
b110 +
#971300000000
0!
0'
#971310000000
1!
b111 %
1'
b111 +
#971320000000
0!
0'
#971330000000
1!
0$
b1000 %
1'
0*
b1000 +
#971340000000
0!
0'
#971350000000
1!
b1001 %
1'
b1001 +
#971360000000
0!
0'
#971370000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#971380000000
0!
0'
#971390000000
1!
1$
b1 %
1'
1*
b1 +
#971400000000
0!
0'
#971410000000
1!
b10 %
1'
b10 +
#971420000000
0!
0'
#971430000000
1!
b11 %
1'
b11 +
#971440000000
0!
0'
#971450000000
1!
b100 %
1'
b100 +
#971460000000
0!
0'
#971470000000
1!
b101 %
1'
b101 +
#971480000000
0!
0'
#971490000000
1!
0$
b110 %
1'
0*
b110 +
#971500000000
0!
0'
#971510000000
1!
b111 %
1'
b111 +
#971520000000
0!
0'
#971530000000
1!
b1000 %
1'
b1000 +
#971540000000
0!
0'
#971550000000
1!
b1001 %
1'
b1001 +
#971560000000
0!
0'
#971570000000
1!
b0 %
1'
b0 +
#971580000000
1"
1(
#971590000000
0!
0"
b100 &
0'
0(
b100 ,
#971600000000
1!
1$
b1 %
1'
1*
b1 +
#971610000000
0!
0'
#971620000000
1!
b10 %
1'
b10 +
#971630000000
0!
0'
#971640000000
1!
b11 %
1'
b11 +
#971650000000
0!
0'
#971660000000
1!
b100 %
1'
b100 +
#971670000000
0!
0'
#971680000000
1!
b101 %
1'
b101 +
#971690000000
0!
0'
#971700000000
1!
b110 %
1'
b110 +
#971710000000
0!
0'
#971720000000
1!
b111 %
1'
b111 +
#971730000000
0!
0'
#971740000000
1!
0$
b1000 %
1'
0*
b1000 +
#971750000000
0!
0'
#971760000000
1!
b1001 %
1'
b1001 +
#971770000000
0!
0'
#971780000000
1!
b0 %
1'
b0 +
#971790000000
0!
0'
#971800000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#971810000000
0!
0'
#971820000000
1!
b10 %
1'
b10 +
#971830000000
0!
0'
#971840000000
1!
b11 %
1'
b11 +
#971850000000
0!
0'
#971860000000
1!
b100 %
1'
b100 +
#971870000000
0!
0'
#971880000000
1!
b101 %
1'
b101 +
#971890000000
0!
0'
#971900000000
1!
0$
b110 %
1'
0*
b110 +
#971910000000
0!
0'
#971920000000
1!
b111 %
1'
b111 +
#971930000000
0!
0'
#971940000000
1!
b1000 %
1'
b1000 +
#971950000000
0!
0'
#971960000000
1!
b1001 %
1'
b1001 +
#971970000000
0!
0'
#971980000000
1!
b0 %
1'
b0 +
#971990000000
0!
0'
#972000000000
1!
1$
b1 %
1'
1*
b1 +
#972010000000
1"
1(
#972020000000
0!
0"
b100 &
0'
0(
b100 ,
#972030000000
1!
b10 %
1'
b10 +
#972040000000
0!
0'
#972050000000
1!
b11 %
1'
b11 +
#972060000000
0!
0'
#972070000000
1!
b100 %
1'
b100 +
#972080000000
0!
0'
#972090000000
1!
b101 %
1'
b101 +
#972100000000
0!
0'
#972110000000
1!
b110 %
1'
b110 +
#972120000000
0!
0'
#972130000000
1!
b111 %
1'
b111 +
#972140000000
0!
0'
#972150000000
1!
0$
b1000 %
1'
0*
b1000 +
#972160000000
0!
0'
#972170000000
1!
b1001 %
1'
b1001 +
#972180000000
0!
0'
#972190000000
1!
b0 %
1'
b0 +
#972200000000
0!
0'
#972210000000
1!
1$
b1 %
1'
1*
b1 +
#972220000000
0!
0'
#972230000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#972240000000
0!
0'
#972250000000
1!
b11 %
1'
b11 +
#972260000000
0!
0'
#972270000000
1!
b100 %
1'
b100 +
#972280000000
0!
0'
#972290000000
1!
b101 %
1'
b101 +
#972300000000
0!
0'
#972310000000
1!
0$
b110 %
1'
0*
b110 +
#972320000000
0!
0'
#972330000000
1!
b111 %
1'
b111 +
#972340000000
0!
0'
#972350000000
1!
b1000 %
1'
b1000 +
#972360000000
0!
0'
#972370000000
1!
b1001 %
1'
b1001 +
#972380000000
0!
0'
#972390000000
1!
b0 %
1'
b0 +
#972400000000
0!
0'
#972410000000
1!
1$
b1 %
1'
1*
b1 +
#972420000000
0!
0'
#972430000000
1!
b10 %
1'
b10 +
#972440000000
1"
1(
#972450000000
0!
0"
b100 &
0'
0(
b100 ,
#972460000000
1!
b11 %
1'
b11 +
#972470000000
0!
0'
#972480000000
1!
b100 %
1'
b100 +
#972490000000
0!
0'
#972500000000
1!
b101 %
1'
b101 +
#972510000000
0!
0'
#972520000000
1!
b110 %
1'
b110 +
#972530000000
0!
0'
#972540000000
1!
b111 %
1'
b111 +
#972550000000
0!
0'
#972560000000
1!
0$
b1000 %
1'
0*
b1000 +
#972570000000
0!
0'
#972580000000
1!
b1001 %
1'
b1001 +
#972590000000
0!
0'
#972600000000
1!
b0 %
1'
b0 +
#972610000000
0!
0'
#972620000000
1!
1$
b1 %
1'
1*
b1 +
#972630000000
0!
0'
#972640000000
1!
b10 %
1'
b10 +
#972650000000
0!
0'
#972660000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#972670000000
0!
0'
#972680000000
1!
b100 %
1'
b100 +
#972690000000
0!
0'
#972700000000
1!
b101 %
1'
b101 +
#972710000000
0!
0'
#972720000000
1!
0$
b110 %
1'
0*
b110 +
#972730000000
0!
0'
#972740000000
1!
b111 %
1'
b111 +
#972750000000
0!
0'
#972760000000
1!
b1000 %
1'
b1000 +
#972770000000
0!
0'
#972780000000
1!
b1001 %
1'
b1001 +
#972790000000
0!
0'
#972800000000
1!
b0 %
1'
b0 +
#972810000000
0!
0'
#972820000000
1!
1$
b1 %
1'
1*
b1 +
#972830000000
0!
0'
#972840000000
1!
b10 %
1'
b10 +
#972850000000
0!
0'
#972860000000
1!
b11 %
1'
b11 +
#972870000000
1"
1(
#972880000000
0!
0"
b100 &
0'
0(
b100 ,
#972890000000
1!
b100 %
1'
b100 +
#972900000000
0!
0'
#972910000000
1!
b101 %
1'
b101 +
#972920000000
0!
0'
#972930000000
1!
b110 %
1'
b110 +
#972940000000
0!
0'
#972950000000
1!
b111 %
1'
b111 +
#972960000000
0!
0'
#972970000000
1!
0$
b1000 %
1'
0*
b1000 +
#972980000000
0!
0'
#972990000000
1!
b1001 %
1'
b1001 +
#973000000000
0!
0'
#973010000000
1!
b0 %
1'
b0 +
#973020000000
0!
0'
#973030000000
1!
1$
b1 %
1'
1*
b1 +
#973040000000
0!
0'
#973050000000
1!
b10 %
1'
b10 +
#973060000000
0!
0'
#973070000000
1!
b11 %
1'
b11 +
#973080000000
0!
0'
#973090000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#973100000000
0!
0'
#973110000000
1!
b101 %
1'
b101 +
#973120000000
0!
0'
#973130000000
1!
0$
b110 %
1'
0*
b110 +
#973140000000
0!
0'
#973150000000
1!
b111 %
1'
b111 +
#973160000000
0!
0'
#973170000000
1!
b1000 %
1'
b1000 +
#973180000000
0!
0'
#973190000000
1!
b1001 %
1'
b1001 +
#973200000000
0!
0'
#973210000000
1!
b0 %
1'
b0 +
#973220000000
0!
0'
#973230000000
1!
1$
b1 %
1'
1*
b1 +
#973240000000
0!
0'
#973250000000
1!
b10 %
1'
b10 +
#973260000000
0!
0'
#973270000000
1!
b11 %
1'
b11 +
#973280000000
0!
0'
#973290000000
1!
b100 %
1'
b100 +
#973300000000
1"
1(
#973310000000
0!
0"
b100 &
0'
0(
b100 ,
#973320000000
1!
b101 %
1'
b101 +
#973330000000
0!
0'
#973340000000
1!
b110 %
1'
b110 +
#973350000000
0!
0'
#973360000000
1!
b111 %
1'
b111 +
#973370000000
0!
0'
#973380000000
1!
0$
b1000 %
1'
0*
b1000 +
#973390000000
0!
0'
#973400000000
1!
b1001 %
1'
b1001 +
#973410000000
0!
0'
#973420000000
1!
b0 %
1'
b0 +
#973430000000
0!
0'
#973440000000
1!
1$
b1 %
1'
1*
b1 +
#973450000000
0!
0'
#973460000000
1!
b10 %
1'
b10 +
#973470000000
0!
0'
#973480000000
1!
b11 %
1'
b11 +
#973490000000
0!
0'
#973500000000
1!
b100 %
1'
b100 +
#973510000000
0!
0'
#973520000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#973530000000
0!
0'
#973540000000
1!
0$
b110 %
1'
0*
b110 +
#973550000000
0!
0'
#973560000000
1!
b111 %
1'
b111 +
#973570000000
0!
0'
#973580000000
1!
b1000 %
1'
b1000 +
#973590000000
0!
0'
#973600000000
1!
b1001 %
1'
b1001 +
#973610000000
0!
0'
#973620000000
1!
b0 %
1'
b0 +
#973630000000
0!
0'
#973640000000
1!
1$
b1 %
1'
1*
b1 +
#973650000000
0!
0'
#973660000000
1!
b10 %
1'
b10 +
#973670000000
0!
0'
#973680000000
1!
b11 %
1'
b11 +
#973690000000
0!
0'
#973700000000
1!
b100 %
1'
b100 +
#973710000000
0!
0'
#973720000000
1!
b101 %
1'
b101 +
#973730000000
1"
1(
#973740000000
0!
0"
b100 &
0'
0(
b100 ,
#973750000000
1!
b110 %
1'
b110 +
#973760000000
0!
0'
#973770000000
1!
b111 %
1'
b111 +
#973780000000
0!
0'
#973790000000
1!
0$
b1000 %
1'
0*
b1000 +
#973800000000
0!
0'
#973810000000
1!
b1001 %
1'
b1001 +
#973820000000
0!
0'
#973830000000
1!
b0 %
1'
b0 +
#973840000000
0!
0'
#973850000000
1!
1$
b1 %
1'
1*
b1 +
#973860000000
0!
0'
#973870000000
1!
b10 %
1'
b10 +
#973880000000
0!
0'
#973890000000
1!
b11 %
1'
b11 +
#973900000000
0!
0'
#973910000000
1!
b100 %
1'
b100 +
#973920000000
0!
0'
#973930000000
1!
b101 %
1'
b101 +
#973940000000
0!
0'
#973950000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#973960000000
0!
0'
#973970000000
1!
b111 %
1'
b111 +
#973980000000
0!
0'
#973990000000
1!
b1000 %
1'
b1000 +
#974000000000
0!
0'
#974010000000
1!
b1001 %
1'
b1001 +
#974020000000
0!
0'
#974030000000
1!
b0 %
1'
b0 +
#974040000000
0!
0'
#974050000000
1!
1$
b1 %
1'
1*
b1 +
#974060000000
0!
0'
#974070000000
1!
b10 %
1'
b10 +
#974080000000
0!
0'
#974090000000
1!
b11 %
1'
b11 +
#974100000000
0!
0'
#974110000000
1!
b100 %
1'
b100 +
#974120000000
0!
0'
#974130000000
1!
b101 %
1'
b101 +
#974140000000
0!
0'
#974150000000
1!
0$
b110 %
1'
0*
b110 +
#974160000000
1"
1(
#974170000000
0!
0"
b100 &
0'
0(
b100 ,
#974180000000
1!
1$
b111 %
1'
1*
b111 +
#974190000000
0!
0'
#974200000000
1!
0$
b1000 %
1'
0*
b1000 +
#974210000000
0!
0'
#974220000000
1!
b1001 %
1'
b1001 +
#974230000000
0!
0'
#974240000000
1!
b0 %
1'
b0 +
#974250000000
0!
0'
#974260000000
1!
1$
b1 %
1'
1*
b1 +
#974270000000
0!
0'
#974280000000
1!
b10 %
1'
b10 +
#974290000000
0!
0'
#974300000000
1!
b11 %
1'
b11 +
#974310000000
0!
0'
#974320000000
1!
b100 %
1'
b100 +
#974330000000
0!
0'
#974340000000
1!
b101 %
1'
b101 +
#974350000000
0!
0'
#974360000000
1!
b110 %
1'
b110 +
#974370000000
0!
0'
#974380000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#974390000000
0!
0'
#974400000000
1!
b1000 %
1'
b1000 +
#974410000000
0!
0'
#974420000000
1!
b1001 %
1'
b1001 +
#974430000000
0!
0'
#974440000000
1!
b0 %
1'
b0 +
#974450000000
0!
0'
#974460000000
1!
1$
b1 %
1'
1*
b1 +
#974470000000
0!
0'
#974480000000
1!
b10 %
1'
b10 +
#974490000000
0!
0'
#974500000000
1!
b11 %
1'
b11 +
#974510000000
0!
0'
#974520000000
1!
b100 %
1'
b100 +
#974530000000
0!
0'
#974540000000
1!
b101 %
1'
b101 +
#974550000000
0!
0'
#974560000000
1!
0$
b110 %
1'
0*
b110 +
#974570000000
0!
0'
#974580000000
1!
b111 %
1'
b111 +
#974590000000
1"
1(
#974600000000
0!
0"
b100 &
0'
0(
b100 ,
#974610000000
1!
b1000 %
1'
b1000 +
#974620000000
0!
0'
#974630000000
1!
b1001 %
1'
b1001 +
#974640000000
0!
0'
#974650000000
1!
b0 %
1'
b0 +
#974660000000
0!
0'
#974670000000
1!
1$
b1 %
1'
1*
b1 +
#974680000000
0!
0'
#974690000000
1!
b10 %
1'
b10 +
#974700000000
0!
0'
#974710000000
1!
b11 %
1'
b11 +
#974720000000
0!
0'
#974730000000
1!
b100 %
1'
b100 +
#974740000000
0!
0'
#974750000000
1!
b101 %
1'
b101 +
#974760000000
0!
0'
#974770000000
1!
b110 %
1'
b110 +
#974780000000
0!
0'
#974790000000
1!
b111 %
1'
b111 +
#974800000000
0!
0'
#974810000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#974820000000
0!
0'
#974830000000
1!
b1001 %
1'
b1001 +
#974840000000
0!
0'
#974850000000
1!
b0 %
1'
b0 +
#974860000000
0!
0'
#974870000000
1!
1$
b1 %
1'
1*
b1 +
#974880000000
0!
0'
#974890000000
1!
b10 %
1'
b10 +
#974900000000
0!
0'
#974910000000
1!
b11 %
1'
b11 +
#974920000000
0!
0'
#974930000000
1!
b100 %
1'
b100 +
#974940000000
0!
0'
#974950000000
1!
b101 %
1'
b101 +
#974960000000
0!
0'
#974970000000
1!
0$
b110 %
1'
0*
b110 +
#974980000000
0!
0'
#974990000000
1!
b111 %
1'
b111 +
#975000000000
0!
0'
#975010000000
1!
b1000 %
1'
b1000 +
#975020000000
1"
1(
#975030000000
0!
0"
b100 &
0'
0(
b100 ,
#975040000000
1!
b1001 %
1'
b1001 +
#975050000000
0!
0'
#975060000000
1!
b0 %
1'
b0 +
#975070000000
0!
0'
#975080000000
1!
1$
b1 %
1'
1*
b1 +
#975090000000
0!
0'
#975100000000
1!
b10 %
1'
b10 +
#975110000000
0!
0'
#975120000000
1!
b11 %
1'
b11 +
#975130000000
0!
0'
#975140000000
1!
b100 %
1'
b100 +
#975150000000
0!
0'
#975160000000
1!
b101 %
1'
b101 +
#975170000000
0!
0'
#975180000000
1!
b110 %
1'
b110 +
#975190000000
0!
0'
#975200000000
1!
b111 %
1'
b111 +
#975210000000
0!
0'
#975220000000
1!
0$
b1000 %
1'
0*
b1000 +
#975230000000
0!
0'
#975240000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#975250000000
0!
0'
#975260000000
1!
b0 %
1'
b0 +
#975270000000
0!
0'
#975280000000
1!
1$
b1 %
1'
1*
b1 +
#975290000000
0!
0'
#975300000000
1!
b10 %
1'
b10 +
#975310000000
0!
0'
#975320000000
1!
b11 %
1'
b11 +
#975330000000
0!
0'
#975340000000
1!
b100 %
1'
b100 +
#975350000000
0!
0'
#975360000000
1!
b101 %
1'
b101 +
#975370000000
0!
0'
#975380000000
1!
0$
b110 %
1'
0*
b110 +
#975390000000
0!
0'
#975400000000
1!
b111 %
1'
b111 +
#975410000000
0!
0'
#975420000000
1!
b1000 %
1'
b1000 +
#975430000000
0!
0'
#975440000000
1!
b1001 %
1'
b1001 +
#975450000000
1"
1(
#975460000000
0!
0"
b100 &
0'
0(
b100 ,
#975470000000
1!
b0 %
1'
b0 +
#975480000000
0!
0'
#975490000000
1!
1$
b1 %
1'
1*
b1 +
#975500000000
0!
0'
#975510000000
1!
b10 %
1'
b10 +
#975520000000
0!
0'
#975530000000
1!
b11 %
1'
b11 +
#975540000000
0!
0'
#975550000000
1!
b100 %
1'
b100 +
#975560000000
0!
0'
#975570000000
1!
b101 %
1'
b101 +
#975580000000
0!
0'
#975590000000
1!
b110 %
1'
b110 +
#975600000000
0!
0'
#975610000000
1!
b111 %
1'
b111 +
#975620000000
0!
0'
#975630000000
1!
0$
b1000 %
1'
0*
b1000 +
#975640000000
0!
0'
#975650000000
1!
b1001 %
1'
b1001 +
#975660000000
0!
0'
#975670000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#975680000000
0!
0'
#975690000000
1!
1$
b1 %
1'
1*
b1 +
#975700000000
0!
0'
#975710000000
1!
b10 %
1'
b10 +
#975720000000
0!
0'
#975730000000
1!
b11 %
1'
b11 +
#975740000000
0!
0'
#975750000000
1!
b100 %
1'
b100 +
#975760000000
0!
0'
#975770000000
1!
b101 %
1'
b101 +
#975780000000
0!
0'
#975790000000
1!
0$
b110 %
1'
0*
b110 +
#975800000000
0!
0'
#975810000000
1!
b111 %
1'
b111 +
#975820000000
0!
0'
#975830000000
1!
b1000 %
1'
b1000 +
#975840000000
0!
0'
#975850000000
1!
b1001 %
1'
b1001 +
#975860000000
0!
0'
#975870000000
1!
b0 %
1'
b0 +
#975880000000
1"
1(
#975890000000
0!
0"
b100 &
0'
0(
b100 ,
#975900000000
1!
1$
b1 %
1'
1*
b1 +
#975910000000
0!
0'
#975920000000
1!
b10 %
1'
b10 +
#975930000000
0!
0'
#975940000000
1!
b11 %
1'
b11 +
#975950000000
0!
0'
#975960000000
1!
b100 %
1'
b100 +
#975970000000
0!
0'
#975980000000
1!
b101 %
1'
b101 +
#975990000000
0!
0'
#976000000000
1!
b110 %
1'
b110 +
#976010000000
0!
0'
#976020000000
1!
b111 %
1'
b111 +
#976030000000
0!
0'
#976040000000
1!
0$
b1000 %
1'
0*
b1000 +
#976050000000
0!
0'
#976060000000
1!
b1001 %
1'
b1001 +
#976070000000
0!
0'
#976080000000
1!
b0 %
1'
b0 +
#976090000000
0!
0'
#976100000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#976110000000
0!
0'
#976120000000
1!
b10 %
1'
b10 +
#976130000000
0!
0'
#976140000000
1!
b11 %
1'
b11 +
#976150000000
0!
0'
#976160000000
1!
b100 %
1'
b100 +
#976170000000
0!
0'
#976180000000
1!
b101 %
1'
b101 +
#976190000000
0!
0'
#976200000000
1!
0$
b110 %
1'
0*
b110 +
#976210000000
0!
0'
#976220000000
1!
b111 %
1'
b111 +
#976230000000
0!
0'
#976240000000
1!
b1000 %
1'
b1000 +
#976250000000
0!
0'
#976260000000
1!
b1001 %
1'
b1001 +
#976270000000
0!
0'
#976280000000
1!
b0 %
1'
b0 +
#976290000000
0!
0'
#976300000000
1!
1$
b1 %
1'
1*
b1 +
#976310000000
1"
1(
#976320000000
0!
0"
b100 &
0'
0(
b100 ,
#976330000000
1!
b10 %
1'
b10 +
#976340000000
0!
0'
#976350000000
1!
b11 %
1'
b11 +
#976360000000
0!
0'
#976370000000
1!
b100 %
1'
b100 +
#976380000000
0!
0'
#976390000000
1!
b101 %
1'
b101 +
#976400000000
0!
0'
#976410000000
1!
b110 %
1'
b110 +
#976420000000
0!
0'
#976430000000
1!
b111 %
1'
b111 +
#976440000000
0!
0'
#976450000000
1!
0$
b1000 %
1'
0*
b1000 +
#976460000000
0!
0'
#976470000000
1!
b1001 %
1'
b1001 +
#976480000000
0!
0'
#976490000000
1!
b0 %
1'
b0 +
#976500000000
0!
0'
#976510000000
1!
1$
b1 %
1'
1*
b1 +
#976520000000
0!
0'
#976530000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#976540000000
0!
0'
#976550000000
1!
b11 %
1'
b11 +
#976560000000
0!
0'
#976570000000
1!
b100 %
1'
b100 +
#976580000000
0!
0'
#976590000000
1!
b101 %
1'
b101 +
#976600000000
0!
0'
#976610000000
1!
0$
b110 %
1'
0*
b110 +
#976620000000
0!
0'
#976630000000
1!
b111 %
1'
b111 +
#976640000000
0!
0'
#976650000000
1!
b1000 %
1'
b1000 +
#976660000000
0!
0'
#976670000000
1!
b1001 %
1'
b1001 +
#976680000000
0!
0'
#976690000000
1!
b0 %
1'
b0 +
#976700000000
0!
0'
#976710000000
1!
1$
b1 %
1'
1*
b1 +
#976720000000
0!
0'
#976730000000
1!
b10 %
1'
b10 +
#976740000000
1"
1(
#976750000000
0!
0"
b100 &
0'
0(
b100 ,
#976760000000
1!
b11 %
1'
b11 +
#976770000000
0!
0'
#976780000000
1!
b100 %
1'
b100 +
#976790000000
0!
0'
#976800000000
1!
b101 %
1'
b101 +
#976810000000
0!
0'
#976820000000
1!
b110 %
1'
b110 +
#976830000000
0!
0'
#976840000000
1!
b111 %
1'
b111 +
#976850000000
0!
0'
#976860000000
1!
0$
b1000 %
1'
0*
b1000 +
#976870000000
0!
0'
#976880000000
1!
b1001 %
1'
b1001 +
#976890000000
0!
0'
#976900000000
1!
b0 %
1'
b0 +
#976910000000
0!
0'
#976920000000
1!
1$
b1 %
1'
1*
b1 +
#976930000000
0!
0'
#976940000000
1!
b10 %
1'
b10 +
#976950000000
0!
0'
#976960000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#976970000000
0!
0'
#976980000000
1!
b100 %
1'
b100 +
#976990000000
0!
0'
#977000000000
1!
b101 %
1'
b101 +
#977010000000
0!
0'
#977020000000
1!
0$
b110 %
1'
0*
b110 +
#977030000000
0!
0'
#977040000000
1!
b111 %
1'
b111 +
#977050000000
0!
0'
#977060000000
1!
b1000 %
1'
b1000 +
#977070000000
0!
0'
#977080000000
1!
b1001 %
1'
b1001 +
#977090000000
0!
0'
#977100000000
1!
b0 %
1'
b0 +
#977110000000
0!
0'
#977120000000
1!
1$
b1 %
1'
1*
b1 +
#977130000000
0!
0'
#977140000000
1!
b10 %
1'
b10 +
#977150000000
0!
0'
#977160000000
1!
b11 %
1'
b11 +
#977170000000
1"
1(
#977180000000
0!
0"
b100 &
0'
0(
b100 ,
#977190000000
1!
b100 %
1'
b100 +
#977200000000
0!
0'
#977210000000
1!
b101 %
1'
b101 +
#977220000000
0!
0'
#977230000000
1!
b110 %
1'
b110 +
#977240000000
0!
0'
#977250000000
1!
b111 %
1'
b111 +
#977260000000
0!
0'
#977270000000
1!
0$
b1000 %
1'
0*
b1000 +
#977280000000
0!
0'
#977290000000
1!
b1001 %
1'
b1001 +
#977300000000
0!
0'
#977310000000
1!
b0 %
1'
b0 +
#977320000000
0!
0'
#977330000000
1!
1$
b1 %
1'
1*
b1 +
#977340000000
0!
0'
#977350000000
1!
b10 %
1'
b10 +
#977360000000
0!
0'
#977370000000
1!
b11 %
1'
b11 +
#977380000000
0!
0'
#977390000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#977400000000
0!
0'
#977410000000
1!
b101 %
1'
b101 +
#977420000000
0!
0'
#977430000000
1!
0$
b110 %
1'
0*
b110 +
#977440000000
0!
0'
#977450000000
1!
b111 %
1'
b111 +
#977460000000
0!
0'
#977470000000
1!
b1000 %
1'
b1000 +
#977480000000
0!
0'
#977490000000
1!
b1001 %
1'
b1001 +
#977500000000
0!
0'
#977510000000
1!
b0 %
1'
b0 +
#977520000000
0!
0'
#977530000000
1!
1$
b1 %
1'
1*
b1 +
#977540000000
0!
0'
#977550000000
1!
b10 %
1'
b10 +
#977560000000
0!
0'
#977570000000
1!
b11 %
1'
b11 +
#977580000000
0!
0'
#977590000000
1!
b100 %
1'
b100 +
#977600000000
1"
1(
#977610000000
0!
0"
b100 &
0'
0(
b100 ,
#977620000000
1!
b101 %
1'
b101 +
#977630000000
0!
0'
#977640000000
1!
b110 %
1'
b110 +
#977650000000
0!
0'
#977660000000
1!
b111 %
1'
b111 +
#977670000000
0!
0'
#977680000000
1!
0$
b1000 %
1'
0*
b1000 +
#977690000000
0!
0'
#977700000000
1!
b1001 %
1'
b1001 +
#977710000000
0!
0'
#977720000000
1!
b0 %
1'
b0 +
#977730000000
0!
0'
#977740000000
1!
1$
b1 %
1'
1*
b1 +
#977750000000
0!
0'
#977760000000
1!
b10 %
1'
b10 +
#977770000000
0!
0'
#977780000000
1!
b11 %
1'
b11 +
#977790000000
0!
0'
#977800000000
1!
b100 %
1'
b100 +
#977810000000
0!
0'
#977820000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#977830000000
0!
0'
#977840000000
1!
0$
b110 %
1'
0*
b110 +
#977850000000
0!
0'
#977860000000
1!
b111 %
1'
b111 +
#977870000000
0!
0'
#977880000000
1!
b1000 %
1'
b1000 +
#977890000000
0!
0'
#977900000000
1!
b1001 %
1'
b1001 +
#977910000000
0!
0'
#977920000000
1!
b0 %
1'
b0 +
#977930000000
0!
0'
#977940000000
1!
1$
b1 %
1'
1*
b1 +
#977950000000
0!
0'
#977960000000
1!
b10 %
1'
b10 +
#977970000000
0!
0'
#977980000000
1!
b11 %
1'
b11 +
#977990000000
0!
0'
#978000000000
1!
b100 %
1'
b100 +
#978010000000
0!
0'
#978020000000
1!
b101 %
1'
b101 +
#978030000000
1"
1(
#978040000000
0!
0"
b100 &
0'
0(
b100 ,
#978050000000
1!
b110 %
1'
b110 +
#978060000000
0!
0'
#978070000000
1!
b111 %
1'
b111 +
#978080000000
0!
0'
#978090000000
1!
0$
b1000 %
1'
0*
b1000 +
#978100000000
0!
0'
#978110000000
1!
b1001 %
1'
b1001 +
#978120000000
0!
0'
#978130000000
1!
b0 %
1'
b0 +
#978140000000
0!
0'
#978150000000
1!
1$
b1 %
1'
1*
b1 +
#978160000000
0!
0'
#978170000000
1!
b10 %
1'
b10 +
#978180000000
0!
0'
#978190000000
1!
b11 %
1'
b11 +
#978200000000
0!
0'
#978210000000
1!
b100 %
1'
b100 +
#978220000000
0!
0'
#978230000000
1!
b101 %
1'
b101 +
#978240000000
0!
0'
#978250000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#978260000000
0!
0'
#978270000000
1!
b111 %
1'
b111 +
#978280000000
0!
0'
#978290000000
1!
b1000 %
1'
b1000 +
#978300000000
0!
0'
#978310000000
1!
b1001 %
1'
b1001 +
#978320000000
0!
0'
#978330000000
1!
b0 %
1'
b0 +
#978340000000
0!
0'
#978350000000
1!
1$
b1 %
1'
1*
b1 +
#978360000000
0!
0'
#978370000000
1!
b10 %
1'
b10 +
#978380000000
0!
0'
#978390000000
1!
b11 %
1'
b11 +
#978400000000
0!
0'
#978410000000
1!
b100 %
1'
b100 +
#978420000000
0!
0'
#978430000000
1!
b101 %
1'
b101 +
#978440000000
0!
0'
#978450000000
1!
0$
b110 %
1'
0*
b110 +
#978460000000
1"
1(
#978470000000
0!
0"
b100 &
0'
0(
b100 ,
#978480000000
1!
1$
b111 %
1'
1*
b111 +
#978490000000
0!
0'
#978500000000
1!
0$
b1000 %
1'
0*
b1000 +
#978510000000
0!
0'
#978520000000
1!
b1001 %
1'
b1001 +
#978530000000
0!
0'
#978540000000
1!
b0 %
1'
b0 +
#978550000000
0!
0'
#978560000000
1!
1$
b1 %
1'
1*
b1 +
#978570000000
0!
0'
#978580000000
1!
b10 %
1'
b10 +
#978590000000
0!
0'
#978600000000
1!
b11 %
1'
b11 +
#978610000000
0!
0'
#978620000000
1!
b100 %
1'
b100 +
#978630000000
0!
0'
#978640000000
1!
b101 %
1'
b101 +
#978650000000
0!
0'
#978660000000
1!
b110 %
1'
b110 +
#978670000000
0!
0'
#978680000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#978690000000
0!
0'
#978700000000
1!
b1000 %
1'
b1000 +
#978710000000
0!
0'
#978720000000
1!
b1001 %
1'
b1001 +
#978730000000
0!
0'
#978740000000
1!
b0 %
1'
b0 +
#978750000000
0!
0'
#978760000000
1!
1$
b1 %
1'
1*
b1 +
#978770000000
0!
0'
#978780000000
1!
b10 %
1'
b10 +
#978790000000
0!
0'
#978800000000
1!
b11 %
1'
b11 +
#978810000000
0!
0'
#978820000000
1!
b100 %
1'
b100 +
#978830000000
0!
0'
#978840000000
1!
b101 %
1'
b101 +
#978850000000
0!
0'
#978860000000
1!
0$
b110 %
1'
0*
b110 +
#978870000000
0!
0'
#978880000000
1!
b111 %
1'
b111 +
#978890000000
1"
1(
#978900000000
0!
0"
b100 &
0'
0(
b100 ,
#978910000000
1!
b1000 %
1'
b1000 +
#978920000000
0!
0'
#978930000000
1!
b1001 %
1'
b1001 +
#978940000000
0!
0'
#978950000000
1!
b0 %
1'
b0 +
#978960000000
0!
0'
#978970000000
1!
1$
b1 %
1'
1*
b1 +
#978980000000
0!
0'
#978990000000
1!
b10 %
1'
b10 +
#979000000000
0!
0'
#979010000000
1!
b11 %
1'
b11 +
#979020000000
0!
0'
#979030000000
1!
b100 %
1'
b100 +
#979040000000
0!
0'
#979050000000
1!
b101 %
1'
b101 +
#979060000000
0!
0'
#979070000000
1!
b110 %
1'
b110 +
#979080000000
0!
0'
#979090000000
1!
b111 %
1'
b111 +
#979100000000
0!
0'
#979110000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#979120000000
0!
0'
#979130000000
1!
b1001 %
1'
b1001 +
#979140000000
0!
0'
#979150000000
1!
b0 %
1'
b0 +
#979160000000
0!
0'
#979170000000
1!
1$
b1 %
1'
1*
b1 +
#979180000000
0!
0'
#979190000000
1!
b10 %
1'
b10 +
#979200000000
0!
0'
#979210000000
1!
b11 %
1'
b11 +
#979220000000
0!
0'
#979230000000
1!
b100 %
1'
b100 +
#979240000000
0!
0'
#979250000000
1!
b101 %
1'
b101 +
#979260000000
0!
0'
#979270000000
1!
0$
b110 %
1'
0*
b110 +
#979280000000
0!
0'
#979290000000
1!
b111 %
1'
b111 +
#979300000000
0!
0'
#979310000000
1!
b1000 %
1'
b1000 +
#979320000000
1"
1(
#979330000000
0!
0"
b100 &
0'
0(
b100 ,
#979340000000
1!
b1001 %
1'
b1001 +
#979350000000
0!
0'
#979360000000
1!
b0 %
1'
b0 +
#979370000000
0!
0'
#979380000000
1!
1$
b1 %
1'
1*
b1 +
#979390000000
0!
0'
#979400000000
1!
b10 %
1'
b10 +
#979410000000
0!
0'
#979420000000
1!
b11 %
1'
b11 +
#979430000000
0!
0'
#979440000000
1!
b100 %
1'
b100 +
#979450000000
0!
0'
#979460000000
1!
b101 %
1'
b101 +
#979470000000
0!
0'
#979480000000
1!
b110 %
1'
b110 +
#979490000000
0!
0'
#979500000000
1!
b111 %
1'
b111 +
#979510000000
0!
0'
#979520000000
1!
0$
b1000 %
1'
0*
b1000 +
#979530000000
0!
0'
#979540000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#979550000000
0!
0'
#979560000000
1!
b0 %
1'
b0 +
#979570000000
0!
0'
#979580000000
1!
1$
b1 %
1'
1*
b1 +
#979590000000
0!
0'
#979600000000
1!
b10 %
1'
b10 +
#979610000000
0!
0'
#979620000000
1!
b11 %
1'
b11 +
#979630000000
0!
0'
#979640000000
1!
b100 %
1'
b100 +
#979650000000
0!
0'
#979660000000
1!
b101 %
1'
b101 +
#979670000000
0!
0'
#979680000000
1!
0$
b110 %
1'
0*
b110 +
#979690000000
0!
0'
#979700000000
1!
b111 %
1'
b111 +
#979710000000
0!
0'
#979720000000
1!
b1000 %
1'
b1000 +
#979730000000
0!
0'
#979740000000
1!
b1001 %
1'
b1001 +
#979750000000
1"
1(
#979760000000
0!
0"
b100 &
0'
0(
b100 ,
#979770000000
1!
b0 %
1'
b0 +
#979780000000
0!
0'
#979790000000
1!
1$
b1 %
1'
1*
b1 +
#979800000000
0!
0'
#979810000000
1!
b10 %
1'
b10 +
#979820000000
0!
0'
#979830000000
1!
b11 %
1'
b11 +
#979840000000
0!
0'
#979850000000
1!
b100 %
1'
b100 +
#979860000000
0!
0'
#979870000000
1!
b101 %
1'
b101 +
#979880000000
0!
0'
#979890000000
1!
b110 %
1'
b110 +
#979900000000
0!
0'
#979910000000
1!
b111 %
1'
b111 +
#979920000000
0!
0'
#979930000000
1!
0$
b1000 %
1'
0*
b1000 +
#979940000000
0!
0'
#979950000000
1!
b1001 %
1'
b1001 +
#979960000000
0!
0'
#979970000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#979980000000
0!
0'
#979990000000
1!
1$
b1 %
1'
1*
b1 +
#980000000000
0!
0'
#980010000000
1!
b10 %
1'
b10 +
#980020000000
0!
0'
#980030000000
1!
b11 %
1'
b11 +
#980040000000
0!
0'
#980050000000
1!
b100 %
1'
b100 +
#980060000000
0!
0'
#980070000000
1!
b101 %
1'
b101 +
#980080000000
0!
0'
#980090000000
1!
0$
b110 %
1'
0*
b110 +
#980100000000
0!
0'
#980110000000
1!
b111 %
1'
b111 +
#980120000000
0!
0'
#980130000000
1!
b1000 %
1'
b1000 +
#980140000000
0!
0'
#980150000000
1!
b1001 %
1'
b1001 +
#980160000000
0!
0'
#980170000000
1!
b0 %
1'
b0 +
#980180000000
1"
1(
#980190000000
0!
0"
b100 &
0'
0(
b100 ,
#980200000000
1!
1$
b1 %
1'
1*
b1 +
#980210000000
0!
0'
#980220000000
1!
b10 %
1'
b10 +
#980230000000
0!
0'
#980240000000
1!
b11 %
1'
b11 +
#980250000000
0!
0'
#980260000000
1!
b100 %
1'
b100 +
#980270000000
0!
0'
#980280000000
1!
b101 %
1'
b101 +
#980290000000
0!
0'
#980300000000
1!
b110 %
1'
b110 +
#980310000000
0!
0'
#980320000000
1!
b111 %
1'
b111 +
#980330000000
0!
0'
#980340000000
1!
0$
b1000 %
1'
0*
b1000 +
#980350000000
0!
0'
#980360000000
1!
b1001 %
1'
b1001 +
#980370000000
0!
0'
#980380000000
1!
b0 %
1'
b0 +
#980390000000
0!
0'
#980400000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#980410000000
0!
0'
#980420000000
1!
b10 %
1'
b10 +
#980430000000
0!
0'
#980440000000
1!
b11 %
1'
b11 +
#980450000000
0!
0'
#980460000000
1!
b100 %
1'
b100 +
#980470000000
0!
0'
#980480000000
1!
b101 %
1'
b101 +
#980490000000
0!
0'
#980500000000
1!
0$
b110 %
1'
0*
b110 +
#980510000000
0!
0'
#980520000000
1!
b111 %
1'
b111 +
#980530000000
0!
0'
#980540000000
1!
b1000 %
1'
b1000 +
#980550000000
0!
0'
#980560000000
1!
b1001 %
1'
b1001 +
#980570000000
0!
0'
#980580000000
1!
b0 %
1'
b0 +
#980590000000
0!
0'
#980600000000
1!
1$
b1 %
1'
1*
b1 +
#980610000000
1"
1(
#980620000000
0!
0"
b100 &
0'
0(
b100 ,
#980630000000
1!
b10 %
1'
b10 +
#980640000000
0!
0'
#980650000000
1!
b11 %
1'
b11 +
#980660000000
0!
0'
#980670000000
1!
b100 %
1'
b100 +
#980680000000
0!
0'
#980690000000
1!
b101 %
1'
b101 +
#980700000000
0!
0'
#980710000000
1!
b110 %
1'
b110 +
#980720000000
0!
0'
#980730000000
1!
b111 %
1'
b111 +
#980740000000
0!
0'
#980750000000
1!
0$
b1000 %
1'
0*
b1000 +
#980760000000
0!
0'
#980770000000
1!
b1001 %
1'
b1001 +
#980780000000
0!
0'
#980790000000
1!
b0 %
1'
b0 +
#980800000000
0!
0'
#980810000000
1!
1$
b1 %
1'
1*
b1 +
#980820000000
0!
0'
#980830000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#980840000000
0!
0'
#980850000000
1!
b11 %
1'
b11 +
#980860000000
0!
0'
#980870000000
1!
b100 %
1'
b100 +
#980880000000
0!
0'
#980890000000
1!
b101 %
1'
b101 +
#980900000000
0!
0'
#980910000000
1!
0$
b110 %
1'
0*
b110 +
#980920000000
0!
0'
#980930000000
1!
b111 %
1'
b111 +
#980940000000
0!
0'
#980950000000
1!
b1000 %
1'
b1000 +
#980960000000
0!
0'
#980970000000
1!
b1001 %
1'
b1001 +
#980980000000
0!
0'
#980990000000
1!
b0 %
1'
b0 +
#981000000000
0!
0'
#981010000000
1!
1$
b1 %
1'
1*
b1 +
#981020000000
0!
0'
#981030000000
1!
b10 %
1'
b10 +
#981040000000
1"
1(
#981050000000
0!
0"
b100 &
0'
0(
b100 ,
#981060000000
1!
b11 %
1'
b11 +
#981070000000
0!
0'
#981080000000
1!
b100 %
1'
b100 +
#981090000000
0!
0'
#981100000000
1!
b101 %
1'
b101 +
#981110000000
0!
0'
#981120000000
1!
b110 %
1'
b110 +
#981130000000
0!
0'
#981140000000
1!
b111 %
1'
b111 +
#981150000000
0!
0'
#981160000000
1!
0$
b1000 %
1'
0*
b1000 +
#981170000000
0!
0'
#981180000000
1!
b1001 %
1'
b1001 +
#981190000000
0!
0'
#981200000000
1!
b0 %
1'
b0 +
#981210000000
0!
0'
#981220000000
1!
1$
b1 %
1'
1*
b1 +
#981230000000
0!
0'
#981240000000
1!
b10 %
1'
b10 +
#981250000000
0!
0'
#981260000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#981270000000
0!
0'
#981280000000
1!
b100 %
1'
b100 +
#981290000000
0!
0'
#981300000000
1!
b101 %
1'
b101 +
#981310000000
0!
0'
#981320000000
1!
0$
b110 %
1'
0*
b110 +
#981330000000
0!
0'
#981340000000
1!
b111 %
1'
b111 +
#981350000000
0!
0'
#981360000000
1!
b1000 %
1'
b1000 +
#981370000000
0!
0'
#981380000000
1!
b1001 %
1'
b1001 +
#981390000000
0!
0'
#981400000000
1!
b0 %
1'
b0 +
#981410000000
0!
0'
#981420000000
1!
1$
b1 %
1'
1*
b1 +
#981430000000
0!
0'
#981440000000
1!
b10 %
1'
b10 +
#981450000000
0!
0'
#981460000000
1!
b11 %
1'
b11 +
#981470000000
1"
1(
#981480000000
0!
0"
b100 &
0'
0(
b100 ,
#981490000000
1!
b100 %
1'
b100 +
#981500000000
0!
0'
#981510000000
1!
b101 %
1'
b101 +
#981520000000
0!
0'
#981530000000
1!
b110 %
1'
b110 +
#981540000000
0!
0'
#981550000000
1!
b111 %
1'
b111 +
#981560000000
0!
0'
#981570000000
1!
0$
b1000 %
1'
0*
b1000 +
#981580000000
0!
0'
#981590000000
1!
b1001 %
1'
b1001 +
#981600000000
0!
0'
#981610000000
1!
b0 %
1'
b0 +
#981620000000
0!
0'
#981630000000
1!
1$
b1 %
1'
1*
b1 +
#981640000000
0!
0'
#981650000000
1!
b10 %
1'
b10 +
#981660000000
0!
0'
#981670000000
1!
b11 %
1'
b11 +
#981680000000
0!
0'
#981690000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#981700000000
0!
0'
#981710000000
1!
b101 %
1'
b101 +
#981720000000
0!
0'
#981730000000
1!
0$
b110 %
1'
0*
b110 +
#981740000000
0!
0'
#981750000000
1!
b111 %
1'
b111 +
#981760000000
0!
0'
#981770000000
1!
b1000 %
1'
b1000 +
#981780000000
0!
0'
#981790000000
1!
b1001 %
1'
b1001 +
#981800000000
0!
0'
#981810000000
1!
b0 %
1'
b0 +
#981820000000
0!
0'
#981830000000
1!
1$
b1 %
1'
1*
b1 +
#981840000000
0!
0'
#981850000000
1!
b10 %
1'
b10 +
#981860000000
0!
0'
#981870000000
1!
b11 %
1'
b11 +
#981880000000
0!
0'
#981890000000
1!
b100 %
1'
b100 +
#981900000000
1"
1(
#981910000000
0!
0"
b100 &
0'
0(
b100 ,
#981920000000
1!
b101 %
1'
b101 +
#981930000000
0!
0'
#981940000000
1!
b110 %
1'
b110 +
#981950000000
0!
0'
#981960000000
1!
b111 %
1'
b111 +
#981970000000
0!
0'
#981980000000
1!
0$
b1000 %
1'
0*
b1000 +
#981990000000
0!
0'
#982000000000
1!
b1001 %
1'
b1001 +
#982010000000
0!
0'
#982020000000
1!
b0 %
1'
b0 +
#982030000000
0!
0'
#982040000000
1!
1$
b1 %
1'
1*
b1 +
#982050000000
0!
0'
#982060000000
1!
b10 %
1'
b10 +
#982070000000
0!
0'
#982080000000
1!
b11 %
1'
b11 +
#982090000000
0!
0'
#982100000000
1!
b100 %
1'
b100 +
#982110000000
0!
0'
#982120000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#982130000000
0!
0'
#982140000000
1!
0$
b110 %
1'
0*
b110 +
#982150000000
0!
0'
#982160000000
1!
b111 %
1'
b111 +
#982170000000
0!
0'
#982180000000
1!
b1000 %
1'
b1000 +
#982190000000
0!
0'
#982200000000
1!
b1001 %
1'
b1001 +
#982210000000
0!
0'
#982220000000
1!
b0 %
1'
b0 +
#982230000000
0!
0'
#982240000000
1!
1$
b1 %
1'
1*
b1 +
#982250000000
0!
0'
#982260000000
1!
b10 %
1'
b10 +
#982270000000
0!
0'
#982280000000
1!
b11 %
1'
b11 +
#982290000000
0!
0'
#982300000000
1!
b100 %
1'
b100 +
#982310000000
0!
0'
#982320000000
1!
b101 %
1'
b101 +
#982330000000
1"
1(
#982340000000
0!
0"
b100 &
0'
0(
b100 ,
#982350000000
1!
b110 %
1'
b110 +
#982360000000
0!
0'
#982370000000
1!
b111 %
1'
b111 +
#982380000000
0!
0'
#982390000000
1!
0$
b1000 %
1'
0*
b1000 +
#982400000000
0!
0'
#982410000000
1!
b1001 %
1'
b1001 +
#982420000000
0!
0'
#982430000000
1!
b0 %
1'
b0 +
#982440000000
0!
0'
#982450000000
1!
1$
b1 %
1'
1*
b1 +
#982460000000
0!
0'
#982470000000
1!
b10 %
1'
b10 +
#982480000000
0!
0'
#982490000000
1!
b11 %
1'
b11 +
#982500000000
0!
0'
#982510000000
1!
b100 %
1'
b100 +
#982520000000
0!
0'
#982530000000
1!
b101 %
1'
b101 +
#982540000000
0!
0'
#982550000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#982560000000
0!
0'
#982570000000
1!
b111 %
1'
b111 +
#982580000000
0!
0'
#982590000000
1!
b1000 %
1'
b1000 +
#982600000000
0!
0'
#982610000000
1!
b1001 %
1'
b1001 +
#982620000000
0!
0'
#982630000000
1!
b0 %
1'
b0 +
#982640000000
0!
0'
#982650000000
1!
1$
b1 %
1'
1*
b1 +
#982660000000
0!
0'
#982670000000
1!
b10 %
1'
b10 +
#982680000000
0!
0'
#982690000000
1!
b11 %
1'
b11 +
#982700000000
0!
0'
#982710000000
1!
b100 %
1'
b100 +
#982720000000
0!
0'
#982730000000
1!
b101 %
1'
b101 +
#982740000000
0!
0'
#982750000000
1!
0$
b110 %
1'
0*
b110 +
#982760000000
1"
1(
#982770000000
0!
0"
b100 &
0'
0(
b100 ,
#982780000000
1!
1$
b111 %
1'
1*
b111 +
#982790000000
0!
0'
#982800000000
1!
0$
b1000 %
1'
0*
b1000 +
#982810000000
0!
0'
#982820000000
1!
b1001 %
1'
b1001 +
#982830000000
0!
0'
#982840000000
1!
b0 %
1'
b0 +
#982850000000
0!
0'
#982860000000
1!
1$
b1 %
1'
1*
b1 +
#982870000000
0!
0'
#982880000000
1!
b10 %
1'
b10 +
#982890000000
0!
0'
#982900000000
1!
b11 %
1'
b11 +
#982910000000
0!
0'
#982920000000
1!
b100 %
1'
b100 +
#982930000000
0!
0'
#982940000000
1!
b101 %
1'
b101 +
#982950000000
0!
0'
#982960000000
1!
b110 %
1'
b110 +
#982970000000
0!
0'
#982980000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#982990000000
0!
0'
#983000000000
1!
b1000 %
1'
b1000 +
#983010000000
0!
0'
#983020000000
1!
b1001 %
1'
b1001 +
#983030000000
0!
0'
#983040000000
1!
b0 %
1'
b0 +
#983050000000
0!
0'
#983060000000
1!
1$
b1 %
1'
1*
b1 +
#983070000000
0!
0'
#983080000000
1!
b10 %
1'
b10 +
#983090000000
0!
0'
#983100000000
1!
b11 %
1'
b11 +
#983110000000
0!
0'
#983120000000
1!
b100 %
1'
b100 +
#983130000000
0!
0'
#983140000000
1!
b101 %
1'
b101 +
#983150000000
0!
0'
#983160000000
1!
0$
b110 %
1'
0*
b110 +
#983170000000
0!
0'
#983180000000
1!
b111 %
1'
b111 +
#983190000000
1"
1(
#983200000000
0!
0"
b100 &
0'
0(
b100 ,
#983210000000
1!
b1000 %
1'
b1000 +
#983220000000
0!
0'
#983230000000
1!
b1001 %
1'
b1001 +
#983240000000
0!
0'
#983250000000
1!
b0 %
1'
b0 +
#983260000000
0!
0'
#983270000000
1!
1$
b1 %
1'
1*
b1 +
#983280000000
0!
0'
#983290000000
1!
b10 %
1'
b10 +
#983300000000
0!
0'
#983310000000
1!
b11 %
1'
b11 +
#983320000000
0!
0'
#983330000000
1!
b100 %
1'
b100 +
#983340000000
0!
0'
#983350000000
1!
b101 %
1'
b101 +
#983360000000
0!
0'
#983370000000
1!
b110 %
1'
b110 +
#983380000000
0!
0'
#983390000000
1!
b111 %
1'
b111 +
#983400000000
0!
0'
#983410000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#983420000000
0!
0'
#983430000000
1!
b1001 %
1'
b1001 +
#983440000000
0!
0'
#983450000000
1!
b0 %
1'
b0 +
#983460000000
0!
0'
#983470000000
1!
1$
b1 %
1'
1*
b1 +
#983480000000
0!
0'
#983490000000
1!
b10 %
1'
b10 +
#983500000000
0!
0'
#983510000000
1!
b11 %
1'
b11 +
#983520000000
0!
0'
#983530000000
1!
b100 %
1'
b100 +
#983540000000
0!
0'
#983550000000
1!
b101 %
1'
b101 +
#983560000000
0!
0'
#983570000000
1!
0$
b110 %
1'
0*
b110 +
#983580000000
0!
0'
#983590000000
1!
b111 %
1'
b111 +
#983600000000
0!
0'
#983610000000
1!
b1000 %
1'
b1000 +
#983620000000
1"
1(
#983630000000
0!
0"
b100 &
0'
0(
b100 ,
#983640000000
1!
b1001 %
1'
b1001 +
#983650000000
0!
0'
#983660000000
1!
b0 %
1'
b0 +
#983670000000
0!
0'
#983680000000
1!
1$
b1 %
1'
1*
b1 +
#983690000000
0!
0'
#983700000000
1!
b10 %
1'
b10 +
#983710000000
0!
0'
#983720000000
1!
b11 %
1'
b11 +
#983730000000
0!
0'
#983740000000
1!
b100 %
1'
b100 +
#983750000000
0!
0'
#983760000000
1!
b101 %
1'
b101 +
#983770000000
0!
0'
#983780000000
1!
b110 %
1'
b110 +
#983790000000
0!
0'
#983800000000
1!
b111 %
1'
b111 +
#983810000000
0!
0'
#983820000000
1!
0$
b1000 %
1'
0*
b1000 +
#983830000000
0!
0'
#983840000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#983850000000
0!
0'
#983860000000
1!
b0 %
1'
b0 +
#983870000000
0!
0'
#983880000000
1!
1$
b1 %
1'
1*
b1 +
#983890000000
0!
0'
#983900000000
1!
b10 %
1'
b10 +
#983910000000
0!
0'
#983920000000
1!
b11 %
1'
b11 +
#983930000000
0!
0'
#983940000000
1!
b100 %
1'
b100 +
#983950000000
0!
0'
#983960000000
1!
b101 %
1'
b101 +
#983970000000
0!
0'
#983980000000
1!
0$
b110 %
1'
0*
b110 +
#983990000000
0!
0'
#984000000000
1!
b111 %
1'
b111 +
#984010000000
0!
0'
#984020000000
1!
b1000 %
1'
b1000 +
#984030000000
0!
0'
#984040000000
1!
b1001 %
1'
b1001 +
#984050000000
1"
1(
#984060000000
0!
0"
b100 &
0'
0(
b100 ,
#984070000000
1!
b0 %
1'
b0 +
#984080000000
0!
0'
#984090000000
1!
1$
b1 %
1'
1*
b1 +
#984100000000
0!
0'
#984110000000
1!
b10 %
1'
b10 +
#984120000000
0!
0'
#984130000000
1!
b11 %
1'
b11 +
#984140000000
0!
0'
#984150000000
1!
b100 %
1'
b100 +
#984160000000
0!
0'
#984170000000
1!
b101 %
1'
b101 +
#984180000000
0!
0'
#984190000000
1!
b110 %
1'
b110 +
#984200000000
0!
0'
#984210000000
1!
b111 %
1'
b111 +
#984220000000
0!
0'
#984230000000
1!
0$
b1000 %
1'
0*
b1000 +
#984240000000
0!
0'
#984250000000
1!
b1001 %
1'
b1001 +
#984260000000
0!
0'
#984270000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#984280000000
0!
0'
#984290000000
1!
1$
b1 %
1'
1*
b1 +
#984300000000
0!
0'
#984310000000
1!
b10 %
1'
b10 +
#984320000000
0!
0'
#984330000000
1!
b11 %
1'
b11 +
#984340000000
0!
0'
#984350000000
1!
b100 %
1'
b100 +
#984360000000
0!
0'
#984370000000
1!
b101 %
1'
b101 +
#984380000000
0!
0'
#984390000000
1!
0$
b110 %
1'
0*
b110 +
#984400000000
0!
0'
#984410000000
1!
b111 %
1'
b111 +
#984420000000
0!
0'
#984430000000
1!
b1000 %
1'
b1000 +
#984440000000
0!
0'
#984450000000
1!
b1001 %
1'
b1001 +
#984460000000
0!
0'
#984470000000
1!
b0 %
1'
b0 +
#984480000000
1"
1(
#984490000000
0!
0"
b100 &
0'
0(
b100 ,
#984500000000
1!
1$
b1 %
1'
1*
b1 +
#984510000000
0!
0'
#984520000000
1!
b10 %
1'
b10 +
#984530000000
0!
0'
#984540000000
1!
b11 %
1'
b11 +
#984550000000
0!
0'
#984560000000
1!
b100 %
1'
b100 +
#984570000000
0!
0'
#984580000000
1!
b101 %
1'
b101 +
#984590000000
0!
0'
#984600000000
1!
b110 %
1'
b110 +
#984610000000
0!
0'
#984620000000
1!
b111 %
1'
b111 +
#984630000000
0!
0'
#984640000000
1!
0$
b1000 %
1'
0*
b1000 +
#984650000000
0!
0'
#984660000000
1!
b1001 %
1'
b1001 +
#984670000000
0!
0'
#984680000000
1!
b0 %
1'
b0 +
#984690000000
0!
0'
#984700000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#984710000000
0!
0'
#984720000000
1!
b10 %
1'
b10 +
#984730000000
0!
0'
#984740000000
1!
b11 %
1'
b11 +
#984750000000
0!
0'
#984760000000
1!
b100 %
1'
b100 +
#984770000000
0!
0'
#984780000000
1!
b101 %
1'
b101 +
#984790000000
0!
0'
#984800000000
1!
0$
b110 %
1'
0*
b110 +
#984810000000
0!
0'
#984820000000
1!
b111 %
1'
b111 +
#984830000000
0!
0'
#984840000000
1!
b1000 %
1'
b1000 +
#984850000000
0!
0'
#984860000000
1!
b1001 %
1'
b1001 +
#984870000000
0!
0'
#984880000000
1!
b0 %
1'
b0 +
#984890000000
0!
0'
#984900000000
1!
1$
b1 %
1'
1*
b1 +
#984910000000
1"
1(
#984920000000
0!
0"
b100 &
0'
0(
b100 ,
#984930000000
1!
b10 %
1'
b10 +
#984940000000
0!
0'
#984950000000
1!
b11 %
1'
b11 +
#984960000000
0!
0'
#984970000000
1!
b100 %
1'
b100 +
#984980000000
0!
0'
#984990000000
1!
b101 %
1'
b101 +
#985000000000
0!
0'
#985010000000
1!
b110 %
1'
b110 +
#985020000000
0!
0'
#985030000000
1!
b111 %
1'
b111 +
#985040000000
0!
0'
#985050000000
1!
0$
b1000 %
1'
0*
b1000 +
#985060000000
0!
0'
#985070000000
1!
b1001 %
1'
b1001 +
#985080000000
0!
0'
#985090000000
1!
b0 %
1'
b0 +
#985100000000
0!
0'
#985110000000
1!
1$
b1 %
1'
1*
b1 +
#985120000000
0!
0'
#985130000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#985140000000
0!
0'
#985150000000
1!
b11 %
1'
b11 +
#985160000000
0!
0'
#985170000000
1!
b100 %
1'
b100 +
#985180000000
0!
0'
#985190000000
1!
b101 %
1'
b101 +
#985200000000
0!
0'
#985210000000
1!
0$
b110 %
1'
0*
b110 +
#985220000000
0!
0'
#985230000000
1!
b111 %
1'
b111 +
#985240000000
0!
0'
#985250000000
1!
b1000 %
1'
b1000 +
#985260000000
0!
0'
#985270000000
1!
b1001 %
1'
b1001 +
#985280000000
0!
0'
#985290000000
1!
b0 %
1'
b0 +
#985300000000
0!
0'
#985310000000
1!
1$
b1 %
1'
1*
b1 +
#985320000000
0!
0'
#985330000000
1!
b10 %
1'
b10 +
#985340000000
1"
1(
#985350000000
0!
0"
b100 &
0'
0(
b100 ,
#985360000000
1!
b11 %
1'
b11 +
#985370000000
0!
0'
#985380000000
1!
b100 %
1'
b100 +
#985390000000
0!
0'
#985400000000
1!
b101 %
1'
b101 +
#985410000000
0!
0'
#985420000000
1!
b110 %
1'
b110 +
#985430000000
0!
0'
#985440000000
1!
b111 %
1'
b111 +
#985450000000
0!
0'
#985460000000
1!
0$
b1000 %
1'
0*
b1000 +
#985470000000
0!
0'
#985480000000
1!
b1001 %
1'
b1001 +
#985490000000
0!
0'
#985500000000
1!
b0 %
1'
b0 +
#985510000000
0!
0'
#985520000000
1!
1$
b1 %
1'
1*
b1 +
#985530000000
0!
0'
#985540000000
1!
b10 %
1'
b10 +
#985550000000
0!
0'
#985560000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#985570000000
0!
0'
#985580000000
1!
b100 %
1'
b100 +
#985590000000
0!
0'
#985600000000
1!
b101 %
1'
b101 +
#985610000000
0!
0'
#985620000000
1!
0$
b110 %
1'
0*
b110 +
#985630000000
0!
0'
#985640000000
1!
b111 %
1'
b111 +
#985650000000
0!
0'
#985660000000
1!
b1000 %
1'
b1000 +
#985670000000
0!
0'
#985680000000
1!
b1001 %
1'
b1001 +
#985690000000
0!
0'
#985700000000
1!
b0 %
1'
b0 +
#985710000000
0!
0'
#985720000000
1!
1$
b1 %
1'
1*
b1 +
#985730000000
0!
0'
#985740000000
1!
b10 %
1'
b10 +
#985750000000
0!
0'
#985760000000
1!
b11 %
1'
b11 +
#985770000000
1"
1(
#985780000000
0!
0"
b100 &
0'
0(
b100 ,
#985790000000
1!
b100 %
1'
b100 +
#985800000000
0!
0'
#985810000000
1!
b101 %
1'
b101 +
#985820000000
0!
0'
#985830000000
1!
b110 %
1'
b110 +
#985840000000
0!
0'
#985850000000
1!
b111 %
1'
b111 +
#985860000000
0!
0'
#985870000000
1!
0$
b1000 %
1'
0*
b1000 +
#985880000000
0!
0'
#985890000000
1!
b1001 %
1'
b1001 +
#985900000000
0!
0'
#985910000000
1!
b0 %
1'
b0 +
#985920000000
0!
0'
#985930000000
1!
1$
b1 %
1'
1*
b1 +
#985940000000
0!
0'
#985950000000
1!
b10 %
1'
b10 +
#985960000000
0!
0'
#985970000000
1!
b11 %
1'
b11 +
#985980000000
0!
0'
#985990000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#986000000000
0!
0'
#986010000000
1!
b101 %
1'
b101 +
#986020000000
0!
0'
#986030000000
1!
0$
b110 %
1'
0*
b110 +
#986040000000
0!
0'
#986050000000
1!
b111 %
1'
b111 +
#986060000000
0!
0'
#986070000000
1!
b1000 %
1'
b1000 +
#986080000000
0!
0'
#986090000000
1!
b1001 %
1'
b1001 +
#986100000000
0!
0'
#986110000000
1!
b0 %
1'
b0 +
#986120000000
0!
0'
#986130000000
1!
1$
b1 %
1'
1*
b1 +
#986140000000
0!
0'
#986150000000
1!
b10 %
1'
b10 +
#986160000000
0!
0'
#986170000000
1!
b11 %
1'
b11 +
#986180000000
0!
0'
#986190000000
1!
b100 %
1'
b100 +
#986200000000
1"
1(
#986210000000
0!
0"
b100 &
0'
0(
b100 ,
#986220000000
1!
b101 %
1'
b101 +
#986230000000
0!
0'
#986240000000
1!
b110 %
1'
b110 +
#986250000000
0!
0'
#986260000000
1!
b111 %
1'
b111 +
#986270000000
0!
0'
#986280000000
1!
0$
b1000 %
1'
0*
b1000 +
#986290000000
0!
0'
#986300000000
1!
b1001 %
1'
b1001 +
#986310000000
0!
0'
#986320000000
1!
b0 %
1'
b0 +
#986330000000
0!
0'
#986340000000
1!
1$
b1 %
1'
1*
b1 +
#986350000000
0!
0'
#986360000000
1!
b10 %
1'
b10 +
#986370000000
0!
0'
#986380000000
1!
b11 %
1'
b11 +
#986390000000
0!
0'
#986400000000
1!
b100 %
1'
b100 +
#986410000000
0!
0'
#986420000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#986430000000
0!
0'
#986440000000
1!
0$
b110 %
1'
0*
b110 +
#986450000000
0!
0'
#986460000000
1!
b111 %
1'
b111 +
#986470000000
0!
0'
#986480000000
1!
b1000 %
1'
b1000 +
#986490000000
0!
0'
#986500000000
1!
b1001 %
1'
b1001 +
#986510000000
0!
0'
#986520000000
1!
b0 %
1'
b0 +
#986530000000
0!
0'
#986540000000
1!
1$
b1 %
1'
1*
b1 +
#986550000000
0!
0'
#986560000000
1!
b10 %
1'
b10 +
#986570000000
0!
0'
#986580000000
1!
b11 %
1'
b11 +
#986590000000
0!
0'
#986600000000
1!
b100 %
1'
b100 +
#986610000000
0!
0'
#986620000000
1!
b101 %
1'
b101 +
#986630000000
1"
1(
#986640000000
0!
0"
b100 &
0'
0(
b100 ,
#986650000000
1!
b110 %
1'
b110 +
#986660000000
0!
0'
#986670000000
1!
b111 %
1'
b111 +
#986680000000
0!
0'
#986690000000
1!
0$
b1000 %
1'
0*
b1000 +
#986700000000
0!
0'
#986710000000
1!
b1001 %
1'
b1001 +
#986720000000
0!
0'
#986730000000
1!
b0 %
1'
b0 +
#986740000000
0!
0'
#986750000000
1!
1$
b1 %
1'
1*
b1 +
#986760000000
0!
0'
#986770000000
1!
b10 %
1'
b10 +
#986780000000
0!
0'
#986790000000
1!
b11 %
1'
b11 +
#986800000000
0!
0'
#986810000000
1!
b100 %
1'
b100 +
#986820000000
0!
0'
#986830000000
1!
b101 %
1'
b101 +
#986840000000
0!
0'
#986850000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#986860000000
0!
0'
#986870000000
1!
b111 %
1'
b111 +
#986880000000
0!
0'
#986890000000
1!
b1000 %
1'
b1000 +
#986900000000
0!
0'
#986910000000
1!
b1001 %
1'
b1001 +
#986920000000
0!
0'
#986930000000
1!
b0 %
1'
b0 +
#986940000000
0!
0'
#986950000000
1!
1$
b1 %
1'
1*
b1 +
#986960000000
0!
0'
#986970000000
1!
b10 %
1'
b10 +
#986980000000
0!
0'
#986990000000
1!
b11 %
1'
b11 +
#987000000000
0!
0'
#987010000000
1!
b100 %
1'
b100 +
#987020000000
0!
0'
#987030000000
1!
b101 %
1'
b101 +
#987040000000
0!
0'
#987050000000
1!
0$
b110 %
1'
0*
b110 +
#987060000000
1"
1(
#987070000000
0!
0"
b100 &
0'
0(
b100 ,
#987080000000
1!
1$
b111 %
1'
1*
b111 +
#987090000000
0!
0'
#987100000000
1!
0$
b1000 %
1'
0*
b1000 +
#987110000000
0!
0'
#987120000000
1!
b1001 %
1'
b1001 +
#987130000000
0!
0'
#987140000000
1!
b0 %
1'
b0 +
#987150000000
0!
0'
#987160000000
1!
1$
b1 %
1'
1*
b1 +
#987170000000
0!
0'
#987180000000
1!
b10 %
1'
b10 +
#987190000000
0!
0'
#987200000000
1!
b11 %
1'
b11 +
#987210000000
0!
0'
#987220000000
1!
b100 %
1'
b100 +
#987230000000
0!
0'
#987240000000
1!
b101 %
1'
b101 +
#987250000000
0!
0'
#987260000000
1!
b110 %
1'
b110 +
#987270000000
0!
0'
#987280000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#987290000000
0!
0'
#987300000000
1!
b1000 %
1'
b1000 +
#987310000000
0!
0'
#987320000000
1!
b1001 %
1'
b1001 +
#987330000000
0!
0'
#987340000000
1!
b0 %
1'
b0 +
#987350000000
0!
0'
#987360000000
1!
1$
b1 %
1'
1*
b1 +
#987370000000
0!
0'
#987380000000
1!
b10 %
1'
b10 +
#987390000000
0!
0'
#987400000000
1!
b11 %
1'
b11 +
#987410000000
0!
0'
#987420000000
1!
b100 %
1'
b100 +
#987430000000
0!
0'
#987440000000
1!
b101 %
1'
b101 +
#987450000000
0!
0'
#987460000000
1!
0$
b110 %
1'
0*
b110 +
#987470000000
0!
0'
#987480000000
1!
b111 %
1'
b111 +
#987490000000
1"
1(
#987500000000
0!
0"
b100 &
0'
0(
b100 ,
#987510000000
1!
b1000 %
1'
b1000 +
#987520000000
0!
0'
#987530000000
1!
b1001 %
1'
b1001 +
#987540000000
0!
0'
#987550000000
1!
b0 %
1'
b0 +
#987560000000
0!
0'
#987570000000
1!
1$
b1 %
1'
1*
b1 +
#987580000000
0!
0'
#987590000000
1!
b10 %
1'
b10 +
#987600000000
0!
0'
#987610000000
1!
b11 %
1'
b11 +
#987620000000
0!
0'
#987630000000
1!
b100 %
1'
b100 +
#987640000000
0!
0'
#987650000000
1!
b101 %
1'
b101 +
#987660000000
0!
0'
#987670000000
1!
b110 %
1'
b110 +
#987680000000
0!
0'
#987690000000
1!
b111 %
1'
b111 +
#987700000000
0!
0'
#987710000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#987720000000
0!
0'
#987730000000
1!
b1001 %
1'
b1001 +
#987740000000
0!
0'
#987750000000
1!
b0 %
1'
b0 +
#987760000000
0!
0'
#987770000000
1!
1$
b1 %
1'
1*
b1 +
#987780000000
0!
0'
#987790000000
1!
b10 %
1'
b10 +
#987800000000
0!
0'
#987810000000
1!
b11 %
1'
b11 +
#987820000000
0!
0'
#987830000000
1!
b100 %
1'
b100 +
#987840000000
0!
0'
#987850000000
1!
b101 %
1'
b101 +
#987860000000
0!
0'
#987870000000
1!
0$
b110 %
1'
0*
b110 +
#987880000000
0!
0'
#987890000000
1!
b111 %
1'
b111 +
#987900000000
0!
0'
#987910000000
1!
b1000 %
1'
b1000 +
#987920000000
1"
1(
#987930000000
0!
0"
b100 &
0'
0(
b100 ,
#987940000000
1!
b1001 %
1'
b1001 +
#987950000000
0!
0'
#987960000000
1!
b0 %
1'
b0 +
#987970000000
0!
0'
#987980000000
1!
1$
b1 %
1'
1*
b1 +
#987990000000
0!
0'
#988000000000
1!
b10 %
1'
b10 +
#988010000000
0!
0'
#988020000000
1!
b11 %
1'
b11 +
#988030000000
0!
0'
#988040000000
1!
b100 %
1'
b100 +
#988050000000
0!
0'
#988060000000
1!
b101 %
1'
b101 +
#988070000000
0!
0'
#988080000000
1!
b110 %
1'
b110 +
#988090000000
0!
0'
#988100000000
1!
b111 %
1'
b111 +
#988110000000
0!
0'
#988120000000
1!
0$
b1000 %
1'
0*
b1000 +
#988130000000
0!
0'
#988140000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#988150000000
0!
0'
#988160000000
1!
b0 %
1'
b0 +
#988170000000
0!
0'
#988180000000
1!
1$
b1 %
1'
1*
b1 +
#988190000000
0!
0'
#988200000000
1!
b10 %
1'
b10 +
#988210000000
0!
0'
#988220000000
1!
b11 %
1'
b11 +
#988230000000
0!
0'
#988240000000
1!
b100 %
1'
b100 +
#988250000000
0!
0'
#988260000000
1!
b101 %
1'
b101 +
#988270000000
0!
0'
#988280000000
1!
0$
b110 %
1'
0*
b110 +
#988290000000
0!
0'
#988300000000
1!
b111 %
1'
b111 +
#988310000000
0!
0'
#988320000000
1!
b1000 %
1'
b1000 +
#988330000000
0!
0'
#988340000000
1!
b1001 %
1'
b1001 +
#988350000000
1"
1(
#988360000000
0!
0"
b100 &
0'
0(
b100 ,
#988370000000
1!
b0 %
1'
b0 +
#988380000000
0!
0'
#988390000000
1!
1$
b1 %
1'
1*
b1 +
#988400000000
0!
0'
#988410000000
1!
b10 %
1'
b10 +
#988420000000
0!
0'
#988430000000
1!
b11 %
1'
b11 +
#988440000000
0!
0'
#988450000000
1!
b100 %
1'
b100 +
#988460000000
0!
0'
#988470000000
1!
b101 %
1'
b101 +
#988480000000
0!
0'
#988490000000
1!
b110 %
1'
b110 +
#988500000000
0!
0'
#988510000000
1!
b111 %
1'
b111 +
#988520000000
0!
0'
#988530000000
1!
0$
b1000 %
1'
0*
b1000 +
#988540000000
0!
0'
#988550000000
1!
b1001 %
1'
b1001 +
#988560000000
0!
0'
#988570000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#988580000000
0!
0'
#988590000000
1!
1$
b1 %
1'
1*
b1 +
#988600000000
0!
0'
#988610000000
1!
b10 %
1'
b10 +
#988620000000
0!
0'
#988630000000
1!
b11 %
1'
b11 +
#988640000000
0!
0'
#988650000000
1!
b100 %
1'
b100 +
#988660000000
0!
0'
#988670000000
1!
b101 %
1'
b101 +
#988680000000
0!
0'
#988690000000
1!
0$
b110 %
1'
0*
b110 +
#988700000000
0!
0'
#988710000000
1!
b111 %
1'
b111 +
#988720000000
0!
0'
#988730000000
1!
b1000 %
1'
b1000 +
#988740000000
0!
0'
#988750000000
1!
b1001 %
1'
b1001 +
#988760000000
0!
0'
#988770000000
1!
b0 %
1'
b0 +
#988780000000
1"
1(
#988790000000
0!
0"
b100 &
0'
0(
b100 ,
#988800000000
1!
1$
b1 %
1'
1*
b1 +
#988810000000
0!
0'
#988820000000
1!
b10 %
1'
b10 +
#988830000000
0!
0'
#988840000000
1!
b11 %
1'
b11 +
#988850000000
0!
0'
#988860000000
1!
b100 %
1'
b100 +
#988870000000
0!
0'
#988880000000
1!
b101 %
1'
b101 +
#988890000000
0!
0'
#988900000000
1!
b110 %
1'
b110 +
#988910000000
0!
0'
#988920000000
1!
b111 %
1'
b111 +
#988930000000
0!
0'
#988940000000
1!
0$
b1000 %
1'
0*
b1000 +
#988950000000
0!
0'
#988960000000
1!
b1001 %
1'
b1001 +
#988970000000
0!
0'
#988980000000
1!
b0 %
1'
b0 +
#988990000000
0!
0'
#989000000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#989010000000
0!
0'
#989020000000
1!
b10 %
1'
b10 +
#989030000000
0!
0'
#989040000000
1!
b11 %
1'
b11 +
#989050000000
0!
0'
#989060000000
1!
b100 %
1'
b100 +
#989070000000
0!
0'
#989080000000
1!
b101 %
1'
b101 +
#989090000000
0!
0'
#989100000000
1!
0$
b110 %
1'
0*
b110 +
#989110000000
0!
0'
#989120000000
1!
b111 %
1'
b111 +
#989130000000
0!
0'
#989140000000
1!
b1000 %
1'
b1000 +
#989150000000
0!
0'
#989160000000
1!
b1001 %
1'
b1001 +
#989170000000
0!
0'
#989180000000
1!
b0 %
1'
b0 +
#989190000000
0!
0'
#989200000000
1!
1$
b1 %
1'
1*
b1 +
#989210000000
1"
1(
#989220000000
0!
0"
b100 &
0'
0(
b100 ,
#989230000000
1!
b10 %
1'
b10 +
#989240000000
0!
0'
#989250000000
1!
b11 %
1'
b11 +
#989260000000
0!
0'
#989270000000
1!
b100 %
1'
b100 +
#989280000000
0!
0'
#989290000000
1!
b101 %
1'
b101 +
#989300000000
0!
0'
#989310000000
1!
b110 %
1'
b110 +
#989320000000
0!
0'
#989330000000
1!
b111 %
1'
b111 +
#989340000000
0!
0'
#989350000000
1!
0$
b1000 %
1'
0*
b1000 +
#989360000000
0!
0'
#989370000000
1!
b1001 %
1'
b1001 +
#989380000000
0!
0'
#989390000000
1!
b0 %
1'
b0 +
#989400000000
0!
0'
#989410000000
1!
1$
b1 %
1'
1*
b1 +
#989420000000
0!
0'
#989430000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#989440000000
0!
0'
#989450000000
1!
b11 %
1'
b11 +
#989460000000
0!
0'
#989470000000
1!
b100 %
1'
b100 +
#989480000000
0!
0'
#989490000000
1!
b101 %
1'
b101 +
#989500000000
0!
0'
#989510000000
1!
0$
b110 %
1'
0*
b110 +
#989520000000
0!
0'
#989530000000
1!
b111 %
1'
b111 +
#989540000000
0!
0'
#989550000000
1!
b1000 %
1'
b1000 +
#989560000000
0!
0'
#989570000000
1!
b1001 %
1'
b1001 +
#989580000000
0!
0'
#989590000000
1!
b0 %
1'
b0 +
#989600000000
0!
0'
#989610000000
1!
1$
b1 %
1'
1*
b1 +
#989620000000
0!
0'
#989630000000
1!
b10 %
1'
b10 +
#989640000000
1"
1(
#989650000000
0!
0"
b100 &
0'
0(
b100 ,
#989660000000
1!
b11 %
1'
b11 +
#989670000000
0!
0'
#989680000000
1!
b100 %
1'
b100 +
#989690000000
0!
0'
#989700000000
1!
b101 %
1'
b101 +
#989710000000
0!
0'
#989720000000
1!
b110 %
1'
b110 +
#989730000000
0!
0'
#989740000000
1!
b111 %
1'
b111 +
#989750000000
0!
0'
#989760000000
1!
0$
b1000 %
1'
0*
b1000 +
#989770000000
0!
0'
#989780000000
1!
b1001 %
1'
b1001 +
#989790000000
0!
0'
#989800000000
1!
b0 %
1'
b0 +
#989810000000
0!
0'
#989820000000
1!
1$
b1 %
1'
1*
b1 +
#989830000000
0!
0'
#989840000000
1!
b10 %
1'
b10 +
#989850000000
0!
0'
#989860000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#989870000000
0!
0'
#989880000000
1!
b100 %
1'
b100 +
#989890000000
0!
0'
#989900000000
1!
b101 %
1'
b101 +
#989910000000
0!
0'
#989920000000
1!
0$
b110 %
1'
0*
b110 +
#989930000000
0!
0'
#989940000000
1!
b111 %
1'
b111 +
#989950000000
0!
0'
#989960000000
1!
b1000 %
1'
b1000 +
#989970000000
0!
0'
#989980000000
1!
b1001 %
1'
b1001 +
#989990000000
0!
0'
#990000000000
1!
b0 %
1'
b0 +
#990010000000
0!
0'
#990020000000
1!
1$
b1 %
1'
1*
b1 +
#990030000000
0!
0'
#990040000000
1!
b10 %
1'
b10 +
#990050000000
0!
0'
#990060000000
1!
b11 %
1'
b11 +
#990070000000
1"
1(
#990080000000
0!
0"
b100 &
0'
0(
b100 ,
#990090000000
1!
b100 %
1'
b100 +
#990100000000
0!
0'
#990110000000
1!
b101 %
1'
b101 +
#990120000000
0!
0'
#990130000000
1!
b110 %
1'
b110 +
#990140000000
0!
0'
#990150000000
1!
b111 %
1'
b111 +
#990160000000
0!
0'
#990170000000
1!
0$
b1000 %
1'
0*
b1000 +
#990180000000
0!
0'
#990190000000
1!
b1001 %
1'
b1001 +
#990200000000
0!
0'
#990210000000
1!
b0 %
1'
b0 +
#990220000000
0!
0'
#990230000000
1!
1$
b1 %
1'
1*
b1 +
#990240000000
0!
0'
#990250000000
1!
b10 %
1'
b10 +
#990260000000
0!
0'
#990270000000
1!
b11 %
1'
b11 +
#990280000000
0!
0'
#990290000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#990300000000
0!
0'
#990310000000
1!
b101 %
1'
b101 +
#990320000000
0!
0'
#990330000000
1!
0$
b110 %
1'
0*
b110 +
#990340000000
0!
0'
#990350000000
1!
b111 %
1'
b111 +
#990360000000
0!
0'
#990370000000
1!
b1000 %
1'
b1000 +
#990380000000
0!
0'
#990390000000
1!
b1001 %
1'
b1001 +
#990400000000
0!
0'
#990410000000
1!
b0 %
1'
b0 +
#990420000000
0!
0'
#990430000000
1!
1$
b1 %
1'
1*
b1 +
#990440000000
0!
0'
#990450000000
1!
b10 %
1'
b10 +
#990460000000
0!
0'
#990470000000
1!
b11 %
1'
b11 +
#990480000000
0!
0'
#990490000000
1!
b100 %
1'
b100 +
#990500000000
1"
1(
#990510000000
0!
0"
b100 &
0'
0(
b100 ,
#990520000000
1!
b101 %
1'
b101 +
#990530000000
0!
0'
#990540000000
1!
b110 %
1'
b110 +
#990550000000
0!
0'
#990560000000
1!
b111 %
1'
b111 +
#990570000000
0!
0'
#990580000000
1!
0$
b1000 %
1'
0*
b1000 +
#990590000000
0!
0'
#990600000000
1!
b1001 %
1'
b1001 +
#990610000000
0!
0'
#990620000000
1!
b0 %
1'
b0 +
#990630000000
0!
0'
#990640000000
1!
1$
b1 %
1'
1*
b1 +
#990650000000
0!
0'
#990660000000
1!
b10 %
1'
b10 +
#990670000000
0!
0'
#990680000000
1!
b11 %
1'
b11 +
#990690000000
0!
0'
#990700000000
1!
b100 %
1'
b100 +
#990710000000
0!
0'
#990720000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#990730000000
0!
0'
#990740000000
1!
0$
b110 %
1'
0*
b110 +
#990750000000
0!
0'
#990760000000
1!
b111 %
1'
b111 +
#990770000000
0!
0'
#990780000000
1!
b1000 %
1'
b1000 +
#990790000000
0!
0'
#990800000000
1!
b1001 %
1'
b1001 +
#990810000000
0!
0'
#990820000000
1!
b0 %
1'
b0 +
#990830000000
0!
0'
#990840000000
1!
1$
b1 %
1'
1*
b1 +
#990850000000
0!
0'
#990860000000
1!
b10 %
1'
b10 +
#990870000000
0!
0'
#990880000000
1!
b11 %
1'
b11 +
#990890000000
0!
0'
#990900000000
1!
b100 %
1'
b100 +
#990910000000
0!
0'
#990920000000
1!
b101 %
1'
b101 +
#990930000000
1"
1(
#990940000000
0!
0"
b100 &
0'
0(
b100 ,
#990950000000
1!
b110 %
1'
b110 +
#990960000000
0!
0'
#990970000000
1!
b111 %
1'
b111 +
#990980000000
0!
0'
#990990000000
1!
0$
b1000 %
1'
0*
b1000 +
#991000000000
0!
0'
#991010000000
1!
b1001 %
1'
b1001 +
#991020000000
0!
0'
#991030000000
1!
b0 %
1'
b0 +
#991040000000
0!
0'
#991050000000
1!
1$
b1 %
1'
1*
b1 +
#991060000000
0!
0'
#991070000000
1!
b10 %
1'
b10 +
#991080000000
0!
0'
#991090000000
1!
b11 %
1'
b11 +
#991100000000
0!
0'
#991110000000
1!
b100 %
1'
b100 +
#991120000000
0!
0'
#991130000000
1!
b101 %
1'
b101 +
#991140000000
0!
0'
#991150000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#991160000000
0!
0'
#991170000000
1!
b111 %
1'
b111 +
#991180000000
0!
0'
#991190000000
1!
b1000 %
1'
b1000 +
#991200000000
0!
0'
#991210000000
1!
b1001 %
1'
b1001 +
#991220000000
0!
0'
#991230000000
1!
b0 %
1'
b0 +
#991240000000
0!
0'
#991250000000
1!
1$
b1 %
1'
1*
b1 +
#991260000000
0!
0'
#991270000000
1!
b10 %
1'
b10 +
#991280000000
0!
0'
#991290000000
1!
b11 %
1'
b11 +
#991300000000
0!
0'
#991310000000
1!
b100 %
1'
b100 +
#991320000000
0!
0'
#991330000000
1!
b101 %
1'
b101 +
#991340000000
0!
0'
#991350000000
1!
0$
b110 %
1'
0*
b110 +
#991360000000
1"
1(
#991370000000
0!
0"
b100 &
0'
0(
b100 ,
#991380000000
1!
1$
b111 %
1'
1*
b111 +
#991390000000
0!
0'
#991400000000
1!
0$
b1000 %
1'
0*
b1000 +
#991410000000
0!
0'
#991420000000
1!
b1001 %
1'
b1001 +
#991430000000
0!
0'
#991440000000
1!
b0 %
1'
b0 +
#991450000000
0!
0'
#991460000000
1!
1$
b1 %
1'
1*
b1 +
#991470000000
0!
0'
#991480000000
1!
b10 %
1'
b10 +
#991490000000
0!
0'
#991500000000
1!
b11 %
1'
b11 +
#991510000000
0!
0'
#991520000000
1!
b100 %
1'
b100 +
#991530000000
0!
0'
#991540000000
1!
b101 %
1'
b101 +
#991550000000
0!
0'
#991560000000
1!
b110 %
1'
b110 +
#991570000000
0!
0'
#991580000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#991590000000
0!
0'
#991600000000
1!
b1000 %
1'
b1000 +
#991610000000
0!
0'
#991620000000
1!
b1001 %
1'
b1001 +
#991630000000
0!
0'
#991640000000
1!
b0 %
1'
b0 +
#991650000000
0!
0'
#991660000000
1!
1$
b1 %
1'
1*
b1 +
#991670000000
0!
0'
#991680000000
1!
b10 %
1'
b10 +
#991690000000
0!
0'
#991700000000
1!
b11 %
1'
b11 +
#991710000000
0!
0'
#991720000000
1!
b100 %
1'
b100 +
#991730000000
0!
0'
#991740000000
1!
b101 %
1'
b101 +
#991750000000
0!
0'
#991760000000
1!
0$
b110 %
1'
0*
b110 +
#991770000000
0!
0'
#991780000000
1!
b111 %
1'
b111 +
#991790000000
1"
1(
#991800000000
0!
0"
b100 &
0'
0(
b100 ,
#991810000000
1!
b1000 %
1'
b1000 +
#991820000000
0!
0'
#991830000000
1!
b1001 %
1'
b1001 +
#991840000000
0!
0'
#991850000000
1!
b0 %
1'
b0 +
#991860000000
0!
0'
#991870000000
1!
1$
b1 %
1'
1*
b1 +
#991880000000
0!
0'
#991890000000
1!
b10 %
1'
b10 +
#991900000000
0!
0'
#991910000000
1!
b11 %
1'
b11 +
#991920000000
0!
0'
#991930000000
1!
b100 %
1'
b100 +
#991940000000
0!
0'
#991950000000
1!
b101 %
1'
b101 +
#991960000000
0!
0'
#991970000000
1!
b110 %
1'
b110 +
#991980000000
0!
0'
#991990000000
1!
b111 %
1'
b111 +
#992000000000
0!
0'
#992010000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#992020000000
0!
0'
#992030000000
1!
b1001 %
1'
b1001 +
#992040000000
0!
0'
#992050000000
1!
b0 %
1'
b0 +
#992060000000
0!
0'
#992070000000
1!
1$
b1 %
1'
1*
b1 +
#992080000000
0!
0'
#992090000000
1!
b10 %
1'
b10 +
#992100000000
0!
0'
#992110000000
1!
b11 %
1'
b11 +
#992120000000
0!
0'
#992130000000
1!
b100 %
1'
b100 +
#992140000000
0!
0'
#992150000000
1!
b101 %
1'
b101 +
#992160000000
0!
0'
#992170000000
1!
0$
b110 %
1'
0*
b110 +
#992180000000
0!
0'
#992190000000
1!
b111 %
1'
b111 +
#992200000000
0!
0'
#992210000000
1!
b1000 %
1'
b1000 +
#992220000000
1"
1(
#992230000000
0!
0"
b100 &
0'
0(
b100 ,
#992240000000
1!
b1001 %
1'
b1001 +
#992250000000
0!
0'
#992260000000
1!
b0 %
1'
b0 +
#992270000000
0!
0'
#992280000000
1!
1$
b1 %
1'
1*
b1 +
#992290000000
0!
0'
#992300000000
1!
b10 %
1'
b10 +
#992310000000
0!
0'
#992320000000
1!
b11 %
1'
b11 +
#992330000000
0!
0'
#992340000000
1!
b100 %
1'
b100 +
#992350000000
0!
0'
#992360000000
1!
b101 %
1'
b101 +
#992370000000
0!
0'
#992380000000
1!
b110 %
1'
b110 +
#992390000000
0!
0'
#992400000000
1!
b111 %
1'
b111 +
#992410000000
0!
0'
#992420000000
1!
0$
b1000 %
1'
0*
b1000 +
#992430000000
0!
0'
#992440000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#992450000000
0!
0'
#992460000000
1!
b0 %
1'
b0 +
#992470000000
0!
0'
#992480000000
1!
1$
b1 %
1'
1*
b1 +
#992490000000
0!
0'
#992500000000
1!
b10 %
1'
b10 +
#992510000000
0!
0'
#992520000000
1!
b11 %
1'
b11 +
#992530000000
0!
0'
#992540000000
1!
b100 %
1'
b100 +
#992550000000
0!
0'
#992560000000
1!
b101 %
1'
b101 +
#992570000000
0!
0'
#992580000000
1!
0$
b110 %
1'
0*
b110 +
#992590000000
0!
0'
#992600000000
1!
b111 %
1'
b111 +
#992610000000
0!
0'
#992620000000
1!
b1000 %
1'
b1000 +
#992630000000
0!
0'
#992640000000
1!
b1001 %
1'
b1001 +
#992650000000
1"
1(
#992660000000
0!
0"
b100 &
0'
0(
b100 ,
#992670000000
1!
b0 %
1'
b0 +
#992680000000
0!
0'
#992690000000
1!
1$
b1 %
1'
1*
b1 +
#992700000000
0!
0'
#992710000000
1!
b10 %
1'
b10 +
#992720000000
0!
0'
#992730000000
1!
b11 %
1'
b11 +
#992740000000
0!
0'
#992750000000
1!
b100 %
1'
b100 +
#992760000000
0!
0'
#992770000000
1!
b101 %
1'
b101 +
#992780000000
0!
0'
#992790000000
1!
b110 %
1'
b110 +
#992800000000
0!
0'
#992810000000
1!
b111 %
1'
b111 +
#992820000000
0!
0'
#992830000000
1!
0$
b1000 %
1'
0*
b1000 +
#992840000000
0!
0'
#992850000000
1!
b1001 %
1'
b1001 +
#992860000000
0!
0'
#992870000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#992880000000
0!
0'
#992890000000
1!
1$
b1 %
1'
1*
b1 +
#992900000000
0!
0'
#992910000000
1!
b10 %
1'
b10 +
#992920000000
0!
0'
#992930000000
1!
b11 %
1'
b11 +
#992940000000
0!
0'
#992950000000
1!
b100 %
1'
b100 +
#992960000000
0!
0'
#992970000000
1!
b101 %
1'
b101 +
#992980000000
0!
0'
#992990000000
1!
0$
b110 %
1'
0*
b110 +
#993000000000
0!
0'
#993010000000
1!
b111 %
1'
b111 +
#993020000000
0!
0'
#993030000000
1!
b1000 %
1'
b1000 +
#993040000000
0!
0'
#993050000000
1!
b1001 %
1'
b1001 +
#993060000000
0!
0'
#993070000000
1!
b0 %
1'
b0 +
#993080000000
1"
1(
#993090000000
0!
0"
b100 &
0'
0(
b100 ,
#993100000000
1!
1$
b1 %
1'
1*
b1 +
#993110000000
0!
0'
#993120000000
1!
b10 %
1'
b10 +
#993130000000
0!
0'
#993140000000
1!
b11 %
1'
b11 +
#993150000000
0!
0'
#993160000000
1!
b100 %
1'
b100 +
#993170000000
0!
0'
#993180000000
1!
b101 %
1'
b101 +
#993190000000
0!
0'
#993200000000
1!
b110 %
1'
b110 +
#993210000000
0!
0'
#993220000000
1!
b111 %
1'
b111 +
#993230000000
0!
0'
#993240000000
1!
0$
b1000 %
1'
0*
b1000 +
#993250000000
0!
0'
#993260000000
1!
b1001 %
1'
b1001 +
#993270000000
0!
0'
#993280000000
1!
b0 %
1'
b0 +
#993290000000
0!
0'
#993300000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#993310000000
0!
0'
#993320000000
1!
b10 %
1'
b10 +
#993330000000
0!
0'
#993340000000
1!
b11 %
1'
b11 +
#993350000000
0!
0'
#993360000000
1!
b100 %
1'
b100 +
#993370000000
0!
0'
#993380000000
1!
b101 %
1'
b101 +
#993390000000
0!
0'
#993400000000
1!
0$
b110 %
1'
0*
b110 +
#993410000000
0!
0'
#993420000000
1!
b111 %
1'
b111 +
#993430000000
0!
0'
#993440000000
1!
b1000 %
1'
b1000 +
#993450000000
0!
0'
#993460000000
1!
b1001 %
1'
b1001 +
#993470000000
0!
0'
#993480000000
1!
b0 %
1'
b0 +
#993490000000
0!
0'
#993500000000
1!
1$
b1 %
1'
1*
b1 +
#993510000000
1"
1(
#993520000000
0!
0"
b100 &
0'
0(
b100 ,
#993530000000
1!
b10 %
1'
b10 +
#993540000000
0!
0'
#993550000000
1!
b11 %
1'
b11 +
#993560000000
0!
0'
#993570000000
1!
b100 %
1'
b100 +
#993580000000
0!
0'
#993590000000
1!
b101 %
1'
b101 +
#993600000000
0!
0'
#993610000000
1!
b110 %
1'
b110 +
#993620000000
0!
0'
#993630000000
1!
b111 %
1'
b111 +
#993640000000
0!
0'
#993650000000
1!
0$
b1000 %
1'
0*
b1000 +
#993660000000
0!
0'
#993670000000
1!
b1001 %
1'
b1001 +
#993680000000
0!
0'
#993690000000
1!
b0 %
1'
b0 +
#993700000000
0!
0'
#993710000000
1!
1$
b1 %
1'
1*
b1 +
#993720000000
0!
0'
#993730000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#993740000000
0!
0'
#993750000000
1!
b11 %
1'
b11 +
#993760000000
0!
0'
#993770000000
1!
b100 %
1'
b100 +
#993780000000
0!
0'
#993790000000
1!
b101 %
1'
b101 +
#993800000000
0!
0'
#993810000000
1!
0$
b110 %
1'
0*
b110 +
#993820000000
0!
0'
#993830000000
1!
b111 %
1'
b111 +
#993840000000
0!
0'
#993850000000
1!
b1000 %
1'
b1000 +
#993860000000
0!
0'
#993870000000
1!
b1001 %
1'
b1001 +
#993880000000
0!
0'
#993890000000
1!
b0 %
1'
b0 +
#993900000000
0!
0'
#993910000000
1!
1$
b1 %
1'
1*
b1 +
#993920000000
0!
0'
#993930000000
1!
b10 %
1'
b10 +
#993940000000
1"
1(
#993950000000
0!
0"
b100 &
0'
0(
b100 ,
#993960000000
1!
b11 %
1'
b11 +
#993970000000
0!
0'
#993980000000
1!
b100 %
1'
b100 +
#993990000000
0!
0'
#994000000000
1!
b101 %
1'
b101 +
#994010000000
0!
0'
#994020000000
1!
b110 %
1'
b110 +
#994030000000
0!
0'
#994040000000
1!
b111 %
1'
b111 +
#994050000000
0!
0'
#994060000000
1!
0$
b1000 %
1'
0*
b1000 +
#994070000000
0!
0'
#994080000000
1!
b1001 %
1'
b1001 +
#994090000000
0!
0'
#994100000000
1!
b0 %
1'
b0 +
#994110000000
0!
0'
#994120000000
1!
1$
b1 %
1'
1*
b1 +
#994130000000
0!
0'
#994140000000
1!
b10 %
1'
b10 +
#994150000000
0!
0'
#994160000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#994170000000
0!
0'
#994180000000
1!
b100 %
1'
b100 +
#994190000000
0!
0'
#994200000000
1!
b101 %
1'
b101 +
#994210000000
0!
0'
#994220000000
1!
0$
b110 %
1'
0*
b110 +
#994230000000
0!
0'
#994240000000
1!
b111 %
1'
b111 +
#994250000000
0!
0'
#994260000000
1!
b1000 %
1'
b1000 +
#994270000000
0!
0'
#994280000000
1!
b1001 %
1'
b1001 +
#994290000000
0!
0'
#994300000000
1!
b0 %
1'
b0 +
#994310000000
0!
0'
#994320000000
1!
1$
b1 %
1'
1*
b1 +
#994330000000
0!
0'
#994340000000
1!
b10 %
1'
b10 +
#994350000000
0!
0'
#994360000000
1!
b11 %
1'
b11 +
#994370000000
1"
1(
#994380000000
0!
0"
b100 &
0'
0(
b100 ,
#994390000000
1!
b100 %
1'
b100 +
#994400000000
0!
0'
#994410000000
1!
b101 %
1'
b101 +
#994420000000
0!
0'
#994430000000
1!
b110 %
1'
b110 +
#994440000000
0!
0'
#994450000000
1!
b111 %
1'
b111 +
#994460000000
0!
0'
#994470000000
1!
0$
b1000 %
1'
0*
b1000 +
#994480000000
0!
0'
#994490000000
1!
b1001 %
1'
b1001 +
#994500000000
0!
0'
#994510000000
1!
b0 %
1'
b0 +
#994520000000
0!
0'
#994530000000
1!
1$
b1 %
1'
1*
b1 +
#994540000000
0!
0'
#994550000000
1!
b10 %
1'
b10 +
#994560000000
0!
0'
#994570000000
1!
b11 %
1'
b11 +
#994580000000
0!
0'
#994590000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#994600000000
0!
0'
#994610000000
1!
b101 %
1'
b101 +
#994620000000
0!
0'
#994630000000
1!
0$
b110 %
1'
0*
b110 +
#994640000000
0!
0'
#994650000000
1!
b111 %
1'
b111 +
#994660000000
0!
0'
#994670000000
1!
b1000 %
1'
b1000 +
#994680000000
0!
0'
#994690000000
1!
b1001 %
1'
b1001 +
#994700000000
0!
0'
#994710000000
1!
b0 %
1'
b0 +
#994720000000
0!
0'
#994730000000
1!
1$
b1 %
1'
1*
b1 +
#994740000000
0!
0'
#994750000000
1!
b10 %
1'
b10 +
#994760000000
0!
0'
#994770000000
1!
b11 %
1'
b11 +
#994780000000
0!
0'
#994790000000
1!
b100 %
1'
b100 +
#994800000000
1"
1(
#994810000000
0!
0"
b100 &
0'
0(
b100 ,
#994820000000
1!
b101 %
1'
b101 +
#994830000000
0!
0'
#994840000000
1!
b110 %
1'
b110 +
#994850000000
0!
0'
#994860000000
1!
b111 %
1'
b111 +
#994870000000
0!
0'
#994880000000
1!
0$
b1000 %
1'
0*
b1000 +
#994890000000
0!
0'
#994900000000
1!
b1001 %
1'
b1001 +
#994910000000
0!
0'
#994920000000
1!
b0 %
1'
b0 +
#994930000000
0!
0'
#994940000000
1!
1$
b1 %
1'
1*
b1 +
#994950000000
0!
0'
#994960000000
1!
b10 %
1'
b10 +
#994970000000
0!
0'
#994980000000
1!
b11 %
1'
b11 +
#994990000000
0!
0'
#995000000000
1!
b100 %
1'
b100 +
#995010000000
0!
0'
#995020000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#995030000000
0!
0'
#995040000000
1!
0$
b110 %
1'
0*
b110 +
#995050000000
0!
0'
#995060000000
1!
b111 %
1'
b111 +
#995070000000
0!
0'
#995080000000
1!
b1000 %
1'
b1000 +
#995090000000
0!
0'
#995100000000
1!
b1001 %
1'
b1001 +
#995110000000
0!
0'
#995120000000
1!
b0 %
1'
b0 +
#995130000000
0!
0'
#995140000000
1!
1$
b1 %
1'
1*
b1 +
#995150000000
0!
0'
#995160000000
1!
b10 %
1'
b10 +
#995170000000
0!
0'
#995180000000
1!
b11 %
1'
b11 +
#995190000000
0!
0'
#995200000000
1!
b100 %
1'
b100 +
#995210000000
0!
0'
#995220000000
1!
b101 %
1'
b101 +
#995230000000
1"
1(
#995240000000
0!
0"
b100 &
0'
0(
b100 ,
#995250000000
1!
b110 %
1'
b110 +
#995260000000
0!
0'
#995270000000
1!
b111 %
1'
b111 +
#995280000000
0!
0'
#995290000000
1!
0$
b1000 %
1'
0*
b1000 +
#995300000000
0!
0'
#995310000000
1!
b1001 %
1'
b1001 +
#995320000000
0!
0'
#995330000000
1!
b0 %
1'
b0 +
#995340000000
0!
0'
#995350000000
1!
1$
b1 %
1'
1*
b1 +
#995360000000
0!
0'
#995370000000
1!
b10 %
1'
b10 +
#995380000000
0!
0'
#995390000000
1!
b11 %
1'
b11 +
#995400000000
0!
0'
#995410000000
1!
b100 %
1'
b100 +
#995420000000
0!
0'
#995430000000
1!
b101 %
1'
b101 +
#995440000000
0!
0'
#995450000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#995460000000
0!
0'
#995470000000
1!
b111 %
1'
b111 +
#995480000000
0!
0'
#995490000000
1!
b1000 %
1'
b1000 +
#995500000000
0!
0'
#995510000000
1!
b1001 %
1'
b1001 +
#995520000000
0!
0'
#995530000000
1!
b0 %
1'
b0 +
#995540000000
0!
0'
#995550000000
1!
1$
b1 %
1'
1*
b1 +
#995560000000
0!
0'
#995570000000
1!
b10 %
1'
b10 +
#995580000000
0!
0'
#995590000000
1!
b11 %
1'
b11 +
#995600000000
0!
0'
#995610000000
1!
b100 %
1'
b100 +
#995620000000
0!
0'
#995630000000
1!
b101 %
1'
b101 +
#995640000000
0!
0'
#995650000000
1!
0$
b110 %
1'
0*
b110 +
#995660000000
1"
1(
#995670000000
0!
0"
b100 &
0'
0(
b100 ,
#995680000000
1!
1$
b111 %
1'
1*
b111 +
#995690000000
0!
0'
#995700000000
1!
0$
b1000 %
1'
0*
b1000 +
#995710000000
0!
0'
#995720000000
1!
b1001 %
1'
b1001 +
#995730000000
0!
0'
#995740000000
1!
b0 %
1'
b0 +
#995750000000
0!
0'
#995760000000
1!
1$
b1 %
1'
1*
b1 +
#995770000000
0!
0'
#995780000000
1!
b10 %
1'
b10 +
#995790000000
0!
0'
#995800000000
1!
b11 %
1'
b11 +
#995810000000
0!
0'
#995820000000
1!
b100 %
1'
b100 +
#995830000000
0!
0'
#995840000000
1!
b101 %
1'
b101 +
#995850000000
0!
0'
#995860000000
1!
b110 %
1'
b110 +
#995870000000
0!
0'
#995880000000
1!
0$
b111 %
b10 &
1'
0*
b111 +
b10 ,
#995890000000
0!
0'
#995900000000
1!
b1000 %
1'
b1000 +
#995910000000
0!
0'
#995920000000
1!
b1001 %
1'
b1001 +
#995930000000
0!
0'
#995940000000
1!
b0 %
1'
b0 +
#995950000000
0!
0'
#995960000000
1!
1$
b1 %
1'
1*
b1 +
#995970000000
0!
0'
#995980000000
1!
b10 %
1'
b10 +
#995990000000
0!
0'
#996000000000
1!
b11 %
1'
b11 +
#996010000000
0!
0'
#996020000000
1!
b100 %
1'
b100 +
#996030000000
0!
0'
#996040000000
1!
b101 %
1'
b101 +
#996050000000
0!
0'
#996060000000
1!
0$
b110 %
1'
0*
b110 +
#996070000000
0!
0'
#996080000000
1!
b111 %
1'
b111 +
#996090000000
1"
1(
#996100000000
0!
0"
b100 &
0'
0(
b100 ,
#996110000000
1!
b1000 %
1'
b1000 +
#996120000000
0!
0'
#996130000000
1!
b1001 %
1'
b1001 +
#996140000000
0!
0'
#996150000000
1!
b0 %
1'
b0 +
#996160000000
0!
0'
#996170000000
1!
1$
b1 %
1'
1*
b1 +
#996180000000
0!
0'
#996190000000
1!
b10 %
1'
b10 +
#996200000000
0!
0'
#996210000000
1!
b11 %
1'
b11 +
#996220000000
0!
0'
#996230000000
1!
b100 %
1'
b100 +
#996240000000
0!
0'
#996250000000
1!
b101 %
1'
b101 +
#996260000000
0!
0'
#996270000000
1!
b110 %
1'
b110 +
#996280000000
0!
0'
#996290000000
1!
b111 %
1'
b111 +
#996300000000
0!
0'
#996310000000
1!
0$
b1000 %
b10 &
1'
0*
b1000 +
b10 ,
#996320000000
0!
0'
#996330000000
1!
b1001 %
1'
b1001 +
#996340000000
0!
0'
#996350000000
1!
b0 %
1'
b0 +
#996360000000
0!
0'
#996370000000
1!
1$
b1 %
1'
1*
b1 +
#996380000000
0!
0'
#996390000000
1!
b10 %
1'
b10 +
#996400000000
0!
0'
#996410000000
1!
b11 %
1'
b11 +
#996420000000
0!
0'
#996430000000
1!
b100 %
1'
b100 +
#996440000000
0!
0'
#996450000000
1!
b101 %
1'
b101 +
#996460000000
0!
0'
#996470000000
1!
0$
b110 %
1'
0*
b110 +
#996480000000
0!
0'
#996490000000
1!
b111 %
1'
b111 +
#996500000000
0!
0'
#996510000000
1!
b1000 %
1'
b1000 +
#996520000000
1"
1(
#996530000000
0!
0"
b100 &
0'
0(
b100 ,
#996540000000
1!
b1001 %
1'
b1001 +
#996550000000
0!
0'
#996560000000
1!
b0 %
1'
b0 +
#996570000000
0!
0'
#996580000000
1!
1$
b1 %
1'
1*
b1 +
#996590000000
0!
0'
#996600000000
1!
b10 %
1'
b10 +
#996610000000
0!
0'
#996620000000
1!
b11 %
1'
b11 +
#996630000000
0!
0'
#996640000000
1!
b100 %
1'
b100 +
#996650000000
0!
0'
#996660000000
1!
b101 %
1'
b101 +
#996670000000
0!
0'
#996680000000
1!
b110 %
1'
b110 +
#996690000000
0!
0'
#996700000000
1!
b111 %
1'
b111 +
#996710000000
0!
0'
#996720000000
1!
0$
b1000 %
1'
0*
b1000 +
#996730000000
0!
0'
#996740000000
1!
b1001 %
b10 &
1'
b1001 +
b10 ,
#996750000000
0!
0'
#996760000000
1!
b0 %
1'
b0 +
#996770000000
0!
0'
#996780000000
1!
1$
b1 %
1'
1*
b1 +
#996790000000
0!
0'
#996800000000
1!
b10 %
1'
b10 +
#996810000000
0!
0'
#996820000000
1!
b11 %
1'
b11 +
#996830000000
0!
0'
#996840000000
1!
b100 %
1'
b100 +
#996850000000
0!
0'
#996860000000
1!
b101 %
1'
b101 +
#996870000000
0!
0'
#996880000000
1!
0$
b110 %
1'
0*
b110 +
#996890000000
0!
0'
#996900000000
1!
b111 %
1'
b111 +
#996910000000
0!
0'
#996920000000
1!
b1000 %
1'
b1000 +
#996930000000
0!
0'
#996940000000
1!
b1001 %
1'
b1001 +
#996950000000
1"
1(
#996960000000
0!
0"
b100 &
0'
0(
b100 ,
#996970000000
1!
b0 %
1'
b0 +
#996980000000
0!
0'
#996990000000
1!
1$
b1 %
1'
1*
b1 +
#997000000000
0!
0'
#997010000000
1!
b10 %
1'
b10 +
#997020000000
0!
0'
#997030000000
1!
b11 %
1'
b11 +
#997040000000
0!
0'
#997050000000
1!
b100 %
1'
b100 +
#997060000000
0!
0'
#997070000000
1!
b101 %
1'
b101 +
#997080000000
0!
0'
#997090000000
1!
b110 %
1'
b110 +
#997100000000
0!
0'
#997110000000
1!
b111 %
1'
b111 +
#997120000000
0!
0'
#997130000000
1!
0$
b1000 %
1'
0*
b1000 +
#997140000000
0!
0'
#997150000000
1!
b1001 %
1'
b1001 +
#997160000000
0!
0'
#997170000000
1!
b0 %
b10 &
1'
b0 +
b10 ,
#997180000000
0!
0'
#997190000000
1!
1$
b1 %
1'
1*
b1 +
#997200000000
0!
0'
#997210000000
1!
b10 %
1'
b10 +
#997220000000
0!
0'
#997230000000
1!
b11 %
1'
b11 +
#997240000000
0!
0'
#997250000000
1!
b100 %
1'
b100 +
#997260000000
0!
0'
#997270000000
1!
b101 %
1'
b101 +
#997280000000
0!
0'
#997290000000
1!
0$
b110 %
1'
0*
b110 +
#997300000000
0!
0'
#997310000000
1!
b111 %
1'
b111 +
#997320000000
0!
0'
#997330000000
1!
b1000 %
1'
b1000 +
#997340000000
0!
0'
#997350000000
1!
b1001 %
1'
b1001 +
#997360000000
0!
0'
#997370000000
1!
b0 %
1'
b0 +
#997380000000
1"
1(
#997390000000
0!
0"
b100 &
0'
0(
b100 ,
#997400000000
1!
1$
b1 %
1'
1*
b1 +
#997410000000
0!
0'
#997420000000
1!
b10 %
1'
b10 +
#997430000000
0!
0'
#997440000000
1!
b11 %
1'
b11 +
#997450000000
0!
0'
#997460000000
1!
b100 %
1'
b100 +
#997470000000
0!
0'
#997480000000
1!
b101 %
1'
b101 +
#997490000000
0!
0'
#997500000000
1!
b110 %
1'
b110 +
#997510000000
0!
0'
#997520000000
1!
b111 %
1'
b111 +
#997530000000
0!
0'
#997540000000
1!
0$
b1000 %
1'
0*
b1000 +
#997550000000
0!
0'
#997560000000
1!
b1001 %
1'
b1001 +
#997570000000
0!
0'
#997580000000
1!
b0 %
1'
b0 +
#997590000000
0!
0'
#997600000000
1!
1$
b1 %
b10 &
1'
1*
b1 +
b10 ,
#997610000000
0!
0'
#997620000000
1!
b10 %
1'
b10 +
#997630000000
0!
0'
#997640000000
1!
b11 %
1'
b11 +
#997650000000
0!
0'
#997660000000
1!
b100 %
1'
b100 +
#997670000000
0!
0'
#997680000000
1!
b101 %
1'
b101 +
#997690000000
0!
0'
#997700000000
1!
0$
b110 %
1'
0*
b110 +
#997710000000
0!
0'
#997720000000
1!
b111 %
1'
b111 +
#997730000000
0!
0'
#997740000000
1!
b1000 %
1'
b1000 +
#997750000000
0!
0'
#997760000000
1!
b1001 %
1'
b1001 +
#997770000000
0!
0'
#997780000000
1!
b0 %
1'
b0 +
#997790000000
0!
0'
#997800000000
1!
1$
b1 %
1'
1*
b1 +
#997810000000
1"
1(
#997820000000
0!
0"
b100 &
0'
0(
b100 ,
#997830000000
1!
b10 %
1'
b10 +
#997840000000
0!
0'
#997850000000
1!
b11 %
1'
b11 +
#997860000000
0!
0'
#997870000000
1!
b100 %
1'
b100 +
#997880000000
0!
0'
#997890000000
1!
b101 %
1'
b101 +
#997900000000
0!
0'
#997910000000
1!
b110 %
1'
b110 +
#997920000000
0!
0'
#997930000000
1!
b111 %
1'
b111 +
#997940000000
0!
0'
#997950000000
1!
0$
b1000 %
1'
0*
b1000 +
#997960000000
0!
0'
#997970000000
1!
b1001 %
1'
b1001 +
#997980000000
0!
0'
#997990000000
1!
b0 %
1'
b0 +
#998000000000
0!
0'
#998010000000
1!
1$
b1 %
1'
1*
b1 +
#998020000000
0!
0'
#998030000000
1!
b10 %
b10 &
1'
b10 +
b10 ,
#998040000000
0!
0'
#998050000000
1!
b11 %
1'
b11 +
#998060000000
0!
0'
#998070000000
1!
b100 %
1'
b100 +
#998080000000
0!
0'
#998090000000
1!
b101 %
1'
b101 +
#998100000000
0!
0'
#998110000000
1!
0$
b110 %
1'
0*
b110 +
#998120000000
0!
0'
#998130000000
1!
b111 %
1'
b111 +
#998140000000
0!
0'
#998150000000
1!
b1000 %
1'
b1000 +
#998160000000
0!
0'
#998170000000
1!
b1001 %
1'
b1001 +
#998180000000
0!
0'
#998190000000
1!
b0 %
1'
b0 +
#998200000000
0!
0'
#998210000000
1!
1$
b1 %
1'
1*
b1 +
#998220000000
0!
0'
#998230000000
1!
b10 %
1'
b10 +
#998240000000
1"
1(
#998250000000
0!
0"
b100 &
0'
0(
b100 ,
#998260000000
1!
b11 %
1'
b11 +
#998270000000
0!
0'
#998280000000
1!
b100 %
1'
b100 +
#998290000000
0!
0'
#998300000000
1!
b101 %
1'
b101 +
#998310000000
0!
0'
#998320000000
1!
b110 %
1'
b110 +
#998330000000
0!
0'
#998340000000
1!
b111 %
1'
b111 +
#998350000000
0!
0'
#998360000000
1!
0$
b1000 %
1'
0*
b1000 +
#998370000000
0!
0'
#998380000000
1!
b1001 %
1'
b1001 +
#998390000000
0!
0'
#998400000000
1!
b0 %
1'
b0 +
#998410000000
0!
0'
#998420000000
1!
1$
b1 %
1'
1*
b1 +
#998430000000
0!
0'
#998440000000
1!
b10 %
1'
b10 +
#998450000000
0!
0'
#998460000000
1!
b11 %
b10 &
1'
b11 +
b10 ,
#998470000000
0!
0'
#998480000000
1!
b100 %
1'
b100 +
#998490000000
0!
0'
#998500000000
1!
b101 %
1'
b101 +
#998510000000
0!
0'
#998520000000
1!
0$
b110 %
1'
0*
b110 +
#998530000000
0!
0'
#998540000000
1!
b111 %
1'
b111 +
#998550000000
0!
0'
#998560000000
1!
b1000 %
1'
b1000 +
#998570000000
0!
0'
#998580000000
1!
b1001 %
1'
b1001 +
#998590000000
0!
0'
#998600000000
1!
b0 %
1'
b0 +
#998610000000
0!
0'
#998620000000
1!
1$
b1 %
1'
1*
b1 +
#998630000000
0!
0'
#998640000000
1!
b10 %
1'
b10 +
#998650000000
0!
0'
#998660000000
1!
b11 %
1'
b11 +
#998670000000
1"
1(
#998680000000
0!
0"
b100 &
0'
0(
b100 ,
#998690000000
1!
b100 %
1'
b100 +
#998700000000
0!
0'
#998710000000
1!
b101 %
1'
b101 +
#998720000000
0!
0'
#998730000000
1!
b110 %
1'
b110 +
#998740000000
0!
0'
#998750000000
1!
b111 %
1'
b111 +
#998760000000
0!
0'
#998770000000
1!
0$
b1000 %
1'
0*
b1000 +
#998780000000
0!
0'
#998790000000
1!
b1001 %
1'
b1001 +
#998800000000
0!
0'
#998810000000
1!
b0 %
1'
b0 +
#998820000000
0!
0'
#998830000000
1!
1$
b1 %
1'
1*
b1 +
#998840000000
0!
0'
#998850000000
1!
b10 %
1'
b10 +
#998860000000
0!
0'
#998870000000
1!
b11 %
1'
b11 +
#998880000000
0!
0'
#998890000000
1!
b100 %
b10 &
1'
b100 +
b10 ,
#998900000000
0!
0'
#998910000000
1!
b101 %
1'
b101 +
#998920000000
0!
0'
#998930000000
1!
0$
b110 %
1'
0*
b110 +
#998940000000
0!
0'
#998950000000
1!
b111 %
1'
b111 +
#998960000000
0!
0'
#998970000000
1!
b1000 %
1'
b1000 +
#998980000000
0!
0'
#998990000000
1!
b1001 %
1'
b1001 +
#999000000000
0!
0'
#999010000000
1!
b0 %
1'
b0 +
#999020000000
0!
0'
#999030000000
1!
1$
b1 %
1'
1*
b1 +
#999040000000
0!
0'
#999050000000
1!
b10 %
1'
b10 +
#999060000000
0!
0'
#999070000000
1!
b11 %
1'
b11 +
#999080000000
0!
0'
#999090000000
1!
b100 %
1'
b100 +
#999100000000
1"
1(
#999110000000
0!
0"
b100 &
0'
0(
b100 ,
#999120000000
1!
b101 %
1'
b101 +
#999130000000
0!
0'
#999140000000
1!
b110 %
1'
b110 +
#999150000000
0!
0'
#999160000000
1!
b111 %
1'
b111 +
#999170000000
0!
0'
#999180000000
1!
0$
b1000 %
1'
0*
b1000 +
#999190000000
0!
0'
#999200000000
1!
b1001 %
1'
b1001 +
#999210000000
0!
0'
#999220000000
1!
b0 %
1'
b0 +
#999230000000
0!
0'
#999240000000
1!
1$
b1 %
1'
1*
b1 +
#999250000000
0!
0'
#999260000000
1!
b10 %
1'
b10 +
#999270000000
0!
0'
#999280000000
1!
b11 %
1'
b11 +
#999290000000
0!
0'
#999300000000
1!
b100 %
1'
b100 +
#999310000000
0!
0'
#999320000000
1!
b101 %
b10 &
1'
b101 +
b10 ,
#999330000000
0!
0'
#999340000000
1!
0$
b110 %
1'
0*
b110 +
#999350000000
0!
0'
#999360000000
1!
b111 %
1'
b111 +
#999370000000
0!
0'
#999380000000
1!
b1000 %
1'
b1000 +
#999390000000
0!
0'
#999400000000
1!
b1001 %
1'
b1001 +
#999410000000
0!
0'
#999420000000
1!
b0 %
1'
b0 +
#999430000000
0!
0'
#999440000000
1!
1$
b1 %
1'
1*
b1 +
#999450000000
0!
0'
#999460000000
1!
b10 %
1'
b10 +
#999470000000
0!
0'
#999480000000
1!
b11 %
1'
b11 +
#999490000000
0!
0'
#999500000000
1!
b100 %
1'
b100 +
#999510000000
0!
0'
#999520000000
1!
b101 %
1'
b101 +
#999530000000
1"
1(
#999540000000
0!
0"
b100 &
0'
0(
b100 ,
#999550000000
1!
b110 %
1'
b110 +
#999560000000
0!
0'
#999570000000
1!
b111 %
1'
b111 +
#999580000000
0!
0'
#999590000000
1!
0$
b1000 %
1'
0*
b1000 +
#999600000000
0!
0'
#999610000000
1!
b1001 %
1'
b1001 +
#999620000000
0!
0'
#999630000000
1!
b0 %
1'
b0 +
#999640000000
0!
0'
#999650000000
1!
1$
b1 %
1'
1*
b1 +
#999660000000
0!
0'
#999670000000
1!
b10 %
1'
b10 +
#999680000000
0!
0'
#999690000000
1!
b11 %
1'
b11 +
#999700000000
0!
0'
#999710000000
1!
b100 %
1'
b100 +
#999720000000
0!
0'
#999730000000
1!
b101 %
1'
b101 +
#999740000000
0!
0'
#999750000000
1!
0$
b110 %
b10 &
1'
0*
b110 +
b10 ,
#999760000000
0!
0'
#999770000000
1!
b111 %
1'
b111 +
#999780000000
0!
0'
#999790000000
1!
b1000 %
1'
b1000 +
#999800000000
0!
0'
#999810000000
1!
b1001 %
1'
b1001 +
#999820000000
0!
0'
#999830000000
1!
b0 %
1'
b0 +
#999840000000
0!
0'
#999850000000
1!
1$
b1 %
1'
1*
b1 +
#999860000000
0!
0'
#999870000000
1!
b10 %
1'
b10 +
#999880000000
0!
0'
#999890000000
1!
b11 %
1'
b11 +
#999900000000
0!
0'
#999910000000
1!
b100 %
1'
b100 +
#999920000000
0!
0'
#999930000000
1!
b101 %
1'
b101 +
#999940000000
0!
0'
#999950000000
1!
0$
b110 %
1'
0*
b110 +
#999960000000
1"
1(
#999970000000
0!
0"
b100 &
0'
0(
b100 ,
#999980000000
1!
1$
b111 %
1'
1*
b111 +
#999990000000
0!
0'
#1000000000000
1!
0$
b1000 %
1'
0*
b1000 +
