$date
  Sat Apr 27 21:01:20 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_tp2_3 $end
$var reg 1 ! clk $end
$var reg 1 " reset $end
$var reg 4 # enable_disp[3:0] $end
$var reg 7 $ segmentos[6:0] $end
$scope module uut $end
$var reg 1 % clk $end
$var reg 1 & reset $end
$var reg 4 ' enable_disp[3:0] $end
$var reg 7 ( segmentos[6:0] $end
$comment state is not handled $end
$var reg 4 ) bcd[3:0] $end
$var integer 32 * cuenta $end
$var reg 1 + debounced_reset $end
$var reg 1 , enable_conta $end
$scope module a $end
$var reg 1 - clk $end
$var reg 1 . key $end
$var reg 1 / debounced_key $end
$var reg 1 0 key_stable $end
$var reg 1 1 last_key $end
$upscope $end
$scope module b $end
$var reg 1 2 clk $end
$var reg 1 3 reset $end
$var reg 1 4 enable $end
$var reg 1 5 cout $end
$var integer 32 6 q $end
$upscope $end
$scope module d0 $end
$var reg 7 7 segmentos[6:0] $end
$var reg 4 8 bcd[3:0] $end
$var reg 1 9 enable $end
$upscope $end
$scope module d1 $end
$var reg 7 : segmentos[6:0] $end
$var reg 4 ; bcd[3:0] $end
$var reg 1 < enable $end
$upscope $end
$scope module d2 $end
$var reg 7 = segmentos[6:0] $end
$var reg 4 > bcd[3:0] $end
$var reg 1 ? enable $end
$upscope $end
$scope module d3 $end
$var reg 7 @ segmentos[6:0] $end
$var reg 4 A bcd[3:0] $end
$var reg 1 B enable $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
U"
b1XXX #
b0110000 $
0%
U&
b1XXX '
b0110000 (
b0001 )
b0 *
U+
1,
0-
U.
U/
U0
U1
02
U3
14
U5
b0 6
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#10000000
1!
1%
1-
12
05
#20000000
0!
0%
b1 *
0-
02
b1 6
#30000000
1!
1%
1-
12
#40000000
0!
0%
b10 *
0-
02
b10 6
#50000000
1!
1%
1-
12
#60000000
0!
0%
b11 *
0-
02
b11 6
#70000000
1!
1%
1-
12
15
#80000000
0!
0%
b100 *
0-
02
b100 6
#90000000
1!
1%
1-
12
#100000000
0!
0%
b101 *
0-
02
b101 6
#110000000
1!
1"
1%
1&
1+
1-
1.
1/
10
11
12
13
#120000000
0!
0%
b110 *
0-
02
b110 6
#130000000
1!
1%
1-
12
05
#140000000
0!
0%
b0 *
0-
02
b0 6
#150000000
1!
1%
1-
12
#160000000
0!
0"
0%
0&
0-
0.
02
#170000000
1!
1%
0+
1-
0/
00
01
12
03
#180000000
0!
0%
0-
02
#190000000
1!
1%
1-
12
#200000000
0!
0%
b1 *
0-
02
b1 6
#210000000
1!
1%
1-
12
#220000000
0!
0%
b10 *
0-
02
b10 6
#230000000
1!
1%
1-
12
#240000000
0!
0%
b11 *
0-
02
b11 6
#250000000
1!
1%
1-
12
15
#260000000
0!
0%
b100 *
0-
02
b100 6
#270000000
1!
1%
1-
12
#280000000
0!
0%
b101 *
0-
02
b101 6
#290000000
1!
1%
1-
12
#300000000
0!
0%
b110 *
0-
02
b110 6
#310000000
1!
1%
1-
12
#320000000
0!
0%
b111 *
0-
02
b111 6
#330000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#340000000
0!
0%
b0 *
0-
02
b0 6
#350000000
1!
1%
1-
12
#360000000
0!
0%
b1 *
0-
02
b1 6
#370000000
1!
1%
1-
12
#380000000
0!
0%
b10 *
0-
02
b10 6
#390000000
1!
1%
1-
12
#400000000
0!
0%
b11 *
0-
02
b11 6
#410000000
1!
1%
1-
12
15
#420000000
0!
0%
b100 *
0-
02
b100 6
#430000000
1!
1%
1-
12
#440000000
0!
0%
b101 *
0-
02
b101 6
#450000000
1!
1%
1-
12
#460000000
0!
0%
b110 *
0-
02
b110 6
#470000000
1!
1%
1-
12
#480000000
0!
0%
b111 *
0-
02
b111 6
#490000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#500000000
0!
0%
b0 *
0-
02
b0 6
#510000000
1!
1%
1-
12
#520000000
0!
0%
b1 *
0-
02
b1 6
#530000000
1!
1%
1-
12
#540000000
0!
0%
b10 *
0-
02
b10 6
#550000000
1!
1%
1-
12
#560000000
0!
0%
b11 *
0-
02
b11 6
#570000000
1!
1%
1-
12
15
#580000000
0!
0%
b100 *
0-
02
b100 6
#590000000
1!
1%
1-
12
#600000000
0!
0%
b101 *
0-
02
b101 6
#610000000
1!
1%
1-
12
#620000000
0!
0%
b110 *
0-
02
b110 6
#630000000
1!
1%
1-
12
#640000000
0!
0%
b111 *
0-
02
b111 6
#650000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#660000000
0!
0%
b0 *
0-
02
b0 6
#670000000
1!
1%
1-
12
#680000000
0!
0%
b1 *
0-
02
b1 6
#690000000
1!
1%
1-
12
#700000000
0!
0%
b10 *
0-
02
b10 6
#710000000
1!
1%
1-
12
#720000000
0!
0%
b11 *
0-
02
b11 6
#730000000
1!
1%
1-
12
15
#740000000
0!
0%
b100 *
0-
02
b100 6
#750000000
1!
1%
1-
12
#760000000
0!
0%
b101 *
0-
02
b101 6
#770000000
1!
1%
1-
12
#780000000
0!
0%
b110 *
0-
02
b110 6
#790000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#800000000
0!
0%
b111 *
0-
02
b111 6
#810000000
1!
1%
1-
12
05
#820000000
0!
0%
b0 *
0-
02
b0 6
#830000000
1!
1%
1-
12
#840000000
0!
0"
0%
0&
0-
0.
02
#850000000
1!
1%
0+
1-
0/
00
01
12
03
#860000000
0!
0%
0-
02
#870000000
1!
1%
1-
12
#880000000
0!
0%
b1 *
0-
02
b1 6
#890000000
1!
1%
1-
12
#900000000
0!
0%
b10 *
0-
02
b10 6
#910000000
1!
1%
1-
12
#920000000
0!
0%
b11 *
0-
02
b11 6
#930000000
1!
1%
1-
12
15
#940000000
0!
0%
b100 *
0-
02
b100 6
#950000000
1!
1%
1-
12
#960000000
0!
0%
b101 *
0-
02
b101 6
#970000000
1!
1%
1-
12
#980000000
0!
0%
b110 *
0-
02
b110 6
#990000000
1!
1%
1-
12
#1000000000
0!
0%
b111 *
0-
02
b111 6
#1010000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#1020000000
0!
0%
b0 *
0-
02
b0 6
#1030000000
1!
1%
1-
12
#1040000000
0!
0%
b1 *
0-
02
b1 6
#1050000000
1!
1%
1-
12
#1060000000
0!
0%
b10 *
0-
02
b10 6
#1070000000
1!
1%
1-
12
#1080000000
0!
0%
b11 *
0-
02
b11 6
#1090000000
1!
1%
1-
12
15
#1100000000
0!
0%
b100 *
0-
02
b100 6
#1110000000
1!
1%
1-
12
#1120000000
0!
0%
b101 *
0-
02
b101 6
#1130000000
1!
1%
1-
12
#1140000000
0!
0%
b110 *
0-
02
b110 6
#1150000000
1!
1%
1-
12
#1160000000
0!
0%
b111 *
0-
02
b111 6
#1170000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#1180000000
0!
0%
b0 *
0-
02
b0 6
#1190000000
1!
1%
1-
12
#1200000000
0!
0%
b1 *
0-
02
b1 6
#1210000000
1!
1%
1-
12
#1220000000
0!
0%
b10 *
0-
02
b10 6
#1230000000
1!
1%
1-
12
#1240000000
0!
0%
b11 *
0-
02
b11 6
#1250000000
1!
1%
1-
12
15
#1260000000
0!
0%
b100 *
0-
02
b100 6
#1270000000
1!
1%
1-
12
#1280000000
0!
0%
b101 *
0-
02
b101 6
#1290000000
1!
1%
1-
12
#1300000000
0!
0%
b110 *
0-
02
b110 6
#1310000000
1!
1%
1-
12
#1320000000
0!
0%
b111 *
0-
02
b111 6
#1330000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#1340000000
0!
0%
b0 *
0-
02
b0 6
#1350000000
1!
1%
1-
12
#1360000000
0!
0%
b1 *
0-
02
b1 6
#1370000000
1!
1%
1-
12
#1380000000
0!
0%
b10 *
0-
02
b10 6
#1390000000
1!
1%
1-
12
#1400000000
0!
0%
b11 *
0-
02
b11 6
#1410000000
1!
1%
1-
12
15
#1420000000
0!
0%
b100 *
0-
02
b100 6
#1430000000
1!
1%
1-
12
#1440000000
0!
0%
b101 *
0-
02
b101 6
#1450000000
1!
1%
1-
12
#1460000000
0!
0%
b110 *
0-
02
b110 6
#1470000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#1480000000
0!
0%
b111 *
0-
02
b111 6
#1490000000
1!
1%
1-
12
05
#1500000000
0!
0%
b0 *
0-
02
b0 6
#1510000000
1!
1%
1-
12
#1520000000
0!
0"
0%
0&
0-
0.
02
#1530000000
1!
1%
0+
1-
0/
00
01
12
03
#1540000000
0!
0%
0-
02
#1550000000
1!
1%
1-
12
#1560000000
0!
0%
b1 *
0-
02
b1 6
#1570000000
1!
1%
1-
12
#1580000000
0!
0%
b10 *
0-
02
b10 6
#1590000000
1!
1%
1-
12
#1600000000
0!
0%
b11 *
0-
02
b11 6
#1610000000
1!
1%
1-
12
15
#1620000000
0!
0%
b100 *
0-
02
b100 6
#1630000000
1!
1%
1-
12
#1640000000
0!
0%
b101 *
0-
02
b101 6
#1650000000
1!
1%
1-
12
#1660000000
0!
0%
b110 *
0-
02
b110 6
#1670000000
1!
1%
1-
12
#1680000000
0!
0%
b111 *
0-
02
b111 6
#1690000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#1700000000
0!
0%
b0 *
0-
02
b0 6
#1710000000
1!
1%
1-
12
#1720000000
0!
0%
b1 *
0-
02
b1 6
#1730000000
1!
1%
1-
12
#1740000000
0!
0%
b10 *
0-
02
b10 6
#1750000000
1!
1%
1-
12
#1760000000
0!
0%
b11 *
0-
02
b11 6
#1770000000
1!
1%
1-
12
15
#1780000000
0!
0%
b100 *
0-
02
b100 6
#1790000000
1!
1%
1-
12
#1800000000
0!
0%
b101 *
0-
02
b101 6
#1810000000
1!
1%
1-
12
#1820000000
0!
0%
b110 *
0-
02
b110 6
#1830000000
1!
1%
1-
12
#1840000000
0!
0%
b111 *
0-
02
b111 6
#1850000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#1860000000
0!
0%
b0 *
0-
02
b0 6
#1870000000
1!
1%
1-
12
#1880000000
0!
0%
b1 *
0-
02
b1 6
#1890000000
1!
1%
1-
12
#1900000000
0!
0%
b10 *
0-
02
b10 6
#1910000000
1!
1%
1-
12
#1920000000
0!
0%
b11 *
0-
02
b11 6
#1930000000
1!
1%
1-
12
15
#1940000000
0!
0%
b100 *
0-
02
b100 6
#1950000000
1!
1%
1-
12
#1960000000
0!
0%
b101 *
0-
02
b101 6
#1970000000
1!
1%
1-
12
#1980000000
0!
0%
b110 *
0-
02
b110 6
#1990000000
1!
1%
1-
12
#2000000000
0!
0%
b111 *
0-
02
b111 6
#2010000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#2020000000
0!
0%
b0 *
0-
02
b0 6
#2030000000
1!
1%
1-
12
#2040000000
0!
0%
b1 *
0-
02
b1 6
#2050000000
1!
1%
1-
12
#2060000000
0!
0%
b10 *
0-
02
b10 6
#2070000000
1!
1%
1-
12
#2080000000
0!
0%
b11 *
0-
02
b11 6
#2090000000
1!
1%
1-
12
15
#2100000000
0!
0%
b100 *
0-
02
b100 6
#2110000000
1!
1%
1-
12
#2120000000
0!
0%
b101 *
0-
02
b101 6
#2130000000
1!
1%
1-
12
#2140000000
0!
0%
b110 *
0-
02
b110 6
#2150000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#2160000000
0!
0%
b111 *
0-
02
b111 6
#2170000000
1!
1%
1-
12
05
#2180000000
0!
0%
b0 *
0-
02
b0 6
#2190000000
1!
1%
1-
12
#2200000000
0!
0"
0%
0&
0-
0.
02
#2210000000
1!
1%
0+
1-
0/
00
01
12
03
#2220000000
0!
0%
0-
02
#2230000000
1!
1%
1-
12
#2240000000
0!
0%
b1 *
0-
02
b1 6
#2250000000
1!
1%
1-
12
#2260000000
0!
0%
b10 *
0-
02
b10 6
#2270000000
1!
1%
1-
12
#2280000000
0!
0%
b11 *
0-
02
b11 6
#2290000000
1!
1%
1-
12
15
#2300000000
0!
0%
b100 *
0-
02
b100 6
#2310000000
1!
1%
1-
12
#2320000000
0!
0%
b101 *
0-
02
b101 6
#2330000000
1!
1%
1-
12
#2340000000
0!
0%
b110 *
0-
02
b110 6
#2350000000
1!
1%
1-
12
#2360000000
0!
0%
b111 *
0-
02
b111 6
#2370000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#2380000000
0!
0%
b0 *
0-
02
b0 6
#2390000000
1!
1%
1-
12
#2400000000
0!
0%
b1 *
0-
02
b1 6
#2410000000
1!
1%
1-
12
#2420000000
0!
0%
b10 *
0-
02
b10 6
#2430000000
1!
1%
1-
12
#2440000000
0!
0%
b11 *
0-
02
b11 6
#2450000000
1!
1%
1-
12
15
#2460000000
0!
0%
b100 *
0-
02
b100 6
#2470000000
1!
1%
1-
12
#2480000000
0!
0%
b101 *
0-
02
b101 6
#2490000000
1!
1%
1-
12
#2500000000
0!
0%
b110 *
0-
02
b110 6
#2510000000
1!
1%
1-
12
#2520000000
0!
0%
b111 *
0-
02
b111 6
#2530000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#2540000000
0!
0%
b0 *
0-
02
b0 6
#2550000000
1!
1%
1-
12
#2560000000
0!
0%
b1 *
0-
02
b1 6
#2570000000
1!
1%
1-
12
#2580000000
0!
0%
b10 *
0-
02
b10 6
#2590000000
1!
1%
1-
12
#2600000000
0!
0%
b11 *
0-
02
b11 6
#2610000000
1!
1%
1-
12
15
#2620000000
0!
0%
b100 *
0-
02
b100 6
#2630000000
1!
1%
1-
12
#2640000000
0!
0%
b101 *
0-
02
b101 6
#2650000000
1!
1%
1-
12
#2660000000
0!
0%
b110 *
0-
02
b110 6
#2670000000
1!
1%
1-
12
#2680000000
0!
0%
b111 *
0-
02
b111 6
#2690000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#2700000000
0!
0%
b0 *
0-
02
b0 6
#2710000000
1!
1%
1-
12
#2720000000
0!
0%
b1 *
0-
02
b1 6
#2730000000
1!
1%
1-
12
#2740000000
0!
0%
b10 *
0-
02
b10 6
#2750000000
1!
1%
1-
12
#2760000000
0!
0%
b11 *
0-
02
b11 6
#2770000000
1!
1%
1-
12
15
#2780000000
0!
0%
b100 *
0-
02
b100 6
#2790000000
1!
1%
1-
12
#2800000000
0!
0%
b101 *
0-
02
b101 6
#2810000000
1!
1%
1-
12
#2820000000
0!
0%
b110 *
0-
02
b110 6
#2830000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#2840000000
0!
0%
b111 *
0-
02
b111 6
#2850000000
1!
1%
1-
12
05
#2860000000
0!
0%
b0 *
0-
02
b0 6
#2870000000
1!
1%
1-
12
#2880000000
0!
0"
0%
0&
0-
0.
02
#2890000000
1!
1%
0+
1-
0/
00
01
12
03
#2900000000
0!
0%
0-
02
#2910000000
1!
1%
1-
12
#2920000000
0!
0%
b1 *
0-
02
b1 6
#2930000000
1!
1%
1-
12
#2940000000
0!
0%
b10 *
0-
02
b10 6
#2950000000
1!
1%
1-
12
#2960000000
0!
0%
b11 *
0-
02
b11 6
#2970000000
1!
1%
1-
12
15
#2980000000
0!
0%
b100 *
0-
02
b100 6
#2990000000
1!
1%
1-
12
#3000000000
0!
0%
b101 *
0-
02
b101 6
#3010000000
1!
1%
1-
12
#3020000000
0!
0%
b110 *
0-
02
b110 6
#3030000000
1!
1%
1-
12
#3040000000
0!
0%
b111 *
0-
02
b111 6
#3050000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#3060000000
0!
0%
b0 *
0-
02
b0 6
#3070000000
1!
1%
1-
12
#3080000000
0!
0%
b1 *
0-
02
b1 6
#3090000000
1!
1%
1-
12
#3100000000
0!
0%
b10 *
0-
02
b10 6
#3110000000
1!
1%
1-
12
#3120000000
0!
0%
b11 *
0-
02
b11 6
#3130000000
1!
1%
1-
12
15
#3140000000
0!
0%
b100 *
0-
02
b100 6
#3150000000
1!
1%
1-
12
#3160000000
0!
0%
b101 *
0-
02
b101 6
#3170000000
1!
1%
1-
12
#3180000000
0!
0%
b110 *
0-
02
b110 6
#3190000000
1!
1%
1-
12
#3200000000
0!
0%
b111 *
0-
02
b111 6
#3210000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#3220000000
0!
0%
b0 *
0-
02
b0 6
#3230000000
1!
1%
1-
12
#3240000000
0!
0%
b1 *
0-
02
b1 6
#3250000000
1!
1%
1-
12
#3260000000
0!
0%
b10 *
0-
02
b10 6
#3270000000
1!
1%
1-
12
#3280000000
0!
0%
b11 *
0-
02
b11 6
#3290000000
1!
1%
1-
12
15
#3300000000
0!
0%
b100 *
0-
02
b100 6
#3310000000
1!
1%
1-
12
#3320000000
0!
0%
b101 *
0-
02
b101 6
#3330000000
1!
1%
1-
12
#3340000000
0!
0%
b110 *
0-
02
b110 6
#3350000000
1!
1%
1-
12
#3360000000
0!
0%
b111 *
0-
02
b111 6
#3370000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#3380000000
0!
0%
b0 *
0-
02
b0 6
#3390000000
1!
1%
1-
12
#3400000000
0!
0%
b1 *
0-
02
b1 6
#3410000000
1!
1%
1-
12
#3420000000
0!
0%
b10 *
0-
02
b10 6
#3430000000
1!
1%
1-
12
#3440000000
0!
0%
b11 *
0-
02
b11 6
#3450000000
1!
1%
1-
12
15
#3460000000
0!
0%
b100 *
0-
02
b100 6
#3470000000
1!
1%
1-
12
#3480000000
0!
0%
b101 *
0-
02
b101 6
#3490000000
1!
1%
1-
12
#3500000000
0!
0%
b110 *
0-
02
b110 6
#3510000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#3520000000
0!
0%
b111 *
0-
02
b111 6
#3530000000
1!
1%
1-
12
05
#3540000000
0!
0%
b0 *
0-
02
b0 6
#3550000000
1!
1%
1-
12
#3560000000
0!
0"
0%
0&
0-
0.
02
#3570000000
1!
1%
0+
1-
0/
00
01
12
03
#3580000000
0!
0%
0-
02
#3590000000
1!
1%
1-
12
#3600000000
0!
0%
b1 *
0-
02
b1 6
#3610000000
1!
1%
1-
12
#3620000000
0!
0%
b10 *
0-
02
b10 6
#3630000000
1!
1%
1-
12
#3640000000
0!
0%
b11 *
0-
02
b11 6
#3650000000
1!
1%
1-
12
15
#3660000000
0!
0%
b100 *
0-
02
b100 6
#3670000000
1!
1%
1-
12
#3680000000
0!
0%
b101 *
0-
02
b101 6
#3690000000
1!
1%
1-
12
#3700000000
0!
0%
b110 *
0-
02
b110 6
#3710000000
1!
1%
1-
12
#3720000000
0!
0%
b111 *
0-
02
b111 6
#3730000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#3740000000
0!
0%
b0 *
0-
02
b0 6
#3750000000
1!
1%
1-
12
#3760000000
0!
0%
b1 *
0-
02
b1 6
#3770000000
1!
1%
1-
12
#3780000000
0!
0%
b10 *
0-
02
b10 6
#3790000000
1!
1%
1-
12
#3800000000
0!
0%
b11 *
0-
02
b11 6
#3810000000
1!
1%
1-
12
15
#3820000000
0!
0%
b100 *
0-
02
b100 6
#3830000000
1!
1%
1-
12
#3840000000
0!
0%
b101 *
0-
02
b101 6
#3850000000
1!
1%
1-
12
#3860000000
0!
0%
b110 *
0-
02
b110 6
#3870000000
1!
1%
1-
12
#3880000000
0!
0%
b111 *
0-
02
b111 6
#3890000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#3900000000
0!
0%
b0 *
0-
02
b0 6
#3910000000
1!
1%
1-
12
#3920000000
0!
0%
b1 *
0-
02
b1 6
#3930000000
1!
1%
1-
12
#3940000000
0!
0%
b10 *
0-
02
b10 6
#3950000000
1!
1%
1-
12
#3960000000
0!
0%
b11 *
0-
02
b11 6
#3970000000
1!
1%
1-
12
15
#3980000000
0!
0%
b100 *
0-
02
b100 6
#3990000000
1!
1%
1-
12
#4000000000
0!
0%
b101 *
0-
02
b101 6
#4010000000
1!
1%
1-
12
#4020000000
0!
0%
b110 *
0-
02
b110 6
#4030000000
1!
1%
1-
12
#4040000000
0!
0%
b111 *
0-
02
b111 6
#4050000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#4060000000
0!
0%
b0 *
0-
02
b0 6
#4070000000
1!
1%
1-
12
#4080000000
0!
0%
b1 *
0-
02
b1 6
#4090000000
1!
1%
1-
12
#4100000000
0!
0%
b10 *
0-
02
b10 6
#4110000000
1!
1%
1-
12
#4120000000
0!
0%
b11 *
0-
02
b11 6
#4130000000
1!
1%
1-
12
15
#4140000000
0!
0%
b100 *
0-
02
b100 6
#4150000000
1!
1%
1-
12
#4160000000
0!
0%
b101 *
0-
02
b101 6
#4170000000
1!
1%
1-
12
#4180000000
0!
0%
b110 *
0-
02
b110 6
#4190000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#4200000000
0!
0%
b111 *
0-
02
b111 6
#4210000000
1!
1%
1-
12
05
#4220000000
0!
0%
b0 *
0-
02
b0 6
#4230000000
1!
1%
1-
12
#4240000000
0!
0"
0%
0&
0-
0.
02
#4250000000
1!
1%
0+
1-
0/
00
01
12
03
#4260000000
0!
0%
0-
02
#4270000000
1!
1%
1-
12
#4280000000
0!
0%
b1 *
0-
02
b1 6
#4290000000
1!
1%
1-
12
#4300000000
0!
0%
b10 *
0-
02
b10 6
#4310000000
1!
1%
1-
12
#4320000000
0!
0%
b11 *
0-
02
b11 6
#4330000000
1!
1%
1-
12
15
#4340000000
0!
0%
b100 *
0-
02
b100 6
#4350000000
1!
1%
1-
12
#4360000000
0!
0%
b101 *
0-
02
b101 6
#4370000000
1!
1%
1-
12
#4380000000
0!
0%
b110 *
0-
02
b110 6
#4390000000
1!
1%
1-
12
#4400000000
0!
0%
b111 *
0-
02
b111 6
#4410000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#4420000000
0!
0%
b0 *
0-
02
b0 6
#4430000000
1!
1%
1-
12
#4440000000
0!
0%
b1 *
0-
02
b1 6
#4450000000
1!
1%
1-
12
#4460000000
0!
0%
b10 *
0-
02
b10 6
#4470000000
1!
1%
1-
12
#4480000000
0!
0%
b11 *
0-
02
b11 6
#4490000000
1!
1%
1-
12
15
#4500000000
0!
0%
b100 *
0-
02
b100 6
#4510000000
1!
1%
1-
12
#4520000000
0!
0%
b101 *
0-
02
b101 6
#4530000000
1!
1%
1-
12
#4540000000
0!
0%
b110 *
0-
02
b110 6
#4550000000
1!
1%
1-
12
#4560000000
0!
0%
b111 *
0-
02
b111 6
#4570000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#4580000000
0!
0%
b0 *
0-
02
b0 6
#4590000000
1!
1%
1-
12
#4600000000
0!
0%
b1 *
0-
02
b1 6
#4610000000
1!
1%
1-
12
#4620000000
0!
0%
b10 *
0-
02
b10 6
#4630000000
1!
1%
1-
12
#4640000000
0!
0%
b11 *
0-
02
b11 6
#4650000000
1!
1%
1-
12
15
#4660000000
0!
0%
b100 *
0-
02
b100 6
#4670000000
1!
1%
1-
12
#4680000000
0!
0%
b101 *
0-
02
b101 6
#4690000000
1!
1%
1-
12
#4700000000
0!
0%
b110 *
0-
02
b110 6
#4710000000
1!
1%
1-
12
#4720000000
0!
0%
b111 *
0-
02
b111 6
#4730000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#4740000000
0!
0%
b0 *
0-
02
b0 6
#4750000000
1!
1%
1-
12
#4760000000
0!
0%
b1 *
0-
02
b1 6
#4770000000
1!
1%
1-
12
#4780000000
0!
0%
b10 *
0-
02
b10 6
#4790000000
1!
1%
1-
12
#4800000000
0!
0%
b11 *
0-
02
b11 6
#4810000000
1!
1%
1-
12
15
#4820000000
0!
0%
b100 *
0-
02
b100 6
#4830000000
1!
1%
1-
12
#4840000000
0!
0%
b101 *
0-
02
b101 6
#4850000000
1!
1%
1-
12
#4860000000
0!
0%
b110 *
0-
02
b110 6
#4870000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#4880000000
0!
0%
b111 *
0-
02
b111 6
#4890000000
1!
1%
1-
12
05
#4900000000
0!
0%
b0 *
0-
02
b0 6
#4910000000
1!
1%
1-
12
#4920000000
0!
0"
0%
0&
0-
0.
02
#4930000000
1!
1%
0+
1-
0/
00
01
12
03
#4940000000
0!
0%
0-
02
#4950000000
1!
1%
1-
12
#4960000000
0!
0%
b1 *
0-
02
b1 6
#4970000000
1!
1%
1-
12
#4980000000
0!
0%
b10 *
0-
02
b10 6
#4990000000
1!
1%
1-
12
#5000000000
0!
0%
b11 *
0-
02
b11 6
#5010000000
1!
1%
1-
12
15
#5020000000
0!
0%
b100 *
0-
02
b100 6
#5030000000
1!
1%
1-
12
#5040000000
0!
0%
b101 *
0-
02
b101 6
#5050000000
1!
1%
1-
12
#5060000000
0!
0%
b110 *
0-
02
b110 6
#5070000000
1!
1%
1-
12
#5080000000
0!
0%
b111 *
0-
02
b111 6
#5090000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#5100000000
0!
0%
b0 *
0-
02
b0 6
#5110000000
1!
1%
1-
12
#5120000000
0!
0%
b1 *
0-
02
b1 6
#5130000000
1!
1%
1-
12
#5140000000
0!
0%
b10 *
0-
02
b10 6
#5150000000
1!
1%
1-
12
#5160000000
0!
0%
b11 *
0-
02
b11 6
#5170000000
1!
1%
1-
12
15
#5180000000
0!
0%
b100 *
0-
02
b100 6
#5190000000
1!
1%
1-
12
#5200000000
0!
0%
b101 *
0-
02
b101 6
#5210000000
1!
1%
1-
12
#5220000000
0!
0%
b110 *
0-
02
b110 6
#5230000000
1!
1%
1-
12
#5240000000
0!
0%
b111 *
0-
02
b111 6
#5250000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#5260000000
0!
0%
b0 *
0-
02
b0 6
#5270000000
1!
1%
1-
12
#5280000000
0!
0%
b1 *
0-
02
b1 6
#5290000000
1!
1%
1-
12
#5300000000
0!
0%
b10 *
0-
02
b10 6
#5310000000
1!
1%
1-
12
#5320000000
0!
0%
b11 *
0-
02
b11 6
#5330000000
1!
1%
1-
12
15
#5340000000
0!
0%
b100 *
0-
02
b100 6
#5350000000
1!
1%
1-
12
#5360000000
0!
0%
b101 *
0-
02
b101 6
#5370000000
1!
1%
1-
12
#5380000000
0!
0%
b110 *
0-
02
b110 6
#5390000000
1!
1%
1-
12
#5400000000
0!
0%
b111 *
0-
02
b111 6
#5410000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#5420000000
0!
0%
b0 *
0-
02
b0 6
#5430000000
1!
1%
1-
12
#5440000000
0!
0%
b1 *
0-
02
b1 6
#5450000000
1!
1%
1-
12
#5460000000
0!
0%
b10 *
0-
02
b10 6
#5470000000
1!
1%
1-
12
#5480000000
0!
0%
b11 *
0-
02
b11 6
#5490000000
1!
1%
1-
12
15
#5500000000
0!
0%
b100 *
0-
02
b100 6
#5510000000
1!
1%
1-
12
#5520000000
0!
0%
b101 *
0-
02
b101 6
#5530000000
1!
1%
1-
12
#5540000000
0!
0%
b110 *
0-
02
b110 6
#5550000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#5560000000
0!
0%
b111 *
0-
02
b111 6
#5570000000
1!
1%
1-
12
05
#5580000000
0!
0%
b0 *
0-
02
b0 6
#5590000000
1!
1%
1-
12
#5600000000
0!
0"
0%
0&
0-
0.
02
#5610000000
1!
1%
0+
1-
0/
00
01
12
03
#5620000000
0!
0%
0-
02
#5630000000
1!
1%
1-
12
#5640000000
0!
0%
b1 *
0-
02
b1 6
#5650000000
1!
1%
1-
12
#5660000000
0!
0%
b10 *
0-
02
b10 6
#5670000000
1!
1%
1-
12
#5680000000
0!
0%
b11 *
0-
02
b11 6
#5690000000
1!
1%
1-
12
15
#5700000000
0!
0%
b100 *
0-
02
b100 6
#5710000000
1!
1%
1-
12
#5720000000
0!
0%
b101 *
0-
02
b101 6
#5730000000
1!
1%
1-
12
#5740000000
0!
0%
b110 *
0-
02
b110 6
#5750000000
1!
1%
1-
12
#5760000000
0!
0%
b111 *
0-
02
b111 6
#5770000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#5780000000
0!
0%
b0 *
0-
02
b0 6
#5790000000
1!
1%
1-
12
#5800000000
0!
0%
b1 *
0-
02
b1 6
#5810000000
1!
1%
1-
12
#5820000000
0!
0%
b10 *
0-
02
b10 6
#5830000000
1!
1%
1-
12
#5840000000
0!
0%
b11 *
0-
02
b11 6
#5850000000
1!
1%
1-
12
15
#5860000000
0!
0%
b100 *
0-
02
b100 6
#5870000000
1!
1%
1-
12
#5880000000
0!
0%
b101 *
0-
02
b101 6
#5890000000
1!
1%
1-
12
#5900000000
0!
0%
b110 *
0-
02
b110 6
#5910000000
1!
1%
1-
12
#5920000000
0!
0%
b111 *
0-
02
b111 6
#5930000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#5940000000
0!
0%
b0 *
0-
02
b0 6
#5950000000
1!
1%
1-
12
#5960000000
0!
0%
b1 *
0-
02
b1 6
#5970000000
1!
1%
1-
12
#5980000000
0!
0%
b10 *
0-
02
b10 6
#5990000000
1!
1%
1-
12
#6000000000
0!
0%
b11 *
0-
02
b11 6
#6010000000
1!
1%
1-
12
15
#6020000000
0!
0%
b100 *
0-
02
b100 6
#6030000000
1!
1%
1-
12
#6040000000
0!
0%
b101 *
0-
02
b101 6
#6050000000
1!
1%
1-
12
#6060000000
0!
0%
b110 *
0-
02
b110 6
#6070000000
1!
1%
1-
12
#6080000000
0!
0%
b111 *
0-
02
b111 6
#6090000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#6100000000
0!
0%
b0 *
0-
02
b0 6
#6110000000
1!
1%
1-
12
#6120000000
0!
0%
b1 *
0-
02
b1 6
#6130000000
1!
1%
1-
12
#6140000000
0!
0%
b10 *
0-
02
b10 6
#6150000000
1!
1%
1-
12
#6160000000
0!
0%
b11 *
0-
02
b11 6
#6170000000
1!
1%
1-
12
15
#6180000000
0!
0%
b100 *
0-
02
b100 6
#6190000000
1!
1%
1-
12
#6200000000
0!
0%
b101 *
0-
02
b101 6
#6210000000
1!
1%
1-
12
#6220000000
0!
0%
b110 *
0-
02
b110 6
#6230000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#6240000000
0!
0%
b111 *
0-
02
b111 6
#6250000000
1!
1%
1-
12
05
#6260000000
0!
0%
b0 *
0-
02
b0 6
#6270000000
1!
1%
1-
12
#6280000000
0!
0"
0%
0&
0-
0.
02
#6290000000
1!
1%
0+
1-
0/
00
01
12
03
#6300000000
0!
0%
0-
02
#6310000000
1!
1%
1-
12
#6320000000
0!
0%
b1 *
0-
02
b1 6
#6330000000
1!
1%
1-
12
#6340000000
0!
0%
b10 *
0-
02
b10 6
#6350000000
1!
1%
1-
12
#6360000000
0!
0%
b11 *
0-
02
b11 6
#6370000000
1!
1%
1-
12
15
#6380000000
0!
0%
b100 *
0-
02
b100 6
#6390000000
1!
1%
1-
12
#6400000000
0!
0%
b101 *
0-
02
b101 6
#6410000000
1!
1%
1-
12
#6420000000
0!
0%
b110 *
0-
02
b110 6
#6430000000
1!
1%
1-
12
#6440000000
0!
0%
b111 *
0-
02
b111 6
#6450000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#6460000000
0!
0%
b0 *
0-
02
b0 6
#6470000000
1!
1%
1-
12
#6480000000
0!
0%
b1 *
0-
02
b1 6
#6490000000
1!
1%
1-
12
#6500000000
0!
0%
b10 *
0-
02
b10 6
#6510000000
1!
1%
1-
12
#6520000000
0!
0%
b11 *
0-
02
b11 6
#6530000000
1!
1%
1-
12
15
#6540000000
0!
0%
b100 *
0-
02
b100 6
#6550000000
1!
1%
1-
12
#6560000000
0!
0%
b101 *
0-
02
b101 6
#6570000000
1!
1%
1-
12
#6580000000
0!
0%
b110 *
0-
02
b110 6
#6590000000
1!
1%
1-
12
#6600000000
0!
0%
b111 *
0-
02
b111 6
#6610000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#6620000000
0!
0%
b0 *
0-
02
b0 6
#6630000000
1!
1%
1-
12
#6640000000
0!
0%
b1 *
0-
02
b1 6
#6650000000
1!
1%
1-
12
#6660000000
0!
0%
b10 *
0-
02
b10 6
#6670000000
1!
1%
1-
12
#6680000000
0!
0%
b11 *
0-
02
b11 6
#6690000000
1!
1%
1-
12
15
#6700000000
0!
0%
b100 *
0-
02
b100 6
#6710000000
1!
1%
1-
12
#6720000000
0!
0%
b101 *
0-
02
b101 6
#6730000000
1!
1%
1-
12
#6740000000
0!
0%
b110 *
0-
02
b110 6
#6750000000
1!
1%
1-
12
#6760000000
0!
0%
b111 *
0-
02
b111 6
#6770000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#6780000000
0!
0%
b0 *
0-
02
b0 6
#6790000000
1!
1%
1-
12
#6800000000
0!
0%
b1 *
0-
02
b1 6
#6810000000
1!
1%
1-
12
#6820000000
0!
0%
b10 *
0-
02
b10 6
#6830000000
1!
1%
1-
12
#6840000000
0!
0%
b11 *
0-
02
b11 6
#6850000000
1!
1%
1-
12
15
#6860000000
0!
0%
b100 *
0-
02
b100 6
#6870000000
1!
1%
1-
12
#6880000000
0!
0%
b101 *
0-
02
b101 6
#6890000000
1!
1%
1-
12
#6900000000
0!
0%
b110 *
0-
02
b110 6
#6910000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#6920000000
0!
0%
b111 *
0-
02
b111 6
#6930000000
1!
1%
1-
12
05
#6940000000
0!
0%
b0 *
0-
02
b0 6
#6950000000
1!
1%
1-
12
#6960000000
0!
0"
0%
0&
0-
0.
02
#6970000000
1!
1%
0+
1-
0/
00
01
12
03
#6980000000
0!
0%
0-
02
#6990000000
1!
1%
1-
12
#7000000000
0!
0%
b1 *
0-
02
b1 6
#7010000000
1!
1%
1-
12
#7020000000
0!
0%
b10 *
0-
02
b10 6
#7030000000
1!
1%
1-
12
#7040000000
0!
0%
b11 *
0-
02
b11 6
#7050000000
1!
1%
1-
12
15
#7060000000
0!
0%
b100 *
0-
02
b100 6
#7070000000
1!
1%
1-
12
#7080000000
0!
0%
b101 *
0-
02
b101 6
#7090000000
1!
1%
1-
12
#7100000000
0!
0%
b110 *
0-
02
b110 6
#7110000000
1!
1%
1-
12
#7120000000
0!
0%
b111 *
0-
02
b111 6
#7130000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#7140000000
0!
0%
b0 *
0-
02
b0 6
#7150000000
1!
1%
1-
12
#7160000000
0!
0%
b1 *
0-
02
b1 6
#7170000000
1!
1%
1-
12
#7180000000
0!
0%
b10 *
0-
02
b10 6
#7190000000
1!
1%
1-
12
#7200000000
0!
0%
b11 *
0-
02
b11 6
#7210000000
1!
1%
1-
12
15
#7220000000
0!
0%
b100 *
0-
02
b100 6
#7230000000
1!
1%
1-
12
#7240000000
0!
0%
b101 *
0-
02
b101 6
#7250000000
1!
1%
1-
12
#7260000000
0!
0%
b110 *
0-
02
b110 6
#7270000000
1!
1%
1-
12
#7280000000
0!
0%
b111 *
0-
02
b111 6
#7290000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#7300000000
0!
0%
b0 *
0-
02
b0 6
#7310000000
1!
1%
1-
12
#7320000000
0!
0%
b1 *
0-
02
b1 6
#7330000000
1!
1%
1-
12
#7340000000
0!
0%
b10 *
0-
02
b10 6
#7350000000
1!
1%
1-
12
#7360000000
0!
0%
b11 *
0-
02
b11 6
#7370000000
1!
1%
1-
12
15
#7380000000
0!
0%
b100 *
0-
02
b100 6
#7390000000
1!
1%
1-
12
#7400000000
0!
0%
b101 *
0-
02
b101 6
#7410000000
1!
1%
1-
12
#7420000000
0!
0%
b110 *
0-
02
b110 6
#7430000000
1!
1%
1-
12
#7440000000
0!
0%
b111 *
0-
02
b111 6
#7450000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#7460000000
0!
0%
b0 *
0-
02
b0 6
#7470000000
1!
1%
1-
12
#7480000000
0!
0%
b1 *
0-
02
b1 6
#7490000000
1!
1%
1-
12
#7500000000
0!
0%
b10 *
0-
02
b10 6
#7510000000
1!
1%
1-
12
#7520000000
0!
0%
b11 *
0-
02
b11 6
#7530000000
1!
1%
1-
12
15
#7540000000
0!
0%
b100 *
0-
02
b100 6
#7550000000
1!
1%
1-
12
#7560000000
0!
0%
b101 *
0-
02
b101 6
#7570000000
1!
1%
1-
12
#7580000000
0!
0%
b110 *
0-
02
b110 6
#7590000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#7600000000
0!
0%
b111 *
0-
02
b111 6
#7610000000
1!
1%
1-
12
05
#7620000000
0!
0%
b0 *
0-
02
b0 6
#7630000000
1!
1%
1-
12
#7640000000
0!
0"
0%
0&
0-
0.
02
#7650000000
1!
1%
0+
1-
0/
00
01
12
03
#7660000000
0!
0%
0-
02
#7670000000
1!
1%
1-
12
#7680000000
0!
0%
b1 *
0-
02
b1 6
#7690000000
1!
1%
1-
12
#7700000000
0!
0%
b10 *
0-
02
b10 6
#7710000000
1!
1%
1-
12
#7720000000
0!
0%
b11 *
0-
02
b11 6
#7730000000
1!
1%
1-
12
15
#7740000000
0!
0%
b100 *
0-
02
b100 6
#7750000000
1!
1%
1-
12
#7760000000
0!
0%
b101 *
0-
02
b101 6
#7770000000
1!
1%
1-
12
#7780000000
0!
0%
b110 *
0-
02
b110 6
#7790000000
1!
1%
1-
12
#7800000000
0!
0%
b111 *
0-
02
b111 6
#7810000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#7820000000
0!
0%
b0 *
0-
02
b0 6
#7830000000
1!
1%
1-
12
#7840000000
0!
0%
b1 *
0-
02
b1 6
#7850000000
1!
1%
1-
12
#7860000000
0!
0%
b10 *
0-
02
b10 6
#7870000000
1!
1%
1-
12
#7880000000
0!
0%
b11 *
0-
02
b11 6
#7890000000
1!
1%
1-
12
15
#7900000000
0!
0%
b100 *
0-
02
b100 6
#7910000000
1!
1%
1-
12
#7920000000
0!
0%
b101 *
0-
02
b101 6
#7930000000
1!
1%
1-
12
#7940000000
0!
0%
b110 *
0-
02
b110 6
#7950000000
1!
1%
1-
12
#7960000000
0!
0%
b111 *
0-
02
b111 6
#7970000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#7980000000
0!
0%
b0 *
0-
02
b0 6
#7990000000
1!
1%
1-
12
#8000000000
0!
0%
b1 *
0-
02
b1 6
#8010000000
1!
1%
1-
12
#8020000000
0!
0%
b10 *
0-
02
b10 6
#8030000000
1!
1%
1-
12
#8040000000
0!
0%
b11 *
0-
02
b11 6
#8050000000
1!
1%
1-
12
15
#8060000000
0!
0%
b100 *
0-
02
b100 6
#8070000000
1!
1%
1-
12
#8080000000
0!
0%
b101 *
0-
02
b101 6
#8090000000
1!
1%
1-
12
#8100000000
0!
0%
b110 *
0-
02
b110 6
#8110000000
1!
1%
1-
12
#8120000000
0!
0%
b111 *
0-
02
b111 6
#8130000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#8140000000
0!
0%
b0 *
0-
02
b0 6
#8150000000
1!
1%
1-
12
#8160000000
0!
0%
b1 *
0-
02
b1 6
#8170000000
1!
1%
1-
12
#8180000000
0!
0%
b10 *
0-
02
b10 6
#8190000000
1!
1%
1-
12
#8200000000
0!
0%
b11 *
0-
02
b11 6
#8210000000
1!
1%
1-
12
15
#8220000000
0!
0%
b100 *
0-
02
b100 6
#8230000000
1!
1%
1-
12
#8240000000
0!
0%
b101 *
0-
02
b101 6
#8250000000
1!
1%
1-
12
#8260000000
0!
0%
b110 *
0-
02
b110 6
#8270000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#8280000000
0!
0%
b111 *
0-
02
b111 6
#8290000000
1!
1%
1-
12
05
#8300000000
0!
0%
b0 *
0-
02
b0 6
#8310000000
1!
1%
1-
12
#8320000000
0!
0"
0%
0&
0-
0.
02
#8330000000
1!
1%
0+
1-
0/
00
01
12
03
#8340000000
0!
0%
0-
02
#8350000000
1!
1%
1-
12
#8360000000
0!
0%
b1 *
0-
02
b1 6
#8370000000
1!
1%
1-
12
#8380000000
0!
0%
b10 *
0-
02
b10 6
#8390000000
1!
1%
1-
12
#8400000000
0!
0%
b11 *
0-
02
b11 6
#8410000000
1!
1%
1-
12
15
#8420000000
0!
0%
b100 *
0-
02
b100 6
#8430000000
1!
1%
1-
12
#8440000000
0!
0%
b101 *
0-
02
b101 6
#8450000000
1!
1%
1-
12
#8460000000
0!
0%
b110 *
0-
02
b110 6
#8470000000
1!
1%
1-
12
#8480000000
0!
0%
b111 *
0-
02
b111 6
#8490000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#8500000000
0!
0%
b0 *
0-
02
b0 6
#8510000000
1!
1%
1-
12
#8520000000
0!
0%
b1 *
0-
02
b1 6
#8530000000
1!
1%
1-
12
#8540000000
0!
0%
b10 *
0-
02
b10 6
#8550000000
1!
1%
1-
12
#8560000000
0!
0%
b11 *
0-
02
b11 6
#8570000000
1!
1%
1-
12
15
#8580000000
0!
0%
b100 *
0-
02
b100 6
#8590000000
1!
1%
1-
12
#8600000000
0!
0%
b101 *
0-
02
b101 6
#8610000000
1!
1%
1-
12
#8620000000
0!
0%
b110 *
0-
02
b110 6
#8630000000
1!
1%
1-
12
#8640000000
0!
0%
b111 *
0-
02
b111 6
#8650000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#8660000000
0!
0%
b0 *
0-
02
b0 6
#8670000000
1!
1%
1-
12
#8680000000
0!
0%
b1 *
0-
02
b1 6
#8690000000
1!
1%
1-
12
#8700000000
0!
0%
b10 *
0-
02
b10 6
#8710000000
1!
1%
1-
12
#8720000000
0!
0%
b11 *
0-
02
b11 6
#8730000000
1!
1%
1-
12
15
#8740000000
0!
0%
b100 *
0-
02
b100 6
#8750000000
1!
1%
1-
12
#8760000000
0!
0%
b101 *
0-
02
b101 6
#8770000000
1!
1%
1-
12
#8780000000
0!
0%
b110 *
0-
02
b110 6
#8790000000
1!
1%
1-
12
#8800000000
0!
0%
b111 *
0-
02
b111 6
#8810000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#8820000000
0!
0%
b0 *
0-
02
b0 6
#8830000000
1!
1%
1-
12
#8840000000
0!
0%
b1 *
0-
02
b1 6
#8850000000
1!
1%
1-
12
#8860000000
0!
0%
b10 *
0-
02
b10 6
#8870000000
1!
1%
1-
12
#8880000000
0!
0%
b11 *
0-
02
b11 6
#8890000000
1!
1%
1-
12
15
#8900000000
0!
0%
b100 *
0-
02
b100 6
#8910000000
1!
1%
1-
12
#8920000000
0!
0%
b101 *
0-
02
b101 6
#8930000000
1!
1%
1-
12
#8940000000
0!
0%
b110 *
0-
02
b110 6
#8950000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#8960000000
0!
0%
b111 *
0-
02
b111 6
#8970000000
1!
1%
1-
12
05
#8980000000
0!
0%
b0 *
0-
02
b0 6
#8990000000
1!
1%
1-
12
#9000000000
0!
0"
0%
0&
0-
0.
02
#9010000000
1!
1%
0+
1-
0/
00
01
12
03
#9020000000
0!
0%
0-
02
#9030000000
1!
1%
1-
12
#9040000000
0!
0%
b1 *
0-
02
b1 6
#9050000000
1!
1%
1-
12
#9060000000
0!
0%
b10 *
0-
02
b10 6
#9070000000
1!
1%
1-
12
#9080000000
0!
0%
b11 *
0-
02
b11 6
#9090000000
1!
1%
1-
12
15
#9100000000
0!
0%
b100 *
0-
02
b100 6
#9110000000
1!
1%
1-
12
#9120000000
0!
0%
b101 *
0-
02
b101 6
#9130000000
1!
1%
1-
12
#9140000000
0!
0%
b110 *
0-
02
b110 6
#9150000000
1!
1%
1-
12
#9160000000
0!
0%
b111 *
0-
02
b111 6
#9170000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#9180000000
0!
0%
b0 *
0-
02
b0 6
#9190000000
1!
1%
1-
12
#9200000000
0!
0%
b1 *
0-
02
b1 6
#9210000000
1!
1%
1-
12
#9220000000
0!
0%
b10 *
0-
02
b10 6
#9230000000
1!
1%
1-
12
#9240000000
0!
0%
b11 *
0-
02
b11 6
#9250000000
1!
1%
1-
12
15
#9260000000
0!
0%
b100 *
0-
02
b100 6
#9270000000
1!
1%
1-
12
#9280000000
0!
0%
b101 *
0-
02
b101 6
#9290000000
1!
1%
1-
12
#9300000000
0!
0%
b110 *
0-
02
b110 6
#9310000000
1!
1%
1-
12
#9320000000
0!
0%
b111 *
0-
02
b111 6
#9330000000
1!
bXX1X #
b1111001 $
1%
bXX1X '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
X9
b1111001 :
b0011 ;
1<
b1111001 =
b0011 >
X?
b1111001 @
b0011 A
XB
#9340000000
0!
0%
b0 *
0-
02
b0 6
#9350000000
1!
1%
1-
12
#9360000000
0!
0%
b1 *
0-
02
b1 6
#9370000000
1!
1%
1-
12
#9380000000
0!
0%
b10 *
0-
02
b10 6
#9390000000
1!
1%
1-
12
#9400000000
0!
0%
b11 *
0-
02
b11 6
#9410000000
1!
1%
1-
12
15
#9420000000
0!
0%
b100 *
0-
02
b100 6
#9430000000
1!
1%
1-
12
#9440000000
0!
0%
b101 *
0-
02
b101 6
#9450000000
1!
1%
1-
12
#9460000000
0!
0%
b110 *
0-
02
b110 6
#9470000000
1!
1%
1-
12
#9480000000
0!
0%
b111 *
0-
02
b111 6
#9490000000
1!
bXXX1 #
b0110011 $
1%
bXXX1 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
19
b0110011 :
b0100 ;
X<
b0110011 =
b0100 >
X?
b0110011 @
b0100 A
XB
#9500000000
0!
0%
b0 *
0-
02
b0 6
#9510000000
1!
1%
1-
12
#9520000000
0!
0%
b1 *
0-
02
b1 6
#9530000000
1!
1%
1-
12
#9540000000
0!
0%
b10 *
0-
02
b10 6
#9550000000
1!
1%
1-
12
#9560000000
0!
0%
b11 *
0-
02
b11 6
#9570000000
1!
1%
1-
12
15
#9580000000
0!
0%
b100 *
0-
02
b100 6
#9590000000
1!
1%
1-
12
#9600000000
0!
0%
b101 *
0-
02
b101 6
#9610000000
1!
1%
1-
12
#9620000000
0!
0%
b110 *
0-
02
b110 6
#9630000000
1!
1"
b1XXX #
b0110000 $
1%
1&
b1XXX '
b0110000 (
b0001 )
1+
1-
1.
1/
10
11
12
13
b0110000 7
b0001 8
X9
b0110000 :
b0001 ;
X<
b0110000 =
b0001 >
X?
b0110000 @
b0001 A
1B
#9640000000
0!
0%
b111 *
0-
02
b111 6
#9650000000
1!
1%
1-
12
05
#9660000000
0!
0%
b0 *
0-
02
b0 6
#9670000000
1!
1%
1-
12
#9680000000
0!
0"
0%
0&
0-
0.
02
#9690000000
1!
1%
0+
1-
0/
00
01
12
03
#9700000000
0!
0%
0-
02
#9710000000
1!
1%
1-
12
#9720000000
0!
0%
b1 *
0-
02
b1 6
#9730000000
1!
1%
1-
12
#9740000000
0!
0%
b10 *
0-
02
b10 6
#9750000000
1!
1%
1-
12
#9760000000
0!
0%
b11 *
0-
02
b11 6
#9770000000
1!
1%
1-
12
15
#9780000000
0!
0%
b100 *
0-
02
b100 6
#9790000000
1!
1%
1-
12
#9800000000
0!
0%
b101 *
0-
02
b101 6
#9810000000
1!
1%
1-
12
#9820000000
0!
0%
b110 *
0-
02
b110 6
#9830000000
1!
1%
1-
12
#9840000000
0!
0%
b111 *
0-
02
b111 6
#9850000000
1!
bX1XX #
b1101101 $
1%
bX1XX '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
X9
b1101101 :
b0010 ;
X<
b1101101 =
b0010 >
1?
b1101101 @
b0010 A
XB
#9860000000
0!
0%
b0 *
0-
02
b0 6
#9870000000
1!
1%
1-
12
#9880000000
0!
0%
b1 *
0-
02
b1 6
#9890000000
1!
1%
1-
12
#9900000000
0!
0%
b10 *
0-
02
b10 6
#9910000000
1!
1%
1-
12
#9920000000
0!
0%
b11 *
0-
02
b11 6
#9930000000
1!
1%
1-
12
15
#9940000000
0!
0%
b100 *
0-
02
b100 6
#9950000000
1!
1%
1-
12
#9960000000
0!
0%
b101 *
0-
02
b101 6
#9970000000
1!
1%
1-
12
#9980000000
0!
0%
b110 *
0-
02
b110 6
#9990000000
1!
1%
1-
12
#10000000000
0!
0%
b111 *
0-
02
b111 6
